
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LSU(
  input          clock,
                 reset,
  output         request_ready,
  input          request_valid,
  input  [2:0]   request_bits_instructionInformation_nf,
  input          request_bits_instructionInformation_mew,
  input  [1:0]   request_bits_instructionInformation_mop,
  input  [4:0]   request_bits_instructionInformation_lumop,
  input  [1:0]   request_bits_instructionInformation_eew,
  input  [4:0]   request_bits_instructionInformation_vs3,
  input          request_bits_instructionInformation_isStore,
                 request_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  request_bits_rs1Data,
                 request_bits_rs2Data,
  input  [2:0]   request_bits_instructionIndex,
  input          v0UpdateVec_0_valid,
  input  [31:0]  v0UpdateVec_0_bits_data,
  input  [7:0]   v0UpdateVec_0_bits_offset,
  input  [3:0]   v0UpdateVec_0_bits_mask,
  input          v0UpdateVec_1_valid,
  input  [31:0]  v0UpdateVec_1_bits_data,
  input  [7:0]   v0UpdateVec_1_bits_offset,
  input  [3:0]   v0UpdateVec_1_bits_mask,
  input          v0UpdateVec_2_valid,
  input  [31:0]  v0UpdateVec_2_bits_data,
  input  [7:0]   v0UpdateVec_2_bits_offset,
  input  [3:0]   v0UpdateVec_2_bits_mask,
  input          v0UpdateVec_3_valid,
  input  [31:0]  v0UpdateVec_3_bits_data,
  input  [7:0]   v0UpdateVec_3_bits_offset,
  input  [3:0]   v0UpdateVec_3_bits_mask,
  input          axi4Port_aw_ready,
  output         axi4Port_aw_valid,
  output [1:0]   axi4Port_aw_bits_id,
  output [31:0]  axi4Port_aw_bits_addr,
  input          axi4Port_w_ready,
  output         axi4Port_w_valid,
  output [127:0] axi4Port_w_bits_data,
  output [15:0]  axi4Port_w_bits_strb,
  input          axi4Port_b_valid,
  input  [1:0]   axi4Port_b_bits_id,
                 axi4Port_b_bits_resp,
  input          axi4Port_ar_ready,
  output         axi4Port_ar_valid,
  output [31:0]  axi4Port_ar_bits_addr,
  output         axi4Port_r_ready,
  input          axi4Port_r_valid,
  input  [1:0]   axi4Port_r_bits_id,
  input  [127:0] axi4Port_r_bits_data,
  input  [1:0]   axi4Port_r_bits_resp,
  input          axi4Port_r_bits_last,
                 simpleAccessPorts_aw_ready,
  output         simpleAccessPorts_aw_valid,
  output [1:0]   simpleAccessPorts_aw_bits_id,
  output [31:0]  simpleAccessPorts_aw_bits_addr,
  output [2:0]   simpleAccessPorts_aw_bits_size,
  input          simpleAccessPorts_w_ready,
  output         simpleAccessPorts_w_valid,
  output [31:0]  simpleAccessPorts_w_bits_data,
  output [3:0]   simpleAccessPorts_w_bits_strb,
  input          simpleAccessPorts_b_valid,
  input  [1:0]   simpleAccessPorts_b_bits_id,
                 simpleAccessPorts_b_bits_resp,
  input          simpleAccessPorts_ar_ready,
  output         simpleAccessPorts_ar_valid,
  output [31:0]  simpleAccessPorts_ar_bits_addr,
  output         simpleAccessPorts_r_ready,
  input          simpleAccessPorts_r_valid,
  input  [1:0]   simpleAccessPorts_r_bits_id,
  input  [31:0]  simpleAccessPorts_r_bits_data,
  input  [1:0]   simpleAccessPorts_r_bits_resp,
  input          simpleAccessPorts_r_bits_last,
                 vrfReadDataPorts_0_ready,
  output         vrfReadDataPorts_0_valid,
  output [4:0]   vrfReadDataPorts_0_bits_vs,
  output [7:0]   vrfReadDataPorts_0_bits_offset,
  output [2:0]   vrfReadDataPorts_0_bits_instructionIndex,
  input          vrfReadDataPorts_1_ready,
  output         vrfReadDataPorts_1_valid,
  output [4:0]   vrfReadDataPorts_1_bits_vs,
  output [7:0]   vrfReadDataPorts_1_bits_offset,
  output [2:0]   vrfReadDataPorts_1_bits_instructionIndex,
  input          vrfReadDataPorts_2_ready,
  output         vrfReadDataPorts_2_valid,
  output [4:0]   vrfReadDataPorts_2_bits_vs,
  output [7:0]   vrfReadDataPorts_2_bits_offset,
  output [2:0]   vrfReadDataPorts_2_bits_instructionIndex,
  input          vrfReadDataPorts_3_ready,
  output         vrfReadDataPorts_3_valid,
  output [4:0]   vrfReadDataPorts_3_bits_vs,
  output [7:0]   vrfReadDataPorts_3_bits_offset,
  output [2:0]   vrfReadDataPorts_3_bits_instructionIndex,
  input          vrfReadResults_0_valid,
  input  [31:0]  vrfReadResults_0_bits,
  input          vrfReadResults_1_valid,
  input  [31:0]  vrfReadResults_1_bits,
  input          vrfReadResults_2_valid,
  input  [31:0]  vrfReadResults_2_bits,
  input          vrfReadResults_3_valid,
  input  [31:0]  vrfReadResults_3_bits,
  input          vrfWritePort_0_ready,
  output         vrfWritePort_0_valid,
  output [4:0]   vrfWritePort_0_bits_vd,
  output [7:0]   vrfWritePort_0_bits_offset,
  output [3:0]   vrfWritePort_0_bits_mask,
  output [31:0]  vrfWritePort_0_bits_data,
  output         vrfWritePort_0_bits_last,
  output [2:0]   vrfWritePort_0_bits_instructionIndex,
  input          vrfWritePort_1_ready,
  output         vrfWritePort_1_valid,
  output [4:0]   vrfWritePort_1_bits_vd,
  output [7:0]   vrfWritePort_1_bits_offset,
  output [3:0]   vrfWritePort_1_bits_mask,
  output [31:0]  vrfWritePort_1_bits_data,
  output         vrfWritePort_1_bits_last,
  output [2:0]   vrfWritePort_1_bits_instructionIndex,
  input          vrfWritePort_2_ready,
  output         vrfWritePort_2_valid,
  output [4:0]   vrfWritePort_2_bits_vd,
  output [7:0]   vrfWritePort_2_bits_offset,
  output [3:0]   vrfWritePort_2_bits_mask,
  output [31:0]  vrfWritePort_2_bits_data,
  output         vrfWritePort_2_bits_last,
  output [2:0]   vrfWritePort_2_bits_instructionIndex,
  input          vrfWritePort_3_ready,
  output         vrfWritePort_3_valid,
  output [4:0]   vrfWritePort_3_bits_vd,
  output [7:0]   vrfWritePort_3_bits_offset,
  output [3:0]   vrfWritePort_3_bits_mask,
  output [31:0]  vrfWritePort_3_bits_data,
  output         vrfWritePort_3_bits_last,
  output [2:0]   vrfWritePort_3_bits_instructionIndex,
  input          writeRelease_0,
                 writeRelease_1,
                 writeRelease_2,
                 writeRelease_3,
  output [7:0]   dataInWriteQueue_0,
                 dataInWriteQueue_1,
                 dataInWriteQueue_2,
                 dataInWriteQueue_3,
  input  [15:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
                 offsetReadResult_0_valid,
  input  [31:0]  offsetReadResult_0_bits,
  input          offsetReadResult_1_valid,
  input  [31:0]  offsetReadResult_1_bits,
  input          offsetReadResult_2_valid,
  input  [31:0]  offsetReadResult_2_bits,
  input          offsetReadResult_3_valid,
  input  [31:0]  offsetReadResult_3_bits,
  output [7:0]   lastReport,
  output [3:0]   tokenIO_offsetGroupRelease
);

  wire                _simpleDataQueue_fifo_empty;
  wire                _simpleDataQueue_fifo_full;
  wire                _simpleDataQueue_fifo_error;
  wire [77:0]         _simpleDataQueue_fifo_data_out;
  wire                _simpleSourceQueue_fifo_empty;
  wire                _simpleSourceQueue_fifo_full;
  wire                _simpleSourceQueue_fifo_error;
  wire                _dataQueue_fifo_empty;
  wire                _dataQueue_fifo_full;
  wire                _dataQueue_fifo_error;
  wire [187:0]        _dataQueue_fifo_data_out;
  wire                _sourceQueue_fifo_empty;
  wire                _sourceQueue_fifo_full;
  wire                _sourceQueue_fifo_error;
  wire                _writeIndexQueue_fifo_3_empty;
  wire                _writeIndexQueue_fifo_3_full;
  wire                _writeIndexQueue_fifo_3_error;
  wire                _writeIndexQueue_fifo_2_empty;
  wire                _writeIndexQueue_fifo_2_full;
  wire                _writeIndexQueue_fifo_2_error;
  wire                _writeIndexQueue_fifo_1_empty;
  wire                _writeIndexQueue_fifo_1_full;
  wire                _writeIndexQueue_fifo_1_error;
  wire                _writeIndexQueue_fifo_empty;
  wire                _writeIndexQueue_fifo_full;
  wire                _writeIndexQueue_fifo_error;
  wire                _otherUnitDataQueueVec_fifo_3_empty;
  wire                _otherUnitDataQueueVec_fifo_3_full;
  wire                _otherUnitDataQueueVec_fifo_3_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_3_data_out;
  wire                _otherUnitDataQueueVec_fifo_2_empty;
  wire                _otherUnitDataQueueVec_fifo_2_full;
  wire                _otherUnitDataQueueVec_fifo_2_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_2_data_out;
  wire                _otherUnitDataQueueVec_fifo_1_empty;
  wire                _otherUnitDataQueueVec_fifo_1_full;
  wire                _otherUnitDataQueueVec_fifo_1_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_1_data_out;
  wire                _otherUnitDataQueueVec_fifo_empty;
  wire                _otherUnitDataQueueVec_fifo_full;
  wire                _otherUnitDataQueueVec_fifo_error;
  wire [31:0]         _otherUnitDataQueueVec_fifo_data_out;
  wire                _otherUnitTargetQueue_fifo_empty;
  wire                _otherUnitTargetQueue_fifo_full;
  wire                _otherUnitTargetQueue_fifo_error;
  wire                _writeQueueVec_fifo_3_empty;
  wire                _writeQueueVec_fifo_3_full;
  wire                _writeQueueVec_fifo_3_error;
  wire [56:0]         _writeQueueVec_fifo_3_data_out;
  wire                _writeQueueVec_fifo_2_empty;
  wire                _writeQueueVec_fifo_2_full;
  wire                _writeQueueVec_fifo_2_error;
  wire [56:0]         _writeQueueVec_fifo_2_data_out;
  wire                _writeQueueVec_fifo_1_empty;
  wire                _writeQueueVec_fifo_1_full;
  wire                _writeQueueVec_fifo_1_error;
  wire [56:0]         _writeQueueVec_fifo_1_data_out;
  wire                _writeQueueVec_fifo_empty;
  wire                _writeQueueVec_fifo_full;
  wire                _writeQueueVec_fifo_error;
  wire [56:0]         _writeQueueVec_fifo_data_out;
  wire                _otherUnit_vrfReadDataPorts_valid;
  wire [4:0]          _otherUnit_vrfReadDataPorts_bits_vs;
  wire [7:0]          _otherUnit_vrfReadDataPorts_bits_offset;
  wire [2:0]          _otherUnit_vrfReadDataPorts_bits_instructionIndex;
  wire                _otherUnit_maskSelect_valid;
  wire [10:0]         _otherUnit_maskSelect_bits;
  wire                _otherUnit_memReadRequest_valid;
  wire                _otherUnit_memWriteRequest_valid;
  wire [7:0]          _otherUnit_memWriteRequest_bits_source;
  wire [31:0]         _otherUnit_memWriteRequest_bits_address;
  wire [1:0]          _otherUnit_memWriteRequest_bits_size;
  wire                _otherUnit_vrfWritePort_valid;
  wire [4:0]          _otherUnit_vrfWritePort_bits_vd;
  wire [7:0]          _otherUnit_vrfWritePort_bits_offset;
  wire [3:0]          _otherUnit_vrfWritePort_bits_mask;
  wire [31:0]         _otherUnit_vrfWritePort_bits_data;
  wire                _otherUnit_vrfWritePort_bits_last;
  wire [2:0]          _otherUnit_vrfWritePort_bits_instructionIndex;
  wire                _otherUnit_status_idle;
  wire                _otherUnit_status_last;
  wire [2:0]          _otherUnit_status_instructionIndex;
  wire [3:0]          _otherUnit_status_targetLane;
  wire                _otherUnit_status_isStore;
  wire                _otherUnit_offsetRelease_0;
  wire                _otherUnit_offsetRelease_1;
  wire                _otherUnit_offsetRelease_2;
  wire                _otherUnit_offsetRelease_3;
  wire                _storeUnit_maskSelect_valid;
  wire [10:0]         _storeUnit_maskSelect_bits;
  wire                _storeUnit_memRequest_valid;
  wire [11:0]         _storeUnit_memRequest_bits_index;
  wire [31:0]         _storeUnit_memRequest_bits_address;
  wire                _storeUnit_status_idle;
  wire                _storeUnit_status_last;
  wire [2:0]          _storeUnit_status_instructionIndex;
  wire [31:0]         _storeUnit_status_startAddress;
  wire [31:0]         _storeUnit_status_endAddress;
  wire                _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [7:0]          _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire                _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [7:0]          _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  wire                _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [7:0]          _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  wire                _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]          _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [7:0]          _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]          _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  wire                _loadUnit_maskSelect_valid;
  wire [10:0]         _loadUnit_maskSelect_bits;
  wire                _loadUnit_memRequest_valid;
  wire                _loadUnit_status_idle;
  wire                _loadUnit_status_last;
  wire [2:0]          _loadUnit_status_instructionIndex;
  wire [31:0]         _loadUnit_status_startAddress;
  wire [31:0]         _loadUnit_status_endAddress;
  wire                _loadUnit_vrfWritePort_0_valid;
  wire [4:0]          _loadUnit_vrfWritePort_0_bits_vd;
  wire [7:0]          _loadUnit_vrfWritePort_0_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_0_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_0_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_0_bits_instructionIndex;
  wire                _loadUnit_vrfWritePort_1_valid;
  wire [4:0]          _loadUnit_vrfWritePort_1_bits_vd;
  wire [7:0]          _loadUnit_vrfWritePort_1_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_1_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_1_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_1_bits_instructionIndex;
  wire                _loadUnit_vrfWritePort_2_valid;
  wire [4:0]          _loadUnit_vrfWritePort_2_bits_vd;
  wire [7:0]          _loadUnit_vrfWritePort_2_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_2_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_2_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_2_bits_instructionIndex;
  wire                _loadUnit_vrfWritePort_3_valid;
  wire [4:0]          _loadUnit_vrfWritePort_3_bits_vd;
  wire [7:0]          _loadUnit_vrfWritePort_3_bits_offset;
  wire [3:0]          _loadUnit_vrfWritePort_3_bits_mask;
  wire [31:0]         _loadUnit_vrfWritePort_3_bits_data;
  wire [2:0]          _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire                simpleDataQueue_almostFull;
  wire                simpleDataQueue_almostEmpty;
  wire                simpleSourceQueue_almostFull;
  wire                simpleSourceQueue_almostEmpty;
  wire                dataQueue_almostFull;
  wire                dataQueue_almostEmpty;
  wire                sourceQueue_almostFull;
  wire                sourceQueue_almostEmpty;
  wire                writeIndexQueue_3_almostFull;
  wire                writeIndexQueue_3_almostEmpty;
  wire                writeIndexQueue_2_almostFull;
  wire                writeIndexQueue_2_almostEmpty;
  wire                writeIndexQueue_1_almostFull;
  wire                writeIndexQueue_1_almostEmpty;
  wire                writeIndexQueue_almostFull;
  wire                writeIndexQueue_almostEmpty;
  wire                otherUnitDataQueueVec_3_almostFull;
  wire                otherUnitDataQueueVec_3_almostEmpty;
  wire                otherUnitDataQueueVec_2_almostFull;
  wire                otherUnitDataQueueVec_2_almostEmpty;
  wire                otherUnitDataQueueVec_1_almostFull;
  wire                otherUnitDataQueueVec_1_almostEmpty;
  wire                otherUnitDataQueueVec_0_almostFull;
  wire                otherUnitDataQueueVec_0_almostEmpty;
  wire                otherUnitTargetQueue_almostFull;
  wire                otherUnitTargetQueue_almostEmpty;
  wire                writeQueueVec_3_almostFull;
  wire                writeQueueVec_3_almostEmpty;
  wire                writeQueueVec_2_almostFull;
  wire                writeQueueVec_2_almostEmpty;
  wire                writeQueueVec_1_almostFull;
  wire                writeQueueVec_1_almostEmpty;
  wire                writeQueueVec_0_almostFull;
  wire                writeQueueVec_0_almostEmpty;
  wire [6:0]          simpleSourceQueue_enq_bits;
  wire [31:0]         simpleAccessPorts_ar_bits_addr_0;
  wire [11:0]         sourceQueue_enq_bits;
  wire [31:0]         axi4Port_ar_bits_addr_0;
  wire                request_valid_0 = request_valid;
  wire [2:0]          request_bits_instructionInformation_nf_0 = request_bits_instructionInformation_nf;
  wire                request_bits_instructionInformation_mew_0 = request_bits_instructionInformation_mew;
  wire [1:0]          request_bits_instructionInformation_mop_0 = request_bits_instructionInformation_mop;
  wire [4:0]          request_bits_instructionInformation_lumop_0 = request_bits_instructionInformation_lumop;
  wire [1:0]          request_bits_instructionInformation_eew_0 = request_bits_instructionInformation_eew;
  wire [4:0]          request_bits_instructionInformation_vs3_0 = request_bits_instructionInformation_vs3;
  wire                request_bits_instructionInformation_isStore_0 = request_bits_instructionInformation_isStore;
  wire                request_bits_instructionInformation_maskedLoadStore_0 = request_bits_instructionInformation_maskedLoadStore;
  wire [31:0]         request_bits_rs1Data_0 = request_bits_rs1Data;
  wire [31:0]         request_bits_rs2Data_0 = request_bits_rs2Data;
  wire [2:0]          request_bits_instructionIndex_0 = request_bits_instructionIndex;
  wire                axi4Port_aw_ready_0 = axi4Port_aw_ready;
  wire                axi4Port_w_ready_0 = axi4Port_w_ready;
  wire                axi4Port_b_valid_0 = axi4Port_b_valid;
  wire [1:0]          axi4Port_b_bits_id_0 = axi4Port_b_bits_id;
  wire [1:0]          axi4Port_b_bits_resp_0 = axi4Port_b_bits_resp;
  wire                axi4Port_ar_ready_0 = axi4Port_ar_ready;
  wire                axi4Port_r_valid_0 = axi4Port_r_valid;
  wire [1:0]          axi4Port_r_bits_id_0 = axi4Port_r_bits_id;
  wire [127:0]        axi4Port_r_bits_data_0 = axi4Port_r_bits_data;
  wire [1:0]          axi4Port_r_bits_resp_0 = axi4Port_r_bits_resp;
  wire                axi4Port_r_bits_last_0 = axi4Port_r_bits_last;
  wire                simpleAccessPorts_aw_ready_0 = simpleAccessPorts_aw_ready;
  wire                simpleAccessPorts_w_ready_0 = simpleAccessPorts_w_ready;
  wire                simpleAccessPorts_b_valid_0 = simpleAccessPorts_b_valid;
  wire [1:0]          simpleAccessPorts_b_bits_id_0 = simpleAccessPorts_b_bits_id;
  wire [1:0]          simpleAccessPorts_b_bits_resp_0 = simpleAccessPorts_b_bits_resp;
  wire                simpleAccessPorts_ar_ready_0 = simpleAccessPorts_ar_ready;
  wire                simpleAccessPorts_r_valid_0 = simpleAccessPorts_r_valid;
  wire [1:0]          simpleAccessPorts_r_bits_id_0 = simpleAccessPorts_r_bits_id;
  wire [31:0]         simpleAccessPorts_r_bits_data_0 = simpleAccessPorts_r_bits_data;
  wire [1:0]          simpleAccessPorts_r_bits_resp_0 = simpleAccessPorts_r_bits_resp;
  wire                simpleAccessPorts_r_bits_last_0 = simpleAccessPorts_r_bits_last;
  wire                vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire                vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire                vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire                vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire                vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire                vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire                vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire                vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire [31:0]         otherUnitDataQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire [31:0]         otherUnitDataQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire [31:0]         otherUnitDataQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire [31:0]         otherUnitDataQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire                writeIndexQueue_deq_ready = writeRelease_0;
  wire                writeIndexQueue_1_deq_ready = writeRelease_1;
  wire                writeIndexQueue_2_deq_ready = writeRelease_2;
  wire                writeIndexQueue_3_deq_ready = writeRelease_3;
  wire [1:0]          vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]          vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]          vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]          vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]          axi4Port_ar_bits_id = 2'h0;
  wire [1:0]          simpleAccessPorts_ar_bits_id = 2'h0;
  wire [1:0]          axi4Port_aw_bits_burst = 2'h1;
  wire [1:0]          axi4Port_ar_bits_burst = 2'h1;
  wire [1:0]          simpleAccessPorts_aw_bits_burst = 2'h1;
  wire [1:0]          simpleAccessPorts_ar_bits_burst = 2'h1;
  wire [3:0]          writeQueueVec_0_enq_bits_targetLane = 4'h1;
  wire [3:0]          writeQueueVec_1_enq_bits_targetLane = 4'h2;
  wire [3:0]          writeQueueVec_2_enq_bits_targetLane = 4'h4;
  wire [3:0]          writeQueueVec_3_enq_bits_targetLane = 4'h8;
  wire [7:0]          axi4Port_aw_bits_len = 8'h0;
  wire [7:0]          axi4Port_ar_bits_len = 8'h0;
  wire [7:0]          simpleAccessPorts_aw_bits_len = 8'h0;
  wire [7:0]          simpleAccessPorts_ar_bits_len = 8'h0;
  wire [2:0]          axi4Port_aw_bits_size = 3'h4;
  wire [2:0]          axi4Port_ar_bits_size = 3'h4;
  wire                axi4Port_aw_bits_lock = 1'h0;
  wire                axi4Port_ar_bits_lock = 1'h0;
  wire                simpleAccessPorts_aw_bits_lock = 1'h0;
  wire                simpleAccessPorts_ar_bits_lock = 1'h0;
  wire [3:0]          axi4Port_aw_bits_cache = 4'h0;
  wire [3:0]          axi4Port_aw_bits_qos = 4'h0;
  wire [3:0]          axi4Port_aw_bits_region = 4'h0;
  wire [3:0]          axi4Port_ar_bits_cache = 4'h0;
  wire [3:0]          axi4Port_ar_bits_qos = 4'h0;
  wire [3:0]          axi4Port_ar_bits_region = 4'h0;
  wire [3:0]          simpleAccessPorts_aw_bits_cache = 4'h0;
  wire [3:0]          simpleAccessPorts_aw_bits_qos = 4'h0;
  wire [3:0]          simpleAccessPorts_aw_bits_region = 4'h0;
  wire [3:0]          simpleAccessPorts_ar_bits_cache = 4'h0;
  wire [3:0]          simpleAccessPorts_ar_bits_qos = 4'h0;
  wire [3:0]          simpleAccessPorts_ar_bits_region = 4'h0;
  wire [2:0]          axi4Port_aw_bits_prot = 3'h0;
  wire [2:0]          axi4Port_ar_bits_prot = 3'h0;
  wire [2:0]          simpleAccessPorts_aw_bits_prot = 3'h0;
  wire [2:0]          simpleAccessPorts_ar_bits_prot = 3'h0;
  wire                axi4Port_w_bits_last = 1'h1;
  wire                axi4Port_b_ready = 1'h1;
  wire                simpleAccessPorts_w_bits_last = 1'h1;
  wire                simpleAccessPorts_b_ready = 1'h1;
  wire [2:0]          simpleAccessPorts_ar_bits_size = 3'h2;
  wire                dataQueue_deq_ready = axi4Port_w_ready_0;
  wire                dataQueue_deq_valid;
  wire [127:0]        dataQueue_deq_bits_data;
  wire [15:0]         dataQueue_deq_bits_mask;
  wire                simpleDataQueue_deq_ready = simpleAccessPorts_w_ready_0;
  wire                simpleDataQueue_deq_valid;
  wire [31:0]         simpleDataQueue_deq_bits_data;
  wire [3:0]          simpleDataQueue_deq_bits_mask;
  wire                writeQueueVec_0_deq_ready = vrfWritePort_0_ready_0;
  wire                writeQueueVec_0_deq_valid;
  wire [4:0]          writeQueueVec_0_deq_bits_data_vd;
  wire [7:0]          writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_0_deq_bits_data_data;
  wire                writeQueueVec_0_deq_bits_data_last;
  wire [2:0]          writeQueueVec_0_deq_bits_data_instructionIndex;
  wire                writeQueueVec_1_deq_ready = vrfWritePort_1_ready_0;
  wire                writeQueueVec_1_deq_valid;
  wire [4:0]          writeQueueVec_1_deq_bits_data_vd;
  wire [7:0]          writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_1_deq_bits_data_data;
  wire                writeQueueVec_1_deq_bits_data_last;
  wire [2:0]          writeQueueVec_1_deq_bits_data_instructionIndex;
  wire                writeQueueVec_2_deq_ready = vrfWritePort_2_ready_0;
  wire                writeQueueVec_2_deq_valid;
  wire [4:0]          writeQueueVec_2_deq_bits_data_vd;
  wire [7:0]          writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_2_deq_bits_data_data;
  wire                writeQueueVec_2_deq_bits_data_last;
  wire [2:0]          writeQueueVec_2_deq_bits_data_instructionIndex;
  wire                writeQueueVec_3_deq_ready = vrfWritePort_3_ready_0;
  wire                writeQueueVec_3_deq_valid;
  wire [4:0]          writeQueueVec_3_deq_bits_data_vd;
  wire [7:0]          writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]          writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]         writeQueueVec_3_deq_bits_data_data;
  wire                writeQueueVec_3_deq_bits_data_last;
  wire [2:0]          writeQueueVec_3_deq_bits_data_instructionIndex;
  reg  [31:0]         v0_0;
  reg  [31:0]         v0_1;
  reg  [31:0]         v0_2;
  reg  [31:0]         v0_3;
  reg  [31:0]         v0_4;
  reg  [31:0]         v0_5;
  reg  [31:0]         v0_6;
  reg  [31:0]         v0_7;
  reg  [31:0]         v0_8;
  reg  [31:0]         v0_9;
  reg  [31:0]         v0_10;
  reg  [31:0]         v0_11;
  reg  [31:0]         v0_12;
  reg  [31:0]         v0_13;
  reg  [31:0]         v0_14;
  reg  [31:0]         v0_15;
  reg  [31:0]         v0_16;
  reg  [31:0]         v0_17;
  reg  [31:0]         v0_18;
  reg  [31:0]         v0_19;
  reg  [31:0]         v0_20;
  reg  [31:0]         v0_21;
  reg  [31:0]         v0_22;
  reg  [31:0]         v0_23;
  reg  [31:0]         v0_24;
  reg  [31:0]         v0_25;
  reg  [31:0]         v0_26;
  reg  [31:0]         v0_27;
  reg  [31:0]         v0_28;
  reg  [31:0]         v0_29;
  reg  [31:0]         v0_30;
  reg  [31:0]         v0_31;
  reg  [31:0]         v0_32;
  reg  [31:0]         v0_33;
  reg  [31:0]         v0_34;
  reg  [31:0]         v0_35;
  reg  [31:0]         v0_36;
  reg  [31:0]         v0_37;
  reg  [31:0]         v0_38;
  reg  [31:0]         v0_39;
  reg  [31:0]         v0_40;
  reg  [31:0]         v0_41;
  reg  [31:0]         v0_42;
  reg  [31:0]         v0_43;
  reg  [31:0]         v0_44;
  reg  [31:0]         v0_45;
  reg  [31:0]         v0_46;
  reg  [31:0]         v0_47;
  reg  [31:0]         v0_48;
  reg  [31:0]         v0_49;
  reg  [31:0]         v0_50;
  reg  [31:0]         v0_51;
  reg  [31:0]         v0_52;
  reg  [31:0]         v0_53;
  reg  [31:0]         v0_54;
  reg  [31:0]         v0_55;
  reg  [31:0]         v0_56;
  reg  [31:0]         v0_57;
  reg  [31:0]         v0_58;
  reg  [31:0]         v0_59;
  reg  [31:0]         v0_60;
  reg  [31:0]         v0_61;
  reg  [31:0]         v0_62;
  reg  [31:0]         v0_63;
  reg  [31:0]         v0_64;
  reg  [31:0]         v0_65;
  reg  [31:0]         v0_66;
  reg  [31:0]         v0_67;
  reg  [31:0]         v0_68;
  reg  [31:0]         v0_69;
  reg  [31:0]         v0_70;
  reg  [31:0]         v0_71;
  reg  [31:0]         v0_72;
  reg  [31:0]         v0_73;
  reg  [31:0]         v0_74;
  reg  [31:0]         v0_75;
  reg  [31:0]         v0_76;
  reg  [31:0]         v0_77;
  reg  [31:0]         v0_78;
  reg  [31:0]         v0_79;
  reg  [31:0]         v0_80;
  reg  [31:0]         v0_81;
  reg  [31:0]         v0_82;
  reg  [31:0]         v0_83;
  reg  [31:0]         v0_84;
  reg  [31:0]         v0_85;
  reg  [31:0]         v0_86;
  reg  [31:0]         v0_87;
  reg  [31:0]         v0_88;
  reg  [31:0]         v0_89;
  reg  [31:0]         v0_90;
  reg  [31:0]         v0_91;
  reg  [31:0]         v0_92;
  reg  [31:0]         v0_93;
  reg  [31:0]         v0_94;
  reg  [31:0]         v0_95;
  reg  [31:0]         v0_96;
  reg  [31:0]         v0_97;
  reg  [31:0]         v0_98;
  reg  [31:0]         v0_99;
  reg  [31:0]         v0_100;
  reg  [31:0]         v0_101;
  reg  [31:0]         v0_102;
  reg  [31:0]         v0_103;
  reg  [31:0]         v0_104;
  reg  [31:0]         v0_105;
  reg  [31:0]         v0_106;
  reg  [31:0]         v0_107;
  reg  [31:0]         v0_108;
  reg  [31:0]         v0_109;
  reg  [31:0]         v0_110;
  reg  [31:0]         v0_111;
  reg  [31:0]         v0_112;
  reg  [31:0]         v0_113;
  reg  [31:0]         v0_114;
  reg  [31:0]         v0_115;
  reg  [31:0]         v0_116;
  reg  [31:0]         v0_117;
  reg  [31:0]         v0_118;
  reg  [31:0]         v0_119;
  reg  [31:0]         v0_120;
  reg  [31:0]         v0_121;
  reg  [31:0]         v0_122;
  reg  [31:0]         v0_123;
  reg  [31:0]         v0_124;
  reg  [31:0]         v0_125;
  reg  [31:0]         v0_126;
  reg  [31:0]         v0_127;
  reg  [31:0]         v0_128;
  reg  [31:0]         v0_129;
  reg  [31:0]         v0_130;
  reg  [31:0]         v0_131;
  reg  [31:0]         v0_132;
  reg  [31:0]         v0_133;
  reg  [31:0]         v0_134;
  reg  [31:0]         v0_135;
  reg  [31:0]         v0_136;
  reg  [31:0]         v0_137;
  reg  [31:0]         v0_138;
  reg  [31:0]         v0_139;
  reg  [31:0]         v0_140;
  reg  [31:0]         v0_141;
  reg  [31:0]         v0_142;
  reg  [31:0]         v0_143;
  reg  [31:0]         v0_144;
  reg  [31:0]         v0_145;
  reg  [31:0]         v0_146;
  reg  [31:0]         v0_147;
  reg  [31:0]         v0_148;
  reg  [31:0]         v0_149;
  reg  [31:0]         v0_150;
  reg  [31:0]         v0_151;
  reg  [31:0]         v0_152;
  reg  [31:0]         v0_153;
  reg  [31:0]         v0_154;
  reg  [31:0]         v0_155;
  reg  [31:0]         v0_156;
  reg  [31:0]         v0_157;
  reg  [31:0]         v0_158;
  reg  [31:0]         v0_159;
  reg  [31:0]         v0_160;
  reg  [31:0]         v0_161;
  reg  [31:0]         v0_162;
  reg  [31:0]         v0_163;
  reg  [31:0]         v0_164;
  reg  [31:0]         v0_165;
  reg  [31:0]         v0_166;
  reg  [31:0]         v0_167;
  reg  [31:0]         v0_168;
  reg  [31:0]         v0_169;
  reg  [31:0]         v0_170;
  reg  [31:0]         v0_171;
  reg  [31:0]         v0_172;
  reg  [31:0]         v0_173;
  reg  [31:0]         v0_174;
  reg  [31:0]         v0_175;
  reg  [31:0]         v0_176;
  reg  [31:0]         v0_177;
  reg  [31:0]         v0_178;
  reg  [31:0]         v0_179;
  reg  [31:0]         v0_180;
  reg  [31:0]         v0_181;
  reg  [31:0]         v0_182;
  reg  [31:0]         v0_183;
  reg  [31:0]         v0_184;
  reg  [31:0]         v0_185;
  reg  [31:0]         v0_186;
  reg  [31:0]         v0_187;
  reg  [31:0]         v0_188;
  reg  [31:0]         v0_189;
  reg  [31:0]         v0_190;
  reg  [31:0]         v0_191;
  reg  [31:0]         v0_192;
  reg  [31:0]         v0_193;
  reg  [31:0]         v0_194;
  reg  [31:0]         v0_195;
  reg  [31:0]         v0_196;
  reg  [31:0]         v0_197;
  reg  [31:0]         v0_198;
  reg  [31:0]         v0_199;
  reg  [31:0]         v0_200;
  reg  [31:0]         v0_201;
  reg  [31:0]         v0_202;
  reg  [31:0]         v0_203;
  reg  [31:0]         v0_204;
  reg  [31:0]         v0_205;
  reg  [31:0]         v0_206;
  reg  [31:0]         v0_207;
  reg  [31:0]         v0_208;
  reg  [31:0]         v0_209;
  reg  [31:0]         v0_210;
  reg  [31:0]         v0_211;
  reg  [31:0]         v0_212;
  reg  [31:0]         v0_213;
  reg  [31:0]         v0_214;
  reg  [31:0]         v0_215;
  reg  [31:0]         v0_216;
  reg  [31:0]         v0_217;
  reg  [31:0]         v0_218;
  reg  [31:0]         v0_219;
  reg  [31:0]         v0_220;
  reg  [31:0]         v0_221;
  reg  [31:0]         v0_222;
  reg  [31:0]         v0_223;
  reg  [31:0]         v0_224;
  reg  [31:0]         v0_225;
  reg  [31:0]         v0_226;
  reg  [31:0]         v0_227;
  reg  [31:0]         v0_228;
  reg  [31:0]         v0_229;
  reg  [31:0]         v0_230;
  reg  [31:0]         v0_231;
  reg  [31:0]         v0_232;
  reg  [31:0]         v0_233;
  reg  [31:0]         v0_234;
  reg  [31:0]         v0_235;
  reg  [31:0]         v0_236;
  reg  [31:0]         v0_237;
  reg  [31:0]         v0_238;
  reg  [31:0]         v0_239;
  reg  [31:0]         v0_240;
  reg  [31:0]         v0_241;
  reg  [31:0]         v0_242;
  reg  [31:0]         v0_243;
  reg  [31:0]         v0_244;
  reg  [31:0]         v0_245;
  reg  [31:0]         v0_246;
  reg  [31:0]         v0_247;
  reg  [31:0]         v0_248;
  reg  [31:0]         v0_249;
  reg  [31:0]         v0_250;
  reg  [31:0]         v0_251;
  reg  [31:0]         v0_252;
  reg  [31:0]         v0_253;
  reg  [31:0]         v0_254;
  reg  [31:0]         v0_255;
  reg  [31:0]         v0_256;
  reg  [31:0]         v0_257;
  reg  [31:0]         v0_258;
  reg  [31:0]         v0_259;
  reg  [31:0]         v0_260;
  reg  [31:0]         v0_261;
  reg  [31:0]         v0_262;
  reg  [31:0]         v0_263;
  reg  [31:0]         v0_264;
  reg  [31:0]         v0_265;
  reg  [31:0]         v0_266;
  reg  [31:0]         v0_267;
  reg  [31:0]         v0_268;
  reg  [31:0]         v0_269;
  reg  [31:0]         v0_270;
  reg  [31:0]         v0_271;
  reg  [31:0]         v0_272;
  reg  [31:0]         v0_273;
  reg  [31:0]         v0_274;
  reg  [31:0]         v0_275;
  reg  [31:0]         v0_276;
  reg  [31:0]         v0_277;
  reg  [31:0]         v0_278;
  reg  [31:0]         v0_279;
  reg  [31:0]         v0_280;
  reg  [31:0]         v0_281;
  reg  [31:0]         v0_282;
  reg  [31:0]         v0_283;
  reg  [31:0]         v0_284;
  reg  [31:0]         v0_285;
  reg  [31:0]         v0_286;
  reg  [31:0]         v0_287;
  reg  [31:0]         v0_288;
  reg  [31:0]         v0_289;
  reg  [31:0]         v0_290;
  reg  [31:0]         v0_291;
  reg  [31:0]         v0_292;
  reg  [31:0]         v0_293;
  reg  [31:0]         v0_294;
  reg  [31:0]         v0_295;
  reg  [31:0]         v0_296;
  reg  [31:0]         v0_297;
  reg  [31:0]         v0_298;
  reg  [31:0]         v0_299;
  reg  [31:0]         v0_300;
  reg  [31:0]         v0_301;
  reg  [31:0]         v0_302;
  reg  [31:0]         v0_303;
  reg  [31:0]         v0_304;
  reg  [31:0]         v0_305;
  reg  [31:0]         v0_306;
  reg  [31:0]         v0_307;
  reg  [31:0]         v0_308;
  reg  [31:0]         v0_309;
  reg  [31:0]         v0_310;
  reg  [31:0]         v0_311;
  reg  [31:0]         v0_312;
  reg  [31:0]         v0_313;
  reg  [31:0]         v0_314;
  reg  [31:0]         v0_315;
  reg  [31:0]         v0_316;
  reg  [31:0]         v0_317;
  reg  [31:0]         v0_318;
  reg  [31:0]         v0_319;
  reg  [31:0]         v0_320;
  reg  [31:0]         v0_321;
  reg  [31:0]         v0_322;
  reg  [31:0]         v0_323;
  reg  [31:0]         v0_324;
  reg  [31:0]         v0_325;
  reg  [31:0]         v0_326;
  reg  [31:0]         v0_327;
  reg  [31:0]         v0_328;
  reg  [31:0]         v0_329;
  reg  [31:0]         v0_330;
  reg  [31:0]         v0_331;
  reg  [31:0]         v0_332;
  reg  [31:0]         v0_333;
  reg  [31:0]         v0_334;
  reg  [31:0]         v0_335;
  reg  [31:0]         v0_336;
  reg  [31:0]         v0_337;
  reg  [31:0]         v0_338;
  reg  [31:0]         v0_339;
  reg  [31:0]         v0_340;
  reg  [31:0]         v0_341;
  reg  [31:0]         v0_342;
  reg  [31:0]         v0_343;
  reg  [31:0]         v0_344;
  reg  [31:0]         v0_345;
  reg  [31:0]         v0_346;
  reg  [31:0]         v0_347;
  reg  [31:0]         v0_348;
  reg  [31:0]         v0_349;
  reg  [31:0]         v0_350;
  reg  [31:0]         v0_351;
  reg  [31:0]         v0_352;
  reg  [31:0]         v0_353;
  reg  [31:0]         v0_354;
  reg  [31:0]         v0_355;
  reg  [31:0]         v0_356;
  reg  [31:0]         v0_357;
  reg  [31:0]         v0_358;
  reg  [31:0]         v0_359;
  reg  [31:0]         v0_360;
  reg  [31:0]         v0_361;
  reg  [31:0]         v0_362;
  reg  [31:0]         v0_363;
  reg  [31:0]         v0_364;
  reg  [31:0]         v0_365;
  reg  [31:0]         v0_366;
  reg  [31:0]         v0_367;
  reg  [31:0]         v0_368;
  reg  [31:0]         v0_369;
  reg  [31:0]         v0_370;
  reg  [31:0]         v0_371;
  reg  [31:0]         v0_372;
  reg  [31:0]         v0_373;
  reg  [31:0]         v0_374;
  reg  [31:0]         v0_375;
  reg  [31:0]         v0_376;
  reg  [31:0]         v0_377;
  reg  [31:0]         v0_378;
  reg  [31:0]         v0_379;
  reg  [31:0]         v0_380;
  reg  [31:0]         v0_381;
  reg  [31:0]         v0_382;
  reg  [31:0]         v0_383;
  reg  [31:0]         v0_384;
  reg  [31:0]         v0_385;
  reg  [31:0]         v0_386;
  reg  [31:0]         v0_387;
  reg  [31:0]         v0_388;
  reg  [31:0]         v0_389;
  reg  [31:0]         v0_390;
  reg  [31:0]         v0_391;
  reg  [31:0]         v0_392;
  reg  [31:0]         v0_393;
  reg  [31:0]         v0_394;
  reg  [31:0]         v0_395;
  reg  [31:0]         v0_396;
  reg  [31:0]         v0_397;
  reg  [31:0]         v0_398;
  reg  [31:0]         v0_399;
  reg  [31:0]         v0_400;
  reg  [31:0]         v0_401;
  reg  [31:0]         v0_402;
  reg  [31:0]         v0_403;
  reg  [31:0]         v0_404;
  reg  [31:0]         v0_405;
  reg  [31:0]         v0_406;
  reg  [31:0]         v0_407;
  reg  [31:0]         v0_408;
  reg  [31:0]         v0_409;
  reg  [31:0]         v0_410;
  reg  [31:0]         v0_411;
  reg  [31:0]         v0_412;
  reg  [31:0]         v0_413;
  reg  [31:0]         v0_414;
  reg  [31:0]         v0_415;
  reg  [31:0]         v0_416;
  reg  [31:0]         v0_417;
  reg  [31:0]         v0_418;
  reg  [31:0]         v0_419;
  reg  [31:0]         v0_420;
  reg  [31:0]         v0_421;
  reg  [31:0]         v0_422;
  reg  [31:0]         v0_423;
  reg  [31:0]         v0_424;
  reg  [31:0]         v0_425;
  reg  [31:0]         v0_426;
  reg  [31:0]         v0_427;
  reg  [31:0]         v0_428;
  reg  [31:0]         v0_429;
  reg  [31:0]         v0_430;
  reg  [31:0]         v0_431;
  reg  [31:0]         v0_432;
  reg  [31:0]         v0_433;
  reg  [31:0]         v0_434;
  reg  [31:0]         v0_435;
  reg  [31:0]         v0_436;
  reg  [31:0]         v0_437;
  reg  [31:0]         v0_438;
  reg  [31:0]         v0_439;
  reg  [31:0]         v0_440;
  reg  [31:0]         v0_441;
  reg  [31:0]         v0_442;
  reg  [31:0]         v0_443;
  reg  [31:0]         v0_444;
  reg  [31:0]         v0_445;
  reg  [31:0]         v0_446;
  reg  [31:0]         v0_447;
  reg  [31:0]         v0_448;
  reg  [31:0]         v0_449;
  reg  [31:0]         v0_450;
  reg  [31:0]         v0_451;
  reg  [31:0]         v0_452;
  reg  [31:0]         v0_453;
  reg  [31:0]         v0_454;
  reg  [31:0]         v0_455;
  reg  [31:0]         v0_456;
  reg  [31:0]         v0_457;
  reg  [31:0]         v0_458;
  reg  [31:0]         v0_459;
  reg  [31:0]         v0_460;
  reg  [31:0]         v0_461;
  reg  [31:0]         v0_462;
  reg  [31:0]         v0_463;
  reg  [31:0]         v0_464;
  reg  [31:0]         v0_465;
  reg  [31:0]         v0_466;
  reg  [31:0]         v0_467;
  reg  [31:0]         v0_468;
  reg  [31:0]         v0_469;
  reg  [31:0]         v0_470;
  reg  [31:0]         v0_471;
  reg  [31:0]         v0_472;
  reg  [31:0]         v0_473;
  reg  [31:0]         v0_474;
  reg  [31:0]         v0_475;
  reg  [31:0]         v0_476;
  reg  [31:0]         v0_477;
  reg  [31:0]         v0_478;
  reg  [31:0]         v0_479;
  reg  [31:0]         v0_480;
  reg  [31:0]         v0_481;
  reg  [31:0]         v0_482;
  reg  [31:0]         v0_483;
  reg  [31:0]         v0_484;
  reg  [31:0]         v0_485;
  reg  [31:0]         v0_486;
  reg  [31:0]         v0_487;
  reg  [31:0]         v0_488;
  reg  [31:0]         v0_489;
  reg  [31:0]         v0_490;
  reg  [31:0]         v0_491;
  reg  [31:0]         v0_492;
  reg  [31:0]         v0_493;
  reg  [31:0]         v0_494;
  reg  [31:0]         v0_495;
  reg  [31:0]         v0_496;
  reg  [31:0]         v0_497;
  reg  [31:0]         v0_498;
  reg  [31:0]         v0_499;
  reg  [31:0]         v0_500;
  reg  [31:0]         v0_501;
  reg  [31:0]         v0_502;
  reg  [31:0]         v0_503;
  reg  [31:0]         v0_504;
  reg  [31:0]         v0_505;
  reg  [31:0]         v0_506;
  reg  [31:0]         v0_507;
  reg  [31:0]         v0_508;
  reg  [31:0]         v0_509;
  reg  [31:0]         v0_510;
  reg  [31:0]         v0_511;
  reg  [31:0]         v0_512;
  reg  [31:0]         v0_513;
  reg  [31:0]         v0_514;
  reg  [31:0]         v0_515;
  reg  [31:0]         v0_516;
  reg  [31:0]         v0_517;
  reg  [31:0]         v0_518;
  reg  [31:0]         v0_519;
  reg  [31:0]         v0_520;
  reg  [31:0]         v0_521;
  reg  [31:0]         v0_522;
  reg  [31:0]         v0_523;
  reg  [31:0]         v0_524;
  reg  [31:0]         v0_525;
  reg  [31:0]         v0_526;
  reg  [31:0]         v0_527;
  reg  [31:0]         v0_528;
  reg  [31:0]         v0_529;
  reg  [31:0]         v0_530;
  reg  [31:0]         v0_531;
  reg  [31:0]         v0_532;
  reg  [31:0]         v0_533;
  reg  [31:0]         v0_534;
  reg  [31:0]         v0_535;
  reg  [31:0]         v0_536;
  reg  [31:0]         v0_537;
  reg  [31:0]         v0_538;
  reg  [31:0]         v0_539;
  reg  [31:0]         v0_540;
  reg  [31:0]         v0_541;
  reg  [31:0]         v0_542;
  reg  [31:0]         v0_543;
  reg  [31:0]         v0_544;
  reg  [31:0]         v0_545;
  reg  [31:0]         v0_546;
  reg  [31:0]         v0_547;
  reg  [31:0]         v0_548;
  reg  [31:0]         v0_549;
  reg  [31:0]         v0_550;
  reg  [31:0]         v0_551;
  reg  [31:0]         v0_552;
  reg  [31:0]         v0_553;
  reg  [31:0]         v0_554;
  reg  [31:0]         v0_555;
  reg  [31:0]         v0_556;
  reg  [31:0]         v0_557;
  reg  [31:0]         v0_558;
  reg  [31:0]         v0_559;
  reg  [31:0]         v0_560;
  reg  [31:0]         v0_561;
  reg  [31:0]         v0_562;
  reg  [31:0]         v0_563;
  reg  [31:0]         v0_564;
  reg  [31:0]         v0_565;
  reg  [31:0]         v0_566;
  reg  [31:0]         v0_567;
  reg  [31:0]         v0_568;
  reg  [31:0]         v0_569;
  reg  [31:0]         v0_570;
  reg  [31:0]         v0_571;
  reg  [31:0]         v0_572;
  reg  [31:0]         v0_573;
  reg  [31:0]         v0_574;
  reg  [31:0]         v0_575;
  reg  [31:0]         v0_576;
  reg  [31:0]         v0_577;
  reg  [31:0]         v0_578;
  reg  [31:0]         v0_579;
  reg  [31:0]         v0_580;
  reg  [31:0]         v0_581;
  reg  [31:0]         v0_582;
  reg  [31:0]         v0_583;
  reg  [31:0]         v0_584;
  reg  [31:0]         v0_585;
  reg  [31:0]         v0_586;
  reg  [31:0]         v0_587;
  reg  [31:0]         v0_588;
  reg  [31:0]         v0_589;
  reg  [31:0]         v0_590;
  reg  [31:0]         v0_591;
  reg  [31:0]         v0_592;
  reg  [31:0]         v0_593;
  reg  [31:0]         v0_594;
  reg  [31:0]         v0_595;
  reg  [31:0]         v0_596;
  reg  [31:0]         v0_597;
  reg  [31:0]         v0_598;
  reg  [31:0]         v0_599;
  reg  [31:0]         v0_600;
  reg  [31:0]         v0_601;
  reg  [31:0]         v0_602;
  reg  [31:0]         v0_603;
  reg  [31:0]         v0_604;
  reg  [31:0]         v0_605;
  reg  [31:0]         v0_606;
  reg  [31:0]         v0_607;
  reg  [31:0]         v0_608;
  reg  [31:0]         v0_609;
  reg  [31:0]         v0_610;
  reg  [31:0]         v0_611;
  reg  [31:0]         v0_612;
  reg  [31:0]         v0_613;
  reg  [31:0]         v0_614;
  reg  [31:0]         v0_615;
  reg  [31:0]         v0_616;
  reg  [31:0]         v0_617;
  reg  [31:0]         v0_618;
  reg  [31:0]         v0_619;
  reg  [31:0]         v0_620;
  reg  [31:0]         v0_621;
  reg  [31:0]         v0_622;
  reg  [31:0]         v0_623;
  reg  [31:0]         v0_624;
  reg  [31:0]         v0_625;
  reg  [31:0]         v0_626;
  reg  [31:0]         v0_627;
  reg  [31:0]         v0_628;
  reg  [31:0]         v0_629;
  reg  [31:0]         v0_630;
  reg  [31:0]         v0_631;
  reg  [31:0]         v0_632;
  reg  [31:0]         v0_633;
  reg  [31:0]         v0_634;
  reg  [31:0]         v0_635;
  reg  [31:0]         v0_636;
  reg  [31:0]         v0_637;
  reg  [31:0]         v0_638;
  reg  [31:0]         v0_639;
  reg  [31:0]         v0_640;
  reg  [31:0]         v0_641;
  reg  [31:0]         v0_642;
  reg  [31:0]         v0_643;
  reg  [31:0]         v0_644;
  reg  [31:0]         v0_645;
  reg  [31:0]         v0_646;
  reg  [31:0]         v0_647;
  reg  [31:0]         v0_648;
  reg  [31:0]         v0_649;
  reg  [31:0]         v0_650;
  reg  [31:0]         v0_651;
  reg  [31:0]         v0_652;
  reg  [31:0]         v0_653;
  reg  [31:0]         v0_654;
  reg  [31:0]         v0_655;
  reg  [31:0]         v0_656;
  reg  [31:0]         v0_657;
  reg  [31:0]         v0_658;
  reg  [31:0]         v0_659;
  reg  [31:0]         v0_660;
  reg  [31:0]         v0_661;
  reg  [31:0]         v0_662;
  reg  [31:0]         v0_663;
  reg  [31:0]         v0_664;
  reg  [31:0]         v0_665;
  reg  [31:0]         v0_666;
  reg  [31:0]         v0_667;
  reg  [31:0]         v0_668;
  reg  [31:0]         v0_669;
  reg  [31:0]         v0_670;
  reg  [31:0]         v0_671;
  reg  [31:0]         v0_672;
  reg  [31:0]         v0_673;
  reg  [31:0]         v0_674;
  reg  [31:0]         v0_675;
  reg  [31:0]         v0_676;
  reg  [31:0]         v0_677;
  reg  [31:0]         v0_678;
  reg  [31:0]         v0_679;
  reg  [31:0]         v0_680;
  reg  [31:0]         v0_681;
  reg  [31:0]         v0_682;
  reg  [31:0]         v0_683;
  reg  [31:0]         v0_684;
  reg  [31:0]         v0_685;
  reg  [31:0]         v0_686;
  reg  [31:0]         v0_687;
  reg  [31:0]         v0_688;
  reg  [31:0]         v0_689;
  reg  [31:0]         v0_690;
  reg  [31:0]         v0_691;
  reg  [31:0]         v0_692;
  reg  [31:0]         v0_693;
  reg  [31:0]         v0_694;
  reg  [31:0]         v0_695;
  reg  [31:0]         v0_696;
  reg  [31:0]         v0_697;
  reg  [31:0]         v0_698;
  reg  [31:0]         v0_699;
  reg  [31:0]         v0_700;
  reg  [31:0]         v0_701;
  reg  [31:0]         v0_702;
  reg  [31:0]         v0_703;
  reg  [31:0]         v0_704;
  reg  [31:0]         v0_705;
  reg  [31:0]         v0_706;
  reg  [31:0]         v0_707;
  reg  [31:0]         v0_708;
  reg  [31:0]         v0_709;
  reg  [31:0]         v0_710;
  reg  [31:0]         v0_711;
  reg  [31:0]         v0_712;
  reg  [31:0]         v0_713;
  reg  [31:0]         v0_714;
  reg  [31:0]         v0_715;
  reg  [31:0]         v0_716;
  reg  [31:0]         v0_717;
  reg  [31:0]         v0_718;
  reg  [31:0]         v0_719;
  reg  [31:0]         v0_720;
  reg  [31:0]         v0_721;
  reg  [31:0]         v0_722;
  reg  [31:0]         v0_723;
  reg  [31:0]         v0_724;
  reg  [31:0]         v0_725;
  reg  [31:0]         v0_726;
  reg  [31:0]         v0_727;
  reg  [31:0]         v0_728;
  reg  [31:0]         v0_729;
  reg  [31:0]         v0_730;
  reg  [31:0]         v0_731;
  reg  [31:0]         v0_732;
  reg  [31:0]         v0_733;
  reg  [31:0]         v0_734;
  reg  [31:0]         v0_735;
  reg  [31:0]         v0_736;
  reg  [31:0]         v0_737;
  reg  [31:0]         v0_738;
  reg  [31:0]         v0_739;
  reg  [31:0]         v0_740;
  reg  [31:0]         v0_741;
  reg  [31:0]         v0_742;
  reg  [31:0]         v0_743;
  reg  [31:0]         v0_744;
  reg  [31:0]         v0_745;
  reg  [31:0]         v0_746;
  reg  [31:0]         v0_747;
  reg  [31:0]         v0_748;
  reg  [31:0]         v0_749;
  reg  [31:0]         v0_750;
  reg  [31:0]         v0_751;
  reg  [31:0]         v0_752;
  reg  [31:0]         v0_753;
  reg  [31:0]         v0_754;
  reg  [31:0]         v0_755;
  reg  [31:0]         v0_756;
  reg  [31:0]         v0_757;
  reg  [31:0]         v0_758;
  reg  [31:0]         v0_759;
  reg  [31:0]         v0_760;
  reg  [31:0]         v0_761;
  reg  [31:0]         v0_762;
  reg  [31:0]         v0_763;
  reg  [31:0]         v0_764;
  reg  [31:0]         v0_765;
  reg  [31:0]         v0_766;
  reg  [31:0]         v0_767;
  reg  [31:0]         v0_768;
  reg  [31:0]         v0_769;
  reg  [31:0]         v0_770;
  reg  [31:0]         v0_771;
  reg  [31:0]         v0_772;
  reg  [31:0]         v0_773;
  reg  [31:0]         v0_774;
  reg  [31:0]         v0_775;
  reg  [31:0]         v0_776;
  reg  [31:0]         v0_777;
  reg  [31:0]         v0_778;
  reg  [31:0]         v0_779;
  reg  [31:0]         v0_780;
  reg  [31:0]         v0_781;
  reg  [31:0]         v0_782;
  reg  [31:0]         v0_783;
  reg  [31:0]         v0_784;
  reg  [31:0]         v0_785;
  reg  [31:0]         v0_786;
  reg  [31:0]         v0_787;
  reg  [31:0]         v0_788;
  reg  [31:0]         v0_789;
  reg  [31:0]         v0_790;
  reg  [31:0]         v0_791;
  reg  [31:0]         v0_792;
  reg  [31:0]         v0_793;
  reg  [31:0]         v0_794;
  reg  [31:0]         v0_795;
  reg  [31:0]         v0_796;
  reg  [31:0]         v0_797;
  reg  [31:0]         v0_798;
  reg  [31:0]         v0_799;
  reg  [31:0]         v0_800;
  reg  [31:0]         v0_801;
  reg  [31:0]         v0_802;
  reg  [31:0]         v0_803;
  reg  [31:0]         v0_804;
  reg  [31:0]         v0_805;
  reg  [31:0]         v0_806;
  reg  [31:0]         v0_807;
  reg  [31:0]         v0_808;
  reg  [31:0]         v0_809;
  reg  [31:0]         v0_810;
  reg  [31:0]         v0_811;
  reg  [31:0]         v0_812;
  reg  [31:0]         v0_813;
  reg  [31:0]         v0_814;
  reg  [31:0]         v0_815;
  reg  [31:0]         v0_816;
  reg  [31:0]         v0_817;
  reg  [31:0]         v0_818;
  reg  [31:0]         v0_819;
  reg  [31:0]         v0_820;
  reg  [31:0]         v0_821;
  reg  [31:0]         v0_822;
  reg  [31:0]         v0_823;
  reg  [31:0]         v0_824;
  reg  [31:0]         v0_825;
  reg  [31:0]         v0_826;
  reg  [31:0]         v0_827;
  reg  [31:0]         v0_828;
  reg  [31:0]         v0_829;
  reg  [31:0]         v0_830;
  reg  [31:0]         v0_831;
  reg  [31:0]         v0_832;
  reg  [31:0]         v0_833;
  reg  [31:0]         v0_834;
  reg  [31:0]         v0_835;
  reg  [31:0]         v0_836;
  reg  [31:0]         v0_837;
  reg  [31:0]         v0_838;
  reg  [31:0]         v0_839;
  reg  [31:0]         v0_840;
  reg  [31:0]         v0_841;
  reg  [31:0]         v0_842;
  reg  [31:0]         v0_843;
  reg  [31:0]         v0_844;
  reg  [31:0]         v0_845;
  reg  [31:0]         v0_846;
  reg  [31:0]         v0_847;
  reg  [31:0]         v0_848;
  reg  [31:0]         v0_849;
  reg  [31:0]         v0_850;
  reg  [31:0]         v0_851;
  reg  [31:0]         v0_852;
  reg  [31:0]         v0_853;
  reg  [31:0]         v0_854;
  reg  [31:0]         v0_855;
  reg  [31:0]         v0_856;
  reg  [31:0]         v0_857;
  reg  [31:0]         v0_858;
  reg  [31:0]         v0_859;
  reg  [31:0]         v0_860;
  reg  [31:0]         v0_861;
  reg  [31:0]         v0_862;
  reg  [31:0]         v0_863;
  reg  [31:0]         v0_864;
  reg  [31:0]         v0_865;
  reg  [31:0]         v0_866;
  reg  [31:0]         v0_867;
  reg  [31:0]         v0_868;
  reg  [31:0]         v0_869;
  reg  [31:0]         v0_870;
  reg  [31:0]         v0_871;
  reg  [31:0]         v0_872;
  reg  [31:0]         v0_873;
  reg  [31:0]         v0_874;
  reg  [31:0]         v0_875;
  reg  [31:0]         v0_876;
  reg  [31:0]         v0_877;
  reg  [31:0]         v0_878;
  reg  [31:0]         v0_879;
  reg  [31:0]         v0_880;
  reg  [31:0]         v0_881;
  reg  [31:0]         v0_882;
  reg  [31:0]         v0_883;
  reg  [31:0]         v0_884;
  reg  [31:0]         v0_885;
  reg  [31:0]         v0_886;
  reg  [31:0]         v0_887;
  reg  [31:0]         v0_888;
  reg  [31:0]         v0_889;
  reg  [31:0]         v0_890;
  reg  [31:0]         v0_891;
  reg  [31:0]         v0_892;
  reg  [31:0]         v0_893;
  reg  [31:0]         v0_894;
  reg  [31:0]         v0_895;
  reg  [31:0]         v0_896;
  reg  [31:0]         v0_897;
  reg  [31:0]         v0_898;
  reg  [31:0]         v0_899;
  reg  [31:0]         v0_900;
  reg  [31:0]         v0_901;
  reg  [31:0]         v0_902;
  reg  [31:0]         v0_903;
  reg  [31:0]         v0_904;
  reg  [31:0]         v0_905;
  reg  [31:0]         v0_906;
  reg  [31:0]         v0_907;
  reg  [31:0]         v0_908;
  reg  [31:0]         v0_909;
  reg  [31:0]         v0_910;
  reg  [31:0]         v0_911;
  reg  [31:0]         v0_912;
  reg  [31:0]         v0_913;
  reg  [31:0]         v0_914;
  reg  [31:0]         v0_915;
  reg  [31:0]         v0_916;
  reg  [31:0]         v0_917;
  reg  [31:0]         v0_918;
  reg  [31:0]         v0_919;
  reg  [31:0]         v0_920;
  reg  [31:0]         v0_921;
  reg  [31:0]         v0_922;
  reg  [31:0]         v0_923;
  reg  [31:0]         v0_924;
  reg  [31:0]         v0_925;
  reg  [31:0]         v0_926;
  reg  [31:0]         v0_927;
  reg  [31:0]         v0_928;
  reg  [31:0]         v0_929;
  reg  [31:0]         v0_930;
  reg  [31:0]         v0_931;
  reg  [31:0]         v0_932;
  reg  [31:0]         v0_933;
  reg  [31:0]         v0_934;
  reg  [31:0]         v0_935;
  reg  [31:0]         v0_936;
  reg  [31:0]         v0_937;
  reg  [31:0]         v0_938;
  reg  [31:0]         v0_939;
  reg  [31:0]         v0_940;
  reg  [31:0]         v0_941;
  reg  [31:0]         v0_942;
  reg  [31:0]         v0_943;
  reg  [31:0]         v0_944;
  reg  [31:0]         v0_945;
  reg  [31:0]         v0_946;
  reg  [31:0]         v0_947;
  reg  [31:0]         v0_948;
  reg  [31:0]         v0_949;
  reg  [31:0]         v0_950;
  reg  [31:0]         v0_951;
  reg  [31:0]         v0_952;
  reg  [31:0]         v0_953;
  reg  [31:0]         v0_954;
  reg  [31:0]         v0_955;
  reg  [31:0]         v0_956;
  reg  [31:0]         v0_957;
  reg  [31:0]         v0_958;
  reg  [31:0]         v0_959;
  reg  [31:0]         v0_960;
  reg  [31:0]         v0_961;
  reg  [31:0]         v0_962;
  reg  [31:0]         v0_963;
  reg  [31:0]         v0_964;
  reg  [31:0]         v0_965;
  reg  [31:0]         v0_966;
  reg  [31:0]         v0_967;
  reg  [31:0]         v0_968;
  reg  [31:0]         v0_969;
  reg  [31:0]         v0_970;
  reg  [31:0]         v0_971;
  reg  [31:0]         v0_972;
  reg  [31:0]         v0_973;
  reg  [31:0]         v0_974;
  reg  [31:0]         v0_975;
  reg  [31:0]         v0_976;
  reg  [31:0]         v0_977;
  reg  [31:0]         v0_978;
  reg  [31:0]         v0_979;
  reg  [31:0]         v0_980;
  reg  [31:0]         v0_981;
  reg  [31:0]         v0_982;
  reg  [31:0]         v0_983;
  reg  [31:0]         v0_984;
  reg  [31:0]         v0_985;
  reg  [31:0]         v0_986;
  reg  [31:0]         v0_987;
  reg  [31:0]         v0_988;
  reg  [31:0]         v0_989;
  reg  [31:0]         v0_990;
  reg  [31:0]         v0_991;
  reg  [31:0]         v0_992;
  reg  [31:0]         v0_993;
  reg  [31:0]         v0_994;
  reg  [31:0]         v0_995;
  reg  [31:0]         v0_996;
  reg  [31:0]         v0_997;
  reg  [31:0]         v0_998;
  reg  [31:0]         v0_999;
  reg  [31:0]         v0_1000;
  reg  [31:0]         v0_1001;
  reg  [31:0]         v0_1002;
  reg  [31:0]         v0_1003;
  reg  [31:0]         v0_1004;
  reg  [31:0]         v0_1005;
  reg  [31:0]         v0_1006;
  reg  [31:0]         v0_1007;
  reg  [31:0]         v0_1008;
  reg  [31:0]         v0_1009;
  reg  [31:0]         v0_1010;
  reg  [31:0]         v0_1011;
  reg  [31:0]         v0_1012;
  reg  [31:0]         v0_1013;
  reg  [31:0]         v0_1014;
  reg  [31:0]         v0_1015;
  reg  [31:0]         v0_1016;
  reg  [31:0]         v0_1017;
  reg  [31:0]         v0_1018;
  reg  [31:0]         v0_1019;
  reg  [31:0]         v0_1020;
  reg  [31:0]         v0_1021;
  reg  [31:0]         v0_1022;
  reg  [31:0]         v0_1023;
  wire [15:0]         maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]         maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]         maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]         maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]         maskExt_lo_4 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_4 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]         maskExt_lo_5 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_5 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]         maskExt_lo_6 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_6 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]         maskExt_lo_7 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_7 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]         maskExt_lo_8 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_8 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]         maskExt_lo_9 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_9 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]         maskExt_lo_10 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_10 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]         maskExt_lo_11 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_11 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]         maskExt_lo_12 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_12 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]         maskExt_lo_13 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_13 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]         maskExt_lo_14 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_14 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]         maskExt_lo_15 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_15 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]         maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]         maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]         maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]         maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]         maskExt_lo_20 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_20 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]         maskExt_lo_21 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_21 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]         maskExt_lo_22 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_22 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]         maskExt_lo_23 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_23 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]         maskExt_lo_24 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_24 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]         maskExt_lo_25 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_25 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]         maskExt_lo_26 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_26 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]         maskExt_lo_27 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_27 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]         maskExt_lo_28 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_28 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]         maskExt_lo_29 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_29 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]         maskExt_lo_30 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_30 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]         maskExt_lo_31 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_31 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [15:0]         maskExt_lo_32 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_32 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_32 = {maskExt_hi_32, maskExt_lo_32};
  wire [15:0]         maskExt_lo_33 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_33 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_33 = {maskExt_hi_33, maskExt_lo_33};
  wire [15:0]         maskExt_lo_34 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_34 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_34 = {maskExt_hi_34, maskExt_lo_34};
  wire [15:0]         maskExt_lo_35 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_35 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_35 = {maskExt_hi_35, maskExt_lo_35};
  wire [15:0]         maskExt_lo_36 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_36 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_36 = {maskExt_hi_36, maskExt_lo_36};
  wire [15:0]         maskExt_lo_37 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_37 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_37 = {maskExt_hi_37, maskExt_lo_37};
  wire [15:0]         maskExt_lo_38 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_38 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_38 = {maskExt_hi_38, maskExt_lo_38};
  wire [15:0]         maskExt_lo_39 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_39 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_39 = {maskExt_hi_39, maskExt_lo_39};
  wire [15:0]         maskExt_lo_40 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_40 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_40 = {maskExt_hi_40, maskExt_lo_40};
  wire [15:0]         maskExt_lo_41 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_41 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_41 = {maskExt_hi_41, maskExt_lo_41};
  wire [15:0]         maskExt_lo_42 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_42 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_42 = {maskExt_hi_42, maskExt_lo_42};
  wire [15:0]         maskExt_lo_43 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_43 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_43 = {maskExt_hi_43, maskExt_lo_43};
  wire [15:0]         maskExt_lo_44 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_44 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_44 = {maskExt_hi_44, maskExt_lo_44};
  wire [15:0]         maskExt_lo_45 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_45 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_45 = {maskExt_hi_45, maskExt_lo_45};
  wire [15:0]         maskExt_lo_46 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_46 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_46 = {maskExt_hi_46, maskExt_lo_46};
  wire [15:0]         maskExt_lo_47 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_47 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_47 = {maskExt_hi_47, maskExt_lo_47};
  wire [15:0]         maskExt_lo_48 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_48 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_48 = {maskExt_hi_48, maskExt_lo_48};
  wire [15:0]         maskExt_lo_49 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_49 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_49 = {maskExt_hi_49, maskExt_lo_49};
  wire [15:0]         maskExt_lo_50 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_50 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_50 = {maskExt_hi_50, maskExt_lo_50};
  wire [15:0]         maskExt_lo_51 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_51 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_51 = {maskExt_hi_51, maskExt_lo_51};
  wire [15:0]         maskExt_lo_52 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_52 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_52 = {maskExt_hi_52, maskExt_lo_52};
  wire [15:0]         maskExt_lo_53 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_53 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_53 = {maskExt_hi_53, maskExt_lo_53};
  wire [15:0]         maskExt_lo_54 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_54 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_54 = {maskExt_hi_54, maskExt_lo_54};
  wire [15:0]         maskExt_lo_55 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_55 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_55 = {maskExt_hi_55, maskExt_lo_55};
  wire [15:0]         maskExt_lo_56 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_56 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_56 = {maskExt_hi_56, maskExt_lo_56};
  wire [15:0]         maskExt_lo_57 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_57 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_57 = {maskExt_hi_57, maskExt_lo_57};
  wire [15:0]         maskExt_lo_58 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_58 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_58 = {maskExt_hi_58, maskExt_lo_58};
  wire [15:0]         maskExt_lo_59 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_59 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_59 = {maskExt_hi_59, maskExt_lo_59};
  wire [15:0]         maskExt_lo_60 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_60 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_60 = {maskExt_hi_60, maskExt_lo_60};
  wire [15:0]         maskExt_lo_61 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_61 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_61 = {maskExt_hi_61, maskExt_lo_61};
  wire [15:0]         maskExt_lo_62 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_62 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_62 = {maskExt_hi_62, maskExt_lo_62};
  wire [15:0]         maskExt_lo_63 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_63 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_63 = {maskExt_hi_63, maskExt_lo_63};
  wire [15:0]         maskExt_lo_64 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_64 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_64 = {maskExt_hi_64, maskExt_lo_64};
  wire [15:0]         maskExt_lo_65 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_65 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_65 = {maskExt_hi_65, maskExt_lo_65};
  wire [15:0]         maskExt_lo_66 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_66 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_66 = {maskExt_hi_66, maskExt_lo_66};
  wire [15:0]         maskExt_lo_67 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_67 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_67 = {maskExt_hi_67, maskExt_lo_67};
  wire [15:0]         maskExt_lo_68 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_68 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_68 = {maskExt_hi_68, maskExt_lo_68};
  wire [15:0]         maskExt_lo_69 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_69 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_69 = {maskExt_hi_69, maskExt_lo_69};
  wire [15:0]         maskExt_lo_70 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_70 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_70 = {maskExt_hi_70, maskExt_lo_70};
  wire [15:0]         maskExt_lo_71 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_71 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_71 = {maskExt_hi_71, maskExt_lo_71};
  wire [15:0]         maskExt_lo_72 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_72 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_72 = {maskExt_hi_72, maskExt_lo_72};
  wire [15:0]         maskExt_lo_73 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_73 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_73 = {maskExt_hi_73, maskExt_lo_73};
  wire [15:0]         maskExt_lo_74 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_74 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_74 = {maskExt_hi_74, maskExt_lo_74};
  wire [15:0]         maskExt_lo_75 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_75 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_75 = {maskExt_hi_75, maskExt_lo_75};
  wire [15:0]         maskExt_lo_76 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_76 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_76 = {maskExt_hi_76, maskExt_lo_76};
  wire [15:0]         maskExt_lo_77 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_77 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_77 = {maskExt_hi_77, maskExt_lo_77};
  wire [15:0]         maskExt_lo_78 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_78 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_78 = {maskExt_hi_78, maskExt_lo_78};
  wire [15:0]         maskExt_lo_79 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_79 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_79 = {maskExt_hi_79, maskExt_lo_79};
  wire [15:0]         maskExt_lo_80 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_80 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_80 = {maskExt_hi_80, maskExt_lo_80};
  wire [15:0]         maskExt_lo_81 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_81 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_81 = {maskExt_hi_81, maskExt_lo_81};
  wire [15:0]         maskExt_lo_82 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_82 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_82 = {maskExt_hi_82, maskExt_lo_82};
  wire [15:0]         maskExt_lo_83 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_83 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_83 = {maskExt_hi_83, maskExt_lo_83};
  wire [15:0]         maskExt_lo_84 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_84 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_84 = {maskExt_hi_84, maskExt_lo_84};
  wire [15:0]         maskExt_lo_85 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_85 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_85 = {maskExt_hi_85, maskExt_lo_85};
  wire [15:0]         maskExt_lo_86 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_86 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_86 = {maskExt_hi_86, maskExt_lo_86};
  wire [15:0]         maskExt_lo_87 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_87 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_87 = {maskExt_hi_87, maskExt_lo_87};
  wire [15:0]         maskExt_lo_88 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_88 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_88 = {maskExt_hi_88, maskExt_lo_88};
  wire [15:0]         maskExt_lo_89 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_89 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_89 = {maskExt_hi_89, maskExt_lo_89};
  wire [15:0]         maskExt_lo_90 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_90 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_90 = {maskExt_hi_90, maskExt_lo_90};
  wire [15:0]         maskExt_lo_91 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_91 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_91 = {maskExt_hi_91, maskExt_lo_91};
  wire [15:0]         maskExt_lo_92 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_92 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_92 = {maskExt_hi_92, maskExt_lo_92};
  wire [15:0]         maskExt_lo_93 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_93 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_93 = {maskExt_hi_93, maskExt_lo_93};
  wire [15:0]         maskExt_lo_94 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_94 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_94 = {maskExt_hi_94, maskExt_lo_94};
  wire [15:0]         maskExt_lo_95 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_95 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_95 = {maskExt_hi_95, maskExt_lo_95};
  wire [15:0]         maskExt_lo_96 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_96 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_96 = {maskExt_hi_96, maskExt_lo_96};
  wire [15:0]         maskExt_lo_97 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_97 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_97 = {maskExt_hi_97, maskExt_lo_97};
  wire [15:0]         maskExt_lo_98 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_98 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_98 = {maskExt_hi_98, maskExt_lo_98};
  wire [15:0]         maskExt_lo_99 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_99 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_99 = {maskExt_hi_99, maskExt_lo_99};
  wire [15:0]         maskExt_lo_100 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_100 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_100 = {maskExt_hi_100, maskExt_lo_100};
  wire [15:0]         maskExt_lo_101 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_101 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_101 = {maskExt_hi_101, maskExt_lo_101};
  wire [15:0]         maskExt_lo_102 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_102 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_102 = {maskExt_hi_102, maskExt_lo_102};
  wire [15:0]         maskExt_lo_103 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_103 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_103 = {maskExt_hi_103, maskExt_lo_103};
  wire [15:0]         maskExt_lo_104 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_104 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_104 = {maskExt_hi_104, maskExt_lo_104};
  wire [15:0]         maskExt_lo_105 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_105 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_105 = {maskExt_hi_105, maskExt_lo_105};
  wire [15:0]         maskExt_lo_106 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_106 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_106 = {maskExt_hi_106, maskExt_lo_106};
  wire [15:0]         maskExt_lo_107 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_107 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_107 = {maskExt_hi_107, maskExt_lo_107};
  wire [15:0]         maskExt_lo_108 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_108 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_108 = {maskExt_hi_108, maskExt_lo_108};
  wire [15:0]         maskExt_lo_109 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_109 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_109 = {maskExt_hi_109, maskExt_lo_109};
  wire [15:0]         maskExt_lo_110 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_110 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_110 = {maskExt_hi_110, maskExt_lo_110};
  wire [15:0]         maskExt_lo_111 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_111 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_111 = {maskExt_hi_111, maskExt_lo_111};
  wire [15:0]         maskExt_lo_112 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_112 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_112 = {maskExt_hi_112, maskExt_lo_112};
  wire [15:0]         maskExt_lo_113 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_113 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_113 = {maskExt_hi_113, maskExt_lo_113};
  wire [15:0]         maskExt_lo_114 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_114 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_114 = {maskExt_hi_114, maskExt_lo_114};
  wire [15:0]         maskExt_lo_115 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_115 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_115 = {maskExt_hi_115, maskExt_lo_115};
  wire [15:0]         maskExt_lo_116 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_116 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_116 = {maskExt_hi_116, maskExt_lo_116};
  wire [15:0]         maskExt_lo_117 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_117 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_117 = {maskExt_hi_117, maskExt_lo_117};
  wire [15:0]         maskExt_lo_118 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_118 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_118 = {maskExt_hi_118, maskExt_lo_118};
  wire [15:0]         maskExt_lo_119 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_119 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_119 = {maskExt_hi_119, maskExt_lo_119};
  wire [15:0]         maskExt_lo_120 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_120 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_120 = {maskExt_hi_120, maskExt_lo_120};
  wire [15:0]         maskExt_lo_121 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_121 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_121 = {maskExt_hi_121, maskExt_lo_121};
  wire [15:0]         maskExt_lo_122 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_122 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_122 = {maskExt_hi_122, maskExt_lo_122};
  wire [15:0]         maskExt_lo_123 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_123 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_123 = {maskExt_hi_123, maskExt_lo_123};
  wire [15:0]         maskExt_lo_124 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_124 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_124 = {maskExt_hi_124, maskExt_lo_124};
  wire [15:0]         maskExt_lo_125 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_125 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_125 = {maskExt_hi_125, maskExt_lo_125};
  wire [15:0]         maskExt_lo_126 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_126 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_126 = {maskExt_hi_126, maskExt_lo_126};
  wire [15:0]         maskExt_lo_127 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_127 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_127 = {maskExt_hi_127, maskExt_lo_127};
  wire [15:0]         maskExt_lo_128 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_128 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_128 = {maskExt_hi_128, maskExt_lo_128};
  wire [15:0]         maskExt_lo_129 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_129 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_129 = {maskExt_hi_129, maskExt_lo_129};
  wire [15:0]         maskExt_lo_130 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_130 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_130 = {maskExt_hi_130, maskExt_lo_130};
  wire [15:0]         maskExt_lo_131 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_131 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_131 = {maskExt_hi_131, maskExt_lo_131};
  wire [15:0]         maskExt_lo_132 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_132 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_132 = {maskExt_hi_132, maskExt_lo_132};
  wire [15:0]         maskExt_lo_133 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_133 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_133 = {maskExt_hi_133, maskExt_lo_133};
  wire [15:0]         maskExt_lo_134 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_134 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_134 = {maskExt_hi_134, maskExt_lo_134};
  wire [15:0]         maskExt_lo_135 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_135 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_135 = {maskExt_hi_135, maskExt_lo_135};
  wire [15:0]         maskExt_lo_136 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_136 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_136 = {maskExt_hi_136, maskExt_lo_136};
  wire [15:0]         maskExt_lo_137 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_137 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_137 = {maskExt_hi_137, maskExt_lo_137};
  wire [15:0]         maskExt_lo_138 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_138 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_138 = {maskExt_hi_138, maskExt_lo_138};
  wire [15:0]         maskExt_lo_139 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_139 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_139 = {maskExt_hi_139, maskExt_lo_139};
  wire [15:0]         maskExt_lo_140 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_140 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_140 = {maskExt_hi_140, maskExt_lo_140};
  wire [15:0]         maskExt_lo_141 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_141 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_141 = {maskExt_hi_141, maskExt_lo_141};
  wire [15:0]         maskExt_lo_142 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_142 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_142 = {maskExt_hi_142, maskExt_lo_142};
  wire [15:0]         maskExt_lo_143 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_143 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_143 = {maskExt_hi_143, maskExt_lo_143};
  wire [15:0]         maskExt_lo_144 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_144 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_144 = {maskExt_hi_144, maskExt_lo_144};
  wire [15:0]         maskExt_lo_145 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_145 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_145 = {maskExt_hi_145, maskExt_lo_145};
  wire [15:0]         maskExt_lo_146 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_146 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_146 = {maskExt_hi_146, maskExt_lo_146};
  wire [15:0]         maskExt_lo_147 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_147 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_147 = {maskExt_hi_147, maskExt_lo_147};
  wire [15:0]         maskExt_lo_148 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_148 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_148 = {maskExt_hi_148, maskExt_lo_148};
  wire [15:0]         maskExt_lo_149 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_149 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_149 = {maskExt_hi_149, maskExt_lo_149};
  wire [15:0]         maskExt_lo_150 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_150 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_150 = {maskExt_hi_150, maskExt_lo_150};
  wire [15:0]         maskExt_lo_151 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_151 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_151 = {maskExt_hi_151, maskExt_lo_151};
  wire [15:0]         maskExt_lo_152 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_152 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_152 = {maskExt_hi_152, maskExt_lo_152};
  wire [15:0]         maskExt_lo_153 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_153 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_153 = {maskExt_hi_153, maskExt_lo_153};
  wire [15:0]         maskExt_lo_154 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_154 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_154 = {maskExt_hi_154, maskExt_lo_154};
  wire [15:0]         maskExt_lo_155 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_155 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_155 = {maskExt_hi_155, maskExt_lo_155};
  wire [15:0]         maskExt_lo_156 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_156 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_156 = {maskExt_hi_156, maskExt_lo_156};
  wire [15:0]         maskExt_lo_157 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_157 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_157 = {maskExt_hi_157, maskExt_lo_157};
  wire [15:0]         maskExt_lo_158 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_158 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_158 = {maskExt_hi_158, maskExt_lo_158};
  wire [15:0]         maskExt_lo_159 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_159 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_159 = {maskExt_hi_159, maskExt_lo_159};
  wire [15:0]         maskExt_lo_160 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_160 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_160 = {maskExt_hi_160, maskExt_lo_160};
  wire [15:0]         maskExt_lo_161 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_161 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_161 = {maskExt_hi_161, maskExt_lo_161};
  wire [15:0]         maskExt_lo_162 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_162 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_162 = {maskExt_hi_162, maskExt_lo_162};
  wire [15:0]         maskExt_lo_163 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_163 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_163 = {maskExt_hi_163, maskExt_lo_163};
  wire [15:0]         maskExt_lo_164 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_164 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_164 = {maskExt_hi_164, maskExt_lo_164};
  wire [15:0]         maskExt_lo_165 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_165 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_165 = {maskExt_hi_165, maskExt_lo_165};
  wire [15:0]         maskExt_lo_166 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_166 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_166 = {maskExt_hi_166, maskExt_lo_166};
  wire [15:0]         maskExt_lo_167 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_167 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_167 = {maskExt_hi_167, maskExt_lo_167};
  wire [15:0]         maskExt_lo_168 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_168 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_168 = {maskExt_hi_168, maskExt_lo_168};
  wire [15:0]         maskExt_lo_169 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_169 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_169 = {maskExt_hi_169, maskExt_lo_169};
  wire [15:0]         maskExt_lo_170 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_170 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_170 = {maskExt_hi_170, maskExt_lo_170};
  wire [15:0]         maskExt_lo_171 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_171 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_171 = {maskExt_hi_171, maskExt_lo_171};
  wire [15:0]         maskExt_lo_172 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_172 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_172 = {maskExt_hi_172, maskExt_lo_172};
  wire [15:0]         maskExt_lo_173 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_173 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_173 = {maskExt_hi_173, maskExt_lo_173};
  wire [15:0]         maskExt_lo_174 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_174 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_174 = {maskExt_hi_174, maskExt_lo_174};
  wire [15:0]         maskExt_lo_175 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_175 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_175 = {maskExt_hi_175, maskExt_lo_175};
  wire [15:0]         maskExt_lo_176 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_176 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_176 = {maskExt_hi_176, maskExt_lo_176};
  wire [15:0]         maskExt_lo_177 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_177 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_177 = {maskExt_hi_177, maskExt_lo_177};
  wire [15:0]         maskExt_lo_178 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_178 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_178 = {maskExt_hi_178, maskExt_lo_178};
  wire [15:0]         maskExt_lo_179 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_179 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_179 = {maskExt_hi_179, maskExt_lo_179};
  wire [15:0]         maskExt_lo_180 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_180 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_180 = {maskExt_hi_180, maskExt_lo_180};
  wire [15:0]         maskExt_lo_181 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_181 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_181 = {maskExt_hi_181, maskExt_lo_181};
  wire [15:0]         maskExt_lo_182 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_182 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_182 = {maskExt_hi_182, maskExt_lo_182};
  wire [15:0]         maskExt_lo_183 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_183 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_183 = {maskExt_hi_183, maskExt_lo_183};
  wire [15:0]         maskExt_lo_184 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_184 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_184 = {maskExt_hi_184, maskExt_lo_184};
  wire [15:0]         maskExt_lo_185 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_185 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_185 = {maskExt_hi_185, maskExt_lo_185};
  wire [15:0]         maskExt_lo_186 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_186 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_186 = {maskExt_hi_186, maskExt_lo_186};
  wire [15:0]         maskExt_lo_187 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_187 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_187 = {maskExt_hi_187, maskExt_lo_187};
  wire [15:0]         maskExt_lo_188 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_188 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_188 = {maskExt_hi_188, maskExt_lo_188};
  wire [15:0]         maskExt_lo_189 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_189 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_189 = {maskExt_hi_189, maskExt_lo_189};
  wire [15:0]         maskExt_lo_190 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_190 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_190 = {maskExt_hi_190, maskExt_lo_190};
  wire [15:0]         maskExt_lo_191 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_191 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_191 = {maskExt_hi_191, maskExt_lo_191};
  wire [15:0]         maskExt_lo_192 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_192 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_192 = {maskExt_hi_192, maskExt_lo_192};
  wire [15:0]         maskExt_lo_193 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_193 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_193 = {maskExt_hi_193, maskExt_lo_193};
  wire [15:0]         maskExt_lo_194 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_194 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_194 = {maskExt_hi_194, maskExt_lo_194};
  wire [15:0]         maskExt_lo_195 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_195 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_195 = {maskExt_hi_195, maskExt_lo_195};
  wire [15:0]         maskExt_lo_196 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_196 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_196 = {maskExt_hi_196, maskExt_lo_196};
  wire [15:0]         maskExt_lo_197 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_197 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_197 = {maskExt_hi_197, maskExt_lo_197};
  wire [15:0]         maskExt_lo_198 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_198 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_198 = {maskExt_hi_198, maskExt_lo_198};
  wire [15:0]         maskExt_lo_199 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_199 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_199 = {maskExt_hi_199, maskExt_lo_199};
  wire [15:0]         maskExt_lo_200 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_200 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_200 = {maskExt_hi_200, maskExt_lo_200};
  wire [15:0]         maskExt_lo_201 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_201 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_201 = {maskExt_hi_201, maskExt_lo_201};
  wire [15:0]         maskExt_lo_202 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_202 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_202 = {maskExt_hi_202, maskExt_lo_202};
  wire [15:0]         maskExt_lo_203 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_203 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_203 = {maskExt_hi_203, maskExt_lo_203};
  wire [15:0]         maskExt_lo_204 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_204 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_204 = {maskExt_hi_204, maskExt_lo_204};
  wire [15:0]         maskExt_lo_205 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_205 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_205 = {maskExt_hi_205, maskExt_lo_205};
  wire [15:0]         maskExt_lo_206 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_206 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_206 = {maskExt_hi_206, maskExt_lo_206};
  wire [15:0]         maskExt_lo_207 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_207 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_207 = {maskExt_hi_207, maskExt_lo_207};
  wire [15:0]         maskExt_lo_208 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_208 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_208 = {maskExt_hi_208, maskExt_lo_208};
  wire [15:0]         maskExt_lo_209 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_209 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_209 = {maskExt_hi_209, maskExt_lo_209};
  wire [15:0]         maskExt_lo_210 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_210 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_210 = {maskExt_hi_210, maskExt_lo_210};
  wire [15:0]         maskExt_lo_211 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_211 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_211 = {maskExt_hi_211, maskExt_lo_211};
  wire [15:0]         maskExt_lo_212 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_212 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_212 = {maskExt_hi_212, maskExt_lo_212};
  wire [15:0]         maskExt_lo_213 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_213 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_213 = {maskExt_hi_213, maskExt_lo_213};
  wire [15:0]         maskExt_lo_214 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_214 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_214 = {maskExt_hi_214, maskExt_lo_214};
  wire [15:0]         maskExt_lo_215 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_215 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_215 = {maskExt_hi_215, maskExt_lo_215};
  wire [15:0]         maskExt_lo_216 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_216 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_216 = {maskExt_hi_216, maskExt_lo_216};
  wire [15:0]         maskExt_lo_217 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_217 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_217 = {maskExt_hi_217, maskExt_lo_217};
  wire [15:0]         maskExt_lo_218 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_218 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_218 = {maskExt_hi_218, maskExt_lo_218};
  wire [15:0]         maskExt_lo_219 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_219 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_219 = {maskExt_hi_219, maskExt_lo_219};
  wire [15:0]         maskExt_lo_220 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_220 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_220 = {maskExt_hi_220, maskExt_lo_220};
  wire [15:0]         maskExt_lo_221 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_221 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_221 = {maskExt_hi_221, maskExt_lo_221};
  wire [15:0]         maskExt_lo_222 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_222 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_222 = {maskExt_hi_222, maskExt_lo_222};
  wire [15:0]         maskExt_lo_223 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_223 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_223 = {maskExt_hi_223, maskExt_lo_223};
  wire [15:0]         maskExt_lo_224 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_224 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_224 = {maskExt_hi_224, maskExt_lo_224};
  wire [15:0]         maskExt_lo_225 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_225 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_225 = {maskExt_hi_225, maskExt_lo_225};
  wire [15:0]         maskExt_lo_226 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_226 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_226 = {maskExt_hi_226, maskExt_lo_226};
  wire [15:0]         maskExt_lo_227 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_227 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_227 = {maskExt_hi_227, maskExt_lo_227};
  wire [15:0]         maskExt_lo_228 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_228 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_228 = {maskExt_hi_228, maskExt_lo_228};
  wire [15:0]         maskExt_lo_229 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_229 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_229 = {maskExt_hi_229, maskExt_lo_229};
  wire [15:0]         maskExt_lo_230 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_230 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_230 = {maskExt_hi_230, maskExt_lo_230};
  wire [15:0]         maskExt_lo_231 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_231 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_231 = {maskExt_hi_231, maskExt_lo_231};
  wire [15:0]         maskExt_lo_232 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_232 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_232 = {maskExt_hi_232, maskExt_lo_232};
  wire [15:0]         maskExt_lo_233 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_233 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_233 = {maskExt_hi_233, maskExt_lo_233};
  wire [15:0]         maskExt_lo_234 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_234 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_234 = {maskExt_hi_234, maskExt_lo_234};
  wire [15:0]         maskExt_lo_235 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_235 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_235 = {maskExt_hi_235, maskExt_lo_235};
  wire [15:0]         maskExt_lo_236 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_236 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_236 = {maskExt_hi_236, maskExt_lo_236};
  wire [15:0]         maskExt_lo_237 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_237 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_237 = {maskExt_hi_237, maskExt_lo_237};
  wire [15:0]         maskExt_lo_238 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_238 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_238 = {maskExt_hi_238, maskExt_lo_238};
  wire [15:0]         maskExt_lo_239 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_239 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_239 = {maskExt_hi_239, maskExt_lo_239};
  wire [15:0]         maskExt_lo_240 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_240 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_240 = {maskExt_hi_240, maskExt_lo_240};
  wire [15:0]         maskExt_lo_241 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_241 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_241 = {maskExt_hi_241, maskExt_lo_241};
  wire [15:0]         maskExt_lo_242 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_242 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_242 = {maskExt_hi_242, maskExt_lo_242};
  wire [15:0]         maskExt_lo_243 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_243 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_243 = {maskExt_hi_243, maskExt_lo_243};
  wire [15:0]         maskExt_lo_244 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_244 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_244 = {maskExt_hi_244, maskExt_lo_244};
  wire [15:0]         maskExt_lo_245 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_245 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_245 = {maskExt_hi_245, maskExt_lo_245};
  wire [15:0]         maskExt_lo_246 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_246 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_246 = {maskExt_hi_246, maskExt_lo_246};
  wire [15:0]         maskExt_lo_247 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_247 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_247 = {maskExt_hi_247, maskExt_lo_247};
  wire [15:0]         maskExt_lo_248 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_248 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_248 = {maskExt_hi_248, maskExt_lo_248};
  wire [15:0]         maskExt_lo_249 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_249 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_249 = {maskExt_hi_249, maskExt_lo_249};
  wire [15:0]         maskExt_lo_250 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_250 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_250 = {maskExt_hi_250, maskExt_lo_250};
  wire [15:0]         maskExt_lo_251 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_251 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_251 = {maskExt_hi_251, maskExt_lo_251};
  wire [15:0]         maskExt_lo_252 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_252 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_252 = {maskExt_hi_252, maskExt_lo_252};
  wire [15:0]         maskExt_lo_253 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_253 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_253 = {maskExt_hi_253, maskExt_lo_253};
  wire [15:0]         maskExt_lo_254 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_254 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_254 = {maskExt_hi_254, maskExt_lo_254};
  wire [15:0]         maskExt_lo_255 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_255 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_255 = {maskExt_hi_255, maskExt_lo_255};
  wire [15:0]         maskExt_lo_256 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_256 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_256 = {maskExt_hi_256, maskExt_lo_256};
  wire [15:0]         maskExt_lo_257 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_257 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_257 = {maskExt_hi_257, maskExt_lo_257};
  wire [15:0]         maskExt_lo_258 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_258 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_258 = {maskExt_hi_258, maskExt_lo_258};
  wire [15:0]         maskExt_lo_259 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_259 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_259 = {maskExt_hi_259, maskExt_lo_259};
  wire [15:0]         maskExt_lo_260 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_260 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_260 = {maskExt_hi_260, maskExt_lo_260};
  wire [15:0]         maskExt_lo_261 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_261 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_261 = {maskExt_hi_261, maskExt_lo_261};
  wire [15:0]         maskExt_lo_262 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_262 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_262 = {maskExt_hi_262, maskExt_lo_262};
  wire [15:0]         maskExt_lo_263 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_263 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_263 = {maskExt_hi_263, maskExt_lo_263};
  wire [15:0]         maskExt_lo_264 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_264 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_264 = {maskExt_hi_264, maskExt_lo_264};
  wire [15:0]         maskExt_lo_265 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_265 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_265 = {maskExt_hi_265, maskExt_lo_265};
  wire [15:0]         maskExt_lo_266 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_266 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_266 = {maskExt_hi_266, maskExt_lo_266};
  wire [15:0]         maskExt_lo_267 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_267 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_267 = {maskExt_hi_267, maskExt_lo_267};
  wire [15:0]         maskExt_lo_268 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_268 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_268 = {maskExt_hi_268, maskExt_lo_268};
  wire [15:0]         maskExt_lo_269 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_269 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_269 = {maskExt_hi_269, maskExt_lo_269};
  wire [15:0]         maskExt_lo_270 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_270 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_270 = {maskExt_hi_270, maskExt_lo_270};
  wire [15:0]         maskExt_lo_271 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_271 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_271 = {maskExt_hi_271, maskExt_lo_271};
  wire [15:0]         maskExt_lo_272 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_272 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_272 = {maskExt_hi_272, maskExt_lo_272};
  wire [15:0]         maskExt_lo_273 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_273 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_273 = {maskExt_hi_273, maskExt_lo_273};
  wire [15:0]         maskExt_lo_274 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_274 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_274 = {maskExt_hi_274, maskExt_lo_274};
  wire [15:0]         maskExt_lo_275 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_275 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_275 = {maskExt_hi_275, maskExt_lo_275};
  wire [15:0]         maskExt_lo_276 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_276 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_276 = {maskExt_hi_276, maskExt_lo_276};
  wire [15:0]         maskExt_lo_277 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_277 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_277 = {maskExt_hi_277, maskExt_lo_277};
  wire [15:0]         maskExt_lo_278 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_278 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_278 = {maskExt_hi_278, maskExt_lo_278};
  wire [15:0]         maskExt_lo_279 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_279 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_279 = {maskExt_hi_279, maskExt_lo_279};
  wire [15:0]         maskExt_lo_280 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_280 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_280 = {maskExt_hi_280, maskExt_lo_280};
  wire [15:0]         maskExt_lo_281 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_281 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_281 = {maskExt_hi_281, maskExt_lo_281};
  wire [15:0]         maskExt_lo_282 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_282 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_282 = {maskExt_hi_282, maskExt_lo_282};
  wire [15:0]         maskExt_lo_283 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_283 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_283 = {maskExt_hi_283, maskExt_lo_283};
  wire [15:0]         maskExt_lo_284 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_284 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_284 = {maskExt_hi_284, maskExt_lo_284};
  wire [15:0]         maskExt_lo_285 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_285 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_285 = {maskExt_hi_285, maskExt_lo_285};
  wire [15:0]         maskExt_lo_286 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_286 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_286 = {maskExt_hi_286, maskExt_lo_286};
  wire [15:0]         maskExt_lo_287 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_287 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_287 = {maskExt_hi_287, maskExt_lo_287};
  wire [15:0]         maskExt_lo_288 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_288 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_288 = {maskExt_hi_288, maskExt_lo_288};
  wire [15:0]         maskExt_lo_289 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_289 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_289 = {maskExt_hi_289, maskExt_lo_289};
  wire [15:0]         maskExt_lo_290 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_290 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_290 = {maskExt_hi_290, maskExt_lo_290};
  wire [15:0]         maskExt_lo_291 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_291 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_291 = {maskExt_hi_291, maskExt_lo_291};
  wire [15:0]         maskExt_lo_292 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_292 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_292 = {maskExt_hi_292, maskExt_lo_292};
  wire [15:0]         maskExt_lo_293 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_293 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_293 = {maskExt_hi_293, maskExt_lo_293};
  wire [15:0]         maskExt_lo_294 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_294 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_294 = {maskExt_hi_294, maskExt_lo_294};
  wire [15:0]         maskExt_lo_295 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_295 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_295 = {maskExt_hi_295, maskExt_lo_295};
  wire [15:0]         maskExt_lo_296 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_296 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_296 = {maskExt_hi_296, maskExt_lo_296};
  wire [15:0]         maskExt_lo_297 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_297 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_297 = {maskExt_hi_297, maskExt_lo_297};
  wire [15:0]         maskExt_lo_298 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_298 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_298 = {maskExt_hi_298, maskExt_lo_298};
  wire [15:0]         maskExt_lo_299 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_299 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_299 = {maskExt_hi_299, maskExt_lo_299};
  wire [15:0]         maskExt_lo_300 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_300 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_300 = {maskExt_hi_300, maskExt_lo_300};
  wire [15:0]         maskExt_lo_301 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_301 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_301 = {maskExt_hi_301, maskExt_lo_301};
  wire [15:0]         maskExt_lo_302 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_302 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_302 = {maskExt_hi_302, maskExt_lo_302};
  wire [15:0]         maskExt_lo_303 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_303 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_303 = {maskExt_hi_303, maskExt_lo_303};
  wire [15:0]         maskExt_lo_304 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_304 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_304 = {maskExt_hi_304, maskExt_lo_304};
  wire [15:0]         maskExt_lo_305 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_305 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_305 = {maskExt_hi_305, maskExt_lo_305};
  wire [15:0]         maskExt_lo_306 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_306 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_306 = {maskExt_hi_306, maskExt_lo_306};
  wire [15:0]         maskExt_lo_307 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_307 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_307 = {maskExt_hi_307, maskExt_lo_307};
  wire [15:0]         maskExt_lo_308 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_308 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_308 = {maskExt_hi_308, maskExt_lo_308};
  wire [15:0]         maskExt_lo_309 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_309 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_309 = {maskExt_hi_309, maskExt_lo_309};
  wire [15:0]         maskExt_lo_310 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_310 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_310 = {maskExt_hi_310, maskExt_lo_310};
  wire [15:0]         maskExt_lo_311 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_311 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_311 = {maskExt_hi_311, maskExt_lo_311};
  wire [15:0]         maskExt_lo_312 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_312 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_312 = {maskExt_hi_312, maskExt_lo_312};
  wire [15:0]         maskExt_lo_313 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_313 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_313 = {maskExt_hi_313, maskExt_lo_313};
  wire [15:0]         maskExt_lo_314 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_314 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_314 = {maskExt_hi_314, maskExt_lo_314};
  wire [15:0]         maskExt_lo_315 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_315 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_315 = {maskExt_hi_315, maskExt_lo_315};
  wire [15:0]         maskExt_lo_316 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_316 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_316 = {maskExt_hi_316, maskExt_lo_316};
  wire [15:0]         maskExt_lo_317 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_317 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_317 = {maskExt_hi_317, maskExt_lo_317};
  wire [15:0]         maskExt_lo_318 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_318 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_318 = {maskExt_hi_318, maskExt_lo_318};
  wire [15:0]         maskExt_lo_319 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_319 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_319 = {maskExt_hi_319, maskExt_lo_319};
  wire [15:0]         maskExt_lo_320 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_320 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_320 = {maskExt_hi_320, maskExt_lo_320};
  wire [15:0]         maskExt_lo_321 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_321 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_321 = {maskExt_hi_321, maskExt_lo_321};
  wire [15:0]         maskExt_lo_322 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_322 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_322 = {maskExt_hi_322, maskExt_lo_322};
  wire [15:0]         maskExt_lo_323 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_323 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_323 = {maskExt_hi_323, maskExt_lo_323};
  wire [15:0]         maskExt_lo_324 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_324 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_324 = {maskExt_hi_324, maskExt_lo_324};
  wire [15:0]         maskExt_lo_325 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_325 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_325 = {maskExt_hi_325, maskExt_lo_325};
  wire [15:0]         maskExt_lo_326 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_326 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_326 = {maskExt_hi_326, maskExt_lo_326};
  wire [15:0]         maskExt_lo_327 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_327 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_327 = {maskExt_hi_327, maskExt_lo_327};
  wire [15:0]         maskExt_lo_328 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_328 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_328 = {maskExt_hi_328, maskExt_lo_328};
  wire [15:0]         maskExt_lo_329 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_329 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_329 = {maskExt_hi_329, maskExt_lo_329};
  wire [15:0]         maskExt_lo_330 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_330 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_330 = {maskExt_hi_330, maskExt_lo_330};
  wire [15:0]         maskExt_lo_331 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_331 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_331 = {maskExt_hi_331, maskExt_lo_331};
  wire [15:0]         maskExt_lo_332 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_332 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_332 = {maskExt_hi_332, maskExt_lo_332};
  wire [15:0]         maskExt_lo_333 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_333 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_333 = {maskExt_hi_333, maskExt_lo_333};
  wire [15:0]         maskExt_lo_334 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_334 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_334 = {maskExt_hi_334, maskExt_lo_334};
  wire [15:0]         maskExt_lo_335 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_335 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_335 = {maskExt_hi_335, maskExt_lo_335};
  wire [15:0]         maskExt_lo_336 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_336 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_336 = {maskExt_hi_336, maskExt_lo_336};
  wire [15:0]         maskExt_lo_337 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_337 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_337 = {maskExt_hi_337, maskExt_lo_337};
  wire [15:0]         maskExt_lo_338 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_338 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_338 = {maskExt_hi_338, maskExt_lo_338};
  wire [15:0]         maskExt_lo_339 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_339 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_339 = {maskExt_hi_339, maskExt_lo_339};
  wire [15:0]         maskExt_lo_340 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_340 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_340 = {maskExt_hi_340, maskExt_lo_340};
  wire [15:0]         maskExt_lo_341 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_341 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_341 = {maskExt_hi_341, maskExt_lo_341};
  wire [15:0]         maskExt_lo_342 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_342 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_342 = {maskExt_hi_342, maskExt_lo_342};
  wire [15:0]         maskExt_lo_343 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_343 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_343 = {maskExt_hi_343, maskExt_lo_343};
  wire [15:0]         maskExt_lo_344 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_344 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_344 = {maskExt_hi_344, maskExt_lo_344};
  wire [15:0]         maskExt_lo_345 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_345 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_345 = {maskExt_hi_345, maskExt_lo_345};
  wire [15:0]         maskExt_lo_346 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_346 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_346 = {maskExt_hi_346, maskExt_lo_346};
  wire [15:0]         maskExt_lo_347 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_347 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_347 = {maskExt_hi_347, maskExt_lo_347};
  wire [15:0]         maskExt_lo_348 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_348 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_348 = {maskExt_hi_348, maskExt_lo_348};
  wire [15:0]         maskExt_lo_349 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_349 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_349 = {maskExt_hi_349, maskExt_lo_349};
  wire [15:0]         maskExt_lo_350 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_350 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_350 = {maskExt_hi_350, maskExt_lo_350};
  wire [15:0]         maskExt_lo_351 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_351 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_351 = {maskExt_hi_351, maskExt_lo_351};
  wire [15:0]         maskExt_lo_352 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_352 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_352 = {maskExt_hi_352, maskExt_lo_352};
  wire [15:0]         maskExt_lo_353 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_353 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_353 = {maskExt_hi_353, maskExt_lo_353};
  wire [15:0]         maskExt_lo_354 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_354 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_354 = {maskExt_hi_354, maskExt_lo_354};
  wire [15:0]         maskExt_lo_355 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_355 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_355 = {maskExt_hi_355, maskExt_lo_355};
  wire [15:0]         maskExt_lo_356 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_356 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_356 = {maskExt_hi_356, maskExt_lo_356};
  wire [15:0]         maskExt_lo_357 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_357 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_357 = {maskExt_hi_357, maskExt_lo_357};
  wire [15:0]         maskExt_lo_358 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_358 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_358 = {maskExt_hi_358, maskExt_lo_358};
  wire [15:0]         maskExt_lo_359 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_359 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_359 = {maskExt_hi_359, maskExt_lo_359};
  wire [15:0]         maskExt_lo_360 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_360 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_360 = {maskExt_hi_360, maskExt_lo_360};
  wire [15:0]         maskExt_lo_361 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_361 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_361 = {maskExt_hi_361, maskExt_lo_361};
  wire [15:0]         maskExt_lo_362 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_362 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_362 = {maskExt_hi_362, maskExt_lo_362};
  wire [15:0]         maskExt_lo_363 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_363 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_363 = {maskExt_hi_363, maskExt_lo_363};
  wire [15:0]         maskExt_lo_364 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_364 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_364 = {maskExt_hi_364, maskExt_lo_364};
  wire [15:0]         maskExt_lo_365 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_365 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_365 = {maskExt_hi_365, maskExt_lo_365};
  wire [15:0]         maskExt_lo_366 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_366 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_366 = {maskExt_hi_366, maskExt_lo_366};
  wire [15:0]         maskExt_lo_367 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_367 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_367 = {maskExt_hi_367, maskExt_lo_367};
  wire [15:0]         maskExt_lo_368 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_368 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_368 = {maskExt_hi_368, maskExt_lo_368};
  wire [15:0]         maskExt_lo_369 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_369 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_369 = {maskExt_hi_369, maskExt_lo_369};
  wire [15:0]         maskExt_lo_370 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_370 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_370 = {maskExt_hi_370, maskExt_lo_370};
  wire [15:0]         maskExt_lo_371 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_371 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_371 = {maskExt_hi_371, maskExt_lo_371};
  wire [15:0]         maskExt_lo_372 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_372 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_372 = {maskExt_hi_372, maskExt_lo_372};
  wire [15:0]         maskExt_lo_373 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_373 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_373 = {maskExt_hi_373, maskExt_lo_373};
  wire [15:0]         maskExt_lo_374 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_374 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_374 = {maskExt_hi_374, maskExt_lo_374};
  wire [15:0]         maskExt_lo_375 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_375 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_375 = {maskExt_hi_375, maskExt_lo_375};
  wire [15:0]         maskExt_lo_376 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_376 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_376 = {maskExt_hi_376, maskExt_lo_376};
  wire [15:0]         maskExt_lo_377 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_377 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_377 = {maskExt_hi_377, maskExt_lo_377};
  wire [15:0]         maskExt_lo_378 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_378 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_378 = {maskExt_hi_378, maskExt_lo_378};
  wire [15:0]         maskExt_lo_379 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_379 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_379 = {maskExt_hi_379, maskExt_lo_379};
  wire [15:0]         maskExt_lo_380 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_380 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_380 = {maskExt_hi_380, maskExt_lo_380};
  wire [15:0]         maskExt_lo_381 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_381 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_381 = {maskExt_hi_381, maskExt_lo_381};
  wire [15:0]         maskExt_lo_382 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_382 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_382 = {maskExt_hi_382, maskExt_lo_382};
  wire [15:0]         maskExt_lo_383 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_383 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_383 = {maskExt_hi_383, maskExt_lo_383};
  wire [15:0]         maskExt_lo_384 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_384 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_384 = {maskExt_hi_384, maskExt_lo_384};
  wire [15:0]         maskExt_lo_385 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_385 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_385 = {maskExt_hi_385, maskExt_lo_385};
  wire [15:0]         maskExt_lo_386 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_386 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_386 = {maskExt_hi_386, maskExt_lo_386};
  wire [15:0]         maskExt_lo_387 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_387 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_387 = {maskExt_hi_387, maskExt_lo_387};
  wire [15:0]         maskExt_lo_388 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_388 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_388 = {maskExt_hi_388, maskExt_lo_388};
  wire [15:0]         maskExt_lo_389 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_389 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_389 = {maskExt_hi_389, maskExt_lo_389};
  wire [15:0]         maskExt_lo_390 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_390 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_390 = {maskExt_hi_390, maskExt_lo_390};
  wire [15:0]         maskExt_lo_391 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_391 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_391 = {maskExt_hi_391, maskExt_lo_391};
  wire [15:0]         maskExt_lo_392 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_392 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_392 = {maskExt_hi_392, maskExt_lo_392};
  wire [15:0]         maskExt_lo_393 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_393 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_393 = {maskExt_hi_393, maskExt_lo_393};
  wire [15:0]         maskExt_lo_394 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_394 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_394 = {maskExt_hi_394, maskExt_lo_394};
  wire [15:0]         maskExt_lo_395 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_395 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_395 = {maskExt_hi_395, maskExt_lo_395};
  wire [15:0]         maskExt_lo_396 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_396 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_396 = {maskExt_hi_396, maskExt_lo_396};
  wire [15:0]         maskExt_lo_397 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_397 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_397 = {maskExt_hi_397, maskExt_lo_397};
  wire [15:0]         maskExt_lo_398 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_398 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_398 = {maskExt_hi_398, maskExt_lo_398};
  wire [15:0]         maskExt_lo_399 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_399 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_399 = {maskExt_hi_399, maskExt_lo_399};
  wire [15:0]         maskExt_lo_400 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_400 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_400 = {maskExt_hi_400, maskExt_lo_400};
  wire [15:0]         maskExt_lo_401 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_401 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_401 = {maskExt_hi_401, maskExt_lo_401};
  wire [15:0]         maskExt_lo_402 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_402 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_402 = {maskExt_hi_402, maskExt_lo_402};
  wire [15:0]         maskExt_lo_403 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_403 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_403 = {maskExt_hi_403, maskExt_lo_403};
  wire [15:0]         maskExt_lo_404 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_404 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_404 = {maskExt_hi_404, maskExt_lo_404};
  wire [15:0]         maskExt_lo_405 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_405 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_405 = {maskExt_hi_405, maskExt_lo_405};
  wire [15:0]         maskExt_lo_406 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_406 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_406 = {maskExt_hi_406, maskExt_lo_406};
  wire [15:0]         maskExt_lo_407 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_407 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_407 = {maskExt_hi_407, maskExt_lo_407};
  wire [15:0]         maskExt_lo_408 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_408 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_408 = {maskExt_hi_408, maskExt_lo_408};
  wire [15:0]         maskExt_lo_409 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_409 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_409 = {maskExt_hi_409, maskExt_lo_409};
  wire [15:0]         maskExt_lo_410 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_410 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_410 = {maskExt_hi_410, maskExt_lo_410};
  wire [15:0]         maskExt_lo_411 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_411 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_411 = {maskExt_hi_411, maskExt_lo_411};
  wire [15:0]         maskExt_lo_412 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_412 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_412 = {maskExt_hi_412, maskExt_lo_412};
  wire [15:0]         maskExt_lo_413 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_413 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_413 = {maskExt_hi_413, maskExt_lo_413};
  wire [15:0]         maskExt_lo_414 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_414 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_414 = {maskExt_hi_414, maskExt_lo_414};
  wire [15:0]         maskExt_lo_415 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_415 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_415 = {maskExt_hi_415, maskExt_lo_415};
  wire [15:0]         maskExt_lo_416 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_416 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_416 = {maskExt_hi_416, maskExt_lo_416};
  wire [15:0]         maskExt_lo_417 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_417 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_417 = {maskExt_hi_417, maskExt_lo_417};
  wire [15:0]         maskExt_lo_418 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_418 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_418 = {maskExt_hi_418, maskExt_lo_418};
  wire [15:0]         maskExt_lo_419 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_419 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_419 = {maskExt_hi_419, maskExt_lo_419};
  wire [15:0]         maskExt_lo_420 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_420 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_420 = {maskExt_hi_420, maskExt_lo_420};
  wire [15:0]         maskExt_lo_421 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_421 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_421 = {maskExt_hi_421, maskExt_lo_421};
  wire [15:0]         maskExt_lo_422 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_422 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_422 = {maskExt_hi_422, maskExt_lo_422};
  wire [15:0]         maskExt_lo_423 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_423 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_423 = {maskExt_hi_423, maskExt_lo_423};
  wire [15:0]         maskExt_lo_424 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_424 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_424 = {maskExt_hi_424, maskExt_lo_424};
  wire [15:0]         maskExt_lo_425 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_425 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_425 = {maskExt_hi_425, maskExt_lo_425};
  wire [15:0]         maskExt_lo_426 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_426 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_426 = {maskExt_hi_426, maskExt_lo_426};
  wire [15:0]         maskExt_lo_427 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_427 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_427 = {maskExt_hi_427, maskExt_lo_427};
  wire [15:0]         maskExt_lo_428 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_428 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_428 = {maskExt_hi_428, maskExt_lo_428};
  wire [15:0]         maskExt_lo_429 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_429 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_429 = {maskExt_hi_429, maskExt_lo_429};
  wire [15:0]         maskExt_lo_430 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_430 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_430 = {maskExt_hi_430, maskExt_lo_430};
  wire [15:0]         maskExt_lo_431 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_431 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_431 = {maskExt_hi_431, maskExt_lo_431};
  wire [15:0]         maskExt_lo_432 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_432 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_432 = {maskExt_hi_432, maskExt_lo_432};
  wire [15:0]         maskExt_lo_433 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_433 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_433 = {maskExt_hi_433, maskExt_lo_433};
  wire [15:0]         maskExt_lo_434 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_434 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_434 = {maskExt_hi_434, maskExt_lo_434};
  wire [15:0]         maskExt_lo_435 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_435 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_435 = {maskExt_hi_435, maskExt_lo_435};
  wire [15:0]         maskExt_lo_436 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_436 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_436 = {maskExt_hi_436, maskExt_lo_436};
  wire [15:0]         maskExt_lo_437 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_437 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_437 = {maskExt_hi_437, maskExt_lo_437};
  wire [15:0]         maskExt_lo_438 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_438 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_438 = {maskExt_hi_438, maskExt_lo_438};
  wire [15:0]         maskExt_lo_439 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_439 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_439 = {maskExt_hi_439, maskExt_lo_439};
  wire [15:0]         maskExt_lo_440 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_440 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_440 = {maskExt_hi_440, maskExt_lo_440};
  wire [15:0]         maskExt_lo_441 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_441 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_441 = {maskExt_hi_441, maskExt_lo_441};
  wire [15:0]         maskExt_lo_442 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_442 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_442 = {maskExt_hi_442, maskExt_lo_442};
  wire [15:0]         maskExt_lo_443 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_443 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_443 = {maskExt_hi_443, maskExt_lo_443};
  wire [15:0]         maskExt_lo_444 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_444 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_444 = {maskExt_hi_444, maskExt_lo_444};
  wire [15:0]         maskExt_lo_445 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_445 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_445 = {maskExt_hi_445, maskExt_lo_445};
  wire [15:0]         maskExt_lo_446 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_446 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_446 = {maskExt_hi_446, maskExt_lo_446};
  wire [15:0]         maskExt_lo_447 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_447 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_447 = {maskExt_hi_447, maskExt_lo_447};
  wire [15:0]         maskExt_lo_448 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_448 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_448 = {maskExt_hi_448, maskExt_lo_448};
  wire [15:0]         maskExt_lo_449 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_449 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_449 = {maskExt_hi_449, maskExt_lo_449};
  wire [15:0]         maskExt_lo_450 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_450 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_450 = {maskExt_hi_450, maskExt_lo_450};
  wire [15:0]         maskExt_lo_451 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_451 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_451 = {maskExt_hi_451, maskExt_lo_451};
  wire [15:0]         maskExt_lo_452 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_452 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_452 = {maskExt_hi_452, maskExt_lo_452};
  wire [15:0]         maskExt_lo_453 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_453 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_453 = {maskExt_hi_453, maskExt_lo_453};
  wire [15:0]         maskExt_lo_454 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_454 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_454 = {maskExt_hi_454, maskExt_lo_454};
  wire [15:0]         maskExt_lo_455 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_455 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_455 = {maskExt_hi_455, maskExt_lo_455};
  wire [15:0]         maskExt_lo_456 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_456 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_456 = {maskExt_hi_456, maskExt_lo_456};
  wire [15:0]         maskExt_lo_457 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_457 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_457 = {maskExt_hi_457, maskExt_lo_457};
  wire [15:0]         maskExt_lo_458 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_458 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_458 = {maskExt_hi_458, maskExt_lo_458};
  wire [15:0]         maskExt_lo_459 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_459 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_459 = {maskExt_hi_459, maskExt_lo_459};
  wire [15:0]         maskExt_lo_460 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_460 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_460 = {maskExt_hi_460, maskExt_lo_460};
  wire [15:0]         maskExt_lo_461 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_461 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_461 = {maskExt_hi_461, maskExt_lo_461};
  wire [15:0]         maskExt_lo_462 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_462 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_462 = {maskExt_hi_462, maskExt_lo_462};
  wire [15:0]         maskExt_lo_463 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_463 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_463 = {maskExt_hi_463, maskExt_lo_463};
  wire [15:0]         maskExt_lo_464 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_464 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_464 = {maskExt_hi_464, maskExt_lo_464};
  wire [15:0]         maskExt_lo_465 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_465 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_465 = {maskExt_hi_465, maskExt_lo_465};
  wire [15:0]         maskExt_lo_466 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_466 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_466 = {maskExt_hi_466, maskExt_lo_466};
  wire [15:0]         maskExt_lo_467 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_467 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_467 = {maskExt_hi_467, maskExt_lo_467};
  wire [15:0]         maskExt_lo_468 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_468 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_468 = {maskExt_hi_468, maskExt_lo_468};
  wire [15:0]         maskExt_lo_469 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_469 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_469 = {maskExt_hi_469, maskExt_lo_469};
  wire [15:0]         maskExt_lo_470 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_470 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_470 = {maskExt_hi_470, maskExt_lo_470};
  wire [15:0]         maskExt_lo_471 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_471 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_471 = {maskExt_hi_471, maskExt_lo_471};
  wire [15:0]         maskExt_lo_472 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_472 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_472 = {maskExt_hi_472, maskExt_lo_472};
  wire [15:0]         maskExt_lo_473 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_473 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_473 = {maskExt_hi_473, maskExt_lo_473};
  wire [15:0]         maskExt_lo_474 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_474 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_474 = {maskExt_hi_474, maskExt_lo_474};
  wire [15:0]         maskExt_lo_475 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_475 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_475 = {maskExt_hi_475, maskExt_lo_475};
  wire [15:0]         maskExt_lo_476 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_476 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_476 = {maskExt_hi_476, maskExt_lo_476};
  wire [15:0]         maskExt_lo_477 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_477 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_477 = {maskExt_hi_477, maskExt_lo_477};
  wire [15:0]         maskExt_lo_478 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_478 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_478 = {maskExt_hi_478, maskExt_lo_478};
  wire [15:0]         maskExt_lo_479 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_479 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_479 = {maskExt_hi_479, maskExt_lo_479};
  wire [15:0]         maskExt_lo_480 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_480 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_480 = {maskExt_hi_480, maskExt_lo_480};
  wire [15:0]         maskExt_lo_481 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_481 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_481 = {maskExt_hi_481, maskExt_lo_481};
  wire [15:0]         maskExt_lo_482 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_482 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_482 = {maskExt_hi_482, maskExt_lo_482};
  wire [15:0]         maskExt_lo_483 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_483 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_483 = {maskExt_hi_483, maskExt_lo_483};
  wire [15:0]         maskExt_lo_484 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_484 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_484 = {maskExt_hi_484, maskExt_lo_484};
  wire [15:0]         maskExt_lo_485 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_485 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_485 = {maskExt_hi_485, maskExt_lo_485};
  wire [15:0]         maskExt_lo_486 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_486 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_486 = {maskExt_hi_486, maskExt_lo_486};
  wire [15:0]         maskExt_lo_487 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_487 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_487 = {maskExt_hi_487, maskExt_lo_487};
  wire [15:0]         maskExt_lo_488 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_488 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_488 = {maskExt_hi_488, maskExt_lo_488};
  wire [15:0]         maskExt_lo_489 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_489 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_489 = {maskExt_hi_489, maskExt_lo_489};
  wire [15:0]         maskExt_lo_490 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_490 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_490 = {maskExt_hi_490, maskExt_lo_490};
  wire [15:0]         maskExt_lo_491 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_491 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_491 = {maskExt_hi_491, maskExt_lo_491};
  wire [15:0]         maskExt_lo_492 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_492 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_492 = {maskExt_hi_492, maskExt_lo_492};
  wire [15:0]         maskExt_lo_493 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_493 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_493 = {maskExt_hi_493, maskExt_lo_493};
  wire [15:0]         maskExt_lo_494 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_494 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_494 = {maskExt_hi_494, maskExt_lo_494};
  wire [15:0]         maskExt_lo_495 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_495 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_495 = {maskExt_hi_495, maskExt_lo_495};
  wire [15:0]         maskExt_lo_496 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_496 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_496 = {maskExt_hi_496, maskExt_lo_496};
  wire [15:0]         maskExt_lo_497 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_497 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_497 = {maskExt_hi_497, maskExt_lo_497};
  wire [15:0]         maskExt_lo_498 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_498 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_498 = {maskExt_hi_498, maskExt_lo_498};
  wire [15:0]         maskExt_lo_499 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_499 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_499 = {maskExt_hi_499, maskExt_lo_499};
  wire [15:0]         maskExt_lo_500 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_500 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_500 = {maskExt_hi_500, maskExt_lo_500};
  wire [15:0]         maskExt_lo_501 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_501 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_501 = {maskExt_hi_501, maskExt_lo_501};
  wire [15:0]         maskExt_lo_502 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_502 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_502 = {maskExt_hi_502, maskExt_lo_502};
  wire [15:0]         maskExt_lo_503 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_503 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_503 = {maskExt_hi_503, maskExt_lo_503};
  wire [15:0]         maskExt_lo_504 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_504 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_504 = {maskExt_hi_504, maskExt_lo_504};
  wire [15:0]         maskExt_lo_505 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_505 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_505 = {maskExt_hi_505, maskExt_lo_505};
  wire [15:0]         maskExt_lo_506 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_506 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_506 = {maskExt_hi_506, maskExt_lo_506};
  wire [15:0]         maskExt_lo_507 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_507 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_507 = {maskExt_hi_507, maskExt_lo_507};
  wire [15:0]         maskExt_lo_508 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_508 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_508 = {maskExt_hi_508, maskExt_lo_508};
  wire [15:0]         maskExt_lo_509 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_509 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_509 = {maskExt_hi_509, maskExt_lo_509};
  wire [15:0]         maskExt_lo_510 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_510 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_510 = {maskExt_hi_510, maskExt_lo_510};
  wire [15:0]         maskExt_lo_511 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_511 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_511 = {maskExt_hi_511, maskExt_lo_511};
  wire [15:0]         maskExt_lo_512 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_512 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_512 = {maskExt_hi_512, maskExt_lo_512};
  wire [15:0]         maskExt_lo_513 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_513 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_513 = {maskExt_hi_513, maskExt_lo_513};
  wire [15:0]         maskExt_lo_514 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_514 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_514 = {maskExt_hi_514, maskExt_lo_514};
  wire [15:0]         maskExt_lo_515 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_515 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_515 = {maskExt_hi_515, maskExt_lo_515};
  wire [15:0]         maskExt_lo_516 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_516 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_516 = {maskExt_hi_516, maskExt_lo_516};
  wire [15:0]         maskExt_lo_517 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_517 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_517 = {maskExt_hi_517, maskExt_lo_517};
  wire [15:0]         maskExt_lo_518 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_518 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_518 = {maskExt_hi_518, maskExt_lo_518};
  wire [15:0]         maskExt_lo_519 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_519 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_519 = {maskExt_hi_519, maskExt_lo_519};
  wire [15:0]         maskExt_lo_520 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_520 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_520 = {maskExt_hi_520, maskExt_lo_520};
  wire [15:0]         maskExt_lo_521 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_521 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_521 = {maskExt_hi_521, maskExt_lo_521};
  wire [15:0]         maskExt_lo_522 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_522 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_522 = {maskExt_hi_522, maskExt_lo_522};
  wire [15:0]         maskExt_lo_523 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_523 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_523 = {maskExt_hi_523, maskExt_lo_523};
  wire [15:0]         maskExt_lo_524 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_524 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_524 = {maskExt_hi_524, maskExt_lo_524};
  wire [15:0]         maskExt_lo_525 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_525 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_525 = {maskExt_hi_525, maskExt_lo_525};
  wire [15:0]         maskExt_lo_526 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_526 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_526 = {maskExt_hi_526, maskExt_lo_526};
  wire [15:0]         maskExt_lo_527 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_527 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_527 = {maskExt_hi_527, maskExt_lo_527};
  wire [15:0]         maskExt_lo_528 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_528 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_528 = {maskExt_hi_528, maskExt_lo_528};
  wire [15:0]         maskExt_lo_529 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_529 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_529 = {maskExt_hi_529, maskExt_lo_529};
  wire [15:0]         maskExt_lo_530 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_530 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_530 = {maskExt_hi_530, maskExt_lo_530};
  wire [15:0]         maskExt_lo_531 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_531 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_531 = {maskExt_hi_531, maskExt_lo_531};
  wire [15:0]         maskExt_lo_532 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_532 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_532 = {maskExt_hi_532, maskExt_lo_532};
  wire [15:0]         maskExt_lo_533 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_533 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_533 = {maskExt_hi_533, maskExt_lo_533};
  wire [15:0]         maskExt_lo_534 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_534 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_534 = {maskExt_hi_534, maskExt_lo_534};
  wire [15:0]         maskExt_lo_535 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_535 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_535 = {maskExt_hi_535, maskExt_lo_535};
  wire [15:0]         maskExt_lo_536 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_536 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_536 = {maskExt_hi_536, maskExt_lo_536};
  wire [15:0]         maskExt_lo_537 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_537 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_537 = {maskExt_hi_537, maskExt_lo_537};
  wire [15:0]         maskExt_lo_538 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_538 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_538 = {maskExt_hi_538, maskExt_lo_538};
  wire [15:0]         maskExt_lo_539 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_539 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_539 = {maskExt_hi_539, maskExt_lo_539};
  wire [15:0]         maskExt_lo_540 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_540 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_540 = {maskExt_hi_540, maskExt_lo_540};
  wire [15:0]         maskExt_lo_541 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_541 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_541 = {maskExt_hi_541, maskExt_lo_541};
  wire [15:0]         maskExt_lo_542 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_542 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_542 = {maskExt_hi_542, maskExt_lo_542};
  wire [15:0]         maskExt_lo_543 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_543 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_543 = {maskExt_hi_543, maskExt_lo_543};
  wire [15:0]         maskExt_lo_544 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_544 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_544 = {maskExt_hi_544, maskExt_lo_544};
  wire [15:0]         maskExt_lo_545 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_545 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_545 = {maskExt_hi_545, maskExt_lo_545};
  wire [15:0]         maskExt_lo_546 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_546 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_546 = {maskExt_hi_546, maskExt_lo_546};
  wire [15:0]         maskExt_lo_547 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_547 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_547 = {maskExt_hi_547, maskExt_lo_547};
  wire [15:0]         maskExt_lo_548 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_548 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_548 = {maskExt_hi_548, maskExt_lo_548};
  wire [15:0]         maskExt_lo_549 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_549 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_549 = {maskExt_hi_549, maskExt_lo_549};
  wire [15:0]         maskExt_lo_550 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_550 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_550 = {maskExt_hi_550, maskExt_lo_550};
  wire [15:0]         maskExt_lo_551 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_551 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_551 = {maskExt_hi_551, maskExt_lo_551};
  wire [15:0]         maskExt_lo_552 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_552 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_552 = {maskExt_hi_552, maskExt_lo_552};
  wire [15:0]         maskExt_lo_553 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_553 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_553 = {maskExt_hi_553, maskExt_lo_553};
  wire [15:0]         maskExt_lo_554 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_554 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_554 = {maskExt_hi_554, maskExt_lo_554};
  wire [15:0]         maskExt_lo_555 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_555 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_555 = {maskExt_hi_555, maskExt_lo_555};
  wire [15:0]         maskExt_lo_556 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_556 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_556 = {maskExt_hi_556, maskExt_lo_556};
  wire [15:0]         maskExt_lo_557 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_557 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_557 = {maskExt_hi_557, maskExt_lo_557};
  wire [15:0]         maskExt_lo_558 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_558 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_558 = {maskExt_hi_558, maskExt_lo_558};
  wire [15:0]         maskExt_lo_559 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_559 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_559 = {maskExt_hi_559, maskExt_lo_559};
  wire [15:0]         maskExt_lo_560 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_560 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_560 = {maskExt_hi_560, maskExt_lo_560};
  wire [15:0]         maskExt_lo_561 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_561 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_561 = {maskExt_hi_561, maskExt_lo_561};
  wire [15:0]         maskExt_lo_562 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_562 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_562 = {maskExt_hi_562, maskExt_lo_562};
  wire [15:0]         maskExt_lo_563 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_563 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_563 = {maskExt_hi_563, maskExt_lo_563};
  wire [15:0]         maskExt_lo_564 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_564 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_564 = {maskExt_hi_564, maskExt_lo_564};
  wire [15:0]         maskExt_lo_565 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_565 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_565 = {maskExt_hi_565, maskExt_lo_565};
  wire [15:0]         maskExt_lo_566 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_566 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_566 = {maskExt_hi_566, maskExt_lo_566};
  wire [15:0]         maskExt_lo_567 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_567 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_567 = {maskExt_hi_567, maskExt_lo_567};
  wire [15:0]         maskExt_lo_568 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_568 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_568 = {maskExt_hi_568, maskExt_lo_568};
  wire [15:0]         maskExt_lo_569 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_569 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_569 = {maskExt_hi_569, maskExt_lo_569};
  wire [15:0]         maskExt_lo_570 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_570 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_570 = {maskExt_hi_570, maskExt_lo_570};
  wire [15:0]         maskExt_lo_571 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_571 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_571 = {maskExt_hi_571, maskExt_lo_571};
  wire [15:0]         maskExt_lo_572 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_572 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_572 = {maskExt_hi_572, maskExt_lo_572};
  wire [15:0]         maskExt_lo_573 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_573 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_573 = {maskExt_hi_573, maskExt_lo_573};
  wire [15:0]         maskExt_lo_574 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_574 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_574 = {maskExt_hi_574, maskExt_lo_574};
  wire [15:0]         maskExt_lo_575 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_575 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_575 = {maskExt_hi_575, maskExt_lo_575};
  wire [15:0]         maskExt_lo_576 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_576 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_576 = {maskExt_hi_576, maskExt_lo_576};
  wire [15:0]         maskExt_lo_577 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_577 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_577 = {maskExt_hi_577, maskExt_lo_577};
  wire [15:0]         maskExt_lo_578 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_578 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_578 = {maskExt_hi_578, maskExt_lo_578};
  wire [15:0]         maskExt_lo_579 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_579 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_579 = {maskExt_hi_579, maskExt_lo_579};
  wire [15:0]         maskExt_lo_580 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_580 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_580 = {maskExt_hi_580, maskExt_lo_580};
  wire [15:0]         maskExt_lo_581 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_581 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_581 = {maskExt_hi_581, maskExt_lo_581};
  wire [15:0]         maskExt_lo_582 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_582 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_582 = {maskExt_hi_582, maskExt_lo_582};
  wire [15:0]         maskExt_lo_583 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_583 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_583 = {maskExt_hi_583, maskExt_lo_583};
  wire [15:0]         maskExt_lo_584 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_584 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_584 = {maskExt_hi_584, maskExt_lo_584};
  wire [15:0]         maskExt_lo_585 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_585 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_585 = {maskExt_hi_585, maskExt_lo_585};
  wire [15:0]         maskExt_lo_586 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_586 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_586 = {maskExt_hi_586, maskExt_lo_586};
  wire [15:0]         maskExt_lo_587 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_587 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_587 = {maskExt_hi_587, maskExt_lo_587};
  wire [15:0]         maskExt_lo_588 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_588 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_588 = {maskExt_hi_588, maskExt_lo_588};
  wire [15:0]         maskExt_lo_589 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_589 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_589 = {maskExt_hi_589, maskExt_lo_589};
  wire [15:0]         maskExt_lo_590 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_590 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_590 = {maskExt_hi_590, maskExt_lo_590};
  wire [15:0]         maskExt_lo_591 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_591 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_591 = {maskExt_hi_591, maskExt_lo_591};
  wire [15:0]         maskExt_lo_592 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_592 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_592 = {maskExt_hi_592, maskExt_lo_592};
  wire [15:0]         maskExt_lo_593 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_593 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_593 = {maskExt_hi_593, maskExt_lo_593};
  wire [15:0]         maskExt_lo_594 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_594 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_594 = {maskExt_hi_594, maskExt_lo_594};
  wire [15:0]         maskExt_lo_595 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_595 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_595 = {maskExt_hi_595, maskExt_lo_595};
  wire [15:0]         maskExt_lo_596 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_596 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_596 = {maskExt_hi_596, maskExt_lo_596};
  wire [15:0]         maskExt_lo_597 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_597 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_597 = {maskExt_hi_597, maskExt_lo_597};
  wire [15:0]         maskExt_lo_598 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_598 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_598 = {maskExt_hi_598, maskExt_lo_598};
  wire [15:0]         maskExt_lo_599 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_599 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_599 = {maskExt_hi_599, maskExt_lo_599};
  wire [15:0]         maskExt_lo_600 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_600 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_600 = {maskExt_hi_600, maskExt_lo_600};
  wire [15:0]         maskExt_lo_601 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_601 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_601 = {maskExt_hi_601, maskExt_lo_601};
  wire [15:0]         maskExt_lo_602 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_602 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_602 = {maskExt_hi_602, maskExt_lo_602};
  wire [15:0]         maskExt_lo_603 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_603 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_603 = {maskExt_hi_603, maskExt_lo_603};
  wire [15:0]         maskExt_lo_604 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_604 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_604 = {maskExt_hi_604, maskExt_lo_604};
  wire [15:0]         maskExt_lo_605 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_605 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_605 = {maskExt_hi_605, maskExt_lo_605};
  wire [15:0]         maskExt_lo_606 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_606 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_606 = {maskExt_hi_606, maskExt_lo_606};
  wire [15:0]         maskExt_lo_607 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_607 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_607 = {maskExt_hi_607, maskExt_lo_607};
  wire [15:0]         maskExt_lo_608 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_608 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_608 = {maskExt_hi_608, maskExt_lo_608};
  wire [15:0]         maskExt_lo_609 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_609 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_609 = {maskExt_hi_609, maskExt_lo_609};
  wire [15:0]         maskExt_lo_610 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_610 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_610 = {maskExt_hi_610, maskExt_lo_610};
  wire [15:0]         maskExt_lo_611 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_611 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_611 = {maskExt_hi_611, maskExt_lo_611};
  wire [15:0]         maskExt_lo_612 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_612 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_612 = {maskExt_hi_612, maskExt_lo_612};
  wire [15:0]         maskExt_lo_613 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_613 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_613 = {maskExt_hi_613, maskExt_lo_613};
  wire [15:0]         maskExt_lo_614 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_614 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_614 = {maskExt_hi_614, maskExt_lo_614};
  wire [15:0]         maskExt_lo_615 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_615 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_615 = {maskExt_hi_615, maskExt_lo_615};
  wire [15:0]         maskExt_lo_616 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_616 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_616 = {maskExt_hi_616, maskExt_lo_616};
  wire [15:0]         maskExt_lo_617 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_617 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_617 = {maskExt_hi_617, maskExt_lo_617};
  wire [15:0]         maskExt_lo_618 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_618 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_618 = {maskExt_hi_618, maskExt_lo_618};
  wire [15:0]         maskExt_lo_619 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_619 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_619 = {maskExt_hi_619, maskExt_lo_619};
  wire [15:0]         maskExt_lo_620 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_620 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_620 = {maskExt_hi_620, maskExt_lo_620};
  wire [15:0]         maskExt_lo_621 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_621 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_621 = {maskExt_hi_621, maskExt_lo_621};
  wire [15:0]         maskExt_lo_622 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_622 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_622 = {maskExt_hi_622, maskExt_lo_622};
  wire [15:0]         maskExt_lo_623 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_623 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_623 = {maskExt_hi_623, maskExt_lo_623};
  wire [15:0]         maskExt_lo_624 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_624 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_624 = {maskExt_hi_624, maskExt_lo_624};
  wire [15:0]         maskExt_lo_625 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_625 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_625 = {maskExt_hi_625, maskExt_lo_625};
  wire [15:0]         maskExt_lo_626 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_626 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_626 = {maskExt_hi_626, maskExt_lo_626};
  wire [15:0]         maskExt_lo_627 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_627 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_627 = {maskExt_hi_627, maskExt_lo_627};
  wire [15:0]         maskExt_lo_628 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_628 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_628 = {maskExt_hi_628, maskExt_lo_628};
  wire [15:0]         maskExt_lo_629 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_629 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_629 = {maskExt_hi_629, maskExt_lo_629};
  wire [15:0]         maskExt_lo_630 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_630 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_630 = {maskExt_hi_630, maskExt_lo_630};
  wire [15:0]         maskExt_lo_631 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_631 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_631 = {maskExt_hi_631, maskExt_lo_631};
  wire [15:0]         maskExt_lo_632 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_632 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_632 = {maskExt_hi_632, maskExt_lo_632};
  wire [15:0]         maskExt_lo_633 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_633 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_633 = {maskExt_hi_633, maskExt_lo_633};
  wire [15:0]         maskExt_lo_634 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_634 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_634 = {maskExt_hi_634, maskExt_lo_634};
  wire [15:0]         maskExt_lo_635 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_635 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_635 = {maskExt_hi_635, maskExt_lo_635};
  wire [15:0]         maskExt_lo_636 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_636 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_636 = {maskExt_hi_636, maskExt_lo_636};
  wire [15:0]         maskExt_lo_637 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_637 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_637 = {maskExt_hi_637, maskExt_lo_637};
  wire [15:0]         maskExt_lo_638 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_638 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_638 = {maskExt_hi_638, maskExt_lo_638};
  wire [15:0]         maskExt_lo_639 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_639 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_639 = {maskExt_hi_639, maskExt_lo_639};
  wire [15:0]         maskExt_lo_640 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_640 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_640 = {maskExt_hi_640, maskExt_lo_640};
  wire [15:0]         maskExt_lo_641 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_641 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_641 = {maskExt_hi_641, maskExt_lo_641};
  wire [15:0]         maskExt_lo_642 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_642 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_642 = {maskExt_hi_642, maskExt_lo_642};
  wire [15:0]         maskExt_lo_643 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_643 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_643 = {maskExt_hi_643, maskExt_lo_643};
  wire [15:0]         maskExt_lo_644 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_644 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_644 = {maskExt_hi_644, maskExt_lo_644};
  wire [15:0]         maskExt_lo_645 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_645 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_645 = {maskExt_hi_645, maskExt_lo_645};
  wire [15:0]         maskExt_lo_646 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_646 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_646 = {maskExt_hi_646, maskExt_lo_646};
  wire [15:0]         maskExt_lo_647 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_647 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_647 = {maskExt_hi_647, maskExt_lo_647};
  wire [15:0]         maskExt_lo_648 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_648 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_648 = {maskExt_hi_648, maskExt_lo_648};
  wire [15:0]         maskExt_lo_649 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_649 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_649 = {maskExt_hi_649, maskExt_lo_649};
  wire [15:0]         maskExt_lo_650 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_650 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_650 = {maskExt_hi_650, maskExt_lo_650};
  wire [15:0]         maskExt_lo_651 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_651 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_651 = {maskExt_hi_651, maskExt_lo_651};
  wire [15:0]         maskExt_lo_652 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_652 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_652 = {maskExt_hi_652, maskExt_lo_652};
  wire [15:0]         maskExt_lo_653 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_653 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_653 = {maskExt_hi_653, maskExt_lo_653};
  wire [15:0]         maskExt_lo_654 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_654 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_654 = {maskExt_hi_654, maskExt_lo_654};
  wire [15:0]         maskExt_lo_655 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_655 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_655 = {maskExt_hi_655, maskExt_lo_655};
  wire [15:0]         maskExt_lo_656 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_656 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_656 = {maskExt_hi_656, maskExt_lo_656};
  wire [15:0]         maskExt_lo_657 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_657 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_657 = {maskExt_hi_657, maskExt_lo_657};
  wire [15:0]         maskExt_lo_658 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_658 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_658 = {maskExt_hi_658, maskExt_lo_658};
  wire [15:0]         maskExt_lo_659 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_659 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_659 = {maskExt_hi_659, maskExt_lo_659};
  wire [15:0]         maskExt_lo_660 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_660 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_660 = {maskExt_hi_660, maskExt_lo_660};
  wire [15:0]         maskExt_lo_661 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_661 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_661 = {maskExt_hi_661, maskExt_lo_661};
  wire [15:0]         maskExt_lo_662 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_662 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_662 = {maskExt_hi_662, maskExt_lo_662};
  wire [15:0]         maskExt_lo_663 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_663 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_663 = {maskExt_hi_663, maskExt_lo_663};
  wire [15:0]         maskExt_lo_664 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_664 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_664 = {maskExt_hi_664, maskExt_lo_664};
  wire [15:0]         maskExt_lo_665 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_665 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_665 = {maskExt_hi_665, maskExt_lo_665};
  wire [15:0]         maskExt_lo_666 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_666 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_666 = {maskExt_hi_666, maskExt_lo_666};
  wire [15:0]         maskExt_lo_667 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_667 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_667 = {maskExt_hi_667, maskExt_lo_667};
  wire [15:0]         maskExt_lo_668 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_668 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_668 = {maskExt_hi_668, maskExt_lo_668};
  wire [15:0]         maskExt_lo_669 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_669 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_669 = {maskExt_hi_669, maskExt_lo_669};
  wire [15:0]         maskExt_lo_670 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_670 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_670 = {maskExt_hi_670, maskExt_lo_670};
  wire [15:0]         maskExt_lo_671 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_671 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_671 = {maskExt_hi_671, maskExt_lo_671};
  wire [15:0]         maskExt_lo_672 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_672 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_672 = {maskExt_hi_672, maskExt_lo_672};
  wire [15:0]         maskExt_lo_673 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_673 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_673 = {maskExt_hi_673, maskExt_lo_673};
  wire [15:0]         maskExt_lo_674 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_674 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_674 = {maskExt_hi_674, maskExt_lo_674};
  wire [15:0]         maskExt_lo_675 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_675 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_675 = {maskExt_hi_675, maskExt_lo_675};
  wire [15:0]         maskExt_lo_676 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_676 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_676 = {maskExt_hi_676, maskExt_lo_676};
  wire [15:0]         maskExt_lo_677 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_677 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_677 = {maskExt_hi_677, maskExt_lo_677};
  wire [15:0]         maskExt_lo_678 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_678 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_678 = {maskExt_hi_678, maskExt_lo_678};
  wire [15:0]         maskExt_lo_679 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_679 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_679 = {maskExt_hi_679, maskExt_lo_679};
  wire [15:0]         maskExt_lo_680 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_680 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_680 = {maskExt_hi_680, maskExt_lo_680};
  wire [15:0]         maskExt_lo_681 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_681 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_681 = {maskExt_hi_681, maskExt_lo_681};
  wire [15:0]         maskExt_lo_682 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_682 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_682 = {maskExt_hi_682, maskExt_lo_682};
  wire [15:0]         maskExt_lo_683 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_683 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_683 = {maskExt_hi_683, maskExt_lo_683};
  wire [15:0]         maskExt_lo_684 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_684 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_684 = {maskExt_hi_684, maskExt_lo_684};
  wire [15:0]         maskExt_lo_685 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_685 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_685 = {maskExt_hi_685, maskExt_lo_685};
  wire [15:0]         maskExt_lo_686 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_686 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_686 = {maskExt_hi_686, maskExt_lo_686};
  wire [15:0]         maskExt_lo_687 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_687 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_687 = {maskExt_hi_687, maskExt_lo_687};
  wire [15:0]         maskExt_lo_688 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_688 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_688 = {maskExt_hi_688, maskExt_lo_688};
  wire [15:0]         maskExt_lo_689 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_689 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_689 = {maskExt_hi_689, maskExt_lo_689};
  wire [15:0]         maskExt_lo_690 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_690 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_690 = {maskExt_hi_690, maskExt_lo_690};
  wire [15:0]         maskExt_lo_691 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_691 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_691 = {maskExt_hi_691, maskExt_lo_691};
  wire [15:0]         maskExt_lo_692 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_692 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_692 = {maskExt_hi_692, maskExt_lo_692};
  wire [15:0]         maskExt_lo_693 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_693 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_693 = {maskExt_hi_693, maskExt_lo_693};
  wire [15:0]         maskExt_lo_694 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_694 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_694 = {maskExt_hi_694, maskExt_lo_694};
  wire [15:0]         maskExt_lo_695 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_695 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_695 = {maskExt_hi_695, maskExt_lo_695};
  wire [15:0]         maskExt_lo_696 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_696 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_696 = {maskExt_hi_696, maskExt_lo_696};
  wire [15:0]         maskExt_lo_697 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_697 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_697 = {maskExt_hi_697, maskExt_lo_697};
  wire [15:0]         maskExt_lo_698 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_698 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_698 = {maskExt_hi_698, maskExt_lo_698};
  wire [15:0]         maskExt_lo_699 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_699 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_699 = {maskExt_hi_699, maskExt_lo_699};
  wire [15:0]         maskExt_lo_700 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_700 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_700 = {maskExt_hi_700, maskExt_lo_700};
  wire [15:0]         maskExt_lo_701 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_701 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_701 = {maskExt_hi_701, maskExt_lo_701};
  wire [15:0]         maskExt_lo_702 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_702 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_702 = {maskExt_hi_702, maskExt_lo_702};
  wire [15:0]         maskExt_lo_703 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_703 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_703 = {maskExt_hi_703, maskExt_lo_703};
  wire [15:0]         maskExt_lo_704 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_704 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_704 = {maskExt_hi_704, maskExt_lo_704};
  wire [15:0]         maskExt_lo_705 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_705 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_705 = {maskExt_hi_705, maskExt_lo_705};
  wire [15:0]         maskExt_lo_706 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_706 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_706 = {maskExt_hi_706, maskExt_lo_706};
  wire [15:0]         maskExt_lo_707 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_707 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_707 = {maskExt_hi_707, maskExt_lo_707};
  wire [15:0]         maskExt_lo_708 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_708 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_708 = {maskExt_hi_708, maskExt_lo_708};
  wire [15:0]         maskExt_lo_709 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_709 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_709 = {maskExt_hi_709, maskExt_lo_709};
  wire [15:0]         maskExt_lo_710 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_710 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_710 = {maskExt_hi_710, maskExt_lo_710};
  wire [15:0]         maskExt_lo_711 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_711 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_711 = {maskExt_hi_711, maskExt_lo_711};
  wire [15:0]         maskExt_lo_712 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_712 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_712 = {maskExt_hi_712, maskExt_lo_712};
  wire [15:0]         maskExt_lo_713 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_713 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_713 = {maskExt_hi_713, maskExt_lo_713};
  wire [15:0]         maskExt_lo_714 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_714 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_714 = {maskExt_hi_714, maskExt_lo_714};
  wire [15:0]         maskExt_lo_715 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_715 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_715 = {maskExt_hi_715, maskExt_lo_715};
  wire [15:0]         maskExt_lo_716 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_716 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_716 = {maskExt_hi_716, maskExt_lo_716};
  wire [15:0]         maskExt_lo_717 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_717 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_717 = {maskExt_hi_717, maskExt_lo_717};
  wire [15:0]         maskExt_lo_718 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_718 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_718 = {maskExt_hi_718, maskExt_lo_718};
  wire [15:0]         maskExt_lo_719 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_719 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_719 = {maskExt_hi_719, maskExt_lo_719};
  wire [15:0]         maskExt_lo_720 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_720 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_720 = {maskExt_hi_720, maskExt_lo_720};
  wire [15:0]         maskExt_lo_721 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_721 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_721 = {maskExt_hi_721, maskExt_lo_721};
  wire [15:0]         maskExt_lo_722 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_722 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_722 = {maskExt_hi_722, maskExt_lo_722};
  wire [15:0]         maskExt_lo_723 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_723 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_723 = {maskExt_hi_723, maskExt_lo_723};
  wire [15:0]         maskExt_lo_724 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_724 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_724 = {maskExt_hi_724, maskExt_lo_724};
  wire [15:0]         maskExt_lo_725 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_725 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_725 = {maskExt_hi_725, maskExt_lo_725};
  wire [15:0]         maskExt_lo_726 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_726 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_726 = {maskExt_hi_726, maskExt_lo_726};
  wire [15:0]         maskExt_lo_727 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_727 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_727 = {maskExt_hi_727, maskExt_lo_727};
  wire [15:0]         maskExt_lo_728 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_728 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_728 = {maskExt_hi_728, maskExt_lo_728};
  wire [15:0]         maskExt_lo_729 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_729 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_729 = {maskExt_hi_729, maskExt_lo_729};
  wire [15:0]         maskExt_lo_730 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_730 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_730 = {maskExt_hi_730, maskExt_lo_730};
  wire [15:0]         maskExt_lo_731 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_731 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_731 = {maskExt_hi_731, maskExt_lo_731};
  wire [15:0]         maskExt_lo_732 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_732 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_732 = {maskExt_hi_732, maskExt_lo_732};
  wire [15:0]         maskExt_lo_733 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_733 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_733 = {maskExt_hi_733, maskExt_lo_733};
  wire [15:0]         maskExt_lo_734 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_734 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_734 = {maskExt_hi_734, maskExt_lo_734};
  wire [15:0]         maskExt_lo_735 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_735 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_735 = {maskExt_hi_735, maskExt_lo_735};
  wire [15:0]         maskExt_lo_736 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_736 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_736 = {maskExt_hi_736, maskExt_lo_736};
  wire [15:0]         maskExt_lo_737 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_737 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_737 = {maskExt_hi_737, maskExt_lo_737};
  wire [15:0]         maskExt_lo_738 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_738 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_738 = {maskExt_hi_738, maskExt_lo_738};
  wire [15:0]         maskExt_lo_739 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_739 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_739 = {maskExt_hi_739, maskExt_lo_739};
  wire [15:0]         maskExt_lo_740 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_740 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_740 = {maskExt_hi_740, maskExt_lo_740};
  wire [15:0]         maskExt_lo_741 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_741 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_741 = {maskExt_hi_741, maskExt_lo_741};
  wire [15:0]         maskExt_lo_742 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_742 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_742 = {maskExt_hi_742, maskExt_lo_742};
  wire [15:0]         maskExt_lo_743 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_743 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_743 = {maskExt_hi_743, maskExt_lo_743};
  wire [15:0]         maskExt_lo_744 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_744 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_744 = {maskExt_hi_744, maskExt_lo_744};
  wire [15:0]         maskExt_lo_745 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_745 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_745 = {maskExt_hi_745, maskExt_lo_745};
  wire [15:0]         maskExt_lo_746 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_746 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_746 = {maskExt_hi_746, maskExt_lo_746};
  wire [15:0]         maskExt_lo_747 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_747 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_747 = {maskExt_hi_747, maskExt_lo_747};
  wire [15:0]         maskExt_lo_748 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_748 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_748 = {maskExt_hi_748, maskExt_lo_748};
  wire [15:0]         maskExt_lo_749 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_749 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_749 = {maskExt_hi_749, maskExt_lo_749};
  wire [15:0]         maskExt_lo_750 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_750 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_750 = {maskExt_hi_750, maskExt_lo_750};
  wire [15:0]         maskExt_lo_751 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_751 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_751 = {maskExt_hi_751, maskExt_lo_751};
  wire [15:0]         maskExt_lo_752 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_752 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_752 = {maskExt_hi_752, maskExt_lo_752};
  wire [15:0]         maskExt_lo_753 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_753 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_753 = {maskExt_hi_753, maskExt_lo_753};
  wire [15:0]         maskExt_lo_754 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_754 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_754 = {maskExt_hi_754, maskExt_lo_754};
  wire [15:0]         maskExt_lo_755 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_755 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_755 = {maskExt_hi_755, maskExt_lo_755};
  wire [15:0]         maskExt_lo_756 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_756 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_756 = {maskExt_hi_756, maskExt_lo_756};
  wire [15:0]         maskExt_lo_757 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_757 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_757 = {maskExt_hi_757, maskExt_lo_757};
  wire [15:0]         maskExt_lo_758 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_758 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_758 = {maskExt_hi_758, maskExt_lo_758};
  wire [15:0]         maskExt_lo_759 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_759 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_759 = {maskExt_hi_759, maskExt_lo_759};
  wire [15:0]         maskExt_lo_760 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_760 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_760 = {maskExt_hi_760, maskExt_lo_760};
  wire [15:0]         maskExt_lo_761 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_761 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_761 = {maskExt_hi_761, maskExt_lo_761};
  wire [15:0]         maskExt_lo_762 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_762 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_762 = {maskExt_hi_762, maskExt_lo_762};
  wire [15:0]         maskExt_lo_763 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_763 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_763 = {maskExt_hi_763, maskExt_lo_763};
  wire [15:0]         maskExt_lo_764 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_764 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_764 = {maskExt_hi_764, maskExt_lo_764};
  wire [15:0]         maskExt_lo_765 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_765 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_765 = {maskExt_hi_765, maskExt_lo_765};
  wire [15:0]         maskExt_lo_766 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_766 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_766 = {maskExt_hi_766, maskExt_lo_766};
  wire [15:0]         maskExt_lo_767 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_767 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_767 = {maskExt_hi_767, maskExt_lo_767};
  wire [15:0]         maskExt_lo_768 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_768 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_768 = {maskExt_hi_768, maskExt_lo_768};
  wire [15:0]         maskExt_lo_769 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_769 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_769 = {maskExt_hi_769, maskExt_lo_769};
  wire [15:0]         maskExt_lo_770 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_770 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_770 = {maskExt_hi_770, maskExt_lo_770};
  wire [15:0]         maskExt_lo_771 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_771 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_771 = {maskExt_hi_771, maskExt_lo_771};
  wire [15:0]         maskExt_lo_772 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_772 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_772 = {maskExt_hi_772, maskExt_lo_772};
  wire [15:0]         maskExt_lo_773 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_773 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_773 = {maskExt_hi_773, maskExt_lo_773};
  wire [15:0]         maskExt_lo_774 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_774 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_774 = {maskExt_hi_774, maskExt_lo_774};
  wire [15:0]         maskExt_lo_775 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_775 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_775 = {maskExt_hi_775, maskExt_lo_775};
  wire [15:0]         maskExt_lo_776 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_776 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_776 = {maskExt_hi_776, maskExt_lo_776};
  wire [15:0]         maskExt_lo_777 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_777 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_777 = {maskExt_hi_777, maskExt_lo_777};
  wire [15:0]         maskExt_lo_778 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_778 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_778 = {maskExt_hi_778, maskExt_lo_778};
  wire [15:0]         maskExt_lo_779 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_779 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_779 = {maskExt_hi_779, maskExt_lo_779};
  wire [15:0]         maskExt_lo_780 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_780 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_780 = {maskExt_hi_780, maskExt_lo_780};
  wire [15:0]         maskExt_lo_781 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_781 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_781 = {maskExt_hi_781, maskExt_lo_781};
  wire [15:0]         maskExt_lo_782 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_782 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_782 = {maskExt_hi_782, maskExt_lo_782};
  wire [15:0]         maskExt_lo_783 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_783 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_783 = {maskExt_hi_783, maskExt_lo_783};
  wire [15:0]         maskExt_lo_784 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_784 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_784 = {maskExt_hi_784, maskExt_lo_784};
  wire [15:0]         maskExt_lo_785 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_785 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_785 = {maskExt_hi_785, maskExt_lo_785};
  wire [15:0]         maskExt_lo_786 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_786 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_786 = {maskExt_hi_786, maskExt_lo_786};
  wire [15:0]         maskExt_lo_787 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_787 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_787 = {maskExt_hi_787, maskExt_lo_787};
  wire [15:0]         maskExt_lo_788 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_788 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_788 = {maskExt_hi_788, maskExt_lo_788};
  wire [15:0]         maskExt_lo_789 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_789 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_789 = {maskExt_hi_789, maskExt_lo_789};
  wire [15:0]         maskExt_lo_790 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_790 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_790 = {maskExt_hi_790, maskExt_lo_790};
  wire [15:0]         maskExt_lo_791 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_791 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_791 = {maskExt_hi_791, maskExt_lo_791};
  wire [15:0]         maskExt_lo_792 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_792 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_792 = {maskExt_hi_792, maskExt_lo_792};
  wire [15:0]         maskExt_lo_793 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_793 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_793 = {maskExt_hi_793, maskExt_lo_793};
  wire [15:0]         maskExt_lo_794 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_794 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_794 = {maskExt_hi_794, maskExt_lo_794};
  wire [15:0]         maskExt_lo_795 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_795 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_795 = {maskExt_hi_795, maskExt_lo_795};
  wire [15:0]         maskExt_lo_796 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_796 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_796 = {maskExt_hi_796, maskExt_lo_796};
  wire [15:0]         maskExt_lo_797 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_797 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_797 = {maskExt_hi_797, maskExt_lo_797};
  wire [15:0]         maskExt_lo_798 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_798 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_798 = {maskExt_hi_798, maskExt_lo_798};
  wire [15:0]         maskExt_lo_799 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_799 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_799 = {maskExt_hi_799, maskExt_lo_799};
  wire [15:0]         maskExt_lo_800 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_800 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_800 = {maskExt_hi_800, maskExt_lo_800};
  wire [15:0]         maskExt_lo_801 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_801 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_801 = {maskExt_hi_801, maskExt_lo_801};
  wire [15:0]         maskExt_lo_802 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_802 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_802 = {maskExt_hi_802, maskExt_lo_802};
  wire [15:0]         maskExt_lo_803 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_803 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_803 = {maskExt_hi_803, maskExt_lo_803};
  wire [15:0]         maskExt_lo_804 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_804 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_804 = {maskExt_hi_804, maskExt_lo_804};
  wire [15:0]         maskExt_lo_805 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_805 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_805 = {maskExt_hi_805, maskExt_lo_805};
  wire [15:0]         maskExt_lo_806 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_806 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_806 = {maskExt_hi_806, maskExt_lo_806};
  wire [15:0]         maskExt_lo_807 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_807 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_807 = {maskExt_hi_807, maskExt_lo_807};
  wire [15:0]         maskExt_lo_808 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_808 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_808 = {maskExt_hi_808, maskExt_lo_808};
  wire [15:0]         maskExt_lo_809 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_809 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_809 = {maskExt_hi_809, maskExt_lo_809};
  wire [15:0]         maskExt_lo_810 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_810 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_810 = {maskExt_hi_810, maskExt_lo_810};
  wire [15:0]         maskExt_lo_811 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_811 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_811 = {maskExt_hi_811, maskExt_lo_811};
  wire [15:0]         maskExt_lo_812 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_812 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_812 = {maskExt_hi_812, maskExt_lo_812};
  wire [15:0]         maskExt_lo_813 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_813 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_813 = {maskExt_hi_813, maskExt_lo_813};
  wire [15:0]         maskExt_lo_814 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_814 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_814 = {maskExt_hi_814, maskExt_lo_814};
  wire [15:0]         maskExt_lo_815 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_815 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_815 = {maskExt_hi_815, maskExt_lo_815};
  wire [15:0]         maskExt_lo_816 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_816 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_816 = {maskExt_hi_816, maskExt_lo_816};
  wire [15:0]         maskExt_lo_817 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_817 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_817 = {maskExt_hi_817, maskExt_lo_817};
  wire [15:0]         maskExt_lo_818 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_818 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_818 = {maskExt_hi_818, maskExt_lo_818};
  wire [15:0]         maskExt_lo_819 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_819 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_819 = {maskExt_hi_819, maskExt_lo_819};
  wire [15:0]         maskExt_lo_820 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_820 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_820 = {maskExt_hi_820, maskExt_lo_820};
  wire [15:0]         maskExt_lo_821 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_821 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_821 = {maskExt_hi_821, maskExt_lo_821};
  wire [15:0]         maskExt_lo_822 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_822 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_822 = {maskExt_hi_822, maskExt_lo_822};
  wire [15:0]         maskExt_lo_823 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_823 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_823 = {maskExt_hi_823, maskExt_lo_823};
  wire [15:0]         maskExt_lo_824 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_824 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_824 = {maskExt_hi_824, maskExt_lo_824};
  wire [15:0]         maskExt_lo_825 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_825 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_825 = {maskExt_hi_825, maskExt_lo_825};
  wire [15:0]         maskExt_lo_826 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_826 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_826 = {maskExt_hi_826, maskExt_lo_826};
  wire [15:0]         maskExt_lo_827 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_827 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_827 = {maskExt_hi_827, maskExt_lo_827};
  wire [15:0]         maskExt_lo_828 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_828 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_828 = {maskExt_hi_828, maskExt_lo_828};
  wire [15:0]         maskExt_lo_829 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_829 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_829 = {maskExt_hi_829, maskExt_lo_829};
  wire [15:0]         maskExt_lo_830 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_830 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_830 = {maskExt_hi_830, maskExt_lo_830};
  wire [15:0]         maskExt_lo_831 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_831 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_831 = {maskExt_hi_831, maskExt_lo_831};
  wire [15:0]         maskExt_lo_832 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_832 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_832 = {maskExt_hi_832, maskExt_lo_832};
  wire [15:0]         maskExt_lo_833 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_833 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_833 = {maskExt_hi_833, maskExt_lo_833};
  wire [15:0]         maskExt_lo_834 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_834 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_834 = {maskExt_hi_834, maskExt_lo_834};
  wire [15:0]         maskExt_lo_835 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_835 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_835 = {maskExt_hi_835, maskExt_lo_835};
  wire [15:0]         maskExt_lo_836 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_836 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_836 = {maskExt_hi_836, maskExt_lo_836};
  wire [15:0]         maskExt_lo_837 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_837 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_837 = {maskExt_hi_837, maskExt_lo_837};
  wire [15:0]         maskExt_lo_838 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_838 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_838 = {maskExt_hi_838, maskExt_lo_838};
  wire [15:0]         maskExt_lo_839 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_839 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_839 = {maskExt_hi_839, maskExt_lo_839};
  wire [15:0]         maskExt_lo_840 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_840 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_840 = {maskExt_hi_840, maskExt_lo_840};
  wire [15:0]         maskExt_lo_841 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_841 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_841 = {maskExt_hi_841, maskExt_lo_841};
  wire [15:0]         maskExt_lo_842 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_842 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_842 = {maskExt_hi_842, maskExt_lo_842};
  wire [15:0]         maskExt_lo_843 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_843 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_843 = {maskExt_hi_843, maskExt_lo_843};
  wire [15:0]         maskExt_lo_844 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_844 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_844 = {maskExt_hi_844, maskExt_lo_844};
  wire [15:0]         maskExt_lo_845 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_845 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_845 = {maskExt_hi_845, maskExt_lo_845};
  wire [15:0]         maskExt_lo_846 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_846 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_846 = {maskExt_hi_846, maskExt_lo_846};
  wire [15:0]         maskExt_lo_847 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_847 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_847 = {maskExt_hi_847, maskExt_lo_847};
  wire [15:0]         maskExt_lo_848 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_848 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_848 = {maskExt_hi_848, maskExt_lo_848};
  wire [15:0]         maskExt_lo_849 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_849 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_849 = {maskExt_hi_849, maskExt_lo_849};
  wire [15:0]         maskExt_lo_850 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_850 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_850 = {maskExt_hi_850, maskExt_lo_850};
  wire [15:0]         maskExt_lo_851 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_851 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_851 = {maskExt_hi_851, maskExt_lo_851};
  wire [15:0]         maskExt_lo_852 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_852 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_852 = {maskExt_hi_852, maskExt_lo_852};
  wire [15:0]         maskExt_lo_853 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_853 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_853 = {maskExt_hi_853, maskExt_lo_853};
  wire [15:0]         maskExt_lo_854 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_854 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_854 = {maskExt_hi_854, maskExt_lo_854};
  wire [15:0]         maskExt_lo_855 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_855 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_855 = {maskExt_hi_855, maskExt_lo_855};
  wire [15:0]         maskExt_lo_856 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_856 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_856 = {maskExt_hi_856, maskExt_lo_856};
  wire [15:0]         maskExt_lo_857 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_857 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_857 = {maskExt_hi_857, maskExt_lo_857};
  wire [15:0]         maskExt_lo_858 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_858 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_858 = {maskExt_hi_858, maskExt_lo_858};
  wire [15:0]         maskExt_lo_859 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_859 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_859 = {maskExt_hi_859, maskExt_lo_859};
  wire [15:0]         maskExt_lo_860 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_860 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_860 = {maskExt_hi_860, maskExt_lo_860};
  wire [15:0]         maskExt_lo_861 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_861 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_861 = {maskExt_hi_861, maskExt_lo_861};
  wire [15:0]         maskExt_lo_862 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_862 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_862 = {maskExt_hi_862, maskExt_lo_862};
  wire [15:0]         maskExt_lo_863 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_863 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_863 = {maskExt_hi_863, maskExt_lo_863};
  wire [15:0]         maskExt_lo_864 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_864 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_864 = {maskExt_hi_864, maskExt_lo_864};
  wire [15:0]         maskExt_lo_865 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_865 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_865 = {maskExt_hi_865, maskExt_lo_865};
  wire [15:0]         maskExt_lo_866 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_866 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_866 = {maskExt_hi_866, maskExt_lo_866};
  wire [15:0]         maskExt_lo_867 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_867 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_867 = {maskExt_hi_867, maskExt_lo_867};
  wire [15:0]         maskExt_lo_868 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_868 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_868 = {maskExt_hi_868, maskExt_lo_868};
  wire [15:0]         maskExt_lo_869 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_869 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_869 = {maskExt_hi_869, maskExt_lo_869};
  wire [15:0]         maskExt_lo_870 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_870 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_870 = {maskExt_hi_870, maskExt_lo_870};
  wire [15:0]         maskExt_lo_871 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_871 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_871 = {maskExt_hi_871, maskExt_lo_871};
  wire [15:0]         maskExt_lo_872 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_872 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_872 = {maskExt_hi_872, maskExt_lo_872};
  wire [15:0]         maskExt_lo_873 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_873 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_873 = {maskExt_hi_873, maskExt_lo_873};
  wire [15:0]         maskExt_lo_874 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_874 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_874 = {maskExt_hi_874, maskExt_lo_874};
  wire [15:0]         maskExt_lo_875 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_875 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_875 = {maskExt_hi_875, maskExt_lo_875};
  wire [15:0]         maskExt_lo_876 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_876 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_876 = {maskExt_hi_876, maskExt_lo_876};
  wire [15:0]         maskExt_lo_877 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_877 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_877 = {maskExt_hi_877, maskExt_lo_877};
  wire [15:0]         maskExt_lo_878 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_878 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_878 = {maskExt_hi_878, maskExt_lo_878};
  wire [15:0]         maskExt_lo_879 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_879 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_879 = {maskExt_hi_879, maskExt_lo_879};
  wire [15:0]         maskExt_lo_880 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_880 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_880 = {maskExt_hi_880, maskExt_lo_880};
  wire [15:0]         maskExt_lo_881 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_881 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_881 = {maskExt_hi_881, maskExt_lo_881};
  wire [15:0]         maskExt_lo_882 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_882 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_882 = {maskExt_hi_882, maskExt_lo_882};
  wire [15:0]         maskExt_lo_883 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_883 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_883 = {maskExt_hi_883, maskExt_lo_883};
  wire [15:0]         maskExt_lo_884 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_884 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_884 = {maskExt_hi_884, maskExt_lo_884};
  wire [15:0]         maskExt_lo_885 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_885 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_885 = {maskExt_hi_885, maskExt_lo_885};
  wire [15:0]         maskExt_lo_886 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_886 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_886 = {maskExt_hi_886, maskExt_lo_886};
  wire [15:0]         maskExt_lo_887 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_887 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_887 = {maskExt_hi_887, maskExt_lo_887};
  wire [15:0]         maskExt_lo_888 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_888 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_888 = {maskExt_hi_888, maskExt_lo_888};
  wire [15:0]         maskExt_lo_889 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_889 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_889 = {maskExt_hi_889, maskExt_lo_889};
  wire [15:0]         maskExt_lo_890 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_890 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_890 = {maskExt_hi_890, maskExt_lo_890};
  wire [15:0]         maskExt_lo_891 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_891 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_891 = {maskExt_hi_891, maskExt_lo_891};
  wire [15:0]         maskExt_lo_892 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_892 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_892 = {maskExt_hi_892, maskExt_lo_892};
  wire [15:0]         maskExt_lo_893 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_893 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_893 = {maskExt_hi_893, maskExt_lo_893};
  wire [15:0]         maskExt_lo_894 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_894 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_894 = {maskExt_hi_894, maskExt_lo_894};
  wire [15:0]         maskExt_lo_895 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_895 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_895 = {maskExt_hi_895, maskExt_lo_895};
  wire [15:0]         maskExt_lo_896 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_896 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_896 = {maskExt_hi_896, maskExt_lo_896};
  wire [15:0]         maskExt_lo_897 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_897 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_897 = {maskExt_hi_897, maskExt_lo_897};
  wire [15:0]         maskExt_lo_898 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_898 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_898 = {maskExt_hi_898, maskExt_lo_898};
  wire [15:0]         maskExt_lo_899 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_899 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_899 = {maskExt_hi_899, maskExt_lo_899};
  wire [15:0]         maskExt_lo_900 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_900 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_900 = {maskExt_hi_900, maskExt_lo_900};
  wire [15:0]         maskExt_lo_901 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_901 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_901 = {maskExt_hi_901, maskExt_lo_901};
  wire [15:0]         maskExt_lo_902 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_902 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_902 = {maskExt_hi_902, maskExt_lo_902};
  wire [15:0]         maskExt_lo_903 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_903 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_903 = {maskExt_hi_903, maskExt_lo_903};
  wire [15:0]         maskExt_lo_904 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_904 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_904 = {maskExt_hi_904, maskExt_lo_904};
  wire [15:0]         maskExt_lo_905 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_905 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_905 = {maskExt_hi_905, maskExt_lo_905};
  wire [15:0]         maskExt_lo_906 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_906 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_906 = {maskExt_hi_906, maskExt_lo_906};
  wire [15:0]         maskExt_lo_907 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_907 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_907 = {maskExt_hi_907, maskExt_lo_907};
  wire [15:0]         maskExt_lo_908 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_908 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_908 = {maskExt_hi_908, maskExt_lo_908};
  wire [15:0]         maskExt_lo_909 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_909 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_909 = {maskExt_hi_909, maskExt_lo_909};
  wire [15:0]         maskExt_lo_910 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_910 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_910 = {maskExt_hi_910, maskExt_lo_910};
  wire [15:0]         maskExt_lo_911 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_911 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_911 = {maskExt_hi_911, maskExt_lo_911};
  wire [15:0]         maskExt_lo_912 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_912 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_912 = {maskExt_hi_912, maskExt_lo_912};
  wire [15:0]         maskExt_lo_913 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_913 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_913 = {maskExt_hi_913, maskExt_lo_913};
  wire [15:0]         maskExt_lo_914 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_914 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_914 = {maskExt_hi_914, maskExt_lo_914};
  wire [15:0]         maskExt_lo_915 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_915 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_915 = {maskExt_hi_915, maskExt_lo_915};
  wire [15:0]         maskExt_lo_916 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_916 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_916 = {maskExt_hi_916, maskExt_lo_916};
  wire [15:0]         maskExt_lo_917 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_917 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_917 = {maskExt_hi_917, maskExt_lo_917};
  wire [15:0]         maskExt_lo_918 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_918 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_918 = {maskExt_hi_918, maskExt_lo_918};
  wire [15:0]         maskExt_lo_919 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_919 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_919 = {maskExt_hi_919, maskExt_lo_919};
  wire [15:0]         maskExt_lo_920 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_920 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_920 = {maskExt_hi_920, maskExt_lo_920};
  wire [15:0]         maskExt_lo_921 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_921 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_921 = {maskExt_hi_921, maskExt_lo_921};
  wire [15:0]         maskExt_lo_922 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_922 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_922 = {maskExt_hi_922, maskExt_lo_922};
  wire [15:0]         maskExt_lo_923 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_923 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_923 = {maskExt_hi_923, maskExt_lo_923};
  wire [15:0]         maskExt_lo_924 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_924 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_924 = {maskExt_hi_924, maskExt_lo_924};
  wire [15:0]         maskExt_lo_925 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_925 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_925 = {maskExt_hi_925, maskExt_lo_925};
  wire [15:0]         maskExt_lo_926 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_926 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_926 = {maskExt_hi_926, maskExt_lo_926};
  wire [15:0]         maskExt_lo_927 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_927 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_927 = {maskExt_hi_927, maskExt_lo_927};
  wire [15:0]         maskExt_lo_928 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_928 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_928 = {maskExt_hi_928, maskExt_lo_928};
  wire [15:0]         maskExt_lo_929 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_929 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_929 = {maskExt_hi_929, maskExt_lo_929};
  wire [15:0]         maskExt_lo_930 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_930 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_930 = {maskExt_hi_930, maskExt_lo_930};
  wire [15:0]         maskExt_lo_931 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_931 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_931 = {maskExt_hi_931, maskExt_lo_931};
  wire [15:0]         maskExt_lo_932 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_932 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_932 = {maskExt_hi_932, maskExt_lo_932};
  wire [15:0]         maskExt_lo_933 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_933 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_933 = {maskExt_hi_933, maskExt_lo_933};
  wire [15:0]         maskExt_lo_934 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_934 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_934 = {maskExt_hi_934, maskExt_lo_934};
  wire [15:0]         maskExt_lo_935 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_935 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_935 = {maskExt_hi_935, maskExt_lo_935};
  wire [15:0]         maskExt_lo_936 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_936 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_936 = {maskExt_hi_936, maskExt_lo_936};
  wire [15:0]         maskExt_lo_937 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_937 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_937 = {maskExt_hi_937, maskExt_lo_937};
  wire [15:0]         maskExt_lo_938 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_938 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_938 = {maskExt_hi_938, maskExt_lo_938};
  wire [15:0]         maskExt_lo_939 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_939 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_939 = {maskExt_hi_939, maskExt_lo_939};
  wire [15:0]         maskExt_lo_940 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_940 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_940 = {maskExt_hi_940, maskExt_lo_940};
  wire [15:0]         maskExt_lo_941 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_941 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_941 = {maskExt_hi_941, maskExt_lo_941};
  wire [15:0]         maskExt_lo_942 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_942 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_942 = {maskExt_hi_942, maskExt_lo_942};
  wire [15:0]         maskExt_lo_943 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_943 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_943 = {maskExt_hi_943, maskExt_lo_943};
  wire [15:0]         maskExt_lo_944 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_944 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_944 = {maskExt_hi_944, maskExt_lo_944};
  wire [15:0]         maskExt_lo_945 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_945 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_945 = {maskExt_hi_945, maskExt_lo_945};
  wire [15:0]         maskExt_lo_946 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_946 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_946 = {maskExt_hi_946, maskExt_lo_946};
  wire [15:0]         maskExt_lo_947 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_947 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_947 = {maskExt_hi_947, maskExt_lo_947};
  wire [15:0]         maskExt_lo_948 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_948 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_948 = {maskExt_hi_948, maskExt_lo_948};
  wire [15:0]         maskExt_lo_949 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_949 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_949 = {maskExt_hi_949, maskExt_lo_949};
  wire [15:0]         maskExt_lo_950 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_950 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_950 = {maskExt_hi_950, maskExt_lo_950};
  wire [15:0]         maskExt_lo_951 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_951 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_951 = {maskExt_hi_951, maskExt_lo_951};
  wire [15:0]         maskExt_lo_952 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_952 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_952 = {maskExt_hi_952, maskExt_lo_952};
  wire [15:0]         maskExt_lo_953 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_953 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_953 = {maskExt_hi_953, maskExt_lo_953};
  wire [15:0]         maskExt_lo_954 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_954 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_954 = {maskExt_hi_954, maskExt_lo_954};
  wire [15:0]         maskExt_lo_955 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_955 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_955 = {maskExt_hi_955, maskExt_lo_955};
  wire [15:0]         maskExt_lo_956 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_956 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_956 = {maskExt_hi_956, maskExt_lo_956};
  wire [15:0]         maskExt_lo_957 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_957 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_957 = {maskExt_hi_957, maskExt_lo_957};
  wire [15:0]         maskExt_lo_958 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_958 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_958 = {maskExt_hi_958, maskExt_lo_958};
  wire [15:0]         maskExt_lo_959 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_959 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_959 = {maskExt_hi_959, maskExt_lo_959};
  wire [15:0]         maskExt_lo_960 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_960 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_960 = {maskExt_hi_960, maskExt_lo_960};
  wire [15:0]         maskExt_lo_961 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_961 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_961 = {maskExt_hi_961, maskExt_lo_961};
  wire [15:0]         maskExt_lo_962 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_962 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_962 = {maskExt_hi_962, maskExt_lo_962};
  wire [15:0]         maskExt_lo_963 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_963 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_963 = {maskExt_hi_963, maskExt_lo_963};
  wire [15:0]         maskExt_lo_964 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_964 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_964 = {maskExt_hi_964, maskExt_lo_964};
  wire [15:0]         maskExt_lo_965 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_965 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_965 = {maskExt_hi_965, maskExt_lo_965};
  wire [15:0]         maskExt_lo_966 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_966 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_966 = {maskExt_hi_966, maskExt_lo_966};
  wire [15:0]         maskExt_lo_967 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_967 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_967 = {maskExt_hi_967, maskExt_lo_967};
  wire [15:0]         maskExt_lo_968 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_968 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_968 = {maskExt_hi_968, maskExt_lo_968};
  wire [15:0]         maskExt_lo_969 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_969 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_969 = {maskExt_hi_969, maskExt_lo_969};
  wire [15:0]         maskExt_lo_970 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_970 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_970 = {maskExt_hi_970, maskExt_lo_970};
  wire [15:0]         maskExt_lo_971 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_971 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_971 = {maskExt_hi_971, maskExt_lo_971};
  wire [15:0]         maskExt_lo_972 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_972 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_972 = {maskExt_hi_972, maskExt_lo_972};
  wire [15:0]         maskExt_lo_973 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_973 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_973 = {maskExt_hi_973, maskExt_lo_973};
  wire [15:0]         maskExt_lo_974 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_974 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_974 = {maskExt_hi_974, maskExt_lo_974};
  wire [15:0]         maskExt_lo_975 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_975 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_975 = {maskExt_hi_975, maskExt_lo_975};
  wire [15:0]         maskExt_lo_976 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_976 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_976 = {maskExt_hi_976, maskExt_lo_976};
  wire [15:0]         maskExt_lo_977 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_977 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_977 = {maskExt_hi_977, maskExt_lo_977};
  wire [15:0]         maskExt_lo_978 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_978 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_978 = {maskExt_hi_978, maskExt_lo_978};
  wire [15:0]         maskExt_lo_979 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_979 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_979 = {maskExt_hi_979, maskExt_lo_979};
  wire [15:0]         maskExt_lo_980 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_980 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_980 = {maskExt_hi_980, maskExt_lo_980};
  wire [15:0]         maskExt_lo_981 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_981 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_981 = {maskExt_hi_981, maskExt_lo_981};
  wire [15:0]         maskExt_lo_982 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_982 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_982 = {maskExt_hi_982, maskExt_lo_982};
  wire [15:0]         maskExt_lo_983 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_983 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_983 = {maskExt_hi_983, maskExt_lo_983};
  wire [15:0]         maskExt_lo_984 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_984 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_984 = {maskExt_hi_984, maskExt_lo_984};
  wire [15:0]         maskExt_lo_985 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_985 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_985 = {maskExt_hi_985, maskExt_lo_985};
  wire [15:0]         maskExt_lo_986 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_986 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_986 = {maskExt_hi_986, maskExt_lo_986};
  wire [15:0]         maskExt_lo_987 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_987 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_987 = {maskExt_hi_987, maskExt_lo_987};
  wire [15:0]         maskExt_lo_988 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_988 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_988 = {maskExt_hi_988, maskExt_lo_988};
  wire [15:0]         maskExt_lo_989 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_989 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_989 = {maskExt_hi_989, maskExt_lo_989};
  wire [15:0]         maskExt_lo_990 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_990 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_990 = {maskExt_hi_990, maskExt_lo_990};
  wire [15:0]         maskExt_lo_991 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_991 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_991 = {maskExt_hi_991, maskExt_lo_991};
  wire [15:0]         maskExt_lo_992 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_992 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_992 = {maskExt_hi_992, maskExt_lo_992};
  wire [15:0]         maskExt_lo_993 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_993 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_993 = {maskExt_hi_993, maskExt_lo_993};
  wire [15:0]         maskExt_lo_994 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_994 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_994 = {maskExt_hi_994, maskExt_lo_994};
  wire [15:0]         maskExt_lo_995 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_995 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_995 = {maskExt_hi_995, maskExt_lo_995};
  wire [15:0]         maskExt_lo_996 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_996 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_996 = {maskExt_hi_996, maskExt_lo_996};
  wire [15:0]         maskExt_lo_997 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_997 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_997 = {maskExt_hi_997, maskExt_lo_997};
  wire [15:0]         maskExt_lo_998 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_998 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_998 = {maskExt_hi_998, maskExt_lo_998};
  wire [15:0]         maskExt_lo_999 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_999 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_999 = {maskExt_hi_999, maskExt_lo_999};
  wire [15:0]         maskExt_lo_1000 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1000 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1000 = {maskExt_hi_1000, maskExt_lo_1000};
  wire [15:0]         maskExt_lo_1001 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1001 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1001 = {maskExt_hi_1001, maskExt_lo_1001};
  wire [15:0]         maskExt_lo_1002 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1002 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1002 = {maskExt_hi_1002, maskExt_lo_1002};
  wire [15:0]         maskExt_lo_1003 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1003 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1003 = {maskExt_hi_1003, maskExt_lo_1003};
  wire [15:0]         maskExt_lo_1004 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1004 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1004 = {maskExt_hi_1004, maskExt_lo_1004};
  wire [15:0]         maskExt_lo_1005 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1005 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1005 = {maskExt_hi_1005, maskExt_lo_1005};
  wire [15:0]         maskExt_lo_1006 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1006 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1006 = {maskExt_hi_1006, maskExt_lo_1006};
  wire [15:0]         maskExt_lo_1007 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1007 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1007 = {maskExt_hi_1007, maskExt_lo_1007};
  wire [15:0]         maskExt_lo_1008 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1008 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1008 = {maskExt_hi_1008, maskExt_lo_1008};
  wire [15:0]         maskExt_lo_1009 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1009 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1009 = {maskExt_hi_1009, maskExt_lo_1009};
  wire [15:0]         maskExt_lo_1010 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1010 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1010 = {maskExt_hi_1010, maskExt_lo_1010};
  wire [15:0]         maskExt_lo_1011 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1011 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1011 = {maskExt_hi_1011, maskExt_lo_1011};
  wire [15:0]         maskExt_lo_1012 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1012 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1012 = {maskExt_hi_1012, maskExt_lo_1012};
  wire [15:0]         maskExt_lo_1013 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1013 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1013 = {maskExt_hi_1013, maskExt_lo_1013};
  wire [15:0]         maskExt_lo_1014 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1014 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1014 = {maskExt_hi_1014, maskExt_lo_1014};
  wire [15:0]         maskExt_lo_1015 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1015 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1015 = {maskExt_hi_1015, maskExt_lo_1015};
  wire [15:0]         maskExt_lo_1016 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1016 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1016 = {maskExt_hi_1016, maskExt_lo_1016};
  wire [15:0]         maskExt_lo_1017 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1017 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1017 = {maskExt_hi_1017, maskExt_lo_1017};
  wire [15:0]         maskExt_lo_1018 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1018 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1018 = {maskExt_hi_1018, maskExt_lo_1018};
  wire [15:0]         maskExt_lo_1019 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1019 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1019 = {maskExt_hi_1019, maskExt_lo_1019};
  wire [15:0]         maskExt_lo_1020 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1020 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]         maskExt_1020 = {maskExt_hi_1020, maskExt_lo_1020};
  wire [15:0]         maskExt_lo_1021 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1021 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]         maskExt_1021 = {maskExt_hi_1021, maskExt_lo_1021};
  wire [15:0]         maskExt_lo_1022 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1022 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]         maskExt_1022 = {maskExt_hi_1022, maskExt_lo_1022};
  wire [15:0]         maskExt_lo_1023 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]         maskExt_hi_1023 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]         maskExt_1023 = {maskExt_hi_1023, maskExt_lo_1023};
  wire                alwaysMerge = {request_bits_instructionInformation_mop_0, request_bits_instructionInformation_lumop_0[2:0], request_bits_instructionInformation_lumop_0[4]} == 6'h0;
  wire                useLoadUnit = alwaysMerge & ~request_bits_instructionInformation_isStore_0;
  wire                useStoreUnit = alwaysMerge & request_bits_instructionInformation_isStore_0;
  wire                useOtherUnit = ~alwaysMerge;
  wire                addressCheck = _otherUnit_status_idle & (~useOtherUnit | _loadUnit_status_idle & _storeUnit_status_idle);
  wire                unitReady = useLoadUnit & _loadUnit_status_idle | useStoreUnit & _storeUnit_status_idle | useOtherUnit & _otherUnit_status_idle;
  wire                request_ready_0 = unitReady & addressCheck;
  wire                requestFire = request_ready_0 & request_valid_0;
  wire                reqEnq_0 = useLoadUnit & requestFire;
  wire                reqEnq_1 = useStoreUnit & requestFire;
  wire                reqEnq_2 = useOtherUnit & requestFire;
  wire [10:0]         maskSelect = _loadUnit_maskSelect_valid ? _loadUnit_maskSelect_bits : 11'h0;
  wire [63:0]         _GEN = {v0_1, v0_0};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]         _GEN_0 = {v0_3, v0_2};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_0;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_1 = {v0_5, v0_4};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]         _GEN_2 = {v0_7, v0_6};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_2;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_3 = {v0_9, v0_8};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]         _GEN_4 = {v0_11, v0_10};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_4;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_5 = {v0_13, v0_12};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]         _GEN_6 = {v0_15, v0_14};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_6;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_7 = {v0_17, v0_16};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]         _GEN_8 = {v0_19, v0_18};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_8;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_9 = {v0_21, v0_20};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]         _GEN_10 = {v0_23, v0_22};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_10;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_11 = {v0_25, v0_24};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]         _GEN_12 = {v0_27, v0_26};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_12;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_13 = {v0_29, v0_28};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]         _GEN_14 = {v0_31, v0_30};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_14;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_15 = {v0_33, v0_32};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]         _GEN_16 = {v0_35, v0_34};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_16;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_17 = {v0_37, v0_36};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]         _GEN_18 = {v0_39, v0_38};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_18;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_19 = {v0_41, v0_40};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]         _GEN_20 = {v0_43, v0_42};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_20;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_21 = {v0_45, v0_44};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]         _GEN_22 = {v0_47, v0_46};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_22;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_23 = {v0_49, v0_48};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]         _GEN_24 = {v0_51, v0_50};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_24;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_25 = {v0_53, v0_52};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]         _GEN_26 = {v0_55, v0_54};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_26;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_27 = {v0_57, v0_56};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]         _GEN_28 = {v0_59, v0_58};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_28;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_29 = {v0_61, v0_60};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]         _GEN_30 = {v0_63, v0_62};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_30;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_31 = {v0_65, v0_64};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_31;
  wire [63:0]         _GEN_32 = {v0_67, v0_66};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_32;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_33 = {v0_69, v0_68};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_33;
  wire [63:0]         _GEN_34 = {v0_71, v0_70};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_34;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_35 = {v0_73, v0_72};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_35;
  wire [63:0]         _GEN_36 = {v0_75, v0_74};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_36;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_37 = {v0_77, v0_76};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_37;
  wire [63:0]         _GEN_38 = {v0_79, v0_78};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_38;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_39 = {v0_81, v0_80};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_39;
  wire [63:0]         _GEN_40 = {v0_83, v0_82};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_40;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_41 = {v0_85, v0_84};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_41;
  wire [63:0]         _GEN_42 = {v0_87, v0_86};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_42;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_43 = {v0_89, v0_88};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_43;
  wire [63:0]         _GEN_44 = {v0_91, v0_90};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_44;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_45 = {v0_93, v0_92};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_45;
  wire [63:0]         _GEN_46 = {v0_95, v0_94};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_46;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_47 = {v0_97, v0_96};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_47;
  wire [63:0]         _GEN_48 = {v0_99, v0_98};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_48;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_49 = {v0_101, v0_100};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_49;
  wire [63:0]         _GEN_50 = {v0_103, v0_102};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_50;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_51 = {v0_105, v0_104};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_51;
  wire [63:0]         _GEN_52 = {v0_107, v0_106};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_52;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_53 = {v0_109, v0_108};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_53;
  wire [63:0]         _GEN_54 = {v0_111, v0_110};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_54;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_55 = {v0_113, v0_112};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_55;
  wire [63:0]         _GEN_56 = {v0_115, v0_114};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_56;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_57 = {v0_117, v0_116};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_57;
  wire [63:0]         _GEN_58 = {v0_119, v0_118};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_58;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_59 = {v0_121, v0_120};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_59;
  wire [63:0]         _GEN_60 = {v0_123, v0_122};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_60;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_61 = {v0_125, v0_124};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_61;
  wire [63:0]         _GEN_62 = {v0_127, v0_126};
  wire [63:0]         loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]         storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [63:0]         otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_62;
  wire [127:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_lo_lo = {loadUnit_maskInput_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_lo_lo};
  wire [63:0]         _GEN_63 = {v0_129, v0_128};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_63;
  wire [63:0]         _GEN_64 = {v0_131, v0_130};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_64;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_65 = {v0_133, v0_132};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_65;
  wire [63:0]         _GEN_66 = {v0_135, v0_134};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_66;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_67 = {v0_137, v0_136};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_67;
  wire [63:0]         _GEN_68 = {v0_139, v0_138};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_68;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_69 = {v0_141, v0_140};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_69;
  wire [63:0]         _GEN_70 = {v0_143, v0_142};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_70;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_71 = {v0_145, v0_144};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_71;
  wire [63:0]         _GEN_72 = {v0_147, v0_146};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_72;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_73 = {v0_149, v0_148};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_73;
  wire [63:0]         _GEN_74 = {v0_151, v0_150};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_74;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_75 = {v0_153, v0_152};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_75;
  wire [63:0]         _GEN_76 = {v0_155, v0_154};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_76;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_77 = {v0_157, v0_156};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_77;
  wire [63:0]         _GEN_78 = {v0_159, v0_158};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_78;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_79 = {v0_161, v0_160};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_79;
  wire [63:0]         _GEN_80 = {v0_163, v0_162};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_80;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_81 = {v0_165, v0_164};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_81;
  wire [63:0]         _GEN_82 = {v0_167, v0_166};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_82;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_83 = {v0_169, v0_168};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_83;
  wire [63:0]         _GEN_84 = {v0_171, v0_170};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_84;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_85 = {v0_173, v0_172};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_85;
  wire [63:0]         _GEN_86 = {v0_175, v0_174};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_86;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_87 = {v0_177, v0_176};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_87;
  wire [63:0]         _GEN_88 = {v0_179, v0_178};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_88;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_89 = {v0_181, v0_180};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_89;
  wire [63:0]         _GEN_90 = {v0_183, v0_182};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_90;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_91 = {v0_185, v0_184};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_91;
  wire [63:0]         _GEN_92 = {v0_187, v0_186};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_92;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_93 = {v0_189, v0_188};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_93;
  wire [63:0]         _GEN_94 = {v0_191, v0_190};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_94;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_95 = {v0_193, v0_192};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_95;
  wire [63:0]         _GEN_96 = {v0_195, v0_194};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_96;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_97 = {v0_197, v0_196};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_97;
  wire [63:0]         _GEN_98 = {v0_199, v0_198};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_98;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_99 = {v0_201, v0_200};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_99;
  wire [63:0]         _GEN_100 = {v0_203, v0_202};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_100;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_101 = {v0_205, v0_204};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_101;
  wire [63:0]         _GEN_102 = {v0_207, v0_206};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_102;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_103 = {v0_209, v0_208};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_103;
  wire [63:0]         _GEN_104 = {v0_211, v0_210};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_104;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_105 = {v0_213, v0_212};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_105;
  wire [63:0]         _GEN_106 = {v0_215, v0_214};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_106;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_107 = {v0_217, v0_216};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_107;
  wire [63:0]         _GEN_108 = {v0_219, v0_218};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_108;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_109 = {v0_221, v0_220};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_109;
  wire [63:0]         _GEN_110 = {v0_223, v0_222};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_110;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_111 = {v0_225, v0_224};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_111;
  wire [63:0]         _GEN_112 = {v0_227, v0_226};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_112;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_113 = {v0_229, v0_228};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_113;
  wire [63:0]         _GEN_114 = {v0_231, v0_230};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_114;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_115 = {v0_233, v0_232};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_115;
  wire [63:0]         _GEN_116 = {v0_235, v0_234};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_116;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_117 = {v0_237, v0_236};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_117;
  wire [63:0]         _GEN_118 = {v0_239, v0_238};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_118;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_119 = {v0_241, v0_240};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_119;
  wire [63:0]         _GEN_120 = {v0_243, v0_242};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_120;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_121 = {v0_245, v0_244};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_121;
  wire [63:0]         _GEN_122 = {v0_247, v0_246};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_122;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_123 = {v0_249, v0_248};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_123;
  wire [63:0]         _GEN_124 = {v0_251, v0_250};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_124;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_125 = {v0_253, v0_252};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_125;
  wire [63:0]         _GEN_126 = {v0_255, v0_254};
  wire [63:0]         loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]         storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [63:0]         otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_126;
  wire [127:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_lo_hi_hi = {loadUnit_maskInput_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_lo_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_lo_hi = {loadUnit_maskInput_lo_lo_hi_hi, loadUnit_maskInput_lo_lo_hi_lo};
  wire [8191:0]       loadUnit_maskInput_lo_lo = {loadUnit_maskInput_lo_lo_hi, loadUnit_maskInput_lo_lo_lo};
  wire [63:0]         _GEN_127 = {v0_257, v0_256};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_127;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_127;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_127;
  wire [63:0]         _GEN_128 = {v0_259, v0_258};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_128;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_128;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_128;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_129 = {v0_261, v0_260};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_129;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_129;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_129;
  wire [63:0]         _GEN_130 = {v0_263, v0_262};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_130;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_130;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_130;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_131 = {v0_265, v0_264};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_131;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_131;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_131;
  wire [63:0]         _GEN_132 = {v0_267, v0_266};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_132;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_132;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_132;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_133 = {v0_269, v0_268};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_133;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_133;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_133;
  wire [63:0]         _GEN_134 = {v0_271, v0_270};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_134;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_134;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_134;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_135 = {v0_273, v0_272};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_135;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_135;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_135;
  wire [63:0]         _GEN_136 = {v0_275, v0_274};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_136;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_136;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_136;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_137 = {v0_277, v0_276};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_137;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_137;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_137;
  wire [63:0]         _GEN_138 = {v0_279, v0_278};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_138;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_138;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_138;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_139 = {v0_281, v0_280};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_139;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_139;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_139;
  wire [63:0]         _GEN_140 = {v0_283, v0_282};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_140;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_140;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_140;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_141 = {v0_285, v0_284};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_141;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_141;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_141;
  wire [63:0]         _GEN_142 = {v0_287, v0_286};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_142;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_142;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_142;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_143 = {v0_289, v0_288};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_143;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_143;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_143;
  wire [63:0]         _GEN_144 = {v0_291, v0_290};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_144;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_144;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_144;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_145 = {v0_293, v0_292};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_145;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_145;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_145;
  wire [63:0]         _GEN_146 = {v0_295, v0_294};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_146;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_146;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_146;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_147 = {v0_297, v0_296};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_147;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_147;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_147;
  wire [63:0]         _GEN_148 = {v0_299, v0_298};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_148;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_148;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_148;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_149 = {v0_301, v0_300};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_149;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_149;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_149;
  wire [63:0]         _GEN_150 = {v0_303, v0_302};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_150;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_150;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_150;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_151 = {v0_305, v0_304};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_151;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_151;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_151;
  wire [63:0]         _GEN_152 = {v0_307, v0_306};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_152;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_152;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_152;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_153 = {v0_309, v0_308};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_153;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_153;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_153;
  wire [63:0]         _GEN_154 = {v0_311, v0_310};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_154;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_154;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_154;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_155 = {v0_313, v0_312};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_155;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_155;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_155;
  wire [63:0]         _GEN_156 = {v0_315, v0_314};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_156;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_156;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_156;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_157 = {v0_317, v0_316};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_157;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_157;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_157;
  wire [63:0]         _GEN_158 = {v0_319, v0_318};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_158;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_158;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_158;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_159 = {v0_321, v0_320};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_159;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_159;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_159;
  wire [63:0]         _GEN_160 = {v0_323, v0_322};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_160;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_160;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_160;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_161 = {v0_325, v0_324};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_161;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_161;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_161;
  wire [63:0]         _GEN_162 = {v0_327, v0_326};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_162;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_162;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_162;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_163 = {v0_329, v0_328};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_163;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_163;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_163;
  wire [63:0]         _GEN_164 = {v0_331, v0_330};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_164;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_164;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_164;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_165 = {v0_333, v0_332};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_165;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_165;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_165;
  wire [63:0]         _GEN_166 = {v0_335, v0_334};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_166;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_166;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_166;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_167 = {v0_337, v0_336};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_167;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_167;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_167;
  wire [63:0]         _GEN_168 = {v0_339, v0_338};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_168;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_168;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_168;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_169 = {v0_341, v0_340};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_169;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_169;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_169;
  wire [63:0]         _GEN_170 = {v0_343, v0_342};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_170;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_170;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_170;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_171 = {v0_345, v0_344};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_171;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_171;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_171;
  wire [63:0]         _GEN_172 = {v0_347, v0_346};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_172;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_172;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_172;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_173 = {v0_349, v0_348};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_173;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_173;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_173;
  wire [63:0]         _GEN_174 = {v0_351, v0_350};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_174;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_174;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_174;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_175 = {v0_353, v0_352};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_175;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_175;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_175;
  wire [63:0]         _GEN_176 = {v0_355, v0_354};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_176;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_176;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_176;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_177 = {v0_357, v0_356};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_177;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_177;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_177;
  wire [63:0]         _GEN_178 = {v0_359, v0_358};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_178;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_178;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_178;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_179 = {v0_361, v0_360};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_179;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_179;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_179;
  wire [63:0]         _GEN_180 = {v0_363, v0_362};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_180;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_180;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_180;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_181 = {v0_365, v0_364};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_181;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_181;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_181;
  wire [63:0]         _GEN_182 = {v0_367, v0_366};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_182;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_182;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_182;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_183 = {v0_369, v0_368};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_183;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_183;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_183;
  wire [63:0]         _GEN_184 = {v0_371, v0_370};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_184;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_184;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_184;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_185 = {v0_373, v0_372};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_185;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_185;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_185;
  wire [63:0]         _GEN_186 = {v0_375, v0_374};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_186;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_186;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_186;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_187 = {v0_377, v0_376};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_187;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_187;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_187;
  wire [63:0]         _GEN_188 = {v0_379, v0_378};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_188;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_188;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_188;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_189 = {v0_381, v0_380};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_189;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_189;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_189;
  wire [63:0]         _GEN_190 = {v0_383, v0_382};
  wire [63:0]         loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_190;
  wire [63:0]         storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_190;
  wire [63:0]         otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_190;
  wire [127:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_hi_lo = {loadUnit_maskInput_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_lo_lo};
  wire [63:0]         _GEN_191 = {v0_385, v0_384};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_191;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_191;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_191;
  wire [63:0]         _GEN_192 = {v0_387, v0_386};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_192;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_192;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_192;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_193 = {v0_389, v0_388};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_193;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_193;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_193;
  wire [63:0]         _GEN_194 = {v0_391, v0_390};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_194;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_194;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_194;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_195 = {v0_393, v0_392};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_195;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_195;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_195;
  wire [63:0]         _GEN_196 = {v0_395, v0_394};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_196;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_196;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_196;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_197 = {v0_397, v0_396};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_197;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_197;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_197;
  wire [63:0]         _GEN_198 = {v0_399, v0_398};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_198;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_198;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_198;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_199 = {v0_401, v0_400};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_199;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_199;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_199;
  wire [63:0]         _GEN_200 = {v0_403, v0_402};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_200;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_200;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_200;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_201 = {v0_405, v0_404};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_201;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_201;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_201;
  wire [63:0]         _GEN_202 = {v0_407, v0_406};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_202;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_202;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_202;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_203 = {v0_409, v0_408};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_203;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_203;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_203;
  wire [63:0]         _GEN_204 = {v0_411, v0_410};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_204;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_204;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_204;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_205 = {v0_413, v0_412};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_205;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_205;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_205;
  wire [63:0]         _GEN_206 = {v0_415, v0_414};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_206;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_206;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_206;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_207 = {v0_417, v0_416};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_207;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_207;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_207;
  wire [63:0]         _GEN_208 = {v0_419, v0_418};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_208;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_208;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_208;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_209 = {v0_421, v0_420};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_209;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_209;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_209;
  wire [63:0]         _GEN_210 = {v0_423, v0_422};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_210;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_210;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_210;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_211 = {v0_425, v0_424};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_211;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_211;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_211;
  wire [63:0]         _GEN_212 = {v0_427, v0_426};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_212;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_212;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_212;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_213 = {v0_429, v0_428};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_213;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_213;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_213;
  wire [63:0]         _GEN_214 = {v0_431, v0_430};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_214;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_214;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_214;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_215 = {v0_433, v0_432};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_215;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_215;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_215;
  wire [63:0]         _GEN_216 = {v0_435, v0_434};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_216;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_216;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_216;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_217 = {v0_437, v0_436};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_217;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_217;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_217;
  wire [63:0]         _GEN_218 = {v0_439, v0_438};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_218;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_218;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_218;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_219 = {v0_441, v0_440};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_219;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_219;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_219;
  wire [63:0]         _GEN_220 = {v0_443, v0_442};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_220;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_220;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_220;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_221 = {v0_445, v0_444};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_221;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_221;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_221;
  wire [63:0]         _GEN_222 = {v0_447, v0_446};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_222;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_222;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_222;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_223 = {v0_449, v0_448};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_223;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_223;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_223;
  wire [63:0]         _GEN_224 = {v0_451, v0_450};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_224;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_224;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_224;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_225 = {v0_453, v0_452};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_225;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_225;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_225;
  wire [63:0]         _GEN_226 = {v0_455, v0_454};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_226;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_226;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_226;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_227 = {v0_457, v0_456};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_227;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_227;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_227;
  wire [63:0]         _GEN_228 = {v0_459, v0_458};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_228;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_228;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_228;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_229 = {v0_461, v0_460};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_229;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_229;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_229;
  wire [63:0]         _GEN_230 = {v0_463, v0_462};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_230;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_230;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_230;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_231 = {v0_465, v0_464};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_231;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_231;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_231;
  wire [63:0]         _GEN_232 = {v0_467, v0_466};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_232;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_232;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_232;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_233 = {v0_469, v0_468};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_233;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_233;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_233;
  wire [63:0]         _GEN_234 = {v0_471, v0_470};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_234;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_234;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_234;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_235 = {v0_473, v0_472};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_235;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_235;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_235;
  wire [63:0]         _GEN_236 = {v0_475, v0_474};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_236;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_236;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_236;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_237 = {v0_477, v0_476};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_237;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_237;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_237;
  wire [63:0]         _GEN_238 = {v0_479, v0_478};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_238;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_238;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_238;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_239 = {v0_481, v0_480};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_239;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_239;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_239;
  wire [63:0]         _GEN_240 = {v0_483, v0_482};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_240;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_240;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_240;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_241 = {v0_485, v0_484};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_241;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_241;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_241;
  wire [63:0]         _GEN_242 = {v0_487, v0_486};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_242;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_242;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_242;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_243 = {v0_489, v0_488};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_243;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_243;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_243;
  wire [63:0]         _GEN_244 = {v0_491, v0_490};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_244;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_244;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_244;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_245 = {v0_493, v0_492};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_245;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_245;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_245;
  wire [63:0]         _GEN_246 = {v0_495, v0_494};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_246;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_246;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_246;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_247 = {v0_497, v0_496};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_247;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_247;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_247;
  wire [63:0]         _GEN_248 = {v0_499, v0_498};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_248;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_248;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_248;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_249 = {v0_501, v0_500};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_249;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_249;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_249;
  wire [63:0]         _GEN_250 = {v0_503, v0_502};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_250;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_250;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_250;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_251 = {v0_505, v0_504};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_251;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_251;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_251;
  wire [63:0]         _GEN_252 = {v0_507, v0_506};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_252;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_252;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_252;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_253 = {v0_509, v0_508};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_253;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_253;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_253;
  wire [63:0]         _GEN_254 = {v0_511, v0_510};
  wire [63:0]         loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_254;
  wire [63:0]         storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_254;
  wire [63:0]         otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_254;
  wire [127:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_lo_hi_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_lo_hi_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_lo_hi_hi = {loadUnit_maskInput_lo_hi_hi_hi, loadUnit_maskInput_lo_hi_hi_lo};
  wire [8191:0]       loadUnit_maskInput_lo_hi = {loadUnit_maskInput_lo_hi_hi, loadUnit_maskInput_lo_hi_lo};
  wire [16383:0]      loadUnit_maskInput_lo = {loadUnit_maskInput_lo_hi, loadUnit_maskInput_lo_lo};
  wire [63:0]         _GEN_255 = {v0_513, v0_512};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_255;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_255;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo = _GEN_255;
  wire [63:0]         _GEN_256 = {v0_515, v0_514};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_256;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_256;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi = _GEN_256;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_257 = {v0_517, v0_516};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_257;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_257;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo = _GEN_257;
  wire [63:0]         _GEN_258 = {v0_519, v0_518};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_258;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_258;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi = _GEN_258;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_259 = {v0_521, v0_520};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_259;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_259;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo = _GEN_259;
  wire [63:0]         _GEN_260 = {v0_523, v0_522};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_260;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_260;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi = _GEN_260;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_261 = {v0_525, v0_524};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_261;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_261;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo = _GEN_261;
  wire [63:0]         _GEN_262 = {v0_527, v0_526};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_262;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_262;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi = _GEN_262;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_263 = {v0_529, v0_528};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_263;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_263;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo = _GEN_263;
  wire [63:0]         _GEN_264 = {v0_531, v0_530};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_264;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_264;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi = _GEN_264;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_265 = {v0_533, v0_532};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_265;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_265;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo = _GEN_265;
  wire [63:0]         _GEN_266 = {v0_535, v0_534};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_266;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_266;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi = _GEN_266;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_267 = {v0_537, v0_536};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_267;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_267;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo = _GEN_267;
  wire [63:0]         _GEN_268 = {v0_539, v0_538};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_268;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_268;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi = _GEN_268;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_269 = {v0_541, v0_540};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_269;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_269;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo = _GEN_269;
  wire [63:0]         _GEN_270 = {v0_543, v0_542};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_270;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_270;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi = _GEN_270;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_271 = {v0_545, v0_544};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_271;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_271;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo = _GEN_271;
  wire [63:0]         _GEN_272 = {v0_547, v0_546};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_272;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_272;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi = _GEN_272;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_273 = {v0_549, v0_548};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_273;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_273;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo = _GEN_273;
  wire [63:0]         _GEN_274 = {v0_551, v0_550};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_274;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_274;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi = _GEN_274;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_275 = {v0_553, v0_552};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_275;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_275;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo = _GEN_275;
  wire [63:0]         _GEN_276 = {v0_555, v0_554};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_276;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_276;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi = _GEN_276;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_277 = {v0_557, v0_556};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_277;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_277;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo = _GEN_277;
  wire [63:0]         _GEN_278 = {v0_559, v0_558};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_278;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_278;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi = _GEN_278;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_279 = {v0_561, v0_560};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_279;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_279;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo = _GEN_279;
  wire [63:0]         _GEN_280 = {v0_563, v0_562};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_280;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_280;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi = _GEN_280;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_281 = {v0_565, v0_564};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_281;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_281;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo = _GEN_281;
  wire [63:0]         _GEN_282 = {v0_567, v0_566};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_282;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_282;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi = _GEN_282;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_283 = {v0_569, v0_568};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_283;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_283;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo = _GEN_283;
  wire [63:0]         _GEN_284 = {v0_571, v0_570};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_284;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_284;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi = _GEN_284;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_285 = {v0_573, v0_572};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_285;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_285;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo = _GEN_285;
  wire [63:0]         _GEN_286 = {v0_575, v0_574};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_286;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_286;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi = _GEN_286;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_287 = {v0_577, v0_576};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_287;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_287;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo = _GEN_287;
  wire [63:0]         _GEN_288 = {v0_579, v0_578};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_288;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_288;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi = _GEN_288;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_289 = {v0_581, v0_580};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_289;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_289;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo = _GEN_289;
  wire [63:0]         _GEN_290 = {v0_583, v0_582};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_290;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_290;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi = _GEN_290;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_291 = {v0_585, v0_584};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_291;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_291;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo = _GEN_291;
  wire [63:0]         _GEN_292 = {v0_587, v0_586};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_292;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_292;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi = _GEN_292;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_293 = {v0_589, v0_588};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_293;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_293;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo = _GEN_293;
  wire [63:0]         _GEN_294 = {v0_591, v0_590};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_294;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_294;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi = _GEN_294;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_295 = {v0_593, v0_592};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_295;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_295;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo = _GEN_295;
  wire [63:0]         _GEN_296 = {v0_595, v0_594};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_296;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_296;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi = _GEN_296;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_297 = {v0_597, v0_596};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_297;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_297;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo = _GEN_297;
  wire [63:0]         _GEN_298 = {v0_599, v0_598};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_298;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_298;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi = _GEN_298;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_299 = {v0_601, v0_600};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_299;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_299;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo = _GEN_299;
  wire [63:0]         _GEN_300 = {v0_603, v0_602};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_300;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_300;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi = _GEN_300;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_301 = {v0_605, v0_604};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_301;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_301;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo = _GEN_301;
  wire [63:0]         _GEN_302 = {v0_607, v0_606};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_302;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_302;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi = _GEN_302;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_303 = {v0_609, v0_608};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_303;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_303;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo = _GEN_303;
  wire [63:0]         _GEN_304 = {v0_611, v0_610};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_304;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_304;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi = _GEN_304;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_305 = {v0_613, v0_612};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_305;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_305;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo = _GEN_305;
  wire [63:0]         _GEN_306 = {v0_615, v0_614};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_306;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_306;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi = _GEN_306;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_307 = {v0_617, v0_616};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_307;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_307;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo = _GEN_307;
  wire [63:0]         _GEN_308 = {v0_619, v0_618};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_308;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_308;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi = _GEN_308;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_309 = {v0_621, v0_620};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_309;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_309;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo = _GEN_309;
  wire [63:0]         _GEN_310 = {v0_623, v0_622};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_310;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_310;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi = _GEN_310;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_311 = {v0_625, v0_624};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_311;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_311;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo = _GEN_311;
  wire [63:0]         _GEN_312 = {v0_627, v0_626};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_312;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_312;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi = _GEN_312;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_313 = {v0_629, v0_628};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_313;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_313;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo = _GEN_313;
  wire [63:0]         _GEN_314 = {v0_631, v0_630};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_314;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_314;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi = _GEN_314;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_315 = {v0_633, v0_632};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_315;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_315;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo = _GEN_315;
  wire [63:0]         _GEN_316 = {v0_635, v0_634};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_316;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_316;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi = _GEN_316;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_317 = {v0_637, v0_636};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_317;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_317;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo = _GEN_317;
  wire [63:0]         _GEN_318 = {v0_639, v0_638};
  wire [63:0]         loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_318;
  wire [63:0]         storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_318;
  wire [63:0]         otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi = _GEN_318;
  wire [127:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_lo_lo = {loadUnit_maskInput_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_lo_lo};
  wire [63:0]         _GEN_319 = {v0_641, v0_640};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_319;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_319;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo = _GEN_319;
  wire [63:0]         _GEN_320 = {v0_643, v0_642};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_320;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_320;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi = _GEN_320;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_321 = {v0_645, v0_644};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_321;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_321;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo = _GEN_321;
  wire [63:0]         _GEN_322 = {v0_647, v0_646};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_322;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_322;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi = _GEN_322;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_323 = {v0_649, v0_648};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_323;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_323;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo = _GEN_323;
  wire [63:0]         _GEN_324 = {v0_651, v0_650};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_324;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_324;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi = _GEN_324;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_325 = {v0_653, v0_652};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_325;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_325;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo = _GEN_325;
  wire [63:0]         _GEN_326 = {v0_655, v0_654};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_326;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_326;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi = _GEN_326;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_327 = {v0_657, v0_656};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_327;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_327;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo = _GEN_327;
  wire [63:0]         _GEN_328 = {v0_659, v0_658};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_328;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_328;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi = _GEN_328;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_329 = {v0_661, v0_660};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_329;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_329;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo = _GEN_329;
  wire [63:0]         _GEN_330 = {v0_663, v0_662};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_330;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_330;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi = _GEN_330;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_331 = {v0_665, v0_664};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_331;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_331;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo = _GEN_331;
  wire [63:0]         _GEN_332 = {v0_667, v0_666};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_332;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_332;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi = _GEN_332;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_333 = {v0_669, v0_668};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_333;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_333;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo = _GEN_333;
  wire [63:0]         _GEN_334 = {v0_671, v0_670};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_334;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_334;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi = _GEN_334;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_335 = {v0_673, v0_672};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_335;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_335;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo = _GEN_335;
  wire [63:0]         _GEN_336 = {v0_675, v0_674};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_336;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_336;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi = _GEN_336;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_337 = {v0_677, v0_676};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_337;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_337;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo = _GEN_337;
  wire [63:0]         _GEN_338 = {v0_679, v0_678};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_338;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_338;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi = _GEN_338;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_339 = {v0_681, v0_680};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_339;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_339;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo = _GEN_339;
  wire [63:0]         _GEN_340 = {v0_683, v0_682};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_340;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_340;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi = _GEN_340;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_341 = {v0_685, v0_684};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_341;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_341;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo = _GEN_341;
  wire [63:0]         _GEN_342 = {v0_687, v0_686};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_342;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_342;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi = _GEN_342;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_343 = {v0_689, v0_688};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_343;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_343;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo = _GEN_343;
  wire [63:0]         _GEN_344 = {v0_691, v0_690};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_344;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_344;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi = _GEN_344;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_345 = {v0_693, v0_692};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_345;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_345;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo = _GEN_345;
  wire [63:0]         _GEN_346 = {v0_695, v0_694};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_346;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_346;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi = _GEN_346;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_347 = {v0_697, v0_696};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_347;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_347;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo = _GEN_347;
  wire [63:0]         _GEN_348 = {v0_699, v0_698};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_348;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_348;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi = _GEN_348;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_349 = {v0_701, v0_700};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_349;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_349;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo = _GEN_349;
  wire [63:0]         _GEN_350 = {v0_703, v0_702};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_350;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_350;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi = _GEN_350;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_351 = {v0_705, v0_704};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_351;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_351;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo = _GEN_351;
  wire [63:0]         _GEN_352 = {v0_707, v0_706};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_352;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_352;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi = _GEN_352;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_353 = {v0_709, v0_708};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_353;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_353;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo = _GEN_353;
  wire [63:0]         _GEN_354 = {v0_711, v0_710};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_354;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_354;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi = _GEN_354;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_355 = {v0_713, v0_712};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_355;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_355;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo = _GEN_355;
  wire [63:0]         _GEN_356 = {v0_715, v0_714};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_356;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_356;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi = _GEN_356;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_357 = {v0_717, v0_716};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_357;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_357;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo = _GEN_357;
  wire [63:0]         _GEN_358 = {v0_719, v0_718};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_358;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_358;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi = _GEN_358;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_359 = {v0_721, v0_720};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_359;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_359;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo = _GEN_359;
  wire [63:0]         _GEN_360 = {v0_723, v0_722};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_360;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_360;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi = _GEN_360;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_361 = {v0_725, v0_724};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_361;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_361;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo = _GEN_361;
  wire [63:0]         _GEN_362 = {v0_727, v0_726};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_362;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_362;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi = _GEN_362;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_363 = {v0_729, v0_728};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_363;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_363;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo = _GEN_363;
  wire [63:0]         _GEN_364 = {v0_731, v0_730};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_364;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_364;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi = _GEN_364;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_365 = {v0_733, v0_732};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_365;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_365;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo = _GEN_365;
  wire [63:0]         _GEN_366 = {v0_735, v0_734};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_366;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_366;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi = _GEN_366;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_367 = {v0_737, v0_736};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_367;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_367;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo = _GEN_367;
  wire [63:0]         _GEN_368 = {v0_739, v0_738};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_368;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_368;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi = _GEN_368;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_369 = {v0_741, v0_740};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_369;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_369;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo = _GEN_369;
  wire [63:0]         _GEN_370 = {v0_743, v0_742};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_370;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_370;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi = _GEN_370;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_371 = {v0_745, v0_744};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_371;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_371;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo = _GEN_371;
  wire [63:0]         _GEN_372 = {v0_747, v0_746};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_372;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_372;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi = _GEN_372;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_373 = {v0_749, v0_748};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_373;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_373;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo = _GEN_373;
  wire [63:0]         _GEN_374 = {v0_751, v0_750};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_374;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_374;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi = _GEN_374;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_375 = {v0_753, v0_752};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_375;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_375;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo = _GEN_375;
  wire [63:0]         _GEN_376 = {v0_755, v0_754};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_376;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_376;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi = _GEN_376;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_377 = {v0_757, v0_756};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_377;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_377;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo = _GEN_377;
  wire [63:0]         _GEN_378 = {v0_759, v0_758};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_378;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_378;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi = _GEN_378;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_379 = {v0_761, v0_760};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_379;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_379;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo = _GEN_379;
  wire [63:0]         _GEN_380 = {v0_763, v0_762};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_380;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_380;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi = _GEN_380;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_381 = {v0_765, v0_764};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_381;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_381;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo = _GEN_381;
  wire [63:0]         _GEN_382 = {v0_767, v0_766};
  wire [63:0]         loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_382;
  wire [63:0]         storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_382;
  wire [63:0]         otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi = _GEN_382;
  wire [127:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_lo_hi_hi = {loadUnit_maskInput_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_lo_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_lo_hi = {loadUnit_maskInput_hi_lo_hi_hi, loadUnit_maskInput_hi_lo_hi_lo};
  wire [8191:0]       loadUnit_maskInput_hi_lo = {loadUnit_maskInput_hi_lo_hi, loadUnit_maskInput_hi_lo_lo};
  wire [63:0]         _GEN_383 = {v0_769, v0_768};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_383;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_383;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo = _GEN_383;
  wire [63:0]         _GEN_384 = {v0_771, v0_770};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_384;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_384;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi = _GEN_384;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_385 = {v0_773, v0_772};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_385;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_385;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo = _GEN_385;
  wire [63:0]         _GEN_386 = {v0_775, v0_774};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_386;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_386;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi = _GEN_386;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_387 = {v0_777, v0_776};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_387;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_387;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo = _GEN_387;
  wire [63:0]         _GEN_388 = {v0_779, v0_778};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_388;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_388;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi = _GEN_388;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_389 = {v0_781, v0_780};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_389;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_389;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo = _GEN_389;
  wire [63:0]         _GEN_390 = {v0_783, v0_782};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_390;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_390;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi = _GEN_390;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_391 = {v0_785, v0_784};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_391;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_391;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo = _GEN_391;
  wire [63:0]         _GEN_392 = {v0_787, v0_786};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_392;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_392;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi = _GEN_392;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_393 = {v0_789, v0_788};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_393;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_393;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo = _GEN_393;
  wire [63:0]         _GEN_394 = {v0_791, v0_790};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_394;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_394;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi = _GEN_394;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_395 = {v0_793, v0_792};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_395;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_395;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo = _GEN_395;
  wire [63:0]         _GEN_396 = {v0_795, v0_794};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_396;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_396;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi = _GEN_396;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_397 = {v0_797, v0_796};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_397;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_397;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo = _GEN_397;
  wire [63:0]         _GEN_398 = {v0_799, v0_798};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_398;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_398;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi = _GEN_398;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_399 = {v0_801, v0_800};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_399;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_399;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo = _GEN_399;
  wire [63:0]         _GEN_400 = {v0_803, v0_802};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_400;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_400;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi = _GEN_400;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_401 = {v0_805, v0_804};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_401;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_401;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo = _GEN_401;
  wire [63:0]         _GEN_402 = {v0_807, v0_806};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_402;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_402;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi = _GEN_402;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_403 = {v0_809, v0_808};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_403;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_403;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo = _GEN_403;
  wire [63:0]         _GEN_404 = {v0_811, v0_810};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_404;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_404;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi = _GEN_404;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_405 = {v0_813, v0_812};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_405;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_405;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo = _GEN_405;
  wire [63:0]         _GEN_406 = {v0_815, v0_814};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_406;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_406;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi = _GEN_406;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_407 = {v0_817, v0_816};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_407;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_407;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo = _GEN_407;
  wire [63:0]         _GEN_408 = {v0_819, v0_818};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_408;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_408;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi = _GEN_408;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_409 = {v0_821, v0_820};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_409;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_409;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo = _GEN_409;
  wire [63:0]         _GEN_410 = {v0_823, v0_822};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_410;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_410;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi = _GEN_410;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_411 = {v0_825, v0_824};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_411;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_411;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo = _GEN_411;
  wire [63:0]         _GEN_412 = {v0_827, v0_826};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_412;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_412;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi = _GEN_412;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_413 = {v0_829, v0_828};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_413;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_413;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo = _GEN_413;
  wire [63:0]         _GEN_414 = {v0_831, v0_830};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_414;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_414;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi = _GEN_414;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_415 = {v0_833, v0_832};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_415;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_415;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo = _GEN_415;
  wire [63:0]         _GEN_416 = {v0_835, v0_834};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_416;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_416;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi = _GEN_416;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_417 = {v0_837, v0_836};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_417;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_417;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo = _GEN_417;
  wire [63:0]         _GEN_418 = {v0_839, v0_838};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_418;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_418;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi = _GEN_418;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_419 = {v0_841, v0_840};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_419;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_419;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo = _GEN_419;
  wire [63:0]         _GEN_420 = {v0_843, v0_842};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_420;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_420;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi = _GEN_420;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_421 = {v0_845, v0_844};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_421;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_421;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo = _GEN_421;
  wire [63:0]         _GEN_422 = {v0_847, v0_846};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_422;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_422;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi = _GEN_422;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_423 = {v0_849, v0_848};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_423;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_423;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo = _GEN_423;
  wire [63:0]         _GEN_424 = {v0_851, v0_850};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_424;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_424;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi = _GEN_424;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_425 = {v0_853, v0_852};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_425;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_425;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo = _GEN_425;
  wire [63:0]         _GEN_426 = {v0_855, v0_854};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_426;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_426;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi = _GEN_426;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_427 = {v0_857, v0_856};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_427;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_427;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo = _GEN_427;
  wire [63:0]         _GEN_428 = {v0_859, v0_858};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_428;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_428;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi = _GEN_428;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_429 = {v0_861, v0_860};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_429;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_429;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo = _GEN_429;
  wire [63:0]         _GEN_430 = {v0_863, v0_862};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_430;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_430;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi = _GEN_430;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_431 = {v0_865, v0_864};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_431;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_431;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo = _GEN_431;
  wire [63:0]         _GEN_432 = {v0_867, v0_866};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_432;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_432;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi = _GEN_432;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_433 = {v0_869, v0_868};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_433;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_433;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo = _GEN_433;
  wire [63:0]         _GEN_434 = {v0_871, v0_870};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_434;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_434;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi = _GEN_434;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_435 = {v0_873, v0_872};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_435;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_435;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo = _GEN_435;
  wire [63:0]         _GEN_436 = {v0_875, v0_874};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_436;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_436;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi = _GEN_436;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_437 = {v0_877, v0_876};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_437;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_437;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo = _GEN_437;
  wire [63:0]         _GEN_438 = {v0_879, v0_878};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_438;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_438;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi = _GEN_438;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_439 = {v0_881, v0_880};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_439;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_439;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo = _GEN_439;
  wire [63:0]         _GEN_440 = {v0_883, v0_882};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_440;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_440;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi = _GEN_440;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_441 = {v0_885, v0_884};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_441;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_441;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo = _GEN_441;
  wire [63:0]         _GEN_442 = {v0_887, v0_886};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_442;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_442;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi = _GEN_442;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_443 = {v0_889, v0_888};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_443;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_443;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo = _GEN_443;
  wire [63:0]         _GEN_444 = {v0_891, v0_890};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_444;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_444;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi = _GEN_444;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_445 = {v0_893, v0_892};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_445;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_445;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo = _GEN_445;
  wire [63:0]         _GEN_446 = {v0_895, v0_894};
  wire [63:0]         loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_446;
  wire [63:0]         storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_446;
  wire [63:0]         otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi = _GEN_446;
  wire [127:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_lo_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_hi_lo = {loadUnit_maskInput_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_lo_lo};
  wire [63:0]         _GEN_447 = {v0_897, v0_896};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_447;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_447;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo = _GEN_447;
  wire [63:0]         _GEN_448 = {v0_899, v0_898};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_448;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_448;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi = _GEN_448;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_449 = {v0_901, v0_900};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_449;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_449;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo = _GEN_449;
  wire [63:0]         _GEN_450 = {v0_903, v0_902};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_450;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_450;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi = _GEN_450;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_451 = {v0_905, v0_904};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_451;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_451;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo = _GEN_451;
  wire [63:0]         _GEN_452 = {v0_907, v0_906};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_452;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_452;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi = _GEN_452;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_453 = {v0_909, v0_908};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_453;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_453;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo = _GEN_453;
  wire [63:0]         _GEN_454 = {v0_911, v0_910};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_454;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_454;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi = _GEN_454;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_455 = {v0_913, v0_912};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_455;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_455;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo = _GEN_455;
  wire [63:0]         _GEN_456 = {v0_915, v0_914};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_456;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_456;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi = _GEN_456;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_457 = {v0_917, v0_916};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_457;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_457;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo = _GEN_457;
  wire [63:0]         _GEN_458 = {v0_919, v0_918};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_458;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_458;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi = _GEN_458;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_459 = {v0_921, v0_920};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_459;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_459;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo = _GEN_459;
  wire [63:0]         _GEN_460 = {v0_923, v0_922};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_460;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_460;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi = _GEN_460;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_461 = {v0_925, v0_924};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_461;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_461;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo = _GEN_461;
  wire [63:0]         _GEN_462 = {v0_927, v0_926};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_462;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_462;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi = _GEN_462;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_463 = {v0_929, v0_928};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_463;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_463;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo = _GEN_463;
  wire [63:0]         _GEN_464 = {v0_931, v0_930};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_464;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_464;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi = _GEN_464;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_465 = {v0_933, v0_932};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_465;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_465;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo = _GEN_465;
  wire [63:0]         _GEN_466 = {v0_935, v0_934};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_466;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_466;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi = _GEN_466;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_467 = {v0_937, v0_936};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_467;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_467;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo = _GEN_467;
  wire [63:0]         _GEN_468 = {v0_939, v0_938};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_468;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_468;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi = _GEN_468;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_469 = {v0_941, v0_940};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_469;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_469;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo = _GEN_469;
  wire [63:0]         _GEN_470 = {v0_943, v0_942};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_470;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_470;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi = _GEN_470;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_471 = {v0_945, v0_944};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_471;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_471;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo = _GEN_471;
  wire [63:0]         _GEN_472 = {v0_947, v0_946};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_472;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_472;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi = _GEN_472;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_473 = {v0_949, v0_948};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_473;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_473;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo = _GEN_473;
  wire [63:0]         _GEN_474 = {v0_951, v0_950};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_474;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_474;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi = _GEN_474;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_475 = {v0_953, v0_952};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_475;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_475;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo = _GEN_475;
  wire [63:0]         _GEN_476 = {v0_955, v0_954};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_476;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_476;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi = _GEN_476;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_477 = {v0_957, v0_956};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_477;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_477;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo = _GEN_477;
  wire [63:0]         _GEN_478 = {v0_959, v0_958};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_478;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_478;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi = _GEN_478;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_479 = {v0_961, v0_960};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_479;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_479;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo = _GEN_479;
  wire [63:0]         _GEN_480 = {v0_963, v0_962};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_480;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_480;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi = _GEN_480;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [63:0]         _GEN_481 = {v0_965, v0_964};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_481;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_481;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo = _GEN_481;
  wire [63:0]         _GEN_482 = {v0_967, v0_966};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_482;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_482;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi = _GEN_482;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_483 = {v0_969, v0_968};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_483;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_483;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo = _GEN_483;
  wire [63:0]         _GEN_484 = {v0_971, v0_970};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_484;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_484;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi = _GEN_484;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [63:0]         _GEN_485 = {v0_973, v0_972};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_485;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_485;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo = _GEN_485;
  wire [63:0]         _GEN_486 = {v0_975, v0_974};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_486;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_486;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi = _GEN_486;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_487 = {v0_977, v0_976};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_487;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_487;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo = _GEN_487;
  wire [63:0]         _GEN_488 = {v0_979, v0_978};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_488;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_488;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi = _GEN_488;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [63:0]         _GEN_489 = {v0_981, v0_980};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_489;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_489;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo = _GEN_489;
  wire [63:0]         _GEN_490 = {v0_983, v0_982};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_490;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_490;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi = _GEN_490;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_491 = {v0_985, v0_984};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_491;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_491;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo = _GEN_491;
  wire [63:0]         _GEN_492 = {v0_987, v0_986};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_492;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_492;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi = _GEN_492;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [63:0]         _GEN_493 = {v0_989, v0_988};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_493;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_493;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo = _GEN_493;
  wire [63:0]         _GEN_494 = {v0_991, v0_990};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_494;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_494;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi = _GEN_494;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_495 = {v0_993, v0_992};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_495;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_495;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo = _GEN_495;
  wire [63:0]         _GEN_496 = {v0_995, v0_994};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_496;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_496;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi = _GEN_496;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [63:0]         _GEN_497 = {v0_997, v0_996};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_497;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_497;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo = _GEN_497;
  wire [63:0]         _GEN_498 = {v0_999, v0_998};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_498;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_498;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi = _GEN_498;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_499 = {v0_1001, v0_1000};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_499;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_499;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo = _GEN_499;
  wire [63:0]         _GEN_500 = {v0_1003, v0_1002};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_500;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_500;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi = _GEN_500;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [63:0]         _GEN_501 = {v0_1005, v0_1004};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_501;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_501;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo = _GEN_501;
  wire [63:0]         _GEN_502 = {v0_1007, v0_1006};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_502;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_502;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi = _GEN_502;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_503 = {v0_1009, v0_1008};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_503;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_503;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo = _GEN_503;
  wire [63:0]         _GEN_504 = {v0_1011, v0_1010};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_504;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_504;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi = _GEN_504;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [63:0]         _GEN_505 = {v0_1013, v0_1012};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_505;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_505;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo = _GEN_505;
  wire [63:0]         _GEN_506 = {v0_1015, v0_1014};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_506;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_506;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi = _GEN_506;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_507 = {v0_1017, v0_1016};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_507;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_507;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo = _GEN_507;
  wire [63:0]         _GEN_508 = {v0_1019, v0_1018};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_508;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_508;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi = _GEN_508;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [63:0]         _GEN_509 = {v0_1021, v0_1020};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_509;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_509;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo = _GEN_509;
  wire [63:0]         _GEN_510 = {v0_1023, v0_1022};
  wire [63:0]         loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_510;
  wire [63:0]         storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_510;
  wire [63:0]         otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi;
  assign otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi = _GEN_510;
  wire [127:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        loadUnit_maskInput_hi_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       loadUnit_maskInput_hi_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       loadUnit_maskInput_hi_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_hi_lo};
  wire [4095:0]       loadUnit_maskInput_hi_hi_hi = {loadUnit_maskInput_hi_hi_hi_hi, loadUnit_maskInput_hi_hi_hi_lo};
  wire [8191:0]       loadUnit_maskInput_hi_hi = {loadUnit_maskInput_hi_hi_hi, loadUnit_maskInput_hi_hi_lo};
  wire [16383:0]      loadUnit_maskInput_hi = {loadUnit_maskInput_hi_hi, loadUnit_maskInput_hi_lo};
  wire [2047:0][15:0] _GEN_511 =
    {{loadUnit_maskInput_hi[16383:16368]},
     {loadUnit_maskInput_hi[16367:16352]},
     {loadUnit_maskInput_hi[16351:16336]},
     {loadUnit_maskInput_hi[16335:16320]},
     {loadUnit_maskInput_hi[16319:16304]},
     {loadUnit_maskInput_hi[16303:16288]},
     {loadUnit_maskInput_hi[16287:16272]},
     {loadUnit_maskInput_hi[16271:16256]},
     {loadUnit_maskInput_hi[16255:16240]},
     {loadUnit_maskInput_hi[16239:16224]},
     {loadUnit_maskInput_hi[16223:16208]},
     {loadUnit_maskInput_hi[16207:16192]},
     {loadUnit_maskInput_hi[16191:16176]},
     {loadUnit_maskInput_hi[16175:16160]},
     {loadUnit_maskInput_hi[16159:16144]},
     {loadUnit_maskInput_hi[16143:16128]},
     {loadUnit_maskInput_hi[16127:16112]},
     {loadUnit_maskInput_hi[16111:16096]},
     {loadUnit_maskInput_hi[16095:16080]},
     {loadUnit_maskInput_hi[16079:16064]},
     {loadUnit_maskInput_hi[16063:16048]},
     {loadUnit_maskInput_hi[16047:16032]},
     {loadUnit_maskInput_hi[16031:16016]},
     {loadUnit_maskInput_hi[16015:16000]},
     {loadUnit_maskInput_hi[15999:15984]},
     {loadUnit_maskInput_hi[15983:15968]},
     {loadUnit_maskInput_hi[15967:15952]},
     {loadUnit_maskInput_hi[15951:15936]},
     {loadUnit_maskInput_hi[15935:15920]},
     {loadUnit_maskInput_hi[15919:15904]},
     {loadUnit_maskInput_hi[15903:15888]},
     {loadUnit_maskInput_hi[15887:15872]},
     {loadUnit_maskInput_hi[15871:15856]},
     {loadUnit_maskInput_hi[15855:15840]},
     {loadUnit_maskInput_hi[15839:15824]},
     {loadUnit_maskInput_hi[15823:15808]},
     {loadUnit_maskInput_hi[15807:15792]},
     {loadUnit_maskInput_hi[15791:15776]},
     {loadUnit_maskInput_hi[15775:15760]},
     {loadUnit_maskInput_hi[15759:15744]},
     {loadUnit_maskInput_hi[15743:15728]},
     {loadUnit_maskInput_hi[15727:15712]},
     {loadUnit_maskInput_hi[15711:15696]},
     {loadUnit_maskInput_hi[15695:15680]},
     {loadUnit_maskInput_hi[15679:15664]},
     {loadUnit_maskInput_hi[15663:15648]},
     {loadUnit_maskInput_hi[15647:15632]},
     {loadUnit_maskInput_hi[15631:15616]},
     {loadUnit_maskInput_hi[15615:15600]},
     {loadUnit_maskInput_hi[15599:15584]},
     {loadUnit_maskInput_hi[15583:15568]},
     {loadUnit_maskInput_hi[15567:15552]},
     {loadUnit_maskInput_hi[15551:15536]},
     {loadUnit_maskInput_hi[15535:15520]},
     {loadUnit_maskInput_hi[15519:15504]},
     {loadUnit_maskInput_hi[15503:15488]},
     {loadUnit_maskInput_hi[15487:15472]},
     {loadUnit_maskInput_hi[15471:15456]},
     {loadUnit_maskInput_hi[15455:15440]},
     {loadUnit_maskInput_hi[15439:15424]},
     {loadUnit_maskInput_hi[15423:15408]},
     {loadUnit_maskInput_hi[15407:15392]},
     {loadUnit_maskInput_hi[15391:15376]},
     {loadUnit_maskInput_hi[15375:15360]},
     {loadUnit_maskInput_hi[15359:15344]},
     {loadUnit_maskInput_hi[15343:15328]},
     {loadUnit_maskInput_hi[15327:15312]},
     {loadUnit_maskInput_hi[15311:15296]},
     {loadUnit_maskInput_hi[15295:15280]},
     {loadUnit_maskInput_hi[15279:15264]},
     {loadUnit_maskInput_hi[15263:15248]},
     {loadUnit_maskInput_hi[15247:15232]},
     {loadUnit_maskInput_hi[15231:15216]},
     {loadUnit_maskInput_hi[15215:15200]},
     {loadUnit_maskInput_hi[15199:15184]},
     {loadUnit_maskInput_hi[15183:15168]},
     {loadUnit_maskInput_hi[15167:15152]},
     {loadUnit_maskInput_hi[15151:15136]},
     {loadUnit_maskInput_hi[15135:15120]},
     {loadUnit_maskInput_hi[15119:15104]},
     {loadUnit_maskInput_hi[15103:15088]},
     {loadUnit_maskInput_hi[15087:15072]},
     {loadUnit_maskInput_hi[15071:15056]},
     {loadUnit_maskInput_hi[15055:15040]},
     {loadUnit_maskInput_hi[15039:15024]},
     {loadUnit_maskInput_hi[15023:15008]},
     {loadUnit_maskInput_hi[15007:14992]},
     {loadUnit_maskInput_hi[14991:14976]},
     {loadUnit_maskInput_hi[14975:14960]},
     {loadUnit_maskInput_hi[14959:14944]},
     {loadUnit_maskInput_hi[14943:14928]},
     {loadUnit_maskInput_hi[14927:14912]},
     {loadUnit_maskInput_hi[14911:14896]},
     {loadUnit_maskInput_hi[14895:14880]},
     {loadUnit_maskInput_hi[14879:14864]},
     {loadUnit_maskInput_hi[14863:14848]},
     {loadUnit_maskInput_hi[14847:14832]},
     {loadUnit_maskInput_hi[14831:14816]},
     {loadUnit_maskInput_hi[14815:14800]},
     {loadUnit_maskInput_hi[14799:14784]},
     {loadUnit_maskInput_hi[14783:14768]},
     {loadUnit_maskInput_hi[14767:14752]},
     {loadUnit_maskInput_hi[14751:14736]},
     {loadUnit_maskInput_hi[14735:14720]},
     {loadUnit_maskInput_hi[14719:14704]},
     {loadUnit_maskInput_hi[14703:14688]},
     {loadUnit_maskInput_hi[14687:14672]},
     {loadUnit_maskInput_hi[14671:14656]},
     {loadUnit_maskInput_hi[14655:14640]},
     {loadUnit_maskInput_hi[14639:14624]},
     {loadUnit_maskInput_hi[14623:14608]},
     {loadUnit_maskInput_hi[14607:14592]},
     {loadUnit_maskInput_hi[14591:14576]},
     {loadUnit_maskInput_hi[14575:14560]},
     {loadUnit_maskInput_hi[14559:14544]},
     {loadUnit_maskInput_hi[14543:14528]},
     {loadUnit_maskInput_hi[14527:14512]},
     {loadUnit_maskInput_hi[14511:14496]},
     {loadUnit_maskInput_hi[14495:14480]},
     {loadUnit_maskInput_hi[14479:14464]},
     {loadUnit_maskInput_hi[14463:14448]},
     {loadUnit_maskInput_hi[14447:14432]},
     {loadUnit_maskInput_hi[14431:14416]},
     {loadUnit_maskInput_hi[14415:14400]},
     {loadUnit_maskInput_hi[14399:14384]},
     {loadUnit_maskInput_hi[14383:14368]},
     {loadUnit_maskInput_hi[14367:14352]},
     {loadUnit_maskInput_hi[14351:14336]},
     {loadUnit_maskInput_hi[14335:14320]},
     {loadUnit_maskInput_hi[14319:14304]},
     {loadUnit_maskInput_hi[14303:14288]},
     {loadUnit_maskInput_hi[14287:14272]},
     {loadUnit_maskInput_hi[14271:14256]},
     {loadUnit_maskInput_hi[14255:14240]},
     {loadUnit_maskInput_hi[14239:14224]},
     {loadUnit_maskInput_hi[14223:14208]},
     {loadUnit_maskInput_hi[14207:14192]},
     {loadUnit_maskInput_hi[14191:14176]},
     {loadUnit_maskInput_hi[14175:14160]},
     {loadUnit_maskInput_hi[14159:14144]},
     {loadUnit_maskInput_hi[14143:14128]},
     {loadUnit_maskInput_hi[14127:14112]},
     {loadUnit_maskInput_hi[14111:14096]},
     {loadUnit_maskInput_hi[14095:14080]},
     {loadUnit_maskInput_hi[14079:14064]},
     {loadUnit_maskInput_hi[14063:14048]},
     {loadUnit_maskInput_hi[14047:14032]},
     {loadUnit_maskInput_hi[14031:14016]},
     {loadUnit_maskInput_hi[14015:14000]},
     {loadUnit_maskInput_hi[13999:13984]},
     {loadUnit_maskInput_hi[13983:13968]},
     {loadUnit_maskInput_hi[13967:13952]},
     {loadUnit_maskInput_hi[13951:13936]},
     {loadUnit_maskInput_hi[13935:13920]},
     {loadUnit_maskInput_hi[13919:13904]},
     {loadUnit_maskInput_hi[13903:13888]},
     {loadUnit_maskInput_hi[13887:13872]},
     {loadUnit_maskInput_hi[13871:13856]},
     {loadUnit_maskInput_hi[13855:13840]},
     {loadUnit_maskInput_hi[13839:13824]},
     {loadUnit_maskInput_hi[13823:13808]},
     {loadUnit_maskInput_hi[13807:13792]},
     {loadUnit_maskInput_hi[13791:13776]},
     {loadUnit_maskInput_hi[13775:13760]},
     {loadUnit_maskInput_hi[13759:13744]},
     {loadUnit_maskInput_hi[13743:13728]},
     {loadUnit_maskInput_hi[13727:13712]},
     {loadUnit_maskInput_hi[13711:13696]},
     {loadUnit_maskInput_hi[13695:13680]},
     {loadUnit_maskInput_hi[13679:13664]},
     {loadUnit_maskInput_hi[13663:13648]},
     {loadUnit_maskInput_hi[13647:13632]},
     {loadUnit_maskInput_hi[13631:13616]},
     {loadUnit_maskInput_hi[13615:13600]},
     {loadUnit_maskInput_hi[13599:13584]},
     {loadUnit_maskInput_hi[13583:13568]},
     {loadUnit_maskInput_hi[13567:13552]},
     {loadUnit_maskInput_hi[13551:13536]},
     {loadUnit_maskInput_hi[13535:13520]},
     {loadUnit_maskInput_hi[13519:13504]},
     {loadUnit_maskInput_hi[13503:13488]},
     {loadUnit_maskInput_hi[13487:13472]},
     {loadUnit_maskInput_hi[13471:13456]},
     {loadUnit_maskInput_hi[13455:13440]},
     {loadUnit_maskInput_hi[13439:13424]},
     {loadUnit_maskInput_hi[13423:13408]},
     {loadUnit_maskInput_hi[13407:13392]},
     {loadUnit_maskInput_hi[13391:13376]},
     {loadUnit_maskInput_hi[13375:13360]},
     {loadUnit_maskInput_hi[13359:13344]},
     {loadUnit_maskInput_hi[13343:13328]},
     {loadUnit_maskInput_hi[13327:13312]},
     {loadUnit_maskInput_hi[13311:13296]},
     {loadUnit_maskInput_hi[13295:13280]},
     {loadUnit_maskInput_hi[13279:13264]},
     {loadUnit_maskInput_hi[13263:13248]},
     {loadUnit_maskInput_hi[13247:13232]},
     {loadUnit_maskInput_hi[13231:13216]},
     {loadUnit_maskInput_hi[13215:13200]},
     {loadUnit_maskInput_hi[13199:13184]},
     {loadUnit_maskInput_hi[13183:13168]},
     {loadUnit_maskInput_hi[13167:13152]},
     {loadUnit_maskInput_hi[13151:13136]},
     {loadUnit_maskInput_hi[13135:13120]},
     {loadUnit_maskInput_hi[13119:13104]},
     {loadUnit_maskInput_hi[13103:13088]},
     {loadUnit_maskInput_hi[13087:13072]},
     {loadUnit_maskInput_hi[13071:13056]},
     {loadUnit_maskInput_hi[13055:13040]},
     {loadUnit_maskInput_hi[13039:13024]},
     {loadUnit_maskInput_hi[13023:13008]},
     {loadUnit_maskInput_hi[13007:12992]},
     {loadUnit_maskInput_hi[12991:12976]},
     {loadUnit_maskInput_hi[12975:12960]},
     {loadUnit_maskInput_hi[12959:12944]},
     {loadUnit_maskInput_hi[12943:12928]},
     {loadUnit_maskInput_hi[12927:12912]},
     {loadUnit_maskInput_hi[12911:12896]},
     {loadUnit_maskInput_hi[12895:12880]},
     {loadUnit_maskInput_hi[12879:12864]},
     {loadUnit_maskInput_hi[12863:12848]},
     {loadUnit_maskInput_hi[12847:12832]},
     {loadUnit_maskInput_hi[12831:12816]},
     {loadUnit_maskInput_hi[12815:12800]},
     {loadUnit_maskInput_hi[12799:12784]},
     {loadUnit_maskInput_hi[12783:12768]},
     {loadUnit_maskInput_hi[12767:12752]},
     {loadUnit_maskInput_hi[12751:12736]},
     {loadUnit_maskInput_hi[12735:12720]},
     {loadUnit_maskInput_hi[12719:12704]},
     {loadUnit_maskInput_hi[12703:12688]},
     {loadUnit_maskInput_hi[12687:12672]},
     {loadUnit_maskInput_hi[12671:12656]},
     {loadUnit_maskInput_hi[12655:12640]},
     {loadUnit_maskInput_hi[12639:12624]},
     {loadUnit_maskInput_hi[12623:12608]},
     {loadUnit_maskInput_hi[12607:12592]},
     {loadUnit_maskInput_hi[12591:12576]},
     {loadUnit_maskInput_hi[12575:12560]},
     {loadUnit_maskInput_hi[12559:12544]},
     {loadUnit_maskInput_hi[12543:12528]},
     {loadUnit_maskInput_hi[12527:12512]},
     {loadUnit_maskInput_hi[12511:12496]},
     {loadUnit_maskInput_hi[12495:12480]},
     {loadUnit_maskInput_hi[12479:12464]},
     {loadUnit_maskInput_hi[12463:12448]},
     {loadUnit_maskInput_hi[12447:12432]},
     {loadUnit_maskInput_hi[12431:12416]},
     {loadUnit_maskInput_hi[12415:12400]},
     {loadUnit_maskInput_hi[12399:12384]},
     {loadUnit_maskInput_hi[12383:12368]},
     {loadUnit_maskInput_hi[12367:12352]},
     {loadUnit_maskInput_hi[12351:12336]},
     {loadUnit_maskInput_hi[12335:12320]},
     {loadUnit_maskInput_hi[12319:12304]},
     {loadUnit_maskInput_hi[12303:12288]},
     {loadUnit_maskInput_hi[12287:12272]},
     {loadUnit_maskInput_hi[12271:12256]},
     {loadUnit_maskInput_hi[12255:12240]},
     {loadUnit_maskInput_hi[12239:12224]},
     {loadUnit_maskInput_hi[12223:12208]},
     {loadUnit_maskInput_hi[12207:12192]},
     {loadUnit_maskInput_hi[12191:12176]},
     {loadUnit_maskInput_hi[12175:12160]},
     {loadUnit_maskInput_hi[12159:12144]},
     {loadUnit_maskInput_hi[12143:12128]},
     {loadUnit_maskInput_hi[12127:12112]},
     {loadUnit_maskInput_hi[12111:12096]},
     {loadUnit_maskInput_hi[12095:12080]},
     {loadUnit_maskInput_hi[12079:12064]},
     {loadUnit_maskInput_hi[12063:12048]},
     {loadUnit_maskInput_hi[12047:12032]},
     {loadUnit_maskInput_hi[12031:12016]},
     {loadUnit_maskInput_hi[12015:12000]},
     {loadUnit_maskInput_hi[11999:11984]},
     {loadUnit_maskInput_hi[11983:11968]},
     {loadUnit_maskInput_hi[11967:11952]},
     {loadUnit_maskInput_hi[11951:11936]},
     {loadUnit_maskInput_hi[11935:11920]},
     {loadUnit_maskInput_hi[11919:11904]},
     {loadUnit_maskInput_hi[11903:11888]},
     {loadUnit_maskInput_hi[11887:11872]},
     {loadUnit_maskInput_hi[11871:11856]},
     {loadUnit_maskInput_hi[11855:11840]},
     {loadUnit_maskInput_hi[11839:11824]},
     {loadUnit_maskInput_hi[11823:11808]},
     {loadUnit_maskInput_hi[11807:11792]},
     {loadUnit_maskInput_hi[11791:11776]},
     {loadUnit_maskInput_hi[11775:11760]},
     {loadUnit_maskInput_hi[11759:11744]},
     {loadUnit_maskInput_hi[11743:11728]},
     {loadUnit_maskInput_hi[11727:11712]},
     {loadUnit_maskInput_hi[11711:11696]},
     {loadUnit_maskInput_hi[11695:11680]},
     {loadUnit_maskInput_hi[11679:11664]},
     {loadUnit_maskInput_hi[11663:11648]},
     {loadUnit_maskInput_hi[11647:11632]},
     {loadUnit_maskInput_hi[11631:11616]},
     {loadUnit_maskInput_hi[11615:11600]},
     {loadUnit_maskInput_hi[11599:11584]},
     {loadUnit_maskInput_hi[11583:11568]},
     {loadUnit_maskInput_hi[11567:11552]},
     {loadUnit_maskInput_hi[11551:11536]},
     {loadUnit_maskInput_hi[11535:11520]},
     {loadUnit_maskInput_hi[11519:11504]},
     {loadUnit_maskInput_hi[11503:11488]},
     {loadUnit_maskInput_hi[11487:11472]},
     {loadUnit_maskInput_hi[11471:11456]},
     {loadUnit_maskInput_hi[11455:11440]},
     {loadUnit_maskInput_hi[11439:11424]},
     {loadUnit_maskInput_hi[11423:11408]},
     {loadUnit_maskInput_hi[11407:11392]},
     {loadUnit_maskInput_hi[11391:11376]},
     {loadUnit_maskInput_hi[11375:11360]},
     {loadUnit_maskInput_hi[11359:11344]},
     {loadUnit_maskInput_hi[11343:11328]},
     {loadUnit_maskInput_hi[11327:11312]},
     {loadUnit_maskInput_hi[11311:11296]},
     {loadUnit_maskInput_hi[11295:11280]},
     {loadUnit_maskInput_hi[11279:11264]},
     {loadUnit_maskInput_hi[11263:11248]},
     {loadUnit_maskInput_hi[11247:11232]},
     {loadUnit_maskInput_hi[11231:11216]},
     {loadUnit_maskInput_hi[11215:11200]},
     {loadUnit_maskInput_hi[11199:11184]},
     {loadUnit_maskInput_hi[11183:11168]},
     {loadUnit_maskInput_hi[11167:11152]},
     {loadUnit_maskInput_hi[11151:11136]},
     {loadUnit_maskInput_hi[11135:11120]},
     {loadUnit_maskInput_hi[11119:11104]},
     {loadUnit_maskInput_hi[11103:11088]},
     {loadUnit_maskInput_hi[11087:11072]},
     {loadUnit_maskInput_hi[11071:11056]},
     {loadUnit_maskInput_hi[11055:11040]},
     {loadUnit_maskInput_hi[11039:11024]},
     {loadUnit_maskInput_hi[11023:11008]},
     {loadUnit_maskInput_hi[11007:10992]},
     {loadUnit_maskInput_hi[10991:10976]},
     {loadUnit_maskInput_hi[10975:10960]},
     {loadUnit_maskInput_hi[10959:10944]},
     {loadUnit_maskInput_hi[10943:10928]},
     {loadUnit_maskInput_hi[10927:10912]},
     {loadUnit_maskInput_hi[10911:10896]},
     {loadUnit_maskInput_hi[10895:10880]},
     {loadUnit_maskInput_hi[10879:10864]},
     {loadUnit_maskInput_hi[10863:10848]},
     {loadUnit_maskInput_hi[10847:10832]},
     {loadUnit_maskInput_hi[10831:10816]},
     {loadUnit_maskInput_hi[10815:10800]},
     {loadUnit_maskInput_hi[10799:10784]},
     {loadUnit_maskInput_hi[10783:10768]},
     {loadUnit_maskInput_hi[10767:10752]},
     {loadUnit_maskInput_hi[10751:10736]},
     {loadUnit_maskInput_hi[10735:10720]},
     {loadUnit_maskInput_hi[10719:10704]},
     {loadUnit_maskInput_hi[10703:10688]},
     {loadUnit_maskInput_hi[10687:10672]},
     {loadUnit_maskInput_hi[10671:10656]},
     {loadUnit_maskInput_hi[10655:10640]},
     {loadUnit_maskInput_hi[10639:10624]},
     {loadUnit_maskInput_hi[10623:10608]},
     {loadUnit_maskInput_hi[10607:10592]},
     {loadUnit_maskInput_hi[10591:10576]},
     {loadUnit_maskInput_hi[10575:10560]},
     {loadUnit_maskInput_hi[10559:10544]},
     {loadUnit_maskInput_hi[10543:10528]},
     {loadUnit_maskInput_hi[10527:10512]},
     {loadUnit_maskInput_hi[10511:10496]},
     {loadUnit_maskInput_hi[10495:10480]},
     {loadUnit_maskInput_hi[10479:10464]},
     {loadUnit_maskInput_hi[10463:10448]},
     {loadUnit_maskInput_hi[10447:10432]},
     {loadUnit_maskInput_hi[10431:10416]},
     {loadUnit_maskInput_hi[10415:10400]},
     {loadUnit_maskInput_hi[10399:10384]},
     {loadUnit_maskInput_hi[10383:10368]},
     {loadUnit_maskInput_hi[10367:10352]},
     {loadUnit_maskInput_hi[10351:10336]},
     {loadUnit_maskInput_hi[10335:10320]},
     {loadUnit_maskInput_hi[10319:10304]},
     {loadUnit_maskInput_hi[10303:10288]},
     {loadUnit_maskInput_hi[10287:10272]},
     {loadUnit_maskInput_hi[10271:10256]},
     {loadUnit_maskInput_hi[10255:10240]},
     {loadUnit_maskInput_hi[10239:10224]},
     {loadUnit_maskInput_hi[10223:10208]},
     {loadUnit_maskInput_hi[10207:10192]},
     {loadUnit_maskInput_hi[10191:10176]},
     {loadUnit_maskInput_hi[10175:10160]},
     {loadUnit_maskInput_hi[10159:10144]},
     {loadUnit_maskInput_hi[10143:10128]},
     {loadUnit_maskInput_hi[10127:10112]},
     {loadUnit_maskInput_hi[10111:10096]},
     {loadUnit_maskInput_hi[10095:10080]},
     {loadUnit_maskInput_hi[10079:10064]},
     {loadUnit_maskInput_hi[10063:10048]},
     {loadUnit_maskInput_hi[10047:10032]},
     {loadUnit_maskInput_hi[10031:10016]},
     {loadUnit_maskInput_hi[10015:10000]},
     {loadUnit_maskInput_hi[9999:9984]},
     {loadUnit_maskInput_hi[9983:9968]},
     {loadUnit_maskInput_hi[9967:9952]},
     {loadUnit_maskInput_hi[9951:9936]},
     {loadUnit_maskInput_hi[9935:9920]},
     {loadUnit_maskInput_hi[9919:9904]},
     {loadUnit_maskInput_hi[9903:9888]},
     {loadUnit_maskInput_hi[9887:9872]},
     {loadUnit_maskInput_hi[9871:9856]},
     {loadUnit_maskInput_hi[9855:9840]},
     {loadUnit_maskInput_hi[9839:9824]},
     {loadUnit_maskInput_hi[9823:9808]},
     {loadUnit_maskInput_hi[9807:9792]},
     {loadUnit_maskInput_hi[9791:9776]},
     {loadUnit_maskInput_hi[9775:9760]},
     {loadUnit_maskInput_hi[9759:9744]},
     {loadUnit_maskInput_hi[9743:9728]},
     {loadUnit_maskInput_hi[9727:9712]},
     {loadUnit_maskInput_hi[9711:9696]},
     {loadUnit_maskInput_hi[9695:9680]},
     {loadUnit_maskInput_hi[9679:9664]},
     {loadUnit_maskInput_hi[9663:9648]},
     {loadUnit_maskInput_hi[9647:9632]},
     {loadUnit_maskInput_hi[9631:9616]},
     {loadUnit_maskInput_hi[9615:9600]},
     {loadUnit_maskInput_hi[9599:9584]},
     {loadUnit_maskInput_hi[9583:9568]},
     {loadUnit_maskInput_hi[9567:9552]},
     {loadUnit_maskInput_hi[9551:9536]},
     {loadUnit_maskInput_hi[9535:9520]},
     {loadUnit_maskInput_hi[9519:9504]},
     {loadUnit_maskInput_hi[9503:9488]},
     {loadUnit_maskInput_hi[9487:9472]},
     {loadUnit_maskInput_hi[9471:9456]},
     {loadUnit_maskInput_hi[9455:9440]},
     {loadUnit_maskInput_hi[9439:9424]},
     {loadUnit_maskInput_hi[9423:9408]},
     {loadUnit_maskInput_hi[9407:9392]},
     {loadUnit_maskInput_hi[9391:9376]},
     {loadUnit_maskInput_hi[9375:9360]},
     {loadUnit_maskInput_hi[9359:9344]},
     {loadUnit_maskInput_hi[9343:9328]},
     {loadUnit_maskInput_hi[9327:9312]},
     {loadUnit_maskInput_hi[9311:9296]},
     {loadUnit_maskInput_hi[9295:9280]},
     {loadUnit_maskInput_hi[9279:9264]},
     {loadUnit_maskInput_hi[9263:9248]},
     {loadUnit_maskInput_hi[9247:9232]},
     {loadUnit_maskInput_hi[9231:9216]},
     {loadUnit_maskInput_hi[9215:9200]},
     {loadUnit_maskInput_hi[9199:9184]},
     {loadUnit_maskInput_hi[9183:9168]},
     {loadUnit_maskInput_hi[9167:9152]},
     {loadUnit_maskInput_hi[9151:9136]},
     {loadUnit_maskInput_hi[9135:9120]},
     {loadUnit_maskInput_hi[9119:9104]},
     {loadUnit_maskInput_hi[9103:9088]},
     {loadUnit_maskInput_hi[9087:9072]},
     {loadUnit_maskInput_hi[9071:9056]},
     {loadUnit_maskInput_hi[9055:9040]},
     {loadUnit_maskInput_hi[9039:9024]},
     {loadUnit_maskInput_hi[9023:9008]},
     {loadUnit_maskInput_hi[9007:8992]},
     {loadUnit_maskInput_hi[8991:8976]},
     {loadUnit_maskInput_hi[8975:8960]},
     {loadUnit_maskInput_hi[8959:8944]},
     {loadUnit_maskInput_hi[8943:8928]},
     {loadUnit_maskInput_hi[8927:8912]},
     {loadUnit_maskInput_hi[8911:8896]},
     {loadUnit_maskInput_hi[8895:8880]},
     {loadUnit_maskInput_hi[8879:8864]},
     {loadUnit_maskInput_hi[8863:8848]},
     {loadUnit_maskInput_hi[8847:8832]},
     {loadUnit_maskInput_hi[8831:8816]},
     {loadUnit_maskInput_hi[8815:8800]},
     {loadUnit_maskInput_hi[8799:8784]},
     {loadUnit_maskInput_hi[8783:8768]},
     {loadUnit_maskInput_hi[8767:8752]},
     {loadUnit_maskInput_hi[8751:8736]},
     {loadUnit_maskInput_hi[8735:8720]},
     {loadUnit_maskInput_hi[8719:8704]},
     {loadUnit_maskInput_hi[8703:8688]},
     {loadUnit_maskInput_hi[8687:8672]},
     {loadUnit_maskInput_hi[8671:8656]},
     {loadUnit_maskInput_hi[8655:8640]},
     {loadUnit_maskInput_hi[8639:8624]},
     {loadUnit_maskInput_hi[8623:8608]},
     {loadUnit_maskInput_hi[8607:8592]},
     {loadUnit_maskInput_hi[8591:8576]},
     {loadUnit_maskInput_hi[8575:8560]},
     {loadUnit_maskInput_hi[8559:8544]},
     {loadUnit_maskInput_hi[8543:8528]},
     {loadUnit_maskInput_hi[8527:8512]},
     {loadUnit_maskInput_hi[8511:8496]},
     {loadUnit_maskInput_hi[8495:8480]},
     {loadUnit_maskInput_hi[8479:8464]},
     {loadUnit_maskInput_hi[8463:8448]},
     {loadUnit_maskInput_hi[8447:8432]},
     {loadUnit_maskInput_hi[8431:8416]},
     {loadUnit_maskInput_hi[8415:8400]},
     {loadUnit_maskInput_hi[8399:8384]},
     {loadUnit_maskInput_hi[8383:8368]},
     {loadUnit_maskInput_hi[8367:8352]},
     {loadUnit_maskInput_hi[8351:8336]},
     {loadUnit_maskInput_hi[8335:8320]},
     {loadUnit_maskInput_hi[8319:8304]},
     {loadUnit_maskInput_hi[8303:8288]},
     {loadUnit_maskInput_hi[8287:8272]},
     {loadUnit_maskInput_hi[8271:8256]},
     {loadUnit_maskInput_hi[8255:8240]},
     {loadUnit_maskInput_hi[8239:8224]},
     {loadUnit_maskInput_hi[8223:8208]},
     {loadUnit_maskInput_hi[8207:8192]},
     {loadUnit_maskInput_hi[8191:8176]},
     {loadUnit_maskInput_hi[8175:8160]},
     {loadUnit_maskInput_hi[8159:8144]},
     {loadUnit_maskInput_hi[8143:8128]},
     {loadUnit_maskInput_hi[8127:8112]},
     {loadUnit_maskInput_hi[8111:8096]},
     {loadUnit_maskInput_hi[8095:8080]},
     {loadUnit_maskInput_hi[8079:8064]},
     {loadUnit_maskInput_hi[8063:8048]},
     {loadUnit_maskInput_hi[8047:8032]},
     {loadUnit_maskInput_hi[8031:8016]},
     {loadUnit_maskInput_hi[8015:8000]},
     {loadUnit_maskInput_hi[7999:7984]},
     {loadUnit_maskInput_hi[7983:7968]},
     {loadUnit_maskInput_hi[7967:7952]},
     {loadUnit_maskInput_hi[7951:7936]},
     {loadUnit_maskInput_hi[7935:7920]},
     {loadUnit_maskInput_hi[7919:7904]},
     {loadUnit_maskInput_hi[7903:7888]},
     {loadUnit_maskInput_hi[7887:7872]},
     {loadUnit_maskInput_hi[7871:7856]},
     {loadUnit_maskInput_hi[7855:7840]},
     {loadUnit_maskInput_hi[7839:7824]},
     {loadUnit_maskInput_hi[7823:7808]},
     {loadUnit_maskInput_hi[7807:7792]},
     {loadUnit_maskInput_hi[7791:7776]},
     {loadUnit_maskInput_hi[7775:7760]},
     {loadUnit_maskInput_hi[7759:7744]},
     {loadUnit_maskInput_hi[7743:7728]},
     {loadUnit_maskInput_hi[7727:7712]},
     {loadUnit_maskInput_hi[7711:7696]},
     {loadUnit_maskInput_hi[7695:7680]},
     {loadUnit_maskInput_hi[7679:7664]},
     {loadUnit_maskInput_hi[7663:7648]},
     {loadUnit_maskInput_hi[7647:7632]},
     {loadUnit_maskInput_hi[7631:7616]},
     {loadUnit_maskInput_hi[7615:7600]},
     {loadUnit_maskInput_hi[7599:7584]},
     {loadUnit_maskInput_hi[7583:7568]},
     {loadUnit_maskInput_hi[7567:7552]},
     {loadUnit_maskInput_hi[7551:7536]},
     {loadUnit_maskInput_hi[7535:7520]},
     {loadUnit_maskInput_hi[7519:7504]},
     {loadUnit_maskInput_hi[7503:7488]},
     {loadUnit_maskInput_hi[7487:7472]},
     {loadUnit_maskInput_hi[7471:7456]},
     {loadUnit_maskInput_hi[7455:7440]},
     {loadUnit_maskInput_hi[7439:7424]},
     {loadUnit_maskInput_hi[7423:7408]},
     {loadUnit_maskInput_hi[7407:7392]},
     {loadUnit_maskInput_hi[7391:7376]},
     {loadUnit_maskInput_hi[7375:7360]},
     {loadUnit_maskInput_hi[7359:7344]},
     {loadUnit_maskInput_hi[7343:7328]},
     {loadUnit_maskInput_hi[7327:7312]},
     {loadUnit_maskInput_hi[7311:7296]},
     {loadUnit_maskInput_hi[7295:7280]},
     {loadUnit_maskInput_hi[7279:7264]},
     {loadUnit_maskInput_hi[7263:7248]},
     {loadUnit_maskInput_hi[7247:7232]},
     {loadUnit_maskInput_hi[7231:7216]},
     {loadUnit_maskInput_hi[7215:7200]},
     {loadUnit_maskInput_hi[7199:7184]},
     {loadUnit_maskInput_hi[7183:7168]},
     {loadUnit_maskInput_hi[7167:7152]},
     {loadUnit_maskInput_hi[7151:7136]},
     {loadUnit_maskInput_hi[7135:7120]},
     {loadUnit_maskInput_hi[7119:7104]},
     {loadUnit_maskInput_hi[7103:7088]},
     {loadUnit_maskInput_hi[7087:7072]},
     {loadUnit_maskInput_hi[7071:7056]},
     {loadUnit_maskInput_hi[7055:7040]},
     {loadUnit_maskInput_hi[7039:7024]},
     {loadUnit_maskInput_hi[7023:7008]},
     {loadUnit_maskInput_hi[7007:6992]},
     {loadUnit_maskInput_hi[6991:6976]},
     {loadUnit_maskInput_hi[6975:6960]},
     {loadUnit_maskInput_hi[6959:6944]},
     {loadUnit_maskInput_hi[6943:6928]},
     {loadUnit_maskInput_hi[6927:6912]},
     {loadUnit_maskInput_hi[6911:6896]},
     {loadUnit_maskInput_hi[6895:6880]},
     {loadUnit_maskInput_hi[6879:6864]},
     {loadUnit_maskInput_hi[6863:6848]},
     {loadUnit_maskInput_hi[6847:6832]},
     {loadUnit_maskInput_hi[6831:6816]},
     {loadUnit_maskInput_hi[6815:6800]},
     {loadUnit_maskInput_hi[6799:6784]},
     {loadUnit_maskInput_hi[6783:6768]},
     {loadUnit_maskInput_hi[6767:6752]},
     {loadUnit_maskInput_hi[6751:6736]},
     {loadUnit_maskInput_hi[6735:6720]},
     {loadUnit_maskInput_hi[6719:6704]},
     {loadUnit_maskInput_hi[6703:6688]},
     {loadUnit_maskInput_hi[6687:6672]},
     {loadUnit_maskInput_hi[6671:6656]},
     {loadUnit_maskInput_hi[6655:6640]},
     {loadUnit_maskInput_hi[6639:6624]},
     {loadUnit_maskInput_hi[6623:6608]},
     {loadUnit_maskInput_hi[6607:6592]},
     {loadUnit_maskInput_hi[6591:6576]},
     {loadUnit_maskInput_hi[6575:6560]},
     {loadUnit_maskInput_hi[6559:6544]},
     {loadUnit_maskInput_hi[6543:6528]},
     {loadUnit_maskInput_hi[6527:6512]},
     {loadUnit_maskInput_hi[6511:6496]},
     {loadUnit_maskInput_hi[6495:6480]},
     {loadUnit_maskInput_hi[6479:6464]},
     {loadUnit_maskInput_hi[6463:6448]},
     {loadUnit_maskInput_hi[6447:6432]},
     {loadUnit_maskInput_hi[6431:6416]},
     {loadUnit_maskInput_hi[6415:6400]},
     {loadUnit_maskInput_hi[6399:6384]},
     {loadUnit_maskInput_hi[6383:6368]},
     {loadUnit_maskInput_hi[6367:6352]},
     {loadUnit_maskInput_hi[6351:6336]},
     {loadUnit_maskInput_hi[6335:6320]},
     {loadUnit_maskInput_hi[6319:6304]},
     {loadUnit_maskInput_hi[6303:6288]},
     {loadUnit_maskInput_hi[6287:6272]},
     {loadUnit_maskInput_hi[6271:6256]},
     {loadUnit_maskInput_hi[6255:6240]},
     {loadUnit_maskInput_hi[6239:6224]},
     {loadUnit_maskInput_hi[6223:6208]},
     {loadUnit_maskInput_hi[6207:6192]},
     {loadUnit_maskInput_hi[6191:6176]},
     {loadUnit_maskInput_hi[6175:6160]},
     {loadUnit_maskInput_hi[6159:6144]},
     {loadUnit_maskInput_hi[6143:6128]},
     {loadUnit_maskInput_hi[6127:6112]},
     {loadUnit_maskInput_hi[6111:6096]},
     {loadUnit_maskInput_hi[6095:6080]},
     {loadUnit_maskInput_hi[6079:6064]},
     {loadUnit_maskInput_hi[6063:6048]},
     {loadUnit_maskInput_hi[6047:6032]},
     {loadUnit_maskInput_hi[6031:6016]},
     {loadUnit_maskInput_hi[6015:6000]},
     {loadUnit_maskInput_hi[5999:5984]},
     {loadUnit_maskInput_hi[5983:5968]},
     {loadUnit_maskInput_hi[5967:5952]},
     {loadUnit_maskInput_hi[5951:5936]},
     {loadUnit_maskInput_hi[5935:5920]},
     {loadUnit_maskInput_hi[5919:5904]},
     {loadUnit_maskInput_hi[5903:5888]},
     {loadUnit_maskInput_hi[5887:5872]},
     {loadUnit_maskInput_hi[5871:5856]},
     {loadUnit_maskInput_hi[5855:5840]},
     {loadUnit_maskInput_hi[5839:5824]},
     {loadUnit_maskInput_hi[5823:5808]},
     {loadUnit_maskInput_hi[5807:5792]},
     {loadUnit_maskInput_hi[5791:5776]},
     {loadUnit_maskInput_hi[5775:5760]},
     {loadUnit_maskInput_hi[5759:5744]},
     {loadUnit_maskInput_hi[5743:5728]},
     {loadUnit_maskInput_hi[5727:5712]},
     {loadUnit_maskInput_hi[5711:5696]},
     {loadUnit_maskInput_hi[5695:5680]},
     {loadUnit_maskInput_hi[5679:5664]},
     {loadUnit_maskInput_hi[5663:5648]},
     {loadUnit_maskInput_hi[5647:5632]},
     {loadUnit_maskInput_hi[5631:5616]},
     {loadUnit_maskInput_hi[5615:5600]},
     {loadUnit_maskInput_hi[5599:5584]},
     {loadUnit_maskInput_hi[5583:5568]},
     {loadUnit_maskInput_hi[5567:5552]},
     {loadUnit_maskInput_hi[5551:5536]},
     {loadUnit_maskInput_hi[5535:5520]},
     {loadUnit_maskInput_hi[5519:5504]},
     {loadUnit_maskInput_hi[5503:5488]},
     {loadUnit_maskInput_hi[5487:5472]},
     {loadUnit_maskInput_hi[5471:5456]},
     {loadUnit_maskInput_hi[5455:5440]},
     {loadUnit_maskInput_hi[5439:5424]},
     {loadUnit_maskInput_hi[5423:5408]},
     {loadUnit_maskInput_hi[5407:5392]},
     {loadUnit_maskInput_hi[5391:5376]},
     {loadUnit_maskInput_hi[5375:5360]},
     {loadUnit_maskInput_hi[5359:5344]},
     {loadUnit_maskInput_hi[5343:5328]},
     {loadUnit_maskInput_hi[5327:5312]},
     {loadUnit_maskInput_hi[5311:5296]},
     {loadUnit_maskInput_hi[5295:5280]},
     {loadUnit_maskInput_hi[5279:5264]},
     {loadUnit_maskInput_hi[5263:5248]},
     {loadUnit_maskInput_hi[5247:5232]},
     {loadUnit_maskInput_hi[5231:5216]},
     {loadUnit_maskInput_hi[5215:5200]},
     {loadUnit_maskInput_hi[5199:5184]},
     {loadUnit_maskInput_hi[5183:5168]},
     {loadUnit_maskInput_hi[5167:5152]},
     {loadUnit_maskInput_hi[5151:5136]},
     {loadUnit_maskInput_hi[5135:5120]},
     {loadUnit_maskInput_hi[5119:5104]},
     {loadUnit_maskInput_hi[5103:5088]},
     {loadUnit_maskInput_hi[5087:5072]},
     {loadUnit_maskInput_hi[5071:5056]},
     {loadUnit_maskInput_hi[5055:5040]},
     {loadUnit_maskInput_hi[5039:5024]},
     {loadUnit_maskInput_hi[5023:5008]},
     {loadUnit_maskInput_hi[5007:4992]},
     {loadUnit_maskInput_hi[4991:4976]},
     {loadUnit_maskInput_hi[4975:4960]},
     {loadUnit_maskInput_hi[4959:4944]},
     {loadUnit_maskInput_hi[4943:4928]},
     {loadUnit_maskInput_hi[4927:4912]},
     {loadUnit_maskInput_hi[4911:4896]},
     {loadUnit_maskInput_hi[4895:4880]},
     {loadUnit_maskInput_hi[4879:4864]},
     {loadUnit_maskInput_hi[4863:4848]},
     {loadUnit_maskInput_hi[4847:4832]},
     {loadUnit_maskInput_hi[4831:4816]},
     {loadUnit_maskInput_hi[4815:4800]},
     {loadUnit_maskInput_hi[4799:4784]},
     {loadUnit_maskInput_hi[4783:4768]},
     {loadUnit_maskInput_hi[4767:4752]},
     {loadUnit_maskInput_hi[4751:4736]},
     {loadUnit_maskInput_hi[4735:4720]},
     {loadUnit_maskInput_hi[4719:4704]},
     {loadUnit_maskInput_hi[4703:4688]},
     {loadUnit_maskInput_hi[4687:4672]},
     {loadUnit_maskInput_hi[4671:4656]},
     {loadUnit_maskInput_hi[4655:4640]},
     {loadUnit_maskInput_hi[4639:4624]},
     {loadUnit_maskInput_hi[4623:4608]},
     {loadUnit_maskInput_hi[4607:4592]},
     {loadUnit_maskInput_hi[4591:4576]},
     {loadUnit_maskInput_hi[4575:4560]},
     {loadUnit_maskInput_hi[4559:4544]},
     {loadUnit_maskInput_hi[4543:4528]},
     {loadUnit_maskInput_hi[4527:4512]},
     {loadUnit_maskInput_hi[4511:4496]},
     {loadUnit_maskInput_hi[4495:4480]},
     {loadUnit_maskInput_hi[4479:4464]},
     {loadUnit_maskInput_hi[4463:4448]},
     {loadUnit_maskInput_hi[4447:4432]},
     {loadUnit_maskInput_hi[4431:4416]},
     {loadUnit_maskInput_hi[4415:4400]},
     {loadUnit_maskInput_hi[4399:4384]},
     {loadUnit_maskInput_hi[4383:4368]},
     {loadUnit_maskInput_hi[4367:4352]},
     {loadUnit_maskInput_hi[4351:4336]},
     {loadUnit_maskInput_hi[4335:4320]},
     {loadUnit_maskInput_hi[4319:4304]},
     {loadUnit_maskInput_hi[4303:4288]},
     {loadUnit_maskInput_hi[4287:4272]},
     {loadUnit_maskInput_hi[4271:4256]},
     {loadUnit_maskInput_hi[4255:4240]},
     {loadUnit_maskInput_hi[4239:4224]},
     {loadUnit_maskInput_hi[4223:4208]},
     {loadUnit_maskInput_hi[4207:4192]},
     {loadUnit_maskInput_hi[4191:4176]},
     {loadUnit_maskInput_hi[4175:4160]},
     {loadUnit_maskInput_hi[4159:4144]},
     {loadUnit_maskInput_hi[4143:4128]},
     {loadUnit_maskInput_hi[4127:4112]},
     {loadUnit_maskInput_hi[4111:4096]},
     {loadUnit_maskInput_hi[4095:4080]},
     {loadUnit_maskInput_hi[4079:4064]},
     {loadUnit_maskInput_hi[4063:4048]},
     {loadUnit_maskInput_hi[4047:4032]},
     {loadUnit_maskInput_hi[4031:4016]},
     {loadUnit_maskInput_hi[4015:4000]},
     {loadUnit_maskInput_hi[3999:3984]},
     {loadUnit_maskInput_hi[3983:3968]},
     {loadUnit_maskInput_hi[3967:3952]},
     {loadUnit_maskInput_hi[3951:3936]},
     {loadUnit_maskInput_hi[3935:3920]},
     {loadUnit_maskInput_hi[3919:3904]},
     {loadUnit_maskInput_hi[3903:3888]},
     {loadUnit_maskInput_hi[3887:3872]},
     {loadUnit_maskInput_hi[3871:3856]},
     {loadUnit_maskInput_hi[3855:3840]},
     {loadUnit_maskInput_hi[3839:3824]},
     {loadUnit_maskInput_hi[3823:3808]},
     {loadUnit_maskInput_hi[3807:3792]},
     {loadUnit_maskInput_hi[3791:3776]},
     {loadUnit_maskInput_hi[3775:3760]},
     {loadUnit_maskInput_hi[3759:3744]},
     {loadUnit_maskInput_hi[3743:3728]},
     {loadUnit_maskInput_hi[3727:3712]},
     {loadUnit_maskInput_hi[3711:3696]},
     {loadUnit_maskInput_hi[3695:3680]},
     {loadUnit_maskInput_hi[3679:3664]},
     {loadUnit_maskInput_hi[3663:3648]},
     {loadUnit_maskInput_hi[3647:3632]},
     {loadUnit_maskInput_hi[3631:3616]},
     {loadUnit_maskInput_hi[3615:3600]},
     {loadUnit_maskInput_hi[3599:3584]},
     {loadUnit_maskInput_hi[3583:3568]},
     {loadUnit_maskInput_hi[3567:3552]},
     {loadUnit_maskInput_hi[3551:3536]},
     {loadUnit_maskInput_hi[3535:3520]},
     {loadUnit_maskInput_hi[3519:3504]},
     {loadUnit_maskInput_hi[3503:3488]},
     {loadUnit_maskInput_hi[3487:3472]},
     {loadUnit_maskInput_hi[3471:3456]},
     {loadUnit_maskInput_hi[3455:3440]},
     {loadUnit_maskInput_hi[3439:3424]},
     {loadUnit_maskInput_hi[3423:3408]},
     {loadUnit_maskInput_hi[3407:3392]},
     {loadUnit_maskInput_hi[3391:3376]},
     {loadUnit_maskInput_hi[3375:3360]},
     {loadUnit_maskInput_hi[3359:3344]},
     {loadUnit_maskInput_hi[3343:3328]},
     {loadUnit_maskInput_hi[3327:3312]},
     {loadUnit_maskInput_hi[3311:3296]},
     {loadUnit_maskInput_hi[3295:3280]},
     {loadUnit_maskInput_hi[3279:3264]},
     {loadUnit_maskInput_hi[3263:3248]},
     {loadUnit_maskInput_hi[3247:3232]},
     {loadUnit_maskInput_hi[3231:3216]},
     {loadUnit_maskInput_hi[3215:3200]},
     {loadUnit_maskInput_hi[3199:3184]},
     {loadUnit_maskInput_hi[3183:3168]},
     {loadUnit_maskInput_hi[3167:3152]},
     {loadUnit_maskInput_hi[3151:3136]},
     {loadUnit_maskInput_hi[3135:3120]},
     {loadUnit_maskInput_hi[3119:3104]},
     {loadUnit_maskInput_hi[3103:3088]},
     {loadUnit_maskInput_hi[3087:3072]},
     {loadUnit_maskInput_hi[3071:3056]},
     {loadUnit_maskInput_hi[3055:3040]},
     {loadUnit_maskInput_hi[3039:3024]},
     {loadUnit_maskInput_hi[3023:3008]},
     {loadUnit_maskInput_hi[3007:2992]},
     {loadUnit_maskInput_hi[2991:2976]},
     {loadUnit_maskInput_hi[2975:2960]},
     {loadUnit_maskInput_hi[2959:2944]},
     {loadUnit_maskInput_hi[2943:2928]},
     {loadUnit_maskInput_hi[2927:2912]},
     {loadUnit_maskInput_hi[2911:2896]},
     {loadUnit_maskInput_hi[2895:2880]},
     {loadUnit_maskInput_hi[2879:2864]},
     {loadUnit_maskInput_hi[2863:2848]},
     {loadUnit_maskInput_hi[2847:2832]},
     {loadUnit_maskInput_hi[2831:2816]},
     {loadUnit_maskInput_hi[2815:2800]},
     {loadUnit_maskInput_hi[2799:2784]},
     {loadUnit_maskInput_hi[2783:2768]},
     {loadUnit_maskInput_hi[2767:2752]},
     {loadUnit_maskInput_hi[2751:2736]},
     {loadUnit_maskInput_hi[2735:2720]},
     {loadUnit_maskInput_hi[2719:2704]},
     {loadUnit_maskInput_hi[2703:2688]},
     {loadUnit_maskInput_hi[2687:2672]},
     {loadUnit_maskInput_hi[2671:2656]},
     {loadUnit_maskInput_hi[2655:2640]},
     {loadUnit_maskInput_hi[2639:2624]},
     {loadUnit_maskInput_hi[2623:2608]},
     {loadUnit_maskInput_hi[2607:2592]},
     {loadUnit_maskInput_hi[2591:2576]},
     {loadUnit_maskInput_hi[2575:2560]},
     {loadUnit_maskInput_hi[2559:2544]},
     {loadUnit_maskInput_hi[2543:2528]},
     {loadUnit_maskInput_hi[2527:2512]},
     {loadUnit_maskInput_hi[2511:2496]},
     {loadUnit_maskInput_hi[2495:2480]},
     {loadUnit_maskInput_hi[2479:2464]},
     {loadUnit_maskInput_hi[2463:2448]},
     {loadUnit_maskInput_hi[2447:2432]},
     {loadUnit_maskInput_hi[2431:2416]},
     {loadUnit_maskInput_hi[2415:2400]},
     {loadUnit_maskInput_hi[2399:2384]},
     {loadUnit_maskInput_hi[2383:2368]},
     {loadUnit_maskInput_hi[2367:2352]},
     {loadUnit_maskInput_hi[2351:2336]},
     {loadUnit_maskInput_hi[2335:2320]},
     {loadUnit_maskInput_hi[2319:2304]},
     {loadUnit_maskInput_hi[2303:2288]},
     {loadUnit_maskInput_hi[2287:2272]},
     {loadUnit_maskInput_hi[2271:2256]},
     {loadUnit_maskInput_hi[2255:2240]},
     {loadUnit_maskInput_hi[2239:2224]},
     {loadUnit_maskInput_hi[2223:2208]},
     {loadUnit_maskInput_hi[2207:2192]},
     {loadUnit_maskInput_hi[2191:2176]},
     {loadUnit_maskInput_hi[2175:2160]},
     {loadUnit_maskInput_hi[2159:2144]},
     {loadUnit_maskInput_hi[2143:2128]},
     {loadUnit_maskInput_hi[2127:2112]},
     {loadUnit_maskInput_hi[2111:2096]},
     {loadUnit_maskInput_hi[2095:2080]},
     {loadUnit_maskInput_hi[2079:2064]},
     {loadUnit_maskInput_hi[2063:2048]},
     {loadUnit_maskInput_hi[2047:2032]},
     {loadUnit_maskInput_hi[2031:2016]},
     {loadUnit_maskInput_hi[2015:2000]},
     {loadUnit_maskInput_hi[1999:1984]},
     {loadUnit_maskInput_hi[1983:1968]},
     {loadUnit_maskInput_hi[1967:1952]},
     {loadUnit_maskInput_hi[1951:1936]},
     {loadUnit_maskInput_hi[1935:1920]},
     {loadUnit_maskInput_hi[1919:1904]},
     {loadUnit_maskInput_hi[1903:1888]},
     {loadUnit_maskInput_hi[1887:1872]},
     {loadUnit_maskInput_hi[1871:1856]},
     {loadUnit_maskInput_hi[1855:1840]},
     {loadUnit_maskInput_hi[1839:1824]},
     {loadUnit_maskInput_hi[1823:1808]},
     {loadUnit_maskInput_hi[1807:1792]},
     {loadUnit_maskInput_hi[1791:1776]},
     {loadUnit_maskInput_hi[1775:1760]},
     {loadUnit_maskInput_hi[1759:1744]},
     {loadUnit_maskInput_hi[1743:1728]},
     {loadUnit_maskInput_hi[1727:1712]},
     {loadUnit_maskInput_hi[1711:1696]},
     {loadUnit_maskInput_hi[1695:1680]},
     {loadUnit_maskInput_hi[1679:1664]},
     {loadUnit_maskInput_hi[1663:1648]},
     {loadUnit_maskInput_hi[1647:1632]},
     {loadUnit_maskInput_hi[1631:1616]},
     {loadUnit_maskInput_hi[1615:1600]},
     {loadUnit_maskInput_hi[1599:1584]},
     {loadUnit_maskInput_hi[1583:1568]},
     {loadUnit_maskInput_hi[1567:1552]},
     {loadUnit_maskInput_hi[1551:1536]},
     {loadUnit_maskInput_hi[1535:1520]},
     {loadUnit_maskInput_hi[1519:1504]},
     {loadUnit_maskInput_hi[1503:1488]},
     {loadUnit_maskInput_hi[1487:1472]},
     {loadUnit_maskInput_hi[1471:1456]},
     {loadUnit_maskInput_hi[1455:1440]},
     {loadUnit_maskInput_hi[1439:1424]},
     {loadUnit_maskInput_hi[1423:1408]},
     {loadUnit_maskInput_hi[1407:1392]},
     {loadUnit_maskInput_hi[1391:1376]},
     {loadUnit_maskInput_hi[1375:1360]},
     {loadUnit_maskInput_hi[1359:1344]},
     {loadUnit_maskInput_hi[1343:1328]},
     {loadUnit_maskInput_hi[1327:1312]},
     {loadUnit_maskInput_hi[1311:1296]},
     {loadUnit_maskInput_hi[1295:1280]},
     {loadUnit_maskInput_hi[1279:1264]},
     {loadUnit_maskInput_hi[1263:1248]},
     {loadUnit_maskInput_hi[1247:1232]},
     {loadUnit_maskInput_hi[1231:1216]},
     {loadUnit_maskInput_hi[1215:1200]},
     {loadUnit_maskInput_hi[1199:1184]},
     {loadUnit_maskInput_hi[1183:1168]},
     {loadUnit_maskInput_hi[1167:1152]},
     {loadUnit_maskInput_hi[1151:1136]},
     {loadUnit_maskInput_hi[1135:1120]},
     {loadUnit_maskInput_hi[1119:1104]},
     {loadUnit_maskInput_hi[1103:1088]},
     {loadUnit_maskInput_hi[1087:1072]},
     {loadUnit_maskInput_hi[1071:1056]},
     {loadUnit_maskInput_hi[1055:1040]},
     {loadUnit_maskInput_hi[1039:1024]},
     {loadUnit_maskInput_hi[1023:1008]},
     {loadUnit_maskInput_hi[1007:992]},
     {loadUnit_maskInput_hi[991:976]},
     {loadUnit_maskInput_hi[975:960]},
     {loadUnit_maskInput_hi[959:944]},
     {loadUnit_maskInput_hi[943:928]},
     {loadUnit_maskInput_hi[927:912]},
     {loadUnit_maskInput_hi[911:896]},
     {loadUnit_maskInput_hi[895:880]},
     {loadUnit_maskInput_hi[879:864]},
     {loadUnit_maskInput_hi[863:848]},
     {loadUnit_maskInput_hi[847:832]},
     {loadUnit_maskInput_hi[831:816]},
     {loadUnit_maskInput_hi[815:800]},
     {loadUnit_maskInput_hi[799:784]},
     {loadUnit_maskInput_hi[783:768]},
     {loadUnit_maskInput_hi[767:752]},
     {loadUnit_maskInput_hi[751:736]},
     {loadUnit_maskInput_hi[735:720]},
     {loadUnit_maskInput_hi[719:704]},
     {loadUnit_maskInput_hi[703:688]},
     {loadUnit_maskInput_hi[687:672]},
     {loadUnit_maskInput_hi[671:656]},
     {loadUnit_maskInput_hi[655:640]},
     {loadUnit_maskInput_hi[639:624]},
     {loadUnit_maskInput_hi[623:608]},
     {loadUnit_maskInput_hi[607:592]},
     {loadUnit_maskInput_hi[591:576]},
     {loadUnit_maskInput_hi[575:560]},
     {loadUnit_maskInput_hi[559:544]},
     {loadUnit_maskInput_hi[543:528]},
     {loadUnit_maskInput_hi[527:512]},
     {loadUnit_maskInput_hi[511:496]},
     {loadUnit_maskInput_hi[495:480]},
     {loadUnit_maskInput_hi[479:464]},
     {loadUnit_maskInput_hi[463:448]},
     {loadUnit_maskInput_hi[447:432]},
     {loadUnit_maskInput_hi[431:416]},
     {loadUnit_maskInput_hi[415:400]},
     {loadUnit_maskInput_hi[399:384]},
     {loadUnit_maskInput_hi[383:368]},
     {loadUnit_maskInput_hi[367:352]},
     {loadUnit_maskInput_hi[351:336]},
     {loadUnit_maskInput_hi[335:320]},
     {loadUnit_maskInput_hi[319:304]},
     {loadUnit_maskInput_hi[303:288]},
     {loadUnit_maskInput_hi[287:272]},
     {loadUnit_maskInput_hi[271:256]},
     {loadUnit_maskInput_hi[255:240]},
     {loadUnit_maskInput_hi[239:224]},
     {loadUnit_maskInput_hi[223:208]},
     {loadUnit_maskInput_hi[207:192]},
     {loadUnit_maskInput_hi[191:176]},
     {loadUnit_maskInput_hi[175:160]},
     {loadUnit_maskInput_hi[159:144]},
     {loadUnit_maskInput_hi[143:128]},
     {loadUnit_maskInput_hi[127:112]},
     {loadUnit_maskInput_hi[111:96]},
     {loadUnit_maskInput_hi[95:80]},
     {loadUnit_maskInput_hi[79:64]},
     {loadUnit_maskInput_hi[63:48]},
     {loadUnit_maskInput_hi[47:32]},
     {loadUnit_maskInput_hi[31:16]},
     {loadUnit_maskInput_hi[15:0]},
     {loadUnit_maskInput_lo[16383:16368]},
     {loadUnit_maskInput_lo[16367:16352]},
     {loadUnit_maskInput_lo[16351:16336]},
     {loadUnit_maskInput_lo[16335:16320]},
     {loadUnit_maskInput_lo[16319:16304]},
     {loadUnit_maskInput_lo[16303:16288]},
     {loadUnit_maskInput_lo[16287:16272]},
     {loadUnit_maskInput_lo[16271:16256]},
     {loadUnit_maskInput_lo[16255:16240]},
     {loadUnit_maskInput_lo[16239:16224]},
     {loadUnit_maskInput_lo[16223:16208]},
     {loadUnit_maskInput_lo[16207:16192]},
     {loadUnit_maskInput_lo[16191:16176]},
     {loadUnit_maskInput_lo[16175:16160]},
     {loadUnit_maskInput_lo[16159:16144]},
     {loadUnit_maskInput_lo[16143:16128]},
     {loadUnit_maskInput_lo[16127:16112]},
     {loadUnit_maskInput_lo[16111:16096]},
     {loadUnit_maskInput_lo[16095:16080]},
     {loadUnit_maskInput_lo[16079:16064]},
     {loadUnit_maskInput_lo[16063:16048]},
     {loadUnit_maskInput_lo[16047:16032]},
     {loadUnit_maskInput_lo[16031:16016]},
     {loadUnit_maskInput_lo[16015:16000]},
     {loadUnit_maskInput_lo[15999:15984]},
     {loadUnit_maskInput_lo[15983:15968]},
     {loadUnit_maskInput_lo[15967:15952]},
     {loadUnit_maskInput_lo[15951:15936]},
     {loadUnit_maskInput_lo[15935:15920]},
     {loadUnit_maskInput_lo[15919:15904]},
     {loadUnit_maskInput_lo[15903:15888]},
     {loadUnit_maskInput_lo[15887:15872]},
     {loadUnit_maskInput_lo[15871:15856]},
     {loadUnit_maskInput_lo[15855:15840]},
     {loadUnit_maskInput_lo[15839:15824]},
     {loadUnit_maskInput_lo[15823:15808]},
     {loadUnit_maskInput_lo[15807:15792]},
     {loadUnit_maskInput_lo[15791:15776]},
     {loadUnit_maskInput_lo[15775:15760]},
     {loadUnit_maskInput_lo[15759:15744]},
     {loadUnit_maskInput_lo[15743:15728]},
     {loadUnit_maskInput_lo[15727:15712]},
     {loadUnit_maskInput_lo[15711:15696]},
     {loadUnit_maskInput_lo[15695:15680]},
     {loadUnit_maskInput_lo[15679:15664]},
     {loadUnit_maskInput_lo[15663:15648]},
     {loadUnit_maskInput_lo[15647:15632]},
     {loadUnit_maskInput_lo[15631:15616]},
     {loadUnit_maskInput_lo[15615:15600]},
     {loadUnit_maskInput_lo[15599:15584]},
     {loadUnit_maskInput_lo[15583:15568]},
     {loadUnit_maskInput_lo[15567:15552]},
     {loadUnit_maskInput_lo[15551:15536]},
     {loadUnit_maskInput_lo[15535:15520]},
     {loadUnit_maskInput_lo[15519:15504]},
     {loadUnit_maskInput_lo[15503:15488]},
     {loadUnit_maskInput_lo[15487:15472]},
     {loadUnit_maskInput_lo[15471:15456]},
     {loadUnit_maskInput_lo[15455:15440]},
     {loadUnit_maskInput_lo[15439:15424]},
     {loadUnit_maskInput_lo[15423:15408]},
     {loadUnit_maskInput_lo[15407:15392]},
     {loadUnit_maskInput_lo[15391:15376]},
     {loadUnit_maskInput_lo[15375:15360]},
     {loadUnit_maskInput_lo[15359:15344]},
     {loadUnit_maskInput_lo[15343:15328]},
     {loadUnit_maskInput_lo[15327:15312]},
     {loadUnit_maskInput_lo[15311:15296]},
     {loadUnit_maskInput_lo[15295:15280]},
     {loadUnit_maskInput_lo[15279:15264]},
     {loadUnit_maskInput_lo[15263:15248]},
     {loadUnit_maskInput_lo[15247:15232]},
     {loadUnit_maskInput_lo[15231:15216]},
     {loadUnit_maskInput_lo[15215:15200]},
     {loadUnit_maskInput_lo[15199:15184]},
     {loadUnit_maskInput_lo[15183:15168]},
     {loadUnit_maskInput_lo[15167:15152]},
     {loadUnit_maskInput_lo[15151:15136]},
     {loadUnit_maskInput_lo[15135:15120]},
     {loadUnit_maskInput_lo[15119:15104]},
     {loadUnit_maskInput_lo[15103:15088]},
     {loadUnit_maskInput_lo[15087:15072]},
     {loadUnit_maskInput_lo[15071:15056]},
     {loadUnit_maskInput_lo[15055:15040]},
     {loadUnit_maskInput_lo[15039:15024]},
     {loadUnit_maskInput_lo[15023:15008]},
     {loadUnit_maskInput_lo[15007:14992]},
     {loadUnit_maskInput_lo[14991:14976]},
     {loadUnit_maskInput_lo[14975:14960]},
     {loadUnit_maskInput_lo[14959:14944]},
     {loadUnit_maskInput_lo[14943:14928]},
     {loadUnit_maskInput_lo[14927:14912]},
     {loadUnit_maskInput_lo[14911:14896]},
     {loadUnit_maskInput_lo[14895:14880]},
     {loadUnit_maskInput_lo[14879:14864]},
     {loadUnit_maskInput_lo[14863:14848]},
     {loadUnit_maskInput_lo[14847:14832]},
     {loadUnit_maskInput_lo[14831:14816]},
     {loadUnit_maskInput_lo[14815:14800]},
     {loadUnit_maskInput_lo[14799:14784]},
     {loadUnit_maskInput_lo[14783:14768]},
     {loadUnit_maskInput_lo[14767:14752]},
     {loadUnit_maskInput_lo[14751:14736]},
     {loadUnit_maskInput_lo[14735:14720]},
     {loadUnit_maskInput_lo[14719:14704]},
     {loadUnit_maskInput_lo[14703:14688]},
     {loadUnit_maskInput_lo[14687:14672]},
     {loadUnit_maskInput_lo[14671:14656]},
     {loadUnit_maskInput_lo[14655:14640]},
     {loadUnit_maskInput_lo[14639:14624]},
     {loadUnit_maskInput_lo[14623:14608]},
     {loadUnit_maskInput_lo[14607:14592]},
     {loadUnit_maskInput_lo[14591:14576]},
     {loadUnit_maskInput_lo[14575:14560]},
     {loadUnit_maskInput_lo[14559:14544]},
     {loadUnit_maskInput_lo[14543:14528]},
     {loadUnit_maskInput_lo[14527:14512]},
     {loadUnit_maskInput_lo[14511:14496]},
     {loadUnit_maskInput_lo[14495:14480]},
     {loadUnit_maskInput_lo[14479:14464]},
     {loadUnit_maskInput_lo[14463:14448]},
     {loadUnit_maskInput_lo[14447:14432]},
     {loadUnit_maskInput_lo[14431:14416]},
     {loadUnit_maskInput_lo[14415:14400]},
     {loadUnit_maskInput_lo[14399:14384]},
     {loadUnit_maskInput_lo[14383:14368]},
     {loadUnit_maskInput_lo[14367:14352]},
     {loadUnit_maskInput_lo[14351:14336]},
     {loadUnit_maskInput_lo[14335:14320]},
     {loadUnit_maskInput_lo[14319:14304]},
     {loadUnit_maskInput_lo[14303:14288]},
     {loadUnit_maskInput_lo[14287:14272]},
     {loadUnit_maskInput_lo[14271:14256]},
     {loadUnit_maskInput_lo[14255:14240]},
     {loadUnit_maskInput_lo[14239:14224]},
     {loadUnit_maskInput_lo[14223:14208]},
     {loadUnit_maskInput_lo[14207:14192]},
     {loadUnit_maskInput_lo[14191:14176]},
     {loadUnit_maskInput_lo[14175:14160]},
     {loadUnit_maskInput_lo[14159:14144]},
     {loadUnit_maskInput_lo[14143:14128]},
     {loadUnit_maskInput_lo[14127:14112]},
     {loadUnit_maskInput_lo[14111:14096]},
     {loadUnit_maskInput_lo[14095:14080]},
     {loadUnit_maskInput_lo[14079:14064]},
     {loadUnit_maskInput_lo[14063:14048]},
     {loadUnit_maskInput_lo[14047:14032]},
     {loadUnit_maskInput_lo[14031:14016]},
     {loadUnit_maskInput_lo[14015:14000]},
     {loadUnit_maskInput_lo[13999:13984]},
     {loadUnit_maskInput_lo[13983:13968]},
     {loadUnit_maskInput_lo[13967:13952]},
     {loadUnit_maskInput_lo[13951:13936]},
     {loadUnit_maskInput_lo[13935:13920]},
     {loadUnit_maskInput_lo[13919:13904]},
     {loadUnit_maskInput_lo[13903:13888]},
     {loadUnit_maskInput_lo[13887:13872]},
     {loadUnit_maskInput_lo[13871:13856]},
     {loadUnit_maskInput_lo[13855:13840]},
     {loadUnit_maskInput_lo[13839:13824]},
     {loadUnit_maskInput_lo[13823:13808]},
     {loadUnit_maskInput_lo[13807:13792]},
     {loadUnit_maskInput_lo[13791:13776]},
     {loadUnit_maskInput_lo[13775:13760]},
     {loadUnit_maskInput_lo[13759:13744]},
     {loadUnit_maskInput_lo[13743:13728]},
     {loadUnit_maskInput_lo[13727:13712]},
     {loadUnit_maskInput_lo[13711:13696]},
     {loadUnit_maskInput_lo[13695:13680]},
     {loadUnit_maskInput_lo[13679:13664]},
     {loadUnit_maskInput_lo[13663:13648]},
     {loadUnit_maskInput_lo[13647:13632]},
     {loadUnit_maskInput_lo[13631:13616]},
     {loadUnit_maskInput_lo[13615:13600]},
     {loadUnit_maskInput_lo[13599:13584]},
     {loadUnit_maskInput_lo[13583:13568]},
     {loadUnit_maskInput_lo[13567:13552]},
     {loadUnit_maskInput_lo[13551:13536]},
     {loadUnit_maskInput_lo[13535:13520]},
     {loadUnit_maskInput_lo[13519:13504]},
     {loadUnit_maskInput_lo[13503:13488]},
     {loadUnit_maskInput_lo[13487:13472]},
     {loadUnit_maskInput_lo[13471:13456]},
     {loadUnit_maskInput_lo[13455:13440]},
     {loadUnit_maskInput_lo[13439:13424]},
     {loadUnit_maskInput_lo[13423:13408]},
     {loadUnit_maskInput_lo[13407:13392]},
     {loadUnit_maskInput_lo[13391:13376]},
     {loadUnit_maskInput_lo[13375:13360]},
     {loadUnit_maskInput_lo[13359:13344]},
     {loadUnit_maskInput_lo[13343:13328]},
     {loadUnit_maskInput_lo[13327:13312]},
     {loadUnit_maskInput_lo[13311:13296]},
     {loadUnit_maskInput_lo[13295:13280]},
     {loadUnit_maskInput_lo[13279:13264]},
     {loadUnit_maskInput_lo[13263:13248]},
     {loadUnit_maskInput_lo[13247:13232]},
     {loadUnit_maskInput_lo[13231:13216]},
     {loadUnit_maskInput_lo[13215:13200]},
     {loadUnit_maskInput_lo[13199:13184]},
     {loadUnit_maskInput_lo[13183:13168]},
     {loadUnit_maskInput_lo[13167:13152]},
     {loadUnit_maskInput_lo[13151:13136]},
     {loadUnit_maskInput_lo[13135:13120]},
     {loadUnit_maskInput_lo[13119:13104]},
     {loadUnit_maskInput_lo[13103:13088]},
     {loadUnit_maskInput_lo[13087:13072]},
     {loadUnit_maskInput_lo[13071:13056]},
     {loadUnit_maskInput_lo[13055:13040]},
     {loadUnit_maskInput_lo[13039:13024]},
     {loadUnit_maskInput_lo[13023:13008]},
     {loadUnit_maskInput_lo[13007:12992]},
     {loadUnit_maskInput_lo[12991:12976]},
     {loadUnit_maskInput_lo[12975:12960]},
     {loadUnit_maskInput_lo[12959:12944]},
     {loadUnit_maskInput_lo[12943:12928]},
     {loadUnit_maskInput_lo[12927:12912]},
     {loadUnit_maskInput_lo[12911:12896]},
     {loadUnit_maskInput_lo[12895:12880]},
     {loadUnit_maskInput_lo[12879:12864]},
     {loadUnit_maskInput_lo[12863:12848]},
     {loadUnit_maskInput_lo[12847:12832]},
     {loadUnit_maskInput_lo[12831:12816]},
     {loadUnit_maskInput_lo[12815:12800]},
     {loadUnit_maskInput_lo[12799:12784]},
     {loadUnit_maskInput_lo[12783:12768]},
     {loadUnit_maskInput_lo[12767:12752]},
     {loadUnit_maskInput_lo[12751:12736]},
     {loadUnit_maskInput_lo[12735:12720]},
     {loadUnit_maskInput_lo[12719:12704]},
     {loadUnit_maskInput_lo[12703:12688]},
     {loadUnit_maskInput_lo[12687:12672]},
     {loadUnit_maskInput_lo[12671:12656]},
     {loadUnit_maskInput_lo[12655:12640]},
     {loadUnit_maskInput_lo[12639:12624]},
     {loadUnit_maskInput_lo[12623:12608]},
     {loadUnit_maskInput_lo[12607:12592]},
     {loadUnit_maskInput_lo[12591:12576]},
     {loadUnit_maskInput_lo[12575:12560]},
     {loadUnit_maskInput_lo[12559:12544]},
     {loadUnit_maskInput_lo[12543:12528]},
     {loadUnit_maskInput_lo[12527:12512]},
     {loadUnit_maskInput_lo[12511:12496]},
     {loadUnit_maskInput_lo[12495:12480]},
     {loadUnit_maskInput_lo[12479:12464]},
     {loadUnit_maskInput_lo[12463:12448]},
     {loadUnit_maskInput_lo[12447:12432]},
     {loadUnit_maskInput_lo[12431:12416]},
     {loadUnit_maskInput_lo[12415:12400]},
     {loadUnit_maskInput_lo[12399:12384]},
     {loadUnit_maskInput_lo[12383:12368]},
     {loadUnit_maskInput_lo[12367:12352]},
     {loadUnit_maskInput_lo[12351:12336]},
     {loadUnit_maskInput_lo[12335:12320]},
     {loadUnit_maskInput_lo[12319:12304]},
     {loadUnit_maskInput_lo[12303:12288]},
     {loadUnit_maskInput_lo[12287:12272]},
     {loadUnit_maskInput_lo[12271:12256]},
     {loadUnit_maskInput_lo[12255:12240]},
     {loadUnit_maskInput_lo[12239:12224]},
     {loadUnit_maskInput_lo[12223:12208]},
     {loadUnit_maskInput_lo[12207:12192]},
     {loadUnit_maskInput_lo[12191:12176]},
     {loadUnit_maskInput_lo[12175:12160]},
     {loadUnit_maskInput_lo[12159:12144]},
     {loadUnit_maskInput_lo[12143:12128]},
     {loadUnit_maskInput_lo[12127:12112]},
     {loadUnit_maskInput_lo[12111:12096]},
     {loadUnit_maskInput_lo[12095:12080]},
     {loadUnit_maskInput_lo[12079:12064]},
     {loadUnit_maskInput_lo[12063:12048]},
     {loadUnit_maskInput_lo[12047:12032]},
     {loadUnit_maskInput_lo[12031:12016]},
     {loadUnit_maskInput_lo[12015:12000]},
     {loadUnit_maskInput_lo[11999:11984]},
     {loadUnit_maskInput_lo[11983:11968]},
     {loadUnit_maskInput_lo[11967:11952]},
     {loadUnit_maskInput_lo[11951:11936]},
     {loadUnit_maskInput_lo[11935:11920]},
     {loadUnit_maskInput_lo[11919:11904]},
     {loadUnit_maskInput_lo[11903:11888]},
     {loadUnit_maskInput_lo[11887:11872]},
     {loadUnit_maskInput_lo[11871:11856]},
     {loadUnit_maskInput_lo[11855:11840]},
     {loadUnit_maskInput_lo[11839:11824]},
     {loadUnit_maskInput_lo[11823:11808]},
     {loadUnit_maskInput_lo[11807:11792]},
     {loadUnit_maskInput_lo[11791:11776]},
     {loadUnit_maskInput_lo[11775:11760]},
     {loadUnit_maskInput_lo[11759:11744]},
     {loadUnit_maskInput_lo[11743:11728]},
     {loadUnit_maskInput_lo[11727:11712]},
     {loadUnit_maskInput_lo[11711:11696]},
     {loadUnit_maskInput_lo[11695:11680]},
     {loadUnit_maskInput_lo[11679:11664]},
     {loadUnit_maskInput_lo[11663:11648]},
     {loadUnit_maskInput_lo[11647:11632]},
     {loadUnit_maskInput_lo[11631:11616]},
     {loadUnit_maskInput_lo[11615:11600]},
     {loadUnit_maskInput_lo[11599:11584]},
     {loadUnit_maskInput_lo[11583:11568]},
     {loadUnit_maskInput_lo[11567:11552]},
     {loadUnit_maskInput_lo[11551:11536]},
     {loadUnit_maskInput_lo[11535:11520]},
     {loadUnit_maskInput_lo[11519:11504]},
     {loadUnit_maskInput_lo[11503:11488]},
     {loadUnit_maskInput_lo[11487:11472]},
     {loadUnit_maskInput_lo[11471:11456]},
     {loadUnit_maskInput_lo[11455:11440]},
     {loadUnit_maskInput_lo[11439:11424]},
     {loadUnit_maskInput_lo[11423:11408]},
     {loadUnit_maskInput_lo[11407:11392]},
     {loadUnit_maskInput_lo[11391:11376]},
     {loadUnit_maskInput_lo[11375:11360]},
     {loadUnit_maskInput_lo[11359:11344]},
     {loadUnit_maskInput_lo[11343:11328]},
     {loadUnit_maskInput_lo[11327:11312]},
     {loadUnit_maskInput_lo[11311:11296]},
     {loadUnit_maskInput_lo[11295:11280]},
     {loadUnit_maskInput_lo[11279:11264]},
     {loadUnit_maskInput_lo[11263:11248]},
     {loadUnit_maskInput_lo[11247:11232]},
     {loadUnit_maskInput_lo[11231:11216]},
     {loadUnit_maskInput_lo[11215:11200]},
     {loadUnit_maskInput_lo[11199:11184]},
     {loadUnit_maskInput_lo[11183:11168]},
     {loadUnit_maskInput_lo[11167:11152]},
     {loadUnit_maskInput_lo[11151:11136]},
     {loadUnit_maskInput_lo[11135:11120]},
     {loadUnit_maskInput_lo[11119:11104]},
     {loadUnit_maskInput_lo[11103:11088]},
     {loadUnit_maskInput_lo[11087:11072]},
     {loadUnit_maskInput_lo[11071:11056]},
     {loadUnit_maskInput_lo[11055:11040]},
     {loadUnit_maskInput_lo[11039:11024]},
     {loadUnit_maskInput_lo[11023:11008]},
     {loadUnit_maskInput_lo[11007:10992]},
     {loadUnit_maskInput_lo[10991:10976]},
     {loadUnit_maskInput_lo[10975:10960]},
     {loadUnit_maskInput_lo[10959:10944]},
     {loadUnit_maskInput_lo[10943:10928]},
     {loadUnit_maskInput_lo[10927:10912]},
     {loadUnit_maskInput_lo[10911:10896]},
     {loadUnit_maskInput_lo[10895:10880]},
     {loadUnit_maskInput_lo[10879:10864]},
     {loadUnit_maskInput_lo[10863:10848]},
     {loadUnit_maskInput_lo[10847:10832]},
     {loadUnit_maskInput_lo[10831:10816]},
     {loadUnit_maskInput_lo[10815:10800]},
     {loadUnit_maskInput_lo[10799:10784]},
     {loadUnit_maskInput_lo[10783:10768]},
     {loadUnit_maskInput_lo[10767:10752]},
     {loadUnit_maskInput_lo[10751:10736]},
     {loadUnit_maskInput_lo[10735:10720]},
     {loadUnit_maskInput_lo[10719:10704]},
     {loadUnit_maskInput_lo[10703:10688]},
     {loadUnit_maskInput_lo[10687:10672]},
     {loadUnit_maskInput_lo[10671:10656]},
     {loadUnit_maskInput_lo[10655:10640]},
     {loadUnit_maskInput_lo[10639:10624]},
     {loadUnit_maskInput_lo[10623:10608]},
     {loadUnit_maskInput_lo[10607:10592]},
     {loadUnit_maskInput_lo[10591:10576]},
     {loadUnit_maskInput_lo[10575:10560]},
     {loadUnit_maskInput_lo[10559:10544]},
     {loadUnit_maskInput_lo[10543:10528]},
     {loadUnit_maskInput_lo[10527:10512]},
     {loadUnit_maskInput_lo[10511:10496]},
     {loadUnit_maskInput_lo[10495:10480]},
     {loadUnit_maskInput_lo[10479:10464]},
     {loadUnit_maskInput_lo[10463:10448]},
     {loadUnit_maskInput_lo[10447:10432]},
     {loadUnit_maskInput_lo[10431:10416]},
     {loadUnit_maskInput_lo[10415:10400]},
     {loadUnit_maskInput_lo[10399:10384]},
     {loadUnit_maskInput_lo[10383:10368]},
     {loadUnit_maskInput_lo[10367:10352]},
     {loadUnit_maskInput_lo[10351:10336]},
     {loadUnit_maskInput_lo[10335:10320]},
     {loadUnit_maskInput_lo[10319:10304]},
     {loadUnit_maskInput_lo[10303:10288]},
     {loadUnit_maskInput_lo[10287:10272]},
     {loadUnit_maskInput_lo[10271:10256]},
     {loadUnit_maskInput_lo[10255:10240]},
     {loadUnit_maskInput_lo[10239:10224]},
     {loadUnit_maskInput_lo[10223:10208]},
     {loadUnit_maskInput_lo[10207:10192]},
     {loadUnit_maskInput_lo[10191:10176]},
     {loadUnit_maskInput_lo[10175:10160]},
     {loadUnit_maskInput_lo[10159:10144]},
     {loadUnit_maskInput_lo[10143:10128]},
     {loadUnit_maskInput_lo[10127:10112]},
     {loadUnit_maskInput_lo[10111:10096]},
     {loadUnit_maskInput_lo[10095:10080]},
     {loadUnit_maskInput_lo[10079:10064]},
     {loadUnit_maskInput_lo[10063:10048]},
     {loadUnit_maskInput_lo[10047:10032]},
     {loadUnit_maskInput_lo[10031:10016]},
     {loadUnit_maskInput_lo[10015:10000]},
     {loadUnit_maskInput_lo[9999:9984]},
     {loadUnit_maskInput_lo[9983:9968]},
     {loadUnit_maskInput_lo[9967:9952]},
     {loadUnit_maskInput_lo[9951:9936]},
     {loadUnit_maskInput_lo[9935:9920]},
     {loadUnit_maskInput_lo[9919:9904]},
     {loadUnit_maskInput_lo[9903:9888]},
     {loadUnit_maskInput_lo[9887:9872]},
     {loadUnit_maskInput_lo[9871:9856]},
     {loadUnit_maskInput_lo[9855:9840]},
     {loadUnit_maskInput_lo[9839:9824]},
     {loadUnit_maskInput_lo[9823:9808]},
     {loadUnit_maskInput_lo[9807:9792]},
     {loadUnit_maskInput_lo[9791:9776]},
     {loadUnit_maskInput_lo[9775:9760]},
     {loadUnit_maskInput_lo[9759:9744]},
     {loadUnit_maskInput_lo[9743:9728]},
     {loadUnit_maskInput_lo[9727:9712]},
     {loadUnit_maskInput_lo[9711:9696]},
     {loadUnit_maskInput_lo[9695:9680]},
     {loadUnit_maskInput_lo[9679:9664]},
     {loadUnit_maskInput_lo[9663:9648]},
     {loadUnit_maskInput_lo[9647:9632]},
     {loadUnit_maskInput_lo[9631:9616]},
     {loadUnit_maskInput_lo[9615:9600]},
     {loadUnit_maskInput_lo[9599:9584]},
     {loadUnit_maskInput_lo[9583:9568]},
     {loadUnit_maskInput_lo[9567:9552]},
     {loadUnit_maskInput_lo[9551:9536]},
     {loadUnit_maskInput_lo[9535:9520]},
     {loadUnit_maskInput_lo[9519:9504]},
     {loadUnit_maskInput_lo[9503:9488]},
     {loadUnit_maskInput_lo[9487:9472]},
     {loadUnit_maskInput_lo[9471:9456]},
     {loadUnit_maskInput_lo[9455:9440]},
     {loadUnit_maskInput_lo[9439:9424]},
     {loadUnit_maskInput_lo[9423:9408]},
     {loadUnit_maskInput_lo[9407:9392]},
     {loadUnit_maskInput_lo[9391:9376]},
     {loadUnit_maskInput_lo[9375:9360]},
     {loadUnit_maskInput_lo[9359:9344]},
     {loadUnit_maskInput_lo[9343:9328]},
     {loadUnit_maskInput_lo[9327:9312]},
     {loadUnit_maskInput_lo[9311:9296]},
     {loadUnit_maskInput_lo[9295:9280]},
     {loadUnit_maskInput_lo[9279:9264]},
     {loadUnit_maskInput_lo[9263:9248]},
     {loadUnit_maskInput_lo[9247:9232]},
     {loadUnit_maskInput_lo[9231:9216]},
     {loadUnit_maskInput_lo[9215:9200]},
     {loadUnit_maskInput_lo[9199:9184]},
     {loadUnit_maskInput_lo[9183:9168]},
     {loadUnit_maskInput_lo[9167:9152]},
     {loadUnit_maskInput_lo[9151:9136]},
     {loadUnit_maskInput_lo[9135:9120]},
     {loadUnit_maskInput_lo[9119:9104]},
     {loadUnit_maskInput_lo[9103:9088]},
     {loadUnit_maskInput_lo[9087:9072]},
     {loadUnit_maskInput_lo[9071:9056]},
     {loadUnit_maskInput_lo[9055:9040]},
     {loadUnit_maskInput_lo[9039:9024]},
     {loadUnit_maskInput_lo[9023:9008]},
     {loadUnit_maskInput_lo[9007:8992]},
     {loadUnit_maskInput_lo[8991:8976]},
     {loadUnit_maskInput_lo[8975:8960]},
     {loadUnit_maskInput_lo[8959:8944]},
     {loadUnit_maskInput_lo[8943:8928]},
     {loadUnit_maskInput_lo[8927:8912]},
     {loadUnit_maskInput_lo[8911:8896]},
     {loadUnit_maskInput_lo[8895:8880]},
     {loadUnit_maskInput_lo[8879:8864]},
     {loadUnit_maskInput_lo[8863:8848]},
     {loadUnit_maskInput_lo[8847:8832]},
     {loadUnit_maskInput_lo[8831:8816]},
     {loadUnit_maskInput_lo[8815:8800]},
     {loadUnit_maskInput_lo[8799:8784]},
     {loadUnit_maskInput_lo[8783:8768]},
     {loadUnit_maskInput_lo[8767:8752]},
     {loadUnit_maskInput_lo[8751:8736]},
     {loadUnit_maskInput_lo[8735:8720]},
     {loadUnit_maskInput_lo[8719:8704]},
     {loadUnit_maskInput_lo[8703:8688]},
     {loadUnit_maskInput_lo[8687:8672]},
     {loadUnit_maskInput_lo[8671:8656]},
     {loadUnit_maskInput_lo[8655:8640]},
     {loadUnit_maskInput_lo[8639:8624]},
     {loadUnit_maskInput_lo[8623:8608]},
     {loadUnit_maskInput_lo[8607:8592]},
     {loadUnit_maskInput_lo[8591:8576]},
     {loadUnit_maskInput_lo[8575:8560]},
     {loadUnit_maskInput_lo[8559:8544]},
     {loadUnit_maskInput_lo[8543:8528]},
     {loadUnit_maskInput_lo[8527:8512]},
     {loadUnit_maskInput_lo[8511:8496]},
     {loadUnit_maskInput_lo[8495:8480]},
     {loadUnit_maskInput_lo[8479:8464]},
     {loadUnit_maskInput_lo[8463:8448]},
     {loadUnit_maskInput_lo[8447:8432]},
     {loadUnit_maskInput_lo[8431:8416]},
     {loadUnit_maskInput_lo[8415:8400]},
     {loadUnit_maskInput_lo[8399:8384]},
     {loadUnit_maskInput_lo[8383:8368]},
     {loadUnit_maskInput_lo[8367:8352]},
     {loadUnit_maskInput_lo[8351:8336]},
     {loadUnit_maskInput_lo[8335:8320]},
     {loadUnit_maskInput_lo[8319:8304]},
     {loadUnit_maskInput_lo[8303:8288]},
     {loadUnit_maskInput_lo[8287:8272]},
     {loadUnit_maskInput_lo[8271:8256]},
     {loadUnit_maskInput_lo[8255:8240]},
     {loadUnit_maskInput_lo[8239:8224]},
     {loadUnit_maskInput_lo[8223:8208]},
     {loadUnit_maskInput_lo[8207:8192]},
     {loadUnit_maskInput_lo[8191:8176]},
     {loadUnit_maskInput_lo[8175:8160]},
     {loadUnit_maskInput_lo[8159:8144]},
     {loadUnit_maskInput_lo[8143:8128]},
     {loadUnit_maskInput_lo[8127:8112]},
     {loadUnit_maskInput_lo[8111:8096]},
     {loadUnit_maskInput_lo[8095:8080]},
     {loadUnit_maskInput_lo[8079:8064]},
     {loadUnit_maskInput_lo[8063:8048]},
     {loadUnit_maskInput_lo[8047:8032]},
     {loadUnit_maskInput_lo[8031:8016]},
     {loadUnit_maskInput_lo[8015:8000]},
     {loadUnit_maskInput_lo[7999:7984]},
     {loadUnit_maskInput_lo[7983:7968]},
     {loadUnit_maskInput_lo[7967:7952]},
     {loadUnit_maskInput_lo[7951:7936]},
     {loadUnit_maskInput_lo[7935:7920]},
     {loadUnit_maskInput_lo[7919:7904]},
     {loadUnit_maskInput_lo[7903:7888]},
     {loadUnit_maskInput_lo[7887:7872]},
     {loadUnit_maskInput_lo[7871:7856]},
     {loadUnit_maskInput_lo[7855:7840]},
     {loadUnit_maskInput_lo[7839:7824]},
     {loadUnit_maskInput_lo[7823:7808]},
     {loadUnit_maskInput_lo[7807:7792]},
     {loadUnit_maskInput_lo[7791:7776]},
     {loadUnit_maskInput_lo[7775:7760]},
     {loadUnit_maskInput_lo[7759:7744]},
     {loadUnit_maskInput_lo[7743:7728]},
     {loadUnit_maskInput_lo[7727:7712]},
     {loadUnit_maskInput_lo[7711:7696]},
     {loadUnit_maskInput_lo[7695:7680]},
     {loadUnit_maskInput_lo[7679:7664]},
     {loadUnit_maskInput_lo[7663:7648]},
     {loadUnit_maskInput_lo[7647:7632]},
     {loadUnit_maskInput_lo[7631:7616]},
     {loadUnit_maskInput_lo[7615:7600]},
     {loadUnit_maskInput_lo[7599:7584]},
     {loadUnit_maskInput_lo[7583:7568]},
     {loadUnit_maskInput_lo[7567:7552]},
     {loadUnit_maskInput_lo[7551:7536]},
     {loadUnit_maskInput_lo[7535:7520]},
     {loadUnit_maskInput_lo[7519:7504]},
     {loadUnit_maskInput_lo[7503:7488]},
     {loadUnit_maskInput_lo[7487:7472]},
     {loadUnit_maskInput_lo[7471:7456]},
     {loadUnit_maskInput_lo[7455:7440]},
     {loadUnit_maskInput_lo[7439:7424]},
     {loadUnit_maskInput_lo[7423:7408]},
     {loadUnit_maskInput_lo[7407:7392]},
     {loadUnit_maskInput_lo[7391:7376]},
     {loadUnit_maskInput_lo[7375:7360]},
     {loadUnit_maskInput_lo[7359:7344]},
     {loadUnit_maskInput_lo[7343:7328]},
     {loadUnit_maskInput_lo[7327:7312]},
     {loadUnit_maskInput_lo[7311:7296]},
     {loadUnit_maskInput_lo[7295:7280]},
     {loadUnit_maskInput_lo[7279:7264]},
     {loadUnit_maskInput_lo[7263:7248]},
     {loadUnit_maskInput_lo[7247:7232]},
     {loadUnit_maskInput_lo[7231:7216]},
     {loadUnit_maskInput_lo[7215:7200]},
     {loadUnit_maskInput_lo[7199:7184]},
     {loadUnit_maskInput_lo[7183:7168]},
     {loadUnit_maskInput_lo[7167:7152]},
     {loadUnit_maskInput_lo[7151:7136]},
     {loadUnit_maskInput_lo[7135:7120]},
     {loadUnit_maskInput_lo[7119:7104]},
     {loadUnit_maskInput_lo[7103:7088]},
     {loadUnit_maskInput_lo[7087:7072]},
     {loadUnit_maskInput_lo[7071:7056]},
     {loadUnit_maskInput_lo[7055:7040]},
     {loadUnit_maskInput_lo[7039:7024]},
     {loadUnit_maskInput_lo[7023:7008]},
     {loadUnit_maskInput_lo[7007:6992]},
     {loadUnit_maskInput_lo[6991:6976]},
     {loadUnit_maskInput_lo[6975:6960]},
     {loadUnit_maskInput_lo[6959:6944]},
     {loadUnit_maskInput_lo[6943:6928]},
     {loadUnit_maskInput_lo[6927:6912]},
     {loadUnit_maskInput_lo[6911:6896]},
     {loadUnit_maskInput_lo[6895:6880]},
     {loadUnit_maskInput_lo[6879:6864]},
     {loadUnit_maskInput_lo[6863:6848]},
     {loadUnit_maskInput_lo[6847:6832]},
     {loadUnit_maskInput_lo[6831:6816]},
     {loadUnit_maskInput_lo[6815:6800]},
     {loadUnit_maskInput_lo[6799:6784]},
     {loadUnit_maskInput_lo[6783:6768]},
     {loadUnit_maskInput_lo[6767:6752]},
     {loadUnit_maskInput_lo[6751:6736]},
     {loadUnit_maskInput_lo[6735:6720]},
     {loadUnit_maskInput_lo[6719:6704]},
     {loadUnit_maskInput_lo[6703:6688]},
     {loadUnit_maskInput_lo[6687:6672]},
     {loadUnit_maskInput_lo[6671:6656]},
     {loadUnit_maskInput_lo[6655:6640]},
     {loadUnit_maskInput_lo[6639:6624]},
     {loadUnit_maskInput_lo[6623:6608]},
     {loadUnit_maskInput_lo[6607:6592]},
     {loadUnit_maskInput_lo[6591:6576]},
     {loadUnit_maskInput_lo[6575:6560]},
     {loadUnit_maskInput_lo[6559:6544]},
     {loadUnit_maskInput_lo[6543:6528]},
     {loadUnit_maskInput_lo[6527:6512]},
     {loadUnit_maskInput_lo[6511:6496]},
     {loadUnit_maskInput_lo[6495:6480]},
     {loadUnit_maskInput_lo[6479:6464]},
     {loadUnit_maskInput_lo[6463:6448]},
     {loadUnit_maskInput_lo[6447:6432]},
     {loadUnit_maskInput_lo[6431:6416]},
     {loadUnit_maskInput_lo[6415:6400]},
     {loadUnit_maskInput_lo[6399:6384]},
     {loadUnit_maskInput_lo[6383:6368]},
     {loadUnit_maskInput_lo[6367:6352]},
     {loadUnit_maskInput_lo[6351:6336]},
     {loadUnit_maskInput_lo[6335:6320]},
     {loadUnit_maskInput_lo[6319:6304]},
     {loadUnit_maskInput_lo[6303:6288]},
     {loadUnit_maskInput_lo[6287:6272]},
     {loadUnit_maskInput_lo[6271:6256]},
     {loadUnit_maskInput_lo[6255:6240]},
     {loadUnit_maskInput_lo[6239:6224]},
     {loadUnit_maskInput_lo[6223:6208]},
     {loadUnit_maskInput_lo[6207:6192]},
     {loadUnit_maskInput_lo[6191:6176]},
     {loadUnit_maskInput_lo[6175:6160]},
     {loadUnit_maskInput_lo[6159:6144]},
     {loadUnit_maskInput_lo[6143:6128]},
     {loadUnit_maskInput_lo[6127:6112]},
     {loadUnit_maskInput_lo[6111:6096]},
     {loadUnit_maskInput_lo[6095:6080]},
     {loadUnit_maskInput_lo[6079:6064]},
     {loadUnit_maskInput_lo[6063:6048]},
     {loadUnit_maskInput_lo[6047:6032]},
     {loadUnit_maskInput_lo[6031:6016]},
     {loadUnit_maskInput_lo[6015:6000]},
     {loadUnit_maskInput_lo[5999:5984]},
     {loadUnit_maskInput_lo[5983:5968]},
     {loadUnit_maskInput_lo[5967:5952]},
     {loadUnit_maskInput_lo[5951:5936]},
     {loadUnit_maskInput_lo[5935:5920]},
     {loadUnit_maskInput_lo[5919:5904]},
     {loadUnit_maskInput_lo[5903:5888]},
     {loadUnit_maskInput_lo[5887:5872]},
     {loadUnit_maskInput_lo[5871:5856]},
     {loadUnit_maskInput_lo[5855:5840]},
     {loadUnit_maskInput_lo[5839:5824]},
     {loadUnit_maskInput_lo[5823:5808]},
     {loadUnit_maskInput_lo[5807:5792]},
     {loadUnit_maskInput_lo[5791:5776]},
     {loadUnit_maskInput_lo[5775:5760]},
     {loadUnit_maskInput_lo[5759:5744]},
     {loadUnit_maskInput_lo[5743:5728]},
     {loadUnit_maskInput_lo[5727:5712]},
     {loadUnit_maskInput_lo[5711:5696]},
     {loadUnit_maskInput_lo[5695:5680]},
     {loadUnit_maskInput_lo[5679:5664]},
     {loadUnit_maskInput_lo[5663:5648]},
     {loadUnit_maskInput_lo[5647:5632]},
     {loadUnit_maskInput_lo[5631:5616]},
     {loadUnit_maskInput_lo[5615:5600]},
     {loadUnit_maskInput_lo[5599:5584]},
     {loadUnit_maskInput_lo[5583:5568]},
     {loadUnit_maskInput_lo[5567:5552]},
     {loadUnit_maskInput_lo[5551:5536]},
     {loadUnit_maskInput_lo[5535:5520]},
     {loadUnit_maskInput_lo[5519:5504]},
     {loadUnit_maskInput_lo[5503:5488]},
     {loadUnit_maskInput_lo[5487:5472]},
     {loadUnit_maskInput_lo[5471:5456]},
     {loadUnit_maskInput_lo[5455:5440]},
     {loadUnit_maskInput_lo[5439:5424]},
     {loadUnit_maskInput_lo[5423:5408]},
     {loadUnit_maskInput_lo[5407:5392]},
     {loadUnit_maskInput_lo[5391:5376]},
     {loadUnit_maskInput_lo[5375:5360]},
     {loadUnit_maskInput_lo[5359:5344]},
     {loadUnit_maskInput_lo[5343:5328]},
     {loadUnit_maskInput_lo[5327:5312]},
     {loadUnit_maskInput_lo[5311:5296]},
     {loadUnit_maskInput_lo[5295:5280]},
     {loadUnit_maskInput_lo[5279:5264]},
     {loadUnit_maskInput_lo[5263:5248]},
     {loadUnit_maskInput_lo[5247:5232]},
     {loadUnit_maskInput_lo[5231:5216]},
     {loadUnit_maskInput_lo[5215:5200]},
     {loadUnit_maskInput_lo[5199:5184]},
     {loadUnit_maskInput_lo[5183:5168]},
     {loadUnit_maskInput_lo[5167:5152]},
     {loadUnit_maskInput_lo[5151:5136]},
     {loadUnit_maskInput_lo[5135:5120]},
     {loadUnit_maskInput_lo[5119:5104]},
     {loadUnit_maskInput_lo[5103:5088]},
     {loadUnit_maskInput_lo[5087:5072]},
     {loadUnit_maskInput_lo[5071:5056]},
     {loadUnit_maskInput_lo[5055:5040]},
     {loadUnit_maskInput_lo[5039:5024]},
     {loadUnit_maskInput_lo[5023:5008]},
     {loadUnit_maskInput_lo[5007:4992]},
     {loadUnit_maskInput_lo[4991:4976]},
     {loadUnit_maskInput_lo[4975:4960]},
     {loadUnit_maskInput_lo[4959:4944]},
     {loadUnit_maskInput_lo[4943:4928]},
     {loadUnit_maskInput_lo[4927:4912]},
     {loadUnit_maskInput_lo[4911:4896]},
     {loadUnit_maskInput_lo[4895:4880]},
     {loadUnit_maskInput_lo[4879:4864]},
     {loadUnit_maskInput_lo[4863:4848]},
     {loadUnit_maskInput_lo[4847:4832]},
     {loadUnit_maskInput_lo[4831:4816]},
     {loadUnit_maskInput_lo[4815:4800]},
     {loadUnit_maskInput_lo[4799:4784]},
     {loadUnit_maskInput_lo[4783:4768]},
     {loadUnit_maskInput_lo[4767:4752]},
     {loadUnit_maskInput_lo[4751:4736]},
     {loadUnit_maskInput_lo[4735:4720]},
     {loadUnit_maskInput_lo[4719:4704]},
     {loadUnit_maskInput_lo[4703:4688]},
     {loadUnit_maskInput_lo[4687:4672]},
     {loadUnit_maskInput_lo[4671:4656]},
     {loadUnit_maskInput_lo[4655:4640]},
     {loadUnit_maskInput_lo[4639:4624]},
     {loadUnit_maskInput_lo[4623:4608]},
     {loadUnit_maskInput_lo[4607:4592]},
     {loadUnit_maskInput_lo[4591:4576]},
     {loadUnit_maskInput_lo[4575:4560]},
     {loadUnit_maskInput_lo[4559:4544]},
     {loadUnit_maskInput_lo[4543:4528]},
     {loadUnit_maskInput_lo[4527:4512]},
     {loadUnit_maskInput_lo[4511:4496]},
     {loadUnit_maskInput_lo[4495:4480]},
     {loadUnit_maskInput_lo[4479:4464]},
     {loadUnit_maskInput_lo[4463:4448]},
     {loadUnit_maskInput_lo[4447:4432]},
     {loadUnit_maskInput_lo[4431:4416]},
     {loadUnit_maskInput_lo[4415:4400]},
     {loadUnit_maskInput_lo[4399:4384]},
     {loadUnit_maskInput_lo[4383:4368]},
     {loadUnit_maskInput_lo[4367:4352]},
     {loadUnit_maskInput_lo[4351:4336]},
     {loadUnit_maskInput_lo[4335:4320]},
     {loadUnit_maskInput_lo[4319:4304]},
     {loadUnit_maskInput_lo[4303:4288]},
     {loadUnit_maskInput_lo[4287:4272]},
     {loadUnit_maskInput_lo[4271:4256]},
     {loadUnit_maskInput_lo[4255:4240]},
     {loadUnit_maskInput_lo[4239:4224]},
     {loadUnit_maskInput_lo[4223:4208]},
     {loadUnit_maskInput_lo[4207:4192]},
     {loadUnit_maskInput_lo[4191:4176]},
     {loadUnit_maskInput_lo[4175:4160]},
     {loadUnit_maskInput_lo[4159:4144]},
     {loadUnit_maskInput_lo[4143:4128]},
     {loadUnit_maskInput_lo[4127:4112]},
     {loadUnit_maskInput_lo[4111:4096]},
     {loadUnit_maskInput_lo[4095:4080]},
     {loadUnit_maskInput_lo[4079:4064]},
     {loadUnit_maskInput_lo[4063:4048]},
     {loadUnit_maskInput_lo[4047:4032]},
     {loadUnit_maskInput_lo[4031:4016]},
     {loadUnit_maskInput_lo[4015:4000]},
     {loadUnit_maskInput_lo[3999:3984]},
     {loadUnit_maskInput_lo[3983:3968]},
     {loadUnit_maskInput_lo[3967:3952]},
     {loadUnit_maskInput_lo[3951:3936]},
     {loadUnit_maskInput_lo[3935:3920]},
     {loadUnit_maskInput_lo[3919:3904]},
     {loadUnit_maskInput_lo[3903:3888]},
     {loadUnit_maskInput_lo[3887:3872]},
     {loadUnit_maskInput_lo[3871:3856]},
     {loadUnit_maskInput_lo[3855:3840]},
     {loadUnit_maskInput_lo[3839:3824]},
     {loadUnit_maskInput_lo[3823:3808]},
     {loadUnit_maskInput_lo[3807:3792]},
     {loadUnit_maskInput_lo[3791:3776]},
     {loadUnit_maskInput_lo[3775:3760]},
     {loadUnit_maskInput_lo[3759:3744]},
     {loadUnit_maskInput_lo[3743:3728]},
     {loadUnit_maskInput_lo[3727:3712]},
     {loadUnit_maskInput_lo[3711:3696]},
     {loadUnit_maskInput_lo[3695:3680]},
     {loadUnit_maskInput_lo[3679:3664]},
     {loadUnit_maskInput_lo[3663:3648]},
     {loadUnit_maskInput_lo[3647:3632]},
     {loadUnit_maskInput_lo[3631:3616]},
     {loadUnit_maskInput_lo[3615:3600]},
     {loadUnit_maskInput_lo[3599:3584]},
     {loadUnit_maskInput_lo[3583:3568]},
     {loadUnit_maskInput_lo[3567:3552]},
     {loadUnit_maskInput_lo[3551:3536]},
     {loadUnit_maskInput_lo[3535:3520]},
     {loadUnit_maskInput_lo[3519:3504]},
     {loadUnit_maskInput_lo[3503:3488]},
     {loadUnit_maskInput_lo[3487:3472]},
     {loadUnit_maskInput_lo[3471:3456]},
     {loadUnit_maskInput_lo[3455:3440]},
     {loadUnit_maskInput_lo[3439:3424]},
     {loadUnit_maskInput_lo[3423:3408]},
     {loadUnit_maskInput_lo[3407:3392]},
     {loadUnit_maskInput_lo[3391:3376]},
     {loadUnit_maskInput_lo[3375:3360]},
     {loadUnit_maskInput_lo[3359:3344]},
     {loadUnit_maskInput_lo[3343:3328]},
     {loadUnit_maskInput_lo[3327:3312]},
     {loadUnit_maskInput_lo[3311:3296]},
     {loadUnit_maskInput_lo[3295:3280]},
     {loadUnit_maskInput_lo[3279:3264]},
     {loadUnit_maskInput_lo[3263:3248]},
     {loadUnit_maskInput_lo[3247:3232]},
     {loadUnit_maskInput_lo[3231:3216]},
     {loadUnit_maskInput_lo[3215:3200]},
     {loadUnit_maskInput_lo[3199:3184]},
     {loadUnit_maskInput_lo[3183:3168]},
     {loadUnit_maskInput_lo[3167:3152]},
     {loadUnit_maskInput_lo[3151:3136]},
     {loadUnit_maskInput_lo[3135:3120]},
     {loadUnit_maskInput_lo[3119:3104]},
     {loadUnit_maskInput_lo[3103:3088]},
     {loadUnit_maskInput_lo[3087:3072]},
     {loadUnit_maskInput_lo[3071:3056]},
     {loadUnit_maskInput_lo[3055:3040]},
     {loadUnit_maskInput_lo[3039:3024]},
     {loadUnit_maskInput_lo[3023:3008]},
     {loadUnit_maskInput_lo[3007:2992]},
     {loadUnit_maskInput_lo[2991:2976]},
     {loadUnit_maskInput_lo[2975:2960]},
     {loadUnit_maskInput_lo[2959:2944]},
     {loadUnit_maskInput_lo[2943:2928]},
     {loadUnit_maskInput_lo[2927:2912]},
     {loadUnit_maskInput_lo[2911:2896]},
     {loadUnit_maskInput_lo[2895:2880]},
     {loadUnit_maskInput_lo[2879:2864]},
     {loadUnit_maskInput_lo[2863:2848]},
     {loadUnit_maskInput_lo[2847:2832]},
     {loadUnit_maskInput_lo[2831:2816]},
     {loadUnit_maskInput_lo[2815:2800]},
     {loadUnit_maskInput_lo[2799:2784]},
     {loadUnit_maskInput_lo[2783:2768]},
     {loadUnit_maskInput_lo[2767:2752]},
     {loadUnit_maskInput_lo[2751:2736]},
     {loadUnit_maskInput_lo[2735:2720]},
     {loadUnit_maskInput_lo[2719:2704]},
     {loadUnit_maskInput_lo[2703:2688]},
     {loadUnit_maskInput_lo[2687:2672]},
     {loadUnit_maskInput_lo[2671:2656]},
     {loadUnit_maskInput_lo[2655:2640]},
     {loadUnit_maskInput_lo[2639:2624]},
     {loadUnit_maskInput_lo[2623:2608]},
     {loadUnit_maskInput_lo[2607:2592]},
     {loadUnit_maskInput_lo[2591:2576]},
     {loadUnit_maskInput_lo[2575:2560]},
     {loadUnit_maskInput_lo[2559:2544]},
     {loadUnit_maskInput_lo[2543:2528]},
     {loadUnit_maskInput_lo[2527:2512]},
     {loadUnit_maskInput_lo[2511:2496]},
     {loadUnit_maskInput_lo[2495:2480]},
     {loadUnit_maskInput_lo[2479:2464]},
     {loadUnit_maskInput_lo[2463:2448]},
     {loadUnit_maskInput_lo[2447:2432]},
     {loadUnit_maskInput_lo[2431:2416]},
     {loadUnit_maskInput_lo[2415:2400]},
     {loadUnit_maskInput_lo[2399:2384]},
     {loadUnit_maskInput_lo[2383:2368]},
     {loadUnit_maskInput_lo[2367:2352]},
     {loadUnit_maskInput_lo[2351:2336]},
     {loadUnit_maskInput_lo[2335:2320]},
     {loadUnit_maskInput_lo[2319:2304]},
     {loadUnit_maskInput_lo[2303:2288]},
     {loadUnit_maskInput_lo[2287:2272]},
     {loadUnit_maskInput_lo[2271:2256]},
     {loadUnit_maskInput_lo[2255:2240]},
     {loadUnit_maskInput_lo[2239:2224]},
     {loadUnit_maskInput_lo[2223:2208]},
     {loadUnit_maskInput_lo[2207:2192]},
     {loadUnit_maskInput_lo[2191:2176]},
     {loadUnit_maskInput_lo[2175:2160]},
     {loadUnit_maskInput_lo[2159:2144]},
     {loadUnit_maskInput_lo[2143:2128]},
     {loadUnit_maskInput_lo[2127:2112]},
     {loadUnit_maskInput_lo[2111:2096]},
     {loadUnit_maskInput_lo[2095:2080]},
     {loadUnit_maskInput_lo[2079:2064]},
     {loadUnit_maskInput_lo[2063:2048]},
     {loadUnit_maskInput_lo[2047:2032]},
     {loadUnit_maskInput_lo[2031:2016]},
     {loadUnit_maskInput_lo[2015:2000]},
     {loadUnit_maskInput_lo[1999:1984]},
     {loadUnit_maskInput_lo[1983:1968]},
     {loadUnit_maskInput_lo[1967:1952]},
     {loadUnit_maskInput_lo[1951:1936]},
     {loadUnit_maskInput_lo[1935:1920]},
     {loadUnit_maskInput_lo[1919:1904]},
     {loadUnit_maskInput_lo[1903:1888]},
     {loadUnit_maskInput_lo[1887:1872]},
     {loadUnit_maskInput_lo[1871:1856]},
     {loadUnit_maskInput_lo[1855:1840]},
     {loadUnit_maskInput_lo[1839:1824]},
     {loadUnit_maskInput_lo[1823:1808]},
     {loadUnit_maskInput_lo[1807:1792]},
     {loadUnit_maskInput_lo[1791:1776]},
     {loadUnit_maskInput_lo[1775:1760]},
     {loadUnit_maskInput_lo[1759:1744]},
     {loadUnit_maskInput_lo[1743:1728]},
     {loadUnit_maskInput_lo[1727:1712]},
     {loadUnit_maskInput_lo[1711:1696]},
     {loadUnit_maskInput_lo[1695:1680]},
     {loadUnit_maskInput_lo[1679:1664]},
     {loadUnit_maskInput_lo[1663:1648]},
     {loadUnit_maskInput_lo[1647:1632]},
     {loadUnit_maskInput_lo[1631:1616]},
     {loadUnit_maskInput_lo[1615:1600]},
     {loadUnit_maskInput_lo[1599:1584]},
     {loadUnit_maskInput_lo[1583:1568]},
     {loadUnit_maskInput_lo[1567:1552]},
     {loadUnit_maskInput_lo[1551:1536]},
     {loadUnit_maskInput_lo[1535:1520]},
     {loadUnit_maskInput_lo[1519:1504]},
     {loadUnit_maskInput_lo[1503:1488]},
     {loadUnit_maskInput_lo[1487:1472]},
     {loadUnit_maskInput_lo[1471:1456]},
     {loadUnit_maskInput_lo[1455:1440]},
     {loadUnit_maskInput_lo[1439:1424]},
     {loadUnit_maskInput_lo[1423:1408]},
     {loadUnit_maskInput_lo[1407:1392]},
     {loadUnit_maskInput_lo[1391:1376]},
     {loadUnit_maskInput_lo[1375:1360]},
     {loadUnit_maskInput_lo[1359:1344]},
     {loadUnit_maskInput_lo[1343:1328]},
     {loadUnit_maskInput_lo[1327:1312]},
     {loadUnit_maskInput_lo[1311:1296]},
     {loadUnit_maskInput_lo[1295:1280]},
     {loadUnit_maskInput_lo[1279:1264]},
     {loadUnit_maskInput_lo[1263:1248]},
     {loadUnit_maskInput_lo[1247:1232]},
     {loadUnit_maskInput_lo[1231:1216]},
     {loadUnit_maskInput_lo[1215:1200]},
     {loadUnit_maskInput_lo[1199:1184]},
     {loadUnit_maskInput_lo[1183:1168]},
     {loadUnit_maskInput_lo[1167:1152]},
     {loadUnit_maskInput_lo[1151:1136]},
     {loadUnit_maskInput_lo[1135:1120]},
     {loadUnit_maskInput_lo[1119:1104]},
     {loadUnit_maskInput_lo[1103:1088]},
     {loadUnit_maskInput_lo[1087:1072]},
     {loadUnit_maskInput_lo[1071:1056]},
     {loadUnit_maskInput_lo[1055:1040]},
     {loadUnit_maskInput_lo[1039:1024]},
     {loadUnit_maskInput_lo[1023:1008]},
     {loadUnit_maskInput_lo[1007:992]},
     {loadUnit_maskInput_lo[991:976]},
     {loadUnit_maskInput_lo[975:960]},
     {loadUnit_maskInput_lo[959:944]},
     {loadUnit_maskInput_lo[943:928]},
     {loadUnit_maskInput_lo[927:912]},
     {loadUnit_maskInput_lo[911:896]},
     {loadUnit_maskInput_lo[895:880]},
     {loadUnit_maskInput_lo[879:864]},
     {loadUnit_maskInput_lo[863:848]},
     {loadUnit_maskInput_lo[847:832]},
     {loadUnit_maskInput_lo[831:816]},
     {loadUnit_maskInput_lo[815:800]},
     {loadUnit_maskInput_lo[799:784]},
     {loadUnit_maskInput_lo[783:768]},
     {loadUnit_maskInput_lo[767:752]},
     {loadUnit_maskInput_lo[751:736]},
     {loadUnit_maskInput_lo[735:720]},
     {loadUnit_maskInput_lo[719:704]},
     {loadUnit_maskInput_lo[703:688]},
     {loadUnit_maskInput_lo[687:672]},
     {loadUnit_maskInput_lo[671:656]},
     {loadUnit_maskInput_lo[655:640]},
     {loadUnit_maskInput_lo[639:624]},
     {loadUnit_maskInput_lo[623:608]},
     {loadUnit_maskInput_lo[607:592]},
     {loadUnit_maskInput_lo[591:576]},
     {loadUnit_maskInput_lo[575:560]},
     {loadUnit_maskInput_lo[559:544]},
     {loadUnit_maskInput_lo[543:528]},
     {loadUnit_maskInput_lo[527:512]},
     {loadUnit_maskInput_lo[511:496]},
     {loadUnit_maskInput_lo[495:480]},
     {loadUnit_maskInput_lo[479:464]},
     {loadUnit_maskInput_lo[463:448]},
     {loadUnit_maskInput_lo[447:432]},
     {loadUnit_maskInput_lo[431:416]},
     {loadUnit_maskInput_lo[415:400]},
     {loadUnit_maskInput_lo[399:384]},
     {loadUnit_maskInput_lo[383:368]},
     {loadUnit_maskInput_lo[367:352]},
     {loadUnit_maskInput_lo[351:336]},
     {loadUnit_maskInput_lo[335:320]},
     {loadUnit_maskInput_lo[319:304]},
     {loadUnit_maskInput_lo[303:288]},
     {loadUnit_maskInput_lo[287:272]},
     {loadUnit_maskInput_lo[271:256]},
     {loadUnit_maskInput_lo[255:240]},
     {loadUnit_maskInput_lo[239:224]},
     {loadUnit_maskInput_lo[223:208]},
     {loadUnit_maskInput_lo[207:192]},
     {loadUnit_maskInput_lo[191:176]},
     {loadUnit_maskInput_lo[175:160]},
     {loadUnit_maskInput_lo[159:144]},
     {loadUnit_maskInput_lo[143:128]},
     {loadUnit_maskInput_lo[127:112]},
     {loadUnit_maskInput_lo[111:96]},
     {loadUnit_maskInput_lo[95:80]},
     {loadUnit_maskInput_lo[79:64]},
     {loadUnit_maskInput_lo[63:48]},
     {loadUnit_maskInput_lo[47:32]},
     {loadUnit_maskInput_lo[31:16]},
     {loadUnit_maskInput_lo[15:0]}};
  wire [10:0]         maskSelect_1 = _storeUnit_maskSelect_valid ? _storeUnit_maskSelect_bits : 11'h0;
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_lo_lo = {storeUnit_maskInput_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_lo_hi_hi = {storeUnit_maskInput_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_lo_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_lo_hi = {storeUnit_maskInput_lo_lo_hi_hi, storeUnit_maskInput_lo_lo_hi_lo};
  wire [8191:0]       storeUnit_maskInput_lo_lo = {storeUnit_maskInput_lo_lo_hi, storeUnit_maskInput_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_hi_lo = {storeUnit_maskInput_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_lo_hi_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_lo_hi_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_lo_hi_hi = {storeUnit_maskInput_lo_hi_hi_hi, storeUnit_maskInput_lo_hi_hi_lo};
  wire [8191:0]       storeUnit_maskInput_lo_hi = {storeUnit_maskInput_lo_hi_hi, storeUnit_maskInput_lo_hi_lo};
  wire [16383:0]      storeUnit_maskInput_lo = {storeUnit_maskInput_lo_hi, storeUnit_maskInput_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_lo_lo = {storeUnit_maskInput_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_lo_hi_hi = {storeUnit_maskInput_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_lo_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_lo_hi = {storeUnit_maskInput_hi_lo_hi_hi, storeUnit_maskInput_hi_lo_hi_lo};
  wire [8191:0]       storeUnit_maskInput_hi_lo = {storeUnit_maskInput_hi_lo_hi, storeUnit_maskInput_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_lo_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_hi_lo = {storeUnit_maskInput_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        storeUnit_maskInput_hi_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       storeUnit_maskInput_hi_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       storeUnit_maskInput_hi_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_hi_lo};
  wire [4095:0]       storeUnit_maskInput_hi_hi_hi = {storeUnit_maskInput_hi_hi_hi_hi, storeUnit_maskInput_hi_hi_hi_lo};
  wire [8191:0]       storeUnit_maskInput_hi_hi = {storeUnit_maskInput_hi_hi_hi, storeUnit_maskInput_hi_hi_lo};
  wire [16383:0]      storeUnit_maskInput_hi = {storeUnit_maskInput_hi_hi, storeUnit_maskInput_hi_lo};
  wire [2047:0][15:0] _GEN_512 =
    {{storeUnit_maskInput_hi[16383:16368]},
     {storeUnit_maskInput_hi[16367:16352]},
     {storeUnit_maskInput_hi[16351:16336]},
     {storeUnit_maskInput_hi[16335:16320]},
     {storeUnit_maskInput_hi[16319:16304]},
     {storeUnit_maskInput_hi[16303:16288]},
     {storeUnit_maskInput_hi[16287:16272]},
     {storeUnit_maskInput_hi[16271:16256]},
     {storeUnit_maskInput_hi[16255:16240]},
     {storeUnit_maskInput_hi[16239:16224]},
     {storeUnit_maskInput_hi[16223:16208]},
     {storeUnit_maskInput_hi[16207:16192]},
     {storeUnit_maskInput_hi[16191:16176]},
     {storeUnit_maskInput_hi[16175:16160]},
     {storeUnit_maskInput_hi[16159:16144]},
     {storeUnit_maskInput_hi[16143:16128]},
     {storeUnit_maskInput_hi[16127:16112]},
     {storeUnit_maskInput_hi[16111:16096]},
     {storeUnit_maskInput_hi[16095:16080]},
     {storeUnit_maskInput_hi[16079:16064]},
     {storeUnit_maskInput_hi[16063:16048]},
     {storeUnit_maskInput_hi[16047:16032]},
     {storeUnit_maskInput_hi[16031:16016]},
     {storeUnit_maskInput_hi[16015:16000]},
     {storeUnit_maskInput_hi[15999:15984]},
     {storeUnit_maskInput_hi[15983:15968]},
     {storeUnit_maskInput_hi[15967:15952]},
     {storeUnit_maskInput_hi[15951:15936]},
     {storeUnit_maskInput_hi[15935:15920]},
     {storeUnit_maskInput_hi[15919:15904]},
     {storeUnit_maskInput_hi[15903:15888]},
     {storeUnit_maskInput_hi[15887:15872]},
     {storeUnit_maskInput_hi[15871:15856]},
     {storeUnit_maskInput_hi[15855:15840]},
     {storeUnit_maskInput_hi[15839:15824]},
     {storeUnit_maskInput_hi[15823:15808]},
     {storeUnit_maskInput_hi[15807:15792]},
     {storeUnit_maskInput_hi[15791:15776]},
     {storeUnit_maskInput_hi[15775:15760]},
     {storeUnit_maskInput_hi[15759:15744]},
     {storeUnit_maskInput_hi[15743:15728]},
     {storeUnit_maskInput_hi[15727:15712]},
     {storeUnit_maskInput_hi[15711:15696]},
     {storeUnit_maskInput_hi[15695:15680]},
     {storeUnit_maskInput_hi[15679:15664]},
     {storeUnit_maskInput_hi[15663:15648]},
     {storeUnit_maskInput_hi[15647:15632]},
     {storeUnit_maskInput_hi[15631:15616]},
     {storeUnit_maskInput_hi[15615:15600]},
     {storeUnit_maskInput_hi[15599:15584]},
     {storeUnit_maskInput_hi[15583:15568]},
     {storeUnit_maskInput_hi[15567:15552]},
     {storeUnit_maskInput_hi[15551:15536]},
     {storeUnit_maskInput_hi[15535:15520]},
     {storeUnit_maskInput_hi[15519:15504]},
     {storeUnit_maskInput_hi[15503:15488]},
     {storeUnit_maskInput_hi[15487:15472]},
     {storeUnit_maskInput_hi[15471:15456]},
     {storeUnit_maskInput_hi[15455:15440]},
     {storeUnit_maskInput_hi[15439:15424]},
     {storeUnit_maskInput_hi[15423:15408]},
     {storeUnit_maskInput_hi[15407:15392]},
     {storeUnit_maskInput_hi[15391:15376]},
     {storeUnit_maskInput_hi[15375:15360]},
     {storeUnit_maskInput_hi[15359:15344]},
     {storeUnit_maskInput_hi[15343:15328]},
     {storeUnit_maskInput_hi[15327:15312]},
     {storeUnit_maskInput_hi[15311:15296]},
     {storeUnit_maskInput_hi[15295:15280]},
     {storeUnit_maskInput_hi[15279:15264]},
     {storeUnit_maskInput_hi[15263:15248]},
     {storeUnit_maskInput_hi[15247:15232]},
     {storeUnit_maskInput_hi[15231:15216]},
     {storeUnit_maskInput_hi[15215:15200]},
     {storeUnit_maskInput_hi[15199:15184]},
     {storeUnit_maskInput_hi[15183:15168]},
     {storeUnit_maskInput_hi[15167:15152]},
     {storeUnit_maskInput_hi[15151:15136]},
     {storeUnit_maskInput_hi[15135:15120]},
     {storeUnit_maskInput_hi[15119:15104]},
     {storeUnit_maskInput_hi[15103:15088]},
     {storeUnit_maskInput_hi[15087:15072]},
     {storeUnit_maskInput_hi[15071:15056]},
     {storeUnit_maskInput_hi[15055:15040]},
     {storeUnit_maskInput_hi[15039:15024]},
     {storeUnit_maskInput_hi[15023:15008]},
     {storeUnit_maskInput_hi[15007:14992]},
     {storeUnit_maskInput_hi[14991:14976]},
     {storeUnit_maskInput_hi[14975:14960]},
     {storeUnit_maskInput_hi[14959:14944]},
     {storeUnit_maskInput_hi[14943:14928]},
     {storeUnit_maskInput_hi[14927:14912]},
     {storeUnit_maskInput_hi[14911:14896]},
     {storeUnit_maskInput_hi[14895:14880]},
     {storeUnit_maskInput_hi[14879:14864]},
     {storeUnit_maskInput_hi[14863:14848]},
     {storeUnit_maskInput_hi[14847:14832]},
     {storeUnit_maskInput_hi[14831:14816]},
     {storeUnit_maskInput_hi[14815:14800]},
     {storeUnit_maskInput_hi[14799:14784]},
     {storeUnit_maskInput_hi[14783:14768]},
     {storeUnit_maskInput_hi[14767:14752]},
     {storeUnit_maskInput_hi[14751:14736]},
     {storeUnit_maskInput_hi[14735:14720]},
     {storeUnit_maskInput_hi[14719:14704]},
     {storeUnit_maskInput_hi[14703:14688]},
     {storeUnit_maskInput_hi[14687:14672]},
     {storeUnit_maskInput_hi[14671:14656]},
     {storeUnit_maskInput_hi[14655:14640]},
     {storeUnit_maskInput_hi[14639:14624]},
     {storeUnit_maskInput_hi[14623:14608]},
     {storeUnit_maskInput_hi[14607:14592]},
     {storeUnit_maskInput_hi[14591:14576]},
     {storeUnit_maskInput_hi[14575:14560]},
     {storeUnit_maskInput_hi[14559:14544]},
     {storeUnit_maskInput_hi[14543:14528]},
     {storeUnit_maskInput_hi[14527:14512]},
     {storeUnit_maskInput_hi[14511:14496]},
     {storeUnit_maskInput_hi[14495:14480]},
     {storeUnit_maskInput_hi[14479:14464]},
     {storeUnit_maskInput_hi[14463:14448]},
     {storeUnit_maskInput_hi[14447:14432]},
     {storeUnit_maskInput_hi[14431:14416]},
     {storeUnit_maskInput_hi[14415:14400]},
     {storeUnit_maskInput_hi[14399:14384]},
     {storeUnit_maskInput_hi[14383:14368]},
     {storeUnit_maskInput_hi[14367:14352]},
     {storeUnit_maskInput_hi[14351:14336]},
     {storeUnit_maskInput_hi[14335:14320]},
     {storeUnit_maskInput_hi[14319:14304]},
     {storeUnit_maskInput_hi[14303:14288]},
     {storeUnit_maskInput_hi[14287:14272]},
     {storeUnit_maskInput_hi[14271:14256]},
     {storeUnit_maskInput_hi[14255:14240]},
     {storeUnit_maskInput_hi[14239:14224]},
     {storeUnit_maskInput_hi[14223:14208]},
     {storeUnit_maskInput_hi[14207:14192]},
     {storeUnit_maskInput_hi[14191:14176]},
     {storeUnit_maskInput_hi[14175:14160]},
     {storeUnit_maskInput_hi[14159:14144]},
     {storeUnit_maskInput_hi[14143:14128]},
     {storeUnit_maskInput_hi[14127:14112]},
     {storeUnit_maskInput_hi[14111:14096]},
     {storeUnit_maskInput_hi[14095:14080]},
     {storeUnit_maskInput_hi[14079:14064]},
     {storeUnit_maskInput_hi[14063:14048]},
     {storeUnit_maskInput_hi[14047:14032]},
     {storeUnit_maskInput_hi[14031:14016]},
     {storeUnit_maskInput_hi[14015:14000]},
     {storeUnit_maskInput_hi[13999:13984]},
     {storeUnit_maskInput_hi[13983:13968]},
     {storeUnit_maskInput_hi[13967:13952]},
     {storeUnit_maskInput_hi[13951:13936]},
     {storeUnit_maskInput_hi[13935:13920]},
     {storeUnit_maskInput_hi[13919:13904]},
     {storeUnit_maskInput_hi[13903:13888]},
     {storeUnit_maskInput_hi[13887:13872]},
     {storeUnit_maskInput_hi[13871:13856]},
     {storeUnit_maskInput_hi[13855:13840]},
     {storeUnit_maskInput_hi[13839:13824]},
     {storeUnit_maskInput_hi[13823:13808]},
     {storeUnit_maskInput_hi[13807:13792]},
     {storeUnit_maskInput_hi[13791:13776]},
     {storeUnit_maskInput_hi[13775:13760]},
     {storeUnit_maskInput_hi[13759:13744]},
     {storeUnit_maskInput_hi[13743:13728]},
     {storeUnit_maskInput_hi[13727:13712]},
     {storeUnit_maskInput_hi[13711:13696]},
     {storeUnit_maskInput_hi[13695:13680]},
     {storeUnit_maskInput_hi[13679:13664]},
     {storeUnit_maskInput_hi[13663:13648]},
     {storeUnit_maskInput_hi[13647:13632]},
     {storeUnit_maskInput_hi[13631:13616]},
     {storeUnit_maskInput_hi[13615:13600]},
     {storeUnit_maskInput_hi[13599:13584]},
     {storeUnit_maskInput_hi[13583:13568]},
     {storeUnit_maskInput_hi[13567:13552]},
     {storeUnit_maskInput_hi[13551:13536]},
     {storeUnit_maskInput_hi[13535:13520]},
     {storeUnit_maskInput_hi[13519:13504]},
     {storeUnit_maskInput_hi[13503:13488]},
     {storeUnit_maskInput_hi[13487:13472]},
     {storeUnit_maskInput_hi[13471:13456]},
     {storeUnit_maskInput_hi[13455:13440]},
     {storeUnit_maskInput_hi[13439:13424]},
     {storeUnit_maskInput_hi[13423:13408]},
     {storeUnit_maskInput_hi[13407:13392]},
     {storeUnit_maskInput_hi[13391:13376]},
     {storeUnit_maskInput_hi[13375:13360]},
     {storeUnit_maskInput_hi[13359:13344]},
     {storeUnit_maskInput_hi[13343:13328]},
     {storeUnit_maskInput_hi[13327:13312]},
     {storeUnit_maskInput_hi[13311:13296]},
     {storeUnit_maskInput_hi[13295:13280]},
     {storeUnit_maskInput_hi[13279:13264]},
     {storeUnit_maskInput_hi[13263:13248]},
     {storeUnit_maskInput_hi[13247:13232]},
     {storeUnit_maskInput_hi[13231:13216]},
     {storeUnit_maskInput_hi[13215:13200]},
     {storeUnit_maskInput_hi[13199:13184]},
     {storeUnit_maskInput_hi[13183:13168]},
     {storeUnit_maskInput_hi[13167:13152]},
     {storeUnit_maskInput_hi[13151:13136]},
     {storeUnit_maskInput_hi[13135:13120]},
     {storeUnit_maskInput_hi[13119:13104]},
     {storeUnit_maskInput_hi[13103:13088]},
     {storeUnit_maskInput_hi[13087:13072]},
     {storeUnit_maskInput_hi[13071:13056]},
     {storeUnit_maskInput_hi[13055:13040]},
     {storeUnit_maskInput_hi[13039:13024]},
     {storeUnit_maskInput_hi[13023:13008]},
     {storeUnit_maskInput_hi[13007:12992]},
     {storeUnit_maskInput_hi[12991:12976]},
     {storeUnit_maskInput_hi[12975:12960]},
     {storeUnit_maskInput_hi[12959:12944]},
     {storeUnit_maskInput_hi[12943:12928]},
     {storeUnit_maskInput_hi[12927:12912]},
     {storeUnit_maskInput_hi[12911:12896]},
     {storeUnit_maskInput_hi[12895:12880]},
     {storeUnit_maskInput_hi[12879:12864]},
     {storeUnit_maskInput_hi[12863:12848]},
     {storeUnit_maskInput_hi[12847:12832]},
     {storeUnit_maskInput_hi[12831:12816]},
     {storeUnit_maskInput_hi[12815:12800]},
     {storeUnit_maskInput_hi[12799:12784]},
     {storeUnit_maskInput_hi[12783:12768]},
     {storeUnit_maskInput_hi[12767:12752]},
     {storeUnit_maskInput_hi[12751:12736]},
     {storeUnit_maskInput_hi[12735:12720]},
     {storeUnit_maskInput_hi[12719:12704]},
     {storeUnit_maskInput_hi[12703:12688]},
     {storeUnit_maskInput_hi[12687:12672]},
     {storeUnit_maskInput_hi[12671:12656]},
     {storeUnit_maskInput_hi[12655:12640]},
     {storeUnit_maskInput_hi[12639:12624]},
     {storeUnit_maskInput_hi[12623:12608]},
     {storeUnit_maskInput_hi[12607:12592]},
     {storeUnit_maskInput_hi[12591:12576]},
     {storeUnit_maskInput_hi[12575:12560]},
     {storeUnit_maskInput_hi[12559:12544]},
     {storeUnit_maskInput_hi[12543:12528]},
     {storeUnit_maskInput_hi[12527:12512]},
     {storeUnit_maskInput_hi[12511:12496]},
     {storeUnit_maskInput_hi[12495:12480]},
     {storeUnit_maskInput_hi[12479:12464]},
     {storeUnit_maskInput_hi[12463:12448]},
     {storeUnit_maskInput_hi[12447:12432]},
     {storeUnit_maskInput_hi[12431:12416]},
     {storeUnit_maskInput_hi[12415:12400]},
     {storeUnit_maskInput_hi[12399:12384]},
     {storeUnit_maskInput_hi[12383:12368]},
     {storeUnit_maskInput_hi[12367:12352]},
     {storeUnit_maskInput_hi[12351:12336]},
     {storeUnit_maskInput_hi[12335:12320]},
     {storeUnit_maskInput_hi[12319:12304]},
     {storeUnit_maskInput_hi[12303:12288]},
     {storeUnit_maskInput_hi[12287:12272]},
     {storeUnit_maskInput_hi[12271:12256]},
     {storeUnit_maskInput_hi[12255:12240]},
     {storeUnit_maskInput_hi[12239:12224]},
     {storeUnit_maskInput_hi[12223:12208]},
     {storeUnit_maskInput_hi[12207:12192]},
     {storeUnit_maskInput_hi[12191:12176]},
     {storeUnit_maskInput_hi[12175:12160]},
     {storeUnit_maskInput_hi[12159:12144]},
     {storeUnit_maskInput_hi[12143:12128]},
     {storeUnit_maskInput_hi[12127:12112]},
     {storeUnit_maskInput_hi[12111:12096]},
     {storeUnit_maskInput_hi[12095:12080]},
     {storeUnit_maskInput_hi[12079:12064]},
     {storeUnit_maskInput_hi[12063:12048]},
     {storeUnit_maskInput_hi[12047:12032]},
     {storeUnit_maskInput_hi[12031:12016]},
     {storeUnit_maskInput_hi[12015:12000]},
     {storeUnit_maskInput_hi[11999:11984]},
     {storeUnit_maskInput_hi[11983:11968]},
     {storeUnit_maskInput_hi[11967:11952]},
     {storeUnit_maskInput_hi[11951:11936]},
     {storeUnit_maskInput_hi[11935:11920]},
     {storeUnit_maskInput_hi[11919:11904]},
     {storeUnit_maskInput_hi[11903:11888]},
     {storeUnit_maskInput_hi[11887:11872]},
     {storeUnit_maskInput_hi[11871:11856]},
     {storeUnit_maskInput_hi[11855:11840]},
     {storeUnit_maskInput_hi[11839:11824]},
     {storeUnit_maskInput_hi[11823:11808]},
     {storeUnit_maskInput_hi[11807:11792]},
     {storeUnit_maskInput_hi[11791:11776]},
     {storeUnit_maskInput_hi[11775:11760]},
     {storeUnit_maskInput_hi[11759:11744]},
     {storeUnit_maskInput_hi[11743:11728]},
     {storeUnit_maskInput_hi[11727:11712]},
     {storeUnit_maskInput_hi[11711:11696]},
     {storeUnit_maskInput_hi[11695:11680]},
     {storeUnit_maskInput_hi[11679:11664]},
     {storeUnit_maskInput_hi[11663:11648]},
     {storeUnit_maskInput_hi[11647:11632]},
     {storeUnit_maskInput_hi[11631:11616]},
     {storeUnit_maskInput_hi[11615:11600]},
     {storeUnit_maskInput_hi[11599:11584]},
     {storeUnit_maskInput_hi[11583:11568]},
     {storeUnit_maskInput_hi[11567:11552]},
     {storeUnit_maskInput_hi[11551:11536]},
     {storeUnit_maskInput_hi[11535:11520]},
     {storeUnit_maskInput_hi[11519:11504]},
     {storeUnit_maskInput_hi[11503:11488]},
     {storeUnit_maskInput_hi[11487:11472]},
     {storeUnit_maskInput_hi[11471:11456]},
     {storeUnit_maskInput_hi[11455:11440]},
     {storeUnit_maskInput_hi[11439:11424]},
     {storeUnit_maskInput_hi[11423:11408]},
     {storeUnit_maskInput_hi[11407:11392]},
     {storeUnit_maskInput_hi[11391:11376]},
     {storeUnit_maskInput_hi[11375:11360]},
     {storeUnit_maskInput_hi[11359:11344]},
     {storeUnit_maskInput_hi[11343:11328]},
     {storeUnit_maskInput_hi[11327:11312]},
     {storeUnit_maskInput_hi[11311:11296]},
     {storeUnit_maskInput_hi[11295:11280]},
     {storeUnit_maskInput_hi[11279:11264]},
     {storeUnit_maskInput_hi[11263:11248]},
     {storeUnit_maskInput_hi[11247:11232]},
     {storeUnit_maskInput_hi[11231:11216]},
     {storeUnit_maskInput_hi[11215:11200]},
     {storeUnit_maskInput_hi[11199:11184]},
     {storeUnit_maskInput_hi[11183:11168]},
     {storeUnit_maskInput_hi[11167:11152]},
     {storeUnit_maskInput_hi[11151:11136]},
     {storeUnit_maskInput_hi[11135:11120]},
     {storeUnit_maskInput_hi[11119:11104]},
     {storeUnit_maskInput_hi[11103:11088]},
     {storeUnit_maskInput_hi[11087:11072]},
     {storeUnit_maskInput_hi[11071:11056]},
     {storeUnit_maskInput_hi[11055:11040]},
     {storeUnit_maskInput_hi[11039:11024]},
     {storeUnit_maskInput_hi[11023:11008]},
     {storeUnit_maskInput_hi[11007:10992]},
     {storeUnit_maskInput_hi[10991:10976]},
     {storeUnit_maskInput_hi[10975:10960]},
     {storeUnit_maskInput_hi[10959:10944]},
     {storeUnit_maskInput_hi[10943:10928]},
     {storeUnit_maskInput_hi[10927:10912]},
     {storeUnit_maskInput_hi[10911:10896]},
     {storeUnit_maskInput_hi[10895:10880]},
     {storeUnit_maskInput_hi[10879:10864]},
     {storeUnit_maskInput_hi[10863:10848]},
     {storeUnit_maskInput_hi[10847:10832]},
     {storeUnit_maskInput_hi[10831:10816]},
     {storeUnit_maskInput_hi[10815:10800]},
     {storeUnit_maskInput_hi[10799:10784]},
     {storeUnit_maskInput_hi[10783:10768]},
     {storeUnit_maskInput_hi[10767:10752]},
     {storeUnit_maskInput_hi[10751:10736]},
     {storeUnit_maskInput_hi[10735:10720]},
     {storeUnit_maskInput_hi[10719:10704]},
     {storeUnit_maskInput_hi[10703:10688]},
     {storeUnit_maskInput_hi[10687:10672]},
     {storeUnit_maskInput_hi[10671:10656]},
     {storeUnit_maskInput_hi[10655:10640]},
     {storeUnit_maskInput_hi[10639:10624]},
     {storeUnit_maskInput_hi[10623:10608]},
     {storeUnit_maskInput_hi[10607:10592]},
     {storeUnit_maskInput_hi[10591:10576]},
     {storeUnit_maskInput_hi[10575:10560]},
     {storeUnit_maskInput_hi[10559:10544]},
     {storeUnit_maskInput_hi[10543:10528]},
     {storeUnit_maskInput_hi[10527:10512]},
     {storeUnit_maskInput_hi[10511:10496]},
     {storeUnit_maskInput_hi[10495:10480]},
     {storeUnit_maskInput_hi[10479:10464]},
     {storeUnit_maskInput_hi[10463:10448]},
     {storeUnit_maskInput_hi[10447:10432]},
     {storeUnit_maskInput_hi[10431:10416]},
     {storeUnit_maskInput_hi[10415:10400]},
     {storeUnit_maskInput_hi[10399:10384]},
     {storeUnit_maskInput_hi[10383:10368]},
     {storeUnit_maskInput_hi[10367:10352]},
     {storeUnit_maskInput_hi[10351:10336]},
     {storeUnit_maskInput_hi[10335:10320]},
     {storeUnit_maskInput_hi[10319:10304]},
     {storeUnit_maskInput_hi[10303:10288]},
     {storeUnit_maskInput_hi[10287:10272]},
     {storeUnit_maskInput_hi[10271:10256]},
     {storeUnit_maskInput_hi[10255:10240]},
     {storeUnit_maskInput_hi[10239:10224]},
     {storeUnit_maskInput_hi[10223:10208]},
     {storeUnit_maskInput_hi[10207:10192]},
     {storeUnit_maskInput_hi[10191:10176]},
     {storeUnit_maskInput_hi[10175:10160]},
     {storeUnit_maskInput_hi[10159:10144]},
     {storeUnit_maskInput_hi[10143:10128]},
     {storeUnit_maskInput_hi[10127:10112]},
     {storeUnit_maskInput_hi[10111:10096]},
     {storeUnit_maskInput_hi[10095:10080]},
     {storeUnit_maskInput_hi[10079:10064]},
     {storeUnit_maskInput_hi[10063:10048]},
     {storeUnit_maskInput_hi[10047:10032]},
     {storeUnit_maskInput_hi[10031:10016]},
     {storeUnit_maskInput_hi[10015:10000]},
     {storeUnit_maskInput_hi[9999:9984]},
     {storeUnit_maskInput_hi[9983:9968]},
     {storeUnit_maskInput_hi[9967:9952]},
     {storeUnit_maskInput_hi[9951:9936]},
     {storeUnit_maskInput_hi[9935:9920]},
     {storeUnit_maskInput_hi[9919:9904]},
     {storeUnit_maskInput_hi[9903:9888]},
     {storeUnit_maskInput_hi[9887:9872]},
     {storeUnit_maskInput_hi[9871:9856]},
     {storeUnit_maskInput_hi[9855:9840]},
     {storeUnit_maskInput_hi[9839:9824]},
     {storeUnit_maskInput_hi[9823:9808]},
     {storeUnit_maskInput_hi[9807:9792]},
     {storeUnit_maskInput_hi[9791:9776]},
     {storeUnit_maskInput_hi[9775:9760]},
     {storeUnit_maskInput_hi[9759:9744]},
     {storeUnit_maskInput_hi[9743:9728]},
     {storeUnit_maskInput_hi[9727:9712]},
     {storeUnit_maskInput_hi[9711:9696]},
     {storeUnit_maskInput_hi[9695:9680]},
     {storeUnit_maskInput_hi[9679:9664]},
     {storeUnit_maskInput_hi[9663:9648]},
     {storeUnit_maskInput_hi[9647:9632]},
     {storeUnit_maskInput_hi[9631:9616]},
     {storeUnit_maskInput_hi[9615:9600]},
     {storeUnit_maskInput_hi[9599:9584]},
     {storeUnit_maskInput_hi[9583:9568]},
     {storeUnit_maskInput_hi[9567:9552]},
     {storeUnit_maskInput_hi[9551:9536]},
     {storeUnit_maskInput_hi[9535:9520]},
     {storeUnit_maskInput_hi[9519:9504]},
     {storeUnit_maskInput_hi[9503:9488]},
     {storeUnit_maskInput_hi[9487:9472]},
     {storeUnit_maskInput_hi[9471:9456]},
     {storeUnit_maskInput_hi[9455:9440]},
     {storeUnit_maskInput_hi[9439:9424]},
     {storeUnit_maskInput_hi[9423:9408]},
     {storeUnit_maskInput_hi[9407:9392]},
     {storeUnit_maskInput_hi[9391:9376]},
     {storeUnit_maskInput_hi[9375:9360]},
     {storeUnit_maskInput_hi[9359:9344]},
     {storeUnit_maskInput_hi[9343:9328]},
     {storeUnit_maskInput_hi[9327:9312]},
     {storeUnit_maskInput_hi[9311:9296]},
     {storeUnit_maskInput_hi[9295:9280]},
     {storeUnit_maskInput_hi[9279:9264]},
     {storeUnit_maskInput_hi[9263:9248]},
     {storeUnit_maskInput_hi[9247:9232]},
     {storeUnit_maskInput_hi[9231:9216]},
     {storeUnit_maskInput_hi[9215:9200]},
     {storeUnit_maskInput_hi[9199:9184]},
     {storeUnit_maskInput_hi[9183:9168]},
     {storeUnit_maskInput_hi[9167:9152]},
     {storeUnit_maskInput_hi[9151:9136]},
     {storeUnit_maskInput_hi[9135:9120]},
     {storeUnit_maskInput_hi[9119:9104]},
     {storeUnit_maskInput_hi[9103:9088]},
     {storeUnit_maskInput_hi[9087:9072]},
     {storeUnit_maskInput_hi[9071:9056]},
     {storeUnit_maskInput_hi[9055:9040]},
     {storeUnit_maskInput_hi[9039:9024]},
     {storeUnit_maskInput_hi[9023:9008]},
     {storeUnit_maskInput_hi[9007:8992]},
     {storeUnit_maskInput_hi[8991:8976]},
     {storeUnit_maskInput_hi[8975:8960]},
     {storeUnit_maskInput_hi[8959:8944]},
     {storeUnit_maskInput_hi[8943:8928]},
     {storeUnit_maskInput_hi[8927:8912]},
     {storeUnit_maskInput_hi[8911:8896]},
     {storeUnit_maskInput_hi[8895:8880]},
     {storeUnit_maskInput_hi[8879:8864]},
     {storeUnit_maskInput_hi[8863:8848]},
     {storeUnit_maskInput_hi[8847:8832]},
     {storeUnit_maskInput_hi[8831:8816]},
     {storeUnit_maskInput_hi[8815:8800]},
     {storeUnit_maskInput_hi[8799:8784]},
     {storeUnit_maskInput_hi[8783:8768]},
     {storeUnit_maskInput_hi[8767:8752]},
     {storeUnit_maskInput_hi[8751:8736]},
     {storeUnit_maskInput_hi[8735:8720]},
     {storeUnit_maskInput_hi[8719:8704]},
     {storeUnit_maskInput_hi[8703:8688]},
     {storeUnit_maskInput_hi[8687:8672]},
     {storeUnit_maskInput_hi[8671:8656]},
     {storeUnit_maskInput_hi[8655:8640]},
     {storeUnit_maskInput_hi[8639:8624]},
     {storeUnit_maskInput_hi[8623:8608]},
     {storeUnit_maskInput_hi[8607:8592]},
     {storeUnit_maskInput_hi[8591:8576]},
     {storeUnit_maskInput_hi[8575:8560]},
     {storeUnit_maskInput_hi[8559:8544]},
     {storeUnit_maskInput_hi[8543:8528]},
     {storeUnit_maskInput_hi[8527:8512]},
     {storeUnit_maskInput_hi[8511:8496]},
     {storeUnit_maskInput_hi[8495:8480]},
     {storeUnit_maskInput_hi[8479:8464]},
     {storeUnit_maskInput_hi[8463:8448]},
     {storeUnit_maskInput_hi[8447:8432]},
     {storeUnit_maskInput_hi[8431:8416]},
     {storeUnit_maskInput_hi[8415:8400]},
     {storeUnit_maskInput_hi[8399:8384]},
     {storeUnit_maskInput_hi[8383:8368]},
     {storeUnit_maskInput_hi[8367:8352]},
     {storeUnit_maskInput_hi[8351:8336]},
     {storeUnit_maskInput_hi[8335:8320]},
     {storeUnit_maskInput_hi[8319:8304]},
     {storeUnit_maskInput_hi[8303:8288]},
     {storeUnit_maskInput_hi[8287:8272]},
     {storeUnit_maskInput_hi[8271:8256]},
     {storeUnit_maskInput_hi[8255:8240]},
     {storeUnit_maskInput_hi[8239:8224]},
     {storeUnit_maskInput_hi[8223:8208]},
     {storeUnit_maskInput_hi[8207:8192]},
     {storeUnit_maskInput_hi[8191:8176]},
     {storeUnit_maskInput_hi[8175:8160]},
     {storeUnit_maskInput_hi[8159:8144]},
     {storeUnit_maskInput_hi[8143:8128]},
     {storeUnit_maskInput_hi[8127:8112]},
     {storeUnit_maskInput_hi[8111:8096]},
     {storeUnit_maskInput_hi[8095:8080]},
     {storeUnit_maskInput_hi[8079:8064]},
     {storeUnit_maskInput_hi[8063:8048]},
     {storeUnit_maskInput_hi[8047:8032]},
     {storeUnit_maskInput_hi[8031:8016]},
     {storeUnit_maskInput_hi[8015:8000]},
     {storeUnit_maskInput_hi[7999:7984]},
     {storeUnit_maskInput_hi[7983:7968]},
     {storeUnit_maskInput_hi[7967:7952]},
     {storeUnit_maskInput_hi[7951:7936]},
     {storeUnit_maskInput_hi[7935:7920]},
     {storeUnit_maskInput_hi[7919:7904]},
     {storeUnit_maskInput_hi[7903:7888]},
     {storeUnit_maskInput_hi[7887:7872]},
     {storeUnit_maskInput_hi[7871:7856]},
     {storeUnit_maskInput_hi[7855:7840]},
     {storeUnit_maskInput_hi[7839:7824]},
     {storeUnit_maskInput_hi[7823:7808]},
     {storeUnit_maskInput_hi[7807:7792]},
     {storeUnit_maskInput_hi[7791:7776]},
     {storeUnit_maskInput_hi[7775:7760]},
     {storeUnit_maskInput_hi[7759:7744]},
     {storeUnit_maskInput_hi[7743:7728]},
     {storeUnit_maskInput_hi[7727:7712]},
     {storeUnit_maskInput_hi[7711:7696]},
     {storeUnit_maskInput_hi[7695:7680]},
     {storeUnit_maskInput_hi[7679:7664]},
     {storeUnit_maskInput_hi[7663:7648]},
     {storeUnit_maskInput_hi[7647:7632]},
     {storeUnit_maskInput_hi[7631:7616]},
     {storeUnit_maskInput_hi[7615:7600]},
     {storeUnit_maskInput_hi[7599:7584]},
     {storeUnit_maskInput_hi[7583:7568]},
     {storeUnit_maskInput_hi[7567:7552]},
     {storeUnit_maskInput_hi[7551:7536]},
     {storeUnit_maskInput_hi[7535:7520]},
     {storeUnit_maskInput_hi[7519:7504]},
     {storeUnit_maskInput_hi[7503:7488]},
     {storeUnit_maskInput_hi[7487:7472]},
     {storeUnit_maskInput_hi[7471:7456]},
     {storeUnit_maskInput_hi[7455:7440]},
     {storeUnit_maskInput_hi[7439:7424]},
     {storeUnit_maskInput_hi[7423:7408]},
     {storeUnit_maskInput_hi[7407:7392]},
     {storeUnit_maskInput_hi[7391:7376]},
     {storeUnit_maskInput_hi[7375:7360]},
     {storeUnit_maskInput_hi[7359:7344]},
     {storeUnit_maskInput_hi[7343:7328]},
     {storeUnit_maskInput_hi[7327:7312]},
     {storeUnit_maskInput_hi[7311:7296]},
     {storeUnit_maskInput_hi[7295:7280]},
     {storeUnit_maskInput_hi[7279:7264]},
     {storeUnit_maskInput_hi[7263:7248]},
     {storeUnit_maskInput_hi[7247:7232]},
     {storeUnit_maskInput_hi[7231:7216]},
     {storeUnit_maskInput_hi[7215:7200]},
     {storeUnit_maskInput_hi[7199:7184]},
     {storeUnit_maskInput_hi[7183:7168]},
     {storeUnit_maskInput_hi[7167:7152]},
     {storeUnit_maskInput_hi[7151:7136]},
     {storeUnit_maskInput_hi[7135:7120]},
     {storeUnit_maskInput_hi[7119:7104]},
     {storeUnit_maskInput_hi[7103:7088]},
     {storeUnit_maskInput_hi[7087:7072]},
     {storeUnit_maskInput_hi[7071:7056]},
     {storeUnit_maskInput_hi[7055:7040]},
     {storeUnit_maskInput_hi[7039:7024]},
     {storeUnit_maskInput_hi[7023:7008]},
     {storeUnit_maskInput_hi[7007:6992]},
     {storeUnit_maskInput_hi[6991:6976]},
     {storeUnit_maskInput_hi[6975:6960]},
     {storeUnit_maskInput_hi[6959:6944]},
     {storeUnit_maskInput_hi[6943:6928]},
     {storeUnit_maskInput_hi[6927:6912]},
     {storeUnit_maskInput_hi[6911:6896]},
     {storeUnit_maskInput_hi[6895:6880]},
     {storeUnit_maskInput_hi[6879:6864]},
     {storeUnit_maskInput_hi[6863:6848]},
     {storeUnit_maskInput_hi[6847:6832]},
     {storeUnit_maskInput_hi[6831:6816]},
     {storeUnit_maskInput_hi[6815:6800]},
     {storeUnit_maskInput_hi[6799:6784]},
     {storeUnit_maskInput_hi[6783:6768]},
     {storeUnit_maskInput_hi[6767:6752]},
     {storeUnit_maskInput_hi[6751:6736]},
     {storeUnit_maskInput_hi[6735:6720]},
     {storeUnit_maskInput_hi[6719:6704]},
     {storeUnit_maskInput_hi[6703:6688]},
     {storeUnit_maskInput_hi[6687:6672]},
     {storeUnit_maskInput_hi[6671:6656]},
     {storeUnit_maskInput_hi[6655:6640]},
     {storeUnit_maskInput_hi[6639:6624]},
     {storeUnit_maskInput_hi[6623:6608]},
     {storeUnit_maskInput_hi[6607:6592]},
     {storeUnit_maskInput_hi[6591:6576]},
     {storeUnit_maskInput_hi[6575:6560]},
     {storeUnit_maskInput_hi[6559:6544]},
     {storeUnit_maskInput_hi[6543:6528]},
     {storeUnit_maskInput_hi[6527:6512]},
     {storeUnit_maskInput_hi[6511:6496]},
     {storeUnit_maskInput_hi[6495:6480]},
     {storeUnit_maskInput_hi[6479:6464]},
     {storeUnit_maskInput_hi[6463:6448]},
     {storeUnit_maskInput_hi[6447:6432]},
     {storeUnit_maskInput_hi[6431:6416]},
     {storeUnit_maskInput_hi[6415:6400]},
     {storeUnit_maskInput_hi[6399:6384]},
     {storeUnit_maskInput_hi[6383:6368]},
     {storeUnit_maskInput_hi[6367:6352]},
     {storeUnit_maskInput_hi[6351:6336]},
     {storeUnit_maskInput_hi[6335:6320]},
     {storeUnit_maskInput_hi[6319:6304]},
     {storeUnit_maskInput_hi[6303:6288]},
     {storeUnit_maskInput_hi[6287:6272]},
     {storeUnit_maskInput_hi[6271:6256]},
     {storeUnit_maskInput_hi[6255:6240]},
     {storeUnit_maskInput_hi[6239:6224]},
     {storeUnit_maskInput_hi[6223:6208]},
     {storeUnit_maskInput_hi[6207:6192]},
     {storeUnit_maskInput_hi[6191:6176]},
     {storeUnit_maskInput_hi[6175:6160]},
     {storeUnit_maskInput_hi[6159:6144]},
     {storeUnit_maskInput_hi[6143:6128]},
     {storeUnit_maskInput_hi[6127:6112]},
     {storeUnit_maskInput_hi[6111:6096]},
     {storeUnit_maskInput_hi[6095:6080]},
     {storeUnit_maskInput_hi[6079:6064]},
     {storeUnit_maskInput_hi[6063:6048]},
     {storeUnit_maskInput_hi[6047:6032]},
     {storeUnit_maskInput_hi[6031:6016]},
     {storeUnit_maskInput_hi[6015:6000]},
     {storeUnit_maskInput_hi[5999:5984]},
     {storeUnit_maskInput_hi[5983:5968]},
     {storeUnit_maskInput_hi[5967:5952]},
     {storeUnit_maskInput_hi[5951:5936]},
     {storeUnit_maskInput_hi[5935:5920]},
     {storeUnit_maskInput_hi[5919:5904]},
     {storeUnit_maskInput_hi[5903:5888]},
     {storeUnit_maskInput_hi[5887:5872]},
     {storeUnit_maskInput_hi[5871:5856]},
     {storeUnit_maskInput_hi[5855:5840]},
     {storeUnit_maskInput_hi[5839:5824]},
     {storeUnit_maskInput_hi[5823:5808]},
     {storeUnit_maskInput_hi[5807:5792]},
     {storeUnit_maskInput_hi[5791:5776]},
     {storeUnit_maskInput_hi[5775:5760]},
     {storeUnit_maskInput_hi[5759:5744]},
     {storeUnit_maskInput_hi[5743:5728]},
     {storeUnit_maskInput_hi[5727:5712]},
     {storeUnit_maskInput_hi[5711:5696]},
     {storeUnit_maskInput_hi[5695:5680]},
     {storeUnit_maskInput_hi[5679:5664]},
     {storeUnit_maskInput_hi[5663:5648]},
     {storeUnit_maskInput_hi[5647:5632]},
     {storeUnit_maskInput_hi[5631:5616]},
     {storeUnit_maskInput_hi[5615:5600]},
     {storeUnit_maskInput_hi[5599:5584]},
     {storeUnit_maskInput_hi[5583:5568]},
     {storeUnit_maskInput_hi[5567:5552]},
     {storeUnit_maskInput_hi[5551:5536]},
     {storeUnit_maskInput_hi[5535:5520]},
     {storeUnit_maskInput_hi[5519:5504]},
     {storeUnit_maskInput_hi[5503:5488]},
     {storeUnit_maskInput_hi[5487:5472]},
     {storeUnit_maskInput_hi[5471:5456]},
     {storeUnit_maskInput_hi[5455:5440]},
     {storeUnit_maskInput_hi[5439:5424]},
     {storeUnit_maskInput_hi[5423:5408]},
     {storeUnit_maskInput_hi[5407:5392]},
     {storeUnit_maskInput_hi[5391:5376]},
     {storeUnit_maskInput_hi[5375:5360]},
     {storeUnit_maskInput_hi[5359:5344]},
     {storeUnit_maskInput_hi[5343:5328]},
     {storeUnit_maskInput_hi[5327:5312]},
     {storeUnit_maskInput_hi[5311:5296]},
     {storeUnit_maskInput_hi[5295:5280]},
     {storeUnit_maskInput_hi[5279:5264]},
     {storeUnit_maskInput_hi[5263:5248]},
     {storeUnit_maskInput_hi[5247:5232]},
     {storeUnit_maskInput_hi[5231:5216]},
     {storeUnit_maskInput_hi[5215:5200]},
     {storeUnit_maskInput_hi[5199:5184]},
     {storeUnit_maskInput_hi[5183:5168]},
     {storeUnit_maskInput_hi[5167:5152]},
     {storeUnit_maskInput_hi[5151:5136]},
     {storeUnit_maskInput_hi[5135:5120]},
     {storeUnit_maskInput_hi[5119:5104]},
     {storeUnit_maskInput_hi[5103:5088]},
     {storeUnit_maskInput_hi[5087:5072]},
     {storeUnit_maskInput_hi[5071:5056]},
     {storeUnit_maskInput_hi[5055:5040]},
     {storeUnit_maskInput_hi[5039:5024]},
     {storeUnit_maskInput_hi[5023:5008]},
     {storeUnit_maskInput_hi[5007:4992]},
     {storeUnit_maskInput_hi[4991:4976]},
     {storeUnit_maskInput_hi[4975:4960]},
     {storeUnit_maskInput_hi[4959:4944]},
     {storeUnit_maskInput_hi[4943:4928]},
     {storeUnit_maskInput_hi[4927:4912]},
     {storeUnit_maskInput_hi[4911:4896]},
     {storeUnit_maskInput_hi[4895:4880]},
     {storeUnit_maskInput_hi[4879:4864]},
     {storeUnit_maskInput_hi[4863:4848]},
     {storeUnit_maskInput_hi[4847:4832]},
     {storeUnit_maskInput_hi[4831:4816]},
     {storeUnit_maskInput_hi[4815:4800]},
     {storeUnit_maskInput_hi[4799:4784]},
     {storeUnit_maskInput_hi[4783:4768]},
     {storeUnit_maskInput_hi[4767:4752]},
     {storeUnit_maskInput_hi[4751:4736]},
     {storeUnit_maskInput_hi[4735:4720]},
     {storeUnit_maskInput_hi[4719:4704]},
     {storeUnit_maskInput_hi[4703:4688]},
     {storeUnit_maskInput_hi[4687:4672]},
     {storeUnit_maskInput_hi[4671:4656]},
     {storeUnit_maskInput_hi[4655:4640]},
     {storeUnit_maskInput_hi[4639:4624]},
     {storeUnit_maskInput_hi[4623:4608]},
     {storeUnit_maskInput_hi[4607:4592]},
     {storeUnit_maskInput_hi[4591:4576]},
     {storeUnit_maskInput_hi[4575:4560]},
     {storeUnit_maskInput_hi[4559:4544]},
     {storeUnit_maskInput_hi[4543:4528]},
     {storeUnit_maskInput_hi[4527:4512]},
     {storeUnit_maskInput_hi[4511:4496]},
     {storeUnit_maskInput_hi[4495:4480]},
     {storeUnit_maskInput_hi[4479:4464]},
     {storeUnit_maskInput_hi[4463:4448]},
     {storeUnit_maskInput_hi[4447:4432]},
     {storeUnit_maskInput_hi[4431:4416]},
     {storeUnit_maskInput_hi[4415:4400]},
     {storeUnit_maskInput_hi[4399:4384]},
     {storeUnit_maskInput_hi[4383:4368]},
     {storeUnit_maskInput_hi[4367:4352]},
     {storeUnit_maskInput_hi[4351:4336]},
     {storeUnit_maskInput_hi[4335:4320]},
     {storeUnit_maskInput_hi[4319:4304]},
     {storeUnit_maskInput_hi[4303:4288]},
     {storeUnit_maskInput_hi[4287:4272]},
     {storeUnit_maskInput_hi[4271:4256]},
     {storeUnit_maskInput_hi[4255:4240]},
     {storeUnit_maskInput_hi[4239:4224]},
     {storeUnit_maskInput_hi[4223:4208]},
     {storeUnit_maskInput_hi[4207:4192]},
     {storeUnit_maskInput_hi[4191:4176]},
     {storeUnit_maskInput_hi[4175:4160]},
     {storeUnit_maskInput_hi[4159:4144]},
     {storeUnit_maskInput_hi[4143:4128]},
     {storeUnit_maskInput_hi[4127:4112]},
     {storeUnit_maskInput_hi[4111:4096]},
     {storeUnit_maskInput_hi[4095:4080]},
     {storeUnit_maskInput_hi[4079:4064]},
     {storeUnit_maskInput_hi[4063:4048]},
     {storeUnit_maskInput_hi[4047:4032]},
     {storeUnit_maskInput_hi[4031:4016]},
     {storeUnit_maskInput_hi[4015:4000]},
     {storeUnit_maskInput_hi[3999:3984]},
     {storeUnit_maskInput_hi[3983:3968]},
     {storeUnit_maskInput_hi[3967:3952]},
     {storeUnit_maskInput_hi[3951:3936]},
     {storeUnit_maskInput_hi[3935:3920]},
     {storeUnit_maskInput_hi[3919:3904]},
     {storeUnit_maskInput_hi[3903:3888]},
     {storeUnit_maskInput_hi[3887:3872]},
     {storeUnit_maskInput_hi[3871:3856]},
     {storeUnit_maskInput_hi[3855:3840]},
     {storeUnit_maskInput_hi[3839:3824]},
     {storeUnit_maskInput_hi[3823:3808]},
     {storeUnit_maskInput_hi[3807:3792]},
     {storeUnit_maskInput_hi[3791:3776]},
     {storeUnit_maskInput_hi[3775:3760]},
     {storeUnit_maskInput_hi[3759:3744]},
     {storeUnit_maskInput_hi[3743:3728]},
     {storeUnit_maskInput_hi[3727:3712]},
     {storeUnit_maskInput_hi[3711:3696]},
     {storeUnit_maskInput_hi[3695:3680]},
     {storeUnit_maskInput_hi[3679:3664]},
     {storeUnit_maskInput_hi[3663:3648]},
     {storeUnit_maskInput_hi[3647:3632]},
     {storeUnit_maskInput_hi[3631:3616]},
     {storeUnit_maskInput_hi[3615:3600]},
     {storeUnit_maskInput_hi[3599:3584]},
     {storeUnit_maskInput_hi[3583:3568]},
     {storeUnit_maskInput_hi[3567:3552]},
     {storeUnit_maskInput_hi[3551:3536]},
     {storeUnit_maskInput_hi[3535:3520]},
     {storeUnit_maskInput_hi[3519:3504]},
     {storeUnit_maskInput_hi[3503:3488]},
     {storeUnit_maskInput_hi[3487:3472]},
     {storeUnit_maskInput_hi[3471:3456]},
     {storeUnit_maskInput_hi[3455:3440]},
     {storeUnit_maskInput_hi[3439:3424]},
     {storeUnit_maskInput_hi[3423:3408]},
     {storeUnit_maskInput_hi[3407:3392]},
     {storeUnit_maskInput_hi[3391:3376]},
     {storeUnit_maskInput_hi[3375:3360]},
     {storeUnit_maskInput_hi[3359:3344]},
     {storeUnit_maskInput_hi[3343:3328]},
     {storeUnit_maskInput_hi[3327:3312]},
     {storeUnit_maskInput_hi[3311:3296]},
     {storeUnit_maskInput_hi[3295:3280]},
     {storeUnit_maskInput_hi[3279:3264]},
     {storeUnit_maskInput_hi[3263:3248]},
     {storeUnit_maskInput_hi[3247:3232]},
     {storeUnit_maskInput_hi[3231:3216]},
     {storeUnit_maskInput_hi[3215:3200]},
     {storeUnit_maskInput_hi[3199:3184]},
     {storeUnit_maskInput_hi[3183:3168]},
     {storeUnit_maskInput_hi[3167:3152]},
     {storeUnit_maskInput_hi[3151:3136]},
     {storeUnit_maskInput_hi[3135:3120]},
     {storeUnit_maskInput_hi[3119:3104]},
     {storeUnit_maskInput_hi[3103:3088]},
     {storeUnit_maskInput_hi[3087:3072]},
     {storeUnit_maskInput_hi[3071:3056]},
     {storeUnit_maskInput_hi[3055:3040]},
     {storeUnit_maskInput_hi[3039:3024]},
     {storeUnit_maskInput_hi[3023:3008]},
     {storeUnit_maskInput_hi[3007:2992]},
     {storeUnit_maskInput_hi[2991:2976]},
     {storeUnit_maskInput_hi[2975:2960]},
     {storeUnit_maskInput_hi[2959:2944]},
     {storeUnit_maskInput_hi[2943:2928]},
     {storeUnit_maskInput_hi[2927:2912]},
     {storeUnit_maskInput_hi[2911:2896]},
     {storeUnit_maskInput_hi[2895:2880]},
     {storeUnit_maskInput_hi[2879:2864]},
     {storeUnit_maskInput_hi[2863:2848]},
     {storeUnit_maskInput_hi[2847:2832]},
     {storeUnit_maskInput_hi[2831:2816]},
     {storeUnit_maskInput_hi[2815:2800]},
     {storeUnit_maskInput_hi[2799:2784]},
     {storeUnit_maskInput_hi[2783:2768]},
     {storeUnit_maskInput_hi[2767:2752]},
     {storeUnit_maskInput_hi[2751:2736]},
     {storeUnit_maskInput_hi[2735:2720]},
     {storeUnit_maskInput_hi[2719:2704]},
     {storeUnit_maskInput_hi[2703:2688]},
     {storeUnit_maskInput_hi[2687:2672]},
     {storeUnit_maskInput_hi[2671:2656]},
     {storeUnit_maskInput_hi[2655:2640]},
     {storeUnit_maskInput_hi[2639:2624]},
     {storeUnit_maskInput_hi[2623:2608]},
     {storeUnit_maskInput_hi[2607:2592]},
     {storeUnit_maskInput_hi[2591:2576]},
     {storeUnit_maskInput_hi[2575:2560]},
     {storeUnit_maskInput_hi[2559:2544]},
     {storeUnit_maskInput_hi[2543:2528]},
     {storeUnit_maskInput_hi[2527:2512]},
     {storeUnit_maskInput_hi[2511:2496]},
     {storeUnit_maskInput_hi[2495:2480]},
     {storeUnit_maskInput_hi[2479:2464]},
     {storeUnit_maskInput_hi[2463:2448]},
     {storeUnit_maskInput_hi[2447:2432]},
     {storeUnit_maskInput_hi[2431:2416]},
     {storeUnit_maskInput_hi[2415:2400]},
     {storeUnit_maskInput_hi[2399:2384]},
     {storeUnit_maskInput_hi[2383:2368]},
     {storeUnit_maskInput_hi[2367:2352]},
     {storeUnit_maskInput_hi[2351:2336]},
     {storeUnit_maskInput_hi[2335:2320]},
     {storeUnit_maskInput_hi[2319:2304]},
     {storeUnit_maskInput_hi[2303:2288]},
     {storeUnit_maskInput_hi[2287:2272]},
     {storeUnit_maskInput_hi[2271:2256]},
     {storeUnit_maskInput_hi[2255:2240]},
     {storeUnit_maskInput_hi[2239:2224]},
     {storeUnit_maskInput_hi[2223:2208]},
     {storeUnit_maskInput_hi[2207:2192]},
     {storeUnit_maskInput_hi[2191:2176]},
     {storeUnit_maskInput_hi[2175:2160]},
     {storeUnit_maskInput_hi[2159:2144]},
     {storeUnit_maskInput_hi[2143:2128]},
     {storeUnit_maskInput_hi[2127:2112]},
     {storeUnit_maskInput_hi[2111:2096]},
     {storeUnit_maskInput_hi[2095:2080]},
     {storeUnit_maskInput_hi[2079:2064]},
     {storeUnit_maskInput_hi[2063:2048]},
     {storeUnit_maskInput_hi[2047:2032]},
     {storeUnit_maskInput_hi[2031:2016]},
     {storeUnit_maskInput_hi[2015:2000]},
     {storeUnit_maskInput_hi[1999:1984]},
     {storeUnit_maskInput_hi[1983:1968]},
     {storeUnit_maskInput_hi[1967:1952]},
     {storeUnit_maskInput_hi[1951:1936]},
     {storeUnit_maskInput_hi[1935:1920]},
     {storeUnit_maskInput_hi[1919:1904]},
     {storeUnit_maskInput_hi[1903:1888]},
     {storeUnit_maskInput_hi[1887:1872]},
     {storeUnit_maskInput_hi[1871:1856]},
     {storeUnit_maskInput_hi[1855:1840]},
     {storeUnit_maskInput_hi[1839:1824]},
     {storeUnit_maskInput_hi[1823:1808]},
     {storeUnit_maskInput_hi[1807:1792]},
     {storeUnit_maskInput_hi[1791:1776]},
     {storeUnit_maskInput_hi[1775:1760]},
     {storeUnit_maskInput_hi[1759:1744]},
     {storeUnit_maskInput_hi[1743:1728]},
     {storeUnit_maskInput_hi[1727:1712]},
     {storeUnit_maskInput_hi[1711:1696]},
     {storeUnit_maskInput_hi[1695:1680]},
     {storeUnit_maskInput_hi[1679:1664]},
     {storeUnit_maskInput_hi[1663:1648]},
     {storeUnit_maskInput_hi[1647:1632]},
     {storeUnit_maskInput_hi[1631:1616]},
     {storeUnit_maskInput_hi[1615:1600]},
     {storeUnit_maskInput_hi[1599:1584]},
     {storeUnit_maskInput_hi[1583:1568]},
     {storeUnit_maskInput_hi[1567:1552]},
     {storeUnit_maskInput_hi[1551:1536]},
     {storeUnit_maskInput_hi[1535:1520]},
     {storeUnit_maskInput_hi[1519:1504]},
     {storeUnit_maskInput_hi[1503:1488]},
     {storeUnit_maskInput_hi[1487:1472]},
     {storeUnit_maskInput_hi[1471:1456]},
     {storeUnit_maskInput_hi[1455:1440]},
     {storeUnit_maskInput_hi[1439:1424]},
     {storeUnit_maskInput_hi[1423:1408]},
     {storeUnit_maskInput_hi[1407:1392]},
     {storeUnit_maskInput_hi[1391:1376]},
     {storeUnit_maskInput_hi[1375:1360]},
     {storeUnit_maskInput_hi[1359:1344]},
     {storeUnit_maskInput_hi[1343:1328]},
     {storeUnit_maskInput_hi[1327:1312]},
     {storeUnit_maskInput_hi[1311:1296]},
     {storeUnit_maskInput_hi[1295:1280]},
     {storeUnit_maskInput_hi[1279:1264]},
     {storeUnit_maskInput_hi[1263:1248]},
     {storeUnit_maskInput_hi[1247:1232]},
     {storeUnit_maskInput_hi[1231:1216]},
     {storeUnit_maskInput_hi[1215:1200]},
     {storeUnit_maskInput_hi[1199:1184]},
     {storeUnit_maskInput_hi[1183:1168]},
     {storeUnit_maskInput_hi[1167:1152]},
     {storeUnit_maskInput_hi[1151:1136]},
     {storeUnit_maskInput_hi[1135:1120]},
     {storeUnit_maskInput_hi[1119:1104]},
     {storeUnit_maskInput_hi[1103:1088]},
     {storeUnit_maskInput_hi[1087:1072]},
     {storeUnit_maskInput_hi[1071:1056]},
     {storeUnit_maskInput_hi[1055:1040]},
     {storeUnit_maskInput_hi[1039:1024]},
     {storeUnit_maskInput_hi[1023:1008]},
     {storeUnit_maskInput_hi[1007:992]},
     {storeUnit_maskInput_hi[991:976]},
     {storeUnit_maskInput_hi[975:960]},
     {storeUnit_maskInput_hi[959:944]},
     {storeUnit_maskInput_hi[943:928]},
     {storeUnit_maskInput_hi[927:912]},
     {storeUnit_maskInput_hi[911:896]},
     {storeUnit_maskInput_hi[895:880]},
     {storeUnit_maskInput_hi[879:864]},
     {storeUnit_maskInput_hi[863:848]},
     {storeUnit_maskInput_hi[847:832]},
     {storeUnit_maskInput_hi[831:816]},
     {storeUnit_maskInput_hi[815:800]},
     {storeUnit_maskInput_hi[799:784]},
     {storeUnit_maskInput_hi[783:768]},
     {storeUnit_maskInput_hi[767:752]},
     {storeUnit_maskInput_hi[751:736]},
     {storeUnit_maskInput_hi[735:720]},
     {storeUnit_maskInput_hi[719:704]},
     {storeUnit_maskInput_hi[703:688]},
     {storeUnit_maskInput_hi[687:672]},
     {storeUnit_maskInput_hi[671:656]},
     {storeUnit_maskInput_hi[655:640]},
     {storeUnit_maskInput_hi[639:624]},
     {storeUnit_maskInput_hi[623:608]},
     {storeUnit_maskInput_hi[607:592]},
     {storeUnit_maskInput_hi[591:576]},
     {storeUnit_maskInput_hi[575:560]},
     {storeUnit_maskInput_hi[559:544]},
     {storeUnit_maskInput_hi[543:528]},
     {storeUnit_maskInput_hi[527:512]},
     {storeUnit_maskInput_hi[511:496]},
     {storeUnit_maskInput_hi[495:480]},
     {storeUnit_maskInput_hi[479:464]},
     {storeUnit_maskInput_hi[463:448]},
     {storeUnit_maskInput_hi[447:432]},
     {storeUnit_maskInput_hi[431:416]},
     {storeUnit_maskInput_hi[415:400]},
     {storeUnit_maskInput_hi[399:384]},
     {storeUnit_maskInput_hi[383:368]},
     {storeUnit_maskInput_hi[367:352]},
     {storeUnit_maskInput_hi[351:336]},
     {storeUnit_maskInput_hi[335:320]},
     {storeUnit_maskInput_hi[319:304]},
     {storeUnit_maskInput_hi[303:288]},
     {storeUnit_maskInput_hi[287:272]},
     {storeUnit_maskInput_hi[271:256]},
     {storeUnit_maskInput_hi[255:240]},
     {storeUnit_maskInput_hi[239:224]},
     {storeUnit_maskInput_hi[223:208]},
     {storeUnit_maskInput_hi[207:192]},
     {storeUnit_maskInput_hi[191:176]},
     {storeUnit_maskInput_hi[175:160]},
     {storeUnit_maskInput_hi[159:144]},
     {storeUnit_maskInput_hi[143:128]},
     {storeUnit_maskInput_hi[127:112]},
     {storeUnit_maskInput_hi[111:96]},
     {storeUnit_maskInput_hi[95:80]},
     {storeUnit_maskInput_hi[79:64]},
     {storeUnit_maskInput_hi[63:48]},
     {storeUnit_maskInput_hi[47:32]},
     {storeUnit_maskInput_hi[31:16]},
     {storeUnit_maskInput_hi[15:0]},
     {storeUnit_maskInput_lo[16383:16368]},
     {storeUnit_maskInput_lo[16367:16352]},
     {storeUnit_maskInput_lo[16351:16336]},
     {storeUnit_maskInput_lo[16335:16320]},
     {storeUnit_maskInput_lo[16319:16304]},
     {storeUnit_maskInput_lo[16303:16288]},
     {storeUnit_maskInput_lo[16287:16272]},
     {storeUnit_maskInput_lo[16271:16256]},
     {storeUnit_maskInput_lo[16255:16240]},
     {storeUnit_maskInput_lo[16239:16224]},
     {storeUnit_maskInput_lo[16223:16208]},
     {storeUnit_maskInput_lo[16207:16192]},
     {storeUnit_maskInput_lo[16191:16176]},
     {storeUnit_maskInput_lo[16175:16160]},
     {storeUnit_maskInput_lo[16159:16144]},
     {storeUnit_maskInput_lo[16143:16128]},
     {storeUnit_maskInput_lo[16127:16112]},
     {storeUnit_maskInput_lo[16111:16096]},
     {storeUnit_maskInput_lo[16095:16080]},
     {storeUnit_maskInput_lo[16079:16064]},
     {storeUnit_maskInput_lo[16063:16048]},
     {storeUnit_maskInput_lo[16047:16032]},
     {storeUnit_maskInput_lo[16031:16016]},
     {storeUnit_maskInput_lo[16015:16000]},
     {storeUnit_maskInput_lo[15999:15984]},
     {storeUnit_maskInput_lo[15983:15968]},
     {storeUnit_maskInput_lo[15967:15952]},
     {storeUnit_maskInput_lo[15951:15936]},
     {storeUnit_maskInput_lo[15935:15920]},
     {storeUnit_maskInput_lo[15919:15904]},
     {storeUnit_maskInput_lo[15903:15888]},
     {storeUnit_maskInput_lo[15887:15872]},
     {storeUnit_maskInput_lo[15871:15856]},
     {storeUnit_maskInput_lo[15855:15840]},
     {storeUnit_maskInput_lo[15839:15824]},
     {storeUnit_maskInput_lo[15823:15808]},
     {storeUnit_maskInput_lo[15807:15792]},
     {storeUnit_maskInput_lo[15791:15776]},
     {storeUnit_maskInput_lo[15775:15760]},
     {storeUnit_maskInput_lo[15759:15744]},
     {storeUnit_maskInput_lo[15743:15728]},
     {storeUnit_maskInput_lo[15727:15712]},
     {storeUnit_maskInput_lo[15711:15696]},
     {storeUnit_maskInput_lo[15695:15680]},
     {storeUnit_maskInput_lo[15679:15664]},
     {storeUnit_maskInput_lo[15663:15648]},
     {storeUnit_maskInput_lo[15647:15632]},
     {storeUnit_maskInput_lo[15631:15616]},
     {storeUnit_maskInput_lo[15615:15600]},
     {storeUnit_maskInput_lo[15599:15584]},
     {storeUnit_maskInput_lo[15583:15568]},
     {storeUnit_maskInput_lo[15567:15552]},
     {storeUnit_maskInput_lo[15551:15536]},
     {storeUnit_maskInput_lo[15535:15520]},
     {storeUnit_maskInput_lo[15519:15504]},
     {storeUnit_maskInput_lo[15503:15488]},
     {storeUnit_maskInput_lo[15487:15472]},
     {storeUnit_maskInput_lo[15471:15456]},
     {storeUnit_maskInput_lo[15455:15440]},
     {storeUnit_maskInput_lo[15439:15424]},
     {storeUnit_maskInput_lo[15423:15408]},
     {storeUnit_maskInput_lo[15407:15392]},
     {storeUnit_maskInput_lo[15391:15376]},
     {storeUnit_maskInput_lo[15375:15360]},
     {storeUnit_maskInput_lo[15359:15344]},
     {storeUnit_maskInput_lo[15343:15328]},
     {storeUnit_maskInput_lo[15327:15312]},
     {storeUnit_maskInput_lo[15311:15296]},
     {storeUnit_maskInput_lo[15295:15280]},
     {storeUnit_maskInput_lo[15279:15264]},
     {storeUnit_maskInput_lo[15263:15248]},
     {storeUnit_maskInput_lo[15247:15232]},
     {storeUnit_maskInput_lo[15231:15216]},
     {storeUnit_maskInput_lo[15215:15200]},
     {storeUnit_maskInput_lo[15199:15184]},
     {storeUnit_maskInput_lo[15183:15168]},
     {storeUnit_maskInput_lo[15167:15152]},
     {storeUnit_maskInput_lo[15151:15136]},
     {storeUnit_maskInput_lo[15135:15120]},
     {storeUnit_maskInput_lo[15119:15104]},
     {storeUnit_maskInput_lo[15103:15088]},
     {storeUnit_maskInput_lo[15087:15072]},
     {storeUnit_maskInput_lo[15071:15056]},
     {storeUnit_maskInput_lo[15055:15040]},
     {storeUnit_maskInput_lo[15039:15024]},
     {storeUnit_maskInput_lo[15023:15008]},
     {storeUnit_maskInput_lo[15007:14992]},
     {storeUnit_maskInput_lo[14991:14976]},
     {storeUnit_maskInput_lo[14975:14960]},
     {storeUnit_maskInput_lo[14959:14944]},
     {storeUnit_maskInput_lo[14943:14928]},
     {storeUnit_maskInput_lo[14927:14912]},
     {storeUnit_maskInput_lo[14911:14896]},
     {storeUnit_maskInput_lo[14895:14880]},
     {storeUnit_maskInput_lo[14879:14864]},
     {storeUnit_maskInput_lo[14863:14848]},
     {storeUnit_maskInput_lo[14847:14832]},
     {storeUnit_maskInput_lo[14831:14816]},
     {storeUnit_maskInput_lo[14815:14800]},
     {storeUnit_maskInput_lo[14799:14784]},
     {storeUnit_maskInput_lo[14783:14768]},
     {storeUnit_maskInput_lo[14767:14752]},
     {storeUnit_maskInput_lo[14751:14736]},
     {storeUnit_maskInput_lo[14735:14720]},
     {storeUnit_maskInput_lo[14719:14704]},
     {storeUnit_maskInput_lo[14703:14688]},
     {storeUnit_maskInput_lo[14687:14672]},
     {storeUnit_maskInput_lo[14671:14656]},
     {storeUnit_maskInput_lo[14655:14640]},
     {storeUnit_maskInput_lo[14639:14624]},
     {storeUnit_maskInput_lo[14623:14608]},
     {storeUnit_maskInput_lo[14607:14592]},
     {storeUnit_maskInput_lo[14591:14576]},
     {storeUnit_maskInput_lo[14575:14560]},
     {storeUnit_maskInput_lo[14559:14544]},
     {storeUnit_maskInput_lo[14543:14528]},
     {storeUnit_maskInput_lo[14527:14512]},
     {storeUnit_maskInput_lo[14511:14496]},
     {storeUnit_maskInput_lo[14495:14480]},
     {storeUnit_maskInput_lo[14479:14464]},
     {storeUnit_maskInput_lo[14463:14448]},
     {storeUnit_maskInput_lo[14447:14432]},
     {storeUnit_maskInput_lo[14431:14416]},
     {storeUnit_maskInput_lo[14415:14400]},
     {storeUnit_maskInput_lo[14399:14384]},
     {storeUnit_maskInput_lo[14383:14368]},
     {storeUnit_maskInput_lo[14367:14352]},
     {storeUnit_maskInput_lo[14351:14336]},
     {storeUnit_maskInput_lo[14335:14320]},
     {storeUnit_maskInput_lo[14319:14304]},
     {storeUnit_maskInput_lo[14303:14288]},
     {storeUnit_maskInput_lo[14287:14272]},
     {storeUnit_maskInput_lo[14271:14256]},
     {storeUnit_maskInput_lo[14255:14240]},
     {storeUnit_maskInput_lo[14239:14224]},
     {storeUnit_maskInput_lo[14223:14208]},
     {storeUnit_maskInput_lo[14207:14192]},
     {storeUnit_maskInput_lo[14191:14176]},
     {storeUnit_maskInput_lo[14175:14160]},
     {storeUnit_maskInput_lo[14159:14144]},
     {storeUnit_maskInput_lo[14143:14128]},
     {storeUnit_maskInput_lo[14127:14112]},
     {storeUnit_maskInput_lo[14111:14096]},
     {storeUnit_maskInput_lo[14095:14080]},
     {storeUnit_maskInput_lo[14079:14064]},
     {storeUnit_maskInput_lo[14063:14048]},
     {storeUnit_maskInput_lo[14047:14032]},
     {storeUnit_maskInput_lo[14031:14016]},
     {storeUnit_maskInput_lo[14015:14000]},
     {storeUnit_maskInput_lo[13999:13984]},
     {storeUnit_maskInput_lo[13983:13968]},
     {storeUnit_maskInput_lo[13967:13952]},
     {storeUnit_maskInput_lo[13951:13936]},
     {storeUnit_maskInput_lo[13935:13920]},
     {storeUnit_maskInput_lo[13919:13904]},
     {storeUnit_maskInput_lo[13903:13888]},
     {storeUnit_maskInput_lo[13887:13872]},
     {storeUnit_maskInput_lo[13871:13856]},
     {storeUnit_maskInput_lo[13855:13840]},
     {storeUnit_maskInput_lo[13839:13824]},
     {storeUnit_maskInput_lo[13823:13808]},
     {storeUnit_maskInput_lo[13807:13792]},
     {storeUnit_maskInput_lo[13791:13776]},
     {storeUnit_maskInput_lo[13775:13760]},
     {storeUnit_maskInput_lo[13759:13744]},
     {storeUnit_maskInput_lo[13743:13728]},
     {storeUnit_maskInput_lo[13727:13712]},
     {storeUnit_maskInput_lo[13711:13696]},
     {storeUnit_maskInput_lo[13695:13680]},
     {storeUnit_maskInput_lo[13679:13664]},
     {storeUnit_maskInput_lo[13663:13648]},
     {storeUnit_maskInput_lo[13647:13632]},
     {storeUnit_maskInput_lo[13631:13616]},
     {storeUnit_maskInput_lo[13615:13600]},
     {storeUnit_maskInput_lo[13599:13584]},
     {storeUnit_maskInput_lo[13583:13568]},
     {storeUnit_maskInput_lo[13567:13552]},
     {storeUnit_maskInput_lo[13551:13536]},
     {storeUnit_maskInput_lo[13535:13520]},
     {storeUnit_maskInput_lo[13519:13504]},
     {storeUnit_maskInput_lo[13503:13488]},
     {storeUnit_maskInput_lo[13487:13472]},
     {storeUnit_maskInput_lo[13471:13456]},
     {storeUnit_maskInput_lo[13455:13440]},
     {storeUnit_maskInput_lo[13439:13424]},
     {storeUnit_maskInput_lo[13423:13408]},
     {storeUnit_maskInput_lo[13407:13392]},
     {storeUnit_maskInput_lo[13391:13376]},
     {storeUnit_maskInput_lo[13375:13360]},
     {storeUnit_maskInput_lo[13359:13344]},
     {storeUnit_maskInput_lo[13343:13328]},
     {storeUnit_maskInput_lo[13327:13312]},
     {storeUnit_maskInput_lo[13311:13296]},
     {storeUnit_maskInput_lo[13295:13280]},
     {storeUnit_maskInput_lo[13279:13264]},
     {storeUnit_maskInput_lo[13263:13248]},
     {storeUnit_maskInput_lo[13247:13232]},
     {storeUnit_maskInput_lo[13231:13216]},
     {storeUnit_maskInput_lo[13215:13200]},
     {storeUnit_maskInput_lo[13199:13184]},
     {storeUnit_maskInput_lo[13183:13168]},
     {storeUnit_maskInput_lo[13167:13152]},
     {storeUnit_maskInput_lo[13151:13136]},
     {storeUnit_maskInput_lo[13135:13120]},
     {storeUnit_maskInput_lo[13119:13104]},
     {storeUnit_maskInput_lo[13103:13088]},
     {storeUnit_maskInput_lo[13087:13072]},
     {storeUnit_maskInput_lo[13071:13056]},
     {storeUnit_maskInput_lo[13055:13040]},
     {storeUnit_maskInput_lo[13039:13024]},
     {storeUnit_maskInput_lo[13023:13008]},
     {storeUnit_maskInput_lo[13007:12992]},
     {storeUnit_maskInput_lo[12991:12976]},
     {storeUnit_maskInput_lo[12975:12960]},
     {storeUnit_maskInput_lo[12959:12944]},
     {storeUnit_maskInput_lo[12943:12928]},
     {storeUnit_maskInput_lo[12927:12912]},
     {storeUnit_maskInput_lo[12911:12896]},
     {storeUnit_maskInput_lo[12895:12880]},
     {storeUnit_maskInput_lo[12879:12864]},
     {storeUnit_maskInput_lo[12863:12848]},
     {storeUnit_maskInput_lo[12847:12832]},
     {storeUnit_maskInput_lo[12831:12816]},
     {storeUnit_maskInput_lo[12815:12800]},
     {storeUnit_maskInput_lo[12799:12784]},
     {storeUnit_maskInput_lo[12783:12768]},
     {storeUnit_maskInput_lo[12767:12752]},
     {storeUnit_maskInput_lo[12751:12736]},
     {storeUnit_maskInput_lo[12735:12720]},
     {storeUnit_maskInput_lo[12719:12704]},
     {storeUnit_maskInput_lo[12703:12688]},
     {storeUnit_maskInput_lo[12687:12672]},
     {storeUnit_maskInput_lo[12671:12656]},
     {storeUnit_maskInput_lo[12655:12640]},
     {storeUnit_maskInput_lo[12639:12624]},
     {storeUnit_maskInput_lo[12623:12608]},
     {storeUnit_maskInput_lo[12607:12592]},
     {storeUnit_maskInput_lo[12591:12576]},
     {storeUnit_maskInput_lo[12575:12560]},
     {storeUnit_maskInput_lo[12559:12544]},
     {storeUnit_maskInput_lo[12543:12528]},
     {storeUnit_maskInput_lo[12527:12512]},
     {storeUnit_maskInput_lo[12511:12496]},
     {storeUnit_maskInput_lo[12495:12480]},
     {storeUnit_maskInput_lo[12479:12464]},
     {storeUnit_maskInput_lo[12463:12448]},
     {storeUnit_maskInput_lo[12447:12432]},
     {storeUnit_maskInput_lo[12431:12416]},
     {storeUnit_maskInput_lo[12415:12400]},
     {storeUnit_maskInput_lo[12399:12384]},
     {storeUnit_maskInput_lo[12383:12368]},
     {storeUnit_maskInput_lo[12367:12352]},
     {storeUnit_maskInput_lo[12351:12336]},
     {storeUnit_maskInput_lo[12335:12320]},
     {storeUnit_maskInput_lo[12319:12304]},
     {storeUnit_maskInput_lo[12303:12288]},
     {storeUnit_maskInput_lo[12287:12272]},
     {storeUnit_maskInput_lo[12271:12256]},
     {storeUnit_maskInput_lo[12255:12240]},
     {storeUnit_maskInput_lo[12239:12224]},
     {storeUnit_maskInput_lo[12223:12208]},
     {storeUnit_maskInput_lo[12207:12192]},
     {storeUnit_maskInput_lo[12191:12176]},
     {storeUnit_maskInput_lo[12175:12160]},
     {storeUnit_maskInput_lo[12159:12144]},
     {storeUnit_maskInput_lo[12143:12128]},
     {storeUnit_maskInput_lo[12127:12112]},
     {storeUnit_maskInput_lo[12111:12096]},
     {storeUnit_maskInput_lo[12095:12080]},
     {storeUnit_maskInput_lo[12079:12064]},
     {storeUnit_maskInput_lo[12063:12048]},
     {storeUnit_maskInput_lo[12047:12032]},
     {storeUnit_maskInput_lo[12031:12016]},
     {storeUnit_maskInput_lo[12015:12000]},
     {storeUnit_maskInput_lo[11999:11984]},
     {storeUnit_maskInput_lo[11983:11968]},
     {storeUnit_maskInput_lo[11967:11952]},
     {storeUnit_maskInput_lo[11951:11936]},
     {storeUnit_maskInput_lo[11935:11920]},
     {storeUnit_maskInput_lo[11919:11904]},
     {storeUnit_maskInput_lo[11903:11888]},
     {storeUnit_maskInput_lo[11887:11872]},
     {storeUnit_maskInput_lo[11871:11856]},
     {storeUnit_maskInput_lo[11855:11840]},
     {storeUnit_maskInput_lo[11839:11824]},
     {storeUnit_maskInput_lo[11823:11808]},
     {storeUnit_maskInput_lo[11807:11792]},
     {storeUnit_maskInput_lo[11791:11776]},
     {storeUnit_maskInput_lo[11775:11760]},
     {storeUnit_maskInput_lo[11759:11744]},
     {storeUnit_maskInput_lo[11743:11728]},
     {storeUnit_maskInput_lo[11727:11712]},
     {storeUnit_maskInput_lo[11711:11696]},
     {storeUnit_maskInput_lo[11695:11680]},
     {storeUnit_maskInput_lo[11679:11664]},
     {storeUnit_maskInput_lo[11663:11648]},
     {storeUnit_maskInput_lo[11647:11632]},
     {storeUnit_maskInput_lo[11631:11616]},
     {storeUnit_maskInput_lo[11615:11600]},
     {storeUnit_maskInput_lo[11599:11584]},
     {storeUnit_maskInput_lo[11583:11568]},
     {storeUnit_maskInput_lo[11567:11552]},
     {storeUnit_maskInput_lo[11551:11536]},
     {storeUnit_maskInput_lo[11535:11520]},
     {storeUnit_maskInput_lo[11519:11504]},
     {storeUnit_maskInput_lo[11503:11488]},
     {storeUnit_maskInput_lo[11487:11472]},
     {storeUnit_maskInput_lo[11471:11456]},
     {storeUnit_maskInput_lo[11455:11440]},
     {storeUnit_maskInput_lo[11439:11424]},
     {storeUnit_maskInput_lo[11423:11408]},
     {storeUnit_maskInput_lo[11407:11392]},
     {storeUnit_maskInput_lo[11391:11376]},
     {storeUnit_maskInput_lo[11375:11360]},
     {storeUnit_maskInput_lo[11359:11344]},
     {storeUnit_maskInput_lo[11343:11328]},
     {storeUnit_maskInput_lo[11327:11312]},
     {storeUnit_maskInput_lo[11311:11296]},
     {storeUnit_maskInput_lo[11295:11280]},
     {storeUnit_maskInput_lo[11279:11264]},
     {storeUnit_maskInput_lo[11263:11248]},
     {storeUnit_maskInput_lo[11247:11232]},
     {storeUnit_maskInput_lo[11231:11216]},
     {storeUnit_maskInput_lo[11215:11200]},
     {storeUnit_maskInput_lo[11199:11184]},
     {storeUnit_maskInput_lo[11183:11168]},
     {storeUnit_maskInput_lo[11167:11152]},
     {storeUnit_maskInput_lo[11151:11136]},
     {storeUnit_maskInput_lo[11135:11120]},
     {storeUnit_maskInput_lo[11119:11104]},
     {storeUnit_maskInput_lo[11103:11088]},
     {storeUnit_maskInput_lo[11087:11072]},
     {storeUnit_maskInput_lo[11071:11056]},
     {storeUnit_maskInput_lo[11055:11040]},
     {storeUnit_maskInput_lo[11039:11024]},
     {storeUnit_maskInput_lo[11023:11008]},
     {storeUnit_maskInput_lo[11007:10992]},
     {storeUnit_maskInput_lo[10991:10976]},
     {storeUnit_maskInput_lo[10975:10960]},
     {storeUnit_maskInput_lo[10959:10944]},
     {storeUnit_maskInput_lo[10943:10928]},
     {storeUnit_maskInput_lo[10927:10912]},
     {storeUnit_maskInput_lo[10911:10896]},
     {storeUnit_maskInput_lo[10895:10880]},
     {storeUnit_maskInput_lo[10879:10864]},
     {storeUnit_maskInput_lo[10863:10848]},
     {storeUnit_maskInput_lo[10847:10832]},
     {storeUnit_maskInput_lo[10831:10816]},
     {storeUnit_maskInput_lo[10815:10800]},
     {storeUnit_maskInput_lo[10799:10784]},
     {storeUnit_maskInput_lo[10783:10768]},
     {storeUnit_maskInput_lo[10767:10752]},
     {storeUnit_maskInput_lo[10751:10736]},
     {storeUnit_maskInput_lo[10735:10720]},
     {storeUnit_maskInput_lo[10719:10704]},
     {storeUnit_maskInput_lo[10703:10688]},
     {storeUnit_maskInput_lo[10687:10672]},
     {storeUnit_maskInput_lo[10671:10656]},
     {storeUnit_maskInput_lo[10655:10640]},
     {storeUnit_maskInput_lo[10639:10624]},
     {storeUnit_maskInput_lo[10623:10608]},
     {storeUnit_maskInput_lo[10607:10592]},
     {storeUnit_maskInput_lo[10591:10576]},
     {storeUnit_maskInput_lo[10575:10560]},
     {storeUnit_maskInput_lo[10559:10544]},
     {storeUnit_maskInput_lo[10543:10528]},
     {storeUnit_maskInput_lo[10527:10512]},
     {storeUnit_maskInput_lo[10511:10496]},
     {storeUnit_maskInput_lo[10495:10480]},
     {storeUnit_maskInput_lo[10479:10464]},
     {storeUnit_maskInput_lo[10463:10448]},
     {storeUnit_maskInput_lo[10447:10432]},
     {storeUnit_maskInput_lo[10431:10416]},
     {storeUnit_maskInput_lo[10415:10400]},
     {storeUnit_maskInput_lo[10399:10384]},
     {storeUnit_maskInput_lo[10383:10368]},
     {storeUnit_maskInput_lo[10367:10352]},
     {storeUnit_maskInput_lo[10351:10336]},
     {storeUnit_maskInput_lo[10335:10320]},
     {storeUnit_maskInput_lo[10319:10304]},
     {storeUnit_maskInput_lo[10303:10288]},
     {storeUnit_maskInput_lo[10287:10272]},
     {storeUnit_maskInput_lo[10271:10256]},
     {storeUnit_maskInput_lo[10255:10240]},
     {storeUnit_maskInput_lo[10239:10224]},
     {storeUnit_maskInput_lo[10223:10208]},
     {storeUnit_maskInput_lo[10207:10192]},
     {storeUnit_maskInput_lo[10191:10176]},
     {storeUnit_maskInput_lo[10175:10160]},
     {storeUnit_maskInput_lo[10159:10144]},
     {storeUnit_maskInput_lo[10143:10128]},
     {storeUnit_maskInput_lo[10127:10112]},
     {storeUnit_maskInput_lo[10111:10096]},
     {storeUnit_maskInput_lo[10095:10080]},
     {storeUnit_maskInput_lo[10079:10064]},
     {storeUnit_maskInput_lo[10063:10048]},
     {storeUnit_maskInput_lo[10047:10032]},
     {storeUnit_maskInput_lo[10031:10016]},
     {storeUnit_maskInput_lo[10015:10000]},
     {storeUnit_maskInput_lo[9999:9984]},
     {storeUnit_maskInput_lo[9983:9968]},
     {storeUnit_maskInput_lo[9967:9952]},
     {storeUnit_maskInput_lo[9951:9936]},
     {storeUnit_maskInput_lo[9935:9920]},
     {storeUnit_maskInput_lo[9919:9904]},
     {storeUnit_maskInput_lo[9903:9888]},
     {storeUnit_maskInput_lo[9887:9872]},
     {storeUnit_maskInput_lo[9871:9856]},
     {storeUnit_maskInput_lo[9855:9840]},
     {storeUnit_maskInput_lo[9839:9824]},
     {storeUnit_maskInput_lo[9823:9808]},
     {storeUnit_maskInput_lo[9807:9792]},
     {storeUnit_maskInput_lo[9791:9776]},
     {storeUnit_maskInput_lo[9775:9760]},
     {storeUnit_maskInput_lo[9759:9744]},
     {storeUnit_maskInput_lo[9743:9728]},
     {storeUnit_maskInput_lo[9727:9712]},
     {storeUnit_maskInput_lo[9711:9696]},
     {storeUnit_maskInput_lo[9695:9680]},
     {storeUnit_maskInput_lo[9679:9664]},
     {storeUnit_maskInput_lo[9663:9648]},
     {storeUnit_maskInput_lo[9647:9632]},
     {storeUnit_maskInput_lo[9631:9616]},
     {storeUnit_maskInput_lo[9615:9600]},
     {storeUnit_maskInput_lo[9599:9584]},
     {storeUnit_maskInput_lo[9583:9568]},
     {storeUnit_maskInput_lo[9567:9552]},
     {storeUnit_maskInput_lo[9551:9536]},
     {storeUnit_maskInput_lo[9535:9520]},
     {storeUnit_maskInput_lo[9519:9504]},
     {storeUnit_maskInput_lo[9503:9488]},
     {storeUnit_maskInput_lo[9487:9472]},
     {storeUnit_maskInput_lo[9471:9456]},
     {storeUnit_maskInput_lo[9455:9440]},
     {storeUnit_maskInput_lo[9439:9424]},
     {storeUnit_maskInput_lo[9423:9408]},
     {storeUnit_maskInput_lo[9407:9392]},
     {storeUnit_maskInput_lo[9391:9376]},
     {storeUnit_maskInput_lo[9375:9360]},
     {storeUnit_maskInput_lo[9359:9344]},
     {storeUnit_maskInput_lo[9343:9328]},
     {storeUnit_maskInput_lo[9327:9312]},
     {storeUnit_maskInput_lo[9311:9296]},
     {storeUnit_maskInput_lo[9295:9280]},
     {storeUnit_maskInput_lo[9279:9264]},
     {storeUnit_maskInput_lo[9263:9248]},
     {storeUnit_maskInput_lo[9247:9232]},
     {storeUnit_maskInput_lo[9231:9216]},
     {storeUnit_maskInput_lo[9215:9200]},
     {storeUnit_maskInput_lo[9199:9184]},
     {storeUnit_maskInput_lo[9183:9168]},
     {storeUnit_maskInput_lo[9167:9152]},
     {storeUnit_maskInput_lo[9151:9136]},
     {storeUnit_maskInput_lo[9135:9120]},
     {storeUnit_maskInput_lo[9119:9104]},
     {storeUnit_maskInput_lo[9103:9088]},
     {storeUnit_maskInput_lo[9087:9072]},
     {storeUnit_maskInput_lo[9071:9056]},
     {storeUnit_maskInput_lo[9055:9040]},
     {storeUnit_maskInput_lo[9039:9024]},
     {storeUnit_maskInput_lo[9023:9008]},
     {storeUnit_maskInput_lo[9007:8992]},
     {storeUnit_maskInput_lo[8991:8976]},
     {storeUnit_maskInput_lo[8975:8960]},
     {storeUnit_maskInput_lo[8959:8944]},
     {storeUnit_maskInput_lo[8943:8928]},
     {storeUnit_maskInput_lo[8927:8912]},
     {storeUnit_maskInput_lo[8911:8896]},
     {storeUnit_maskInput_lo[8895:8880]},
     {storeUnit_maskInput_lo[8879:8864]},
     {storeUnit_maskInput_lo[8863:8848]},
     {storeUnit_maskInput_lo[8847:8832]},
     {storeUnit_maskInput_lo[8831:8816]},
     {storeUnit_maskInput_lo[8815:8800]},
     {storeUnit_maskInput_lo[8799:8784]},
     {storeUnit_maskInput_lo[8783:8768]},
     {storeUnit_maskInput_lo[8767:8752]},
     {storeUnit_maskInput_lo[8751:8736]},
     {storeUnit_maskInput_lo[8735:8720]},
     {storeUnit_maskInput_lo[8719:8704]},
     {storeUnit_maskInput_lo[8703:8688]},
     {storeUnit_maskInput_lo[8687:8672]},
     {storeUnit_maskInput_lo[8671:8656]},
     {storeUnit_maskInput_lo[8655:8640]},
     {storeUnit_maskInput_lo[8639:8624]},
     {storeUnit_maskInput_lo[8623:8608]},
     {storeUnit_maskInput_lo[8607:8592]},
     {storeUnit_maskInput_lo[8591:8576]},
     {storeUnit_maskInput_lo[8575:8560]},
     {storeUnit_maskInput_lo[8559:8544]},
     {storeUnit_maskInput_lo[8543:8528]},
     {storeUnit_maskInput_lo[8527:8512]},
     {storeUnit_maskInput_lo[8511:8496]},
     {storeUnit_maskInput_lo[8495:8480]},
     {storeUnit_maskInput_lo[8479:8464]},
     {storeUnit_maskInput_lo[8463:8448]},
     {storeUnit_maskInput_lo[8447:8432]},
     {storeUnit_maskInput_lo[8431:8416]},
     {storeUnit_maskInput_lo[8415:8400]},
     {storeUnit_maskInput_lo[8399:8384]},
     {storeUnit_maskInput_lo[8383:8368]},
     {storeUnit_maskInput_lo[8367:8352]},
     {storeUnit_maskInput_lo[8351:8336]},
     {storeUnit_maskInput_lo[8335:8320]},
     {storeUnit_maskInput_lo[8319:8304]},
     {storeUnit_maskInput_lo[8303:8288]},
     {storeUnit_maskInput_lo[8287:8272]},
     {storeUnit_maskInput_lo[8271:8256]},
     {storeUnit_maskInput_lo[8255:8240]},
     {storeUnit_maskInput_lo[8239:8224]},
     {storeUnit_maskInput_lo[8223:8208]},
     {storeUnit_maskInput_lo[8207:8192]},
     {storeUnit_maskInput_lo[8191:8176]},
     {storeUnit_maskInput_lo[8175:8160]},
     {storeUnit_maskInput_lo[8159:8144]},
     {storeUnit_maskInput_lo[8143:8128]},
     {storeUnit_maskInput_lo[8127:8112]},
     {storeUnit_maskInput_lo[8111:8096]},
     {storeUnit_maskInput_lo[8095:8080]},
     {storeUnit_maskInput_lo[8079:8064]},
     {storeUnit_maskInput_lo[8063:8048]},
     {storeUnit_maskInput_lo[8047:8032]},
     {storeUnit_maskInput_lo[8031:8016]},
     {storeUnit_maskInput_lo[8015:8000]},
     {storeUnit_maskInput_lo[7999:7984]},
     {storeUnit_maskInput_lo[7983:7968]},
     {storeUnit_maskInput_lo[7967:7952]},
     {storeUnit_maskInput_lo[7951:7936]},
     {storeUnit_maskInput_lo[7935:7920]},
     {storeUnit_maskInput_lo[7919:7904]},
     {storeUnit_maskInput_lo[7903:7888]},
     {storeUnit_maskInput_lo[7887:7872]},
     {storeUnit_maskInput_lo[7871:7856]},
     {storeUnit_maskInput_lo[7855:7840]},
     {storeUnit_maskInput_lo[7839:7824]},
     {storeUnit_maskInput_lo[7823:7808]},
     {storeUnit_maskInput_lo[7807:7792]},
     {storeUnit_maskInput_lo[7791:7776]},
     {storeUnit_maskInput_lo[7775:7760]},
     {storeUnit_maskInput_lo[7759:7744]},
     {storeUnit_maskInput_lo[7743:7728]},
     {storeUnit_maskInput_lo[7727:7712]},
     {storeUnit_maskInput_lo[7711:7696]},
     {storeUnit_maskInput_lo[7695:7680]},
     {storeUnit_maskInput_lo[7679:7664]},
     {storeUnit_maskInput_lo[7663:7648]},
     {storeUnit_maskInput_lo[7647:7632]},
     {storeUnit_maskInput_lo[7631:7616]},
     {storeUnit_maskInput_lo[7615:7600]},
     {storeUnit_maskInput_lo[7599:7584]},
     {storeUnit_maskInput_lo[7583:7568]},
     {storeUnit_maskInput_lo[7567:7552]},
     {storeUnit_maskInput_lo[7551:7536]},
     {storeUnit_maskInput_lo[7535:7520]},
     {storeUnit_maskInput_lo[7519:7504]},
     {storeUnit_maskInput_lo[7503:7488]},
     {storeUnit_maskInput_lo[7487:7472]},
     {storeUnit_maskInput_lo[7471:7456]},
     {storeUnit_maskInput_lo[7455:7440]},
     {storeUnit_maskInput_lo[7439:7424]},
     {storeUnit_maskInput_lo[7423:7408]},
     {storeUnit_maskInput_lo[7407:7392]},
     {storeUnit_maskInput_lo[7391:7376]},
     {storeUnit_maskInput_lo[7375:7360]},
     {storeUnit_maskInput_lo[7359:7344]},
     {storeUnit_maskInput_lo[7343:7328]},
     {storeUnit_maskInput_lo[7327:7312]},
     {storeUnit_maskInput_lo[7311:7296]},
     {storeUnit_maskInput_lo[7295:7280]},
     {storeUnit_maskInput_lo[7279:7264]},
     {storeUnit_maskInput_lo[7263:7248]},
     {storeUnit_maskInput_lo[7247:7232]},
     {storeUnit_maskInput_lo[7231:7216]},
     {storeUnit_maskInput_lo[7215:7200]},
     {storeUnit_maskInput_lo[7199:7184]},
     {storeUnit_maskInput_lo[7183:7168]},
     {storeUnit_maskInput_lo[7167:7152]},
     {storeUnit_maskInput_lo[7151:7136]},
     {storeUnit_maskInput_lo[7135:7120]},
     {storeUnit_maskInput_lo[7119:7104]},
     {storeUnit_maskInput_lo[7103:7088]},
     {storeUnit_maskInput_lo[7087:7072]},
     {storeUnit_maskInput_lo[7071:7056]},
     {storeUnit_maskInput_lo[7055:7040]},
     {storeUnit_maskInput_lo[7039:7024]},
     {storeUnit_maskInput_lo[7023:7008]},
     {storeUnit_maskInput_lo[7007:6992]},
     {storeUnit_maskInput_lo[6991:6976]},
     {storeUnit_maskInput_lo[6975:6960]},
     {storeUnit_maskInput_lo[6959:6944]},
     {storeUnit_maskInput_lo[6943:6928]},
     {storeUnit_maskInput_lo[6927:6912]},
     {storeUnit_maskInput_lo[6911:6896]},
     {storeUnit_maskInput_lo[6895:6880]},
     {storeUnit_maskInput_lo[6879:6864]},
     {storeUnit_maskInput_lo[6863:6848]},
     {storeUnit_maskInput_lo[6847:6832]},
     {storeUnit_maskInput_lo[6831:6816]},
     {storeUnit_maskInput_lo[6815:6800]},
     {storeUnit_maskInput_lo[6799:6784]},
     {storeUnit_maskInput_lo[6783:6768]},
     {storeUnit_maskInput_lo[6767:6752]},
     {storeUnit_maskInput_lo[6751:6736]},
     {storeUnit_maskInput_lo[6735:6720]},
     {storeUnit_maskInput_lo[6719:6704]},
     {storeUnit_maskInput_lo[6703:6688]},
     {storeUnit_maskInput_lo[6687:6672]},
     {storeUnit_maskInput_lo[6671:6656]},
     {storeUnit_maskInput_lo[6655:6640]},
     {storeUnit_maskInput_lo[6639:6624]},
     {storeUnit_maskInput_lo[6623:6608]},
     {storeUnit_maskInput_lo[6607:6592]},
     {storeUnit_maskInput_lo[6591:6576]},
     {storeUnit_maskInput_lo[6575:6560]},
     {storeUnit_maskInput_lo[6559:6544]},
     {storeUnit_maskInput_lo[6543:6528]},
     {storeUnit_maskInput_lo[6527:6512]},
     {storeUnit_maskInput_lo[6511:6496]},
     {storeUnit_maskInput_lo[6495:6480]},
     {storeUnit_maskInput_lo[6479:6464]},
     {storeUnit_maskInput_lo[6463:6448]},
     {storeUnit_maskInput_lo[6447:6432]},
     {storeUnit_maskInput_lo[6431:6416]},
     {storeUnit_maskInput_lo[6415:6400]},
     {storeUnit_maskInput_lo[6399:6384]},
     {storeUnit_maskInput_lo[6383:6368]},
     {storeUnit_maskInput_lo[6367:6352]},
     {storeUnit_maskInput_lo[6351:6336]},
     {storeUnit_maskInput_lo[6335:6320]},
     {storeUnit_maskInput_lo[6319:6304]},
     {storeUnit_maskInput_lo[6303:6288]},
     {storeUnit_maskInput_lo[6287:6272]},
     {storeUnit_maskInput_lo[6271:6256]},
     {storeUnit_maskInput_lo[6255:6240]},
     {storeUnit_maskInput_lo[6239:6224]},
     {storeUnit_maskInput_lo[6223:6208]},
     {storeUnit_maskInput_lo[6207:6192]},
     {storeUnit_maskInput_lo[6191:6176]},
     {storeUnit_maskInput_lo[6175:6160]},
     {storeUnit_maskInput_lo[6159:6144]},
     {storeUnit_maskInput_lo[6143:6128]},
     {storeUnit_maskInput_lo[6127:6112]},
     {storeUnit_maskInput_lo[6111:6096]},
     {storeUnit_maskInput_lo[6095:6080]},
     {storeUnit_maskInput_lo[6079:6064]},
     {storeUnit_maskInput_lo[6063:6048]},
     {storeUnit_maskInput_lo[6047:6032]},
     {storeUnit_maskInput_lo[6031:6016]},
     {storeUnit_maskInput_lo[6015:6000]},
     {storeUnit_maskInput_lo[5999:5984]},
     {storeUnit_maskInput_lo[5983:5968]},
     {storeUnit_maskInput_lo[5967:5952]},
     {storeUnit_maskInput_lo[5951:5936]},
     {storeUnit_maskInput_lo[5935:5920]},
     {storeUnit_maskInput_lo[5919:5904]},
     {storeUnit_maskInput_lo[5903:5888]},
     {storeUnit_maskInput_lo[5887:5872]},
     {storeUnit_maskInput_lo[5871:5856]},
     {storeUnit_maskInput_lo[5855:5840]},
     {storeUnit_maskInput_lo[5839:5824]},
     {storeUnit_maskInput_lo[5823:5808]},
     {storeUnit_maskInput_lo[5807:5792]},
     {storeUnit_maskInput_lo[5791:5776]},
     {storeUnit_maskInput_lo[5775:5760]},
     {storeUnit_maskInput_lo[5759:5744]},
     {storeUnit_maskInput_lo[5743:5728]},
     {storeUnit_maskInput_lo[5727:5712]},
     {storeUnit_maskInput_lo[5711:5696]},
     {storeUnit_maskInput_lo[5695:5680]},
     {storeUnit_maskInput_lo[5679:5664]},
     {storeUnit_maskInput_lo[5663:5648]},
     {storeUnit_maskInput_lo[5647:5632]},
     {storeUnit_maskInput_lo[5631:5616]},
     {storeUnit_maskInput_lo[5615:5600]},
     {storeUnit_maskInput_lo[5599:5584]},
     {storeUnit_maskInput_lo[5583:5568]},
     {storeUnit_maskInput_lo[5567:5552]},
     {storeUnit_maskInput_lo[5551:5536]},
     {storeUnit_maskInput_lo[5535:5520]},
     {storeUnit_maskInput_lo[5519:5504]},
     {storeUnit_maskInput_lo[5503:5488]},
     {storeUnit_maskInput_lo[5487:5472]},
     {storeUnit_maskInput_lo[5471:5456]},
     {storeUnit_maskInput_lo[5455:5440]},
     {storeUnit_maskInput_lo[5439:5424]},
     {storeUnit_maskInput_lo[5423:5408]},
     {storeUnit_maskInput_lo[5407:5392]},
     {storeUnit_maskInput_lo[5391:5376]},
     {storeUnit_maskInput_lo[5375:5360]},
     {storeUnit_maskInput_lo[5359:5344]},
     {storeUnit_maskInput_lo[5343:5328]},
     {storeUnit_maskInput_lo[5327:5312]},
     {storeUnit_maskInput_lo[5311:5296]},
     {storeUnit_maskInput_lo[5295:5280]},
     {storeUnit_maskInput_lo[5279:5264]},
     {storeUnit_maskInput_lo[5263:5248]},
     {storeUnit_maskInput_lo[5247:5232]},
     {storeUnit_maskInput_lo[5231:5216]},
     {storeUnit_maskInput_lo[5215:5200]},
     {storeUnit_maskInput_lo[5199:5184]},
     {storeUnit_maskInput_lo[5183:5168]},
     {storeUnit_maskInput_lo[5167:5152]},
     {storeUnit_maskInput_lo[5151:5136]},
     {storeUnit_maskInput_lo[5135:5120]},
     {storeUnit_maskInput_lo[5119:5104]},
     {storeUnit_maskInput_lo[5103:5088]},
     {storeUnit_maskInput_lo[5087:5072]},
     {storeUnit_maskInput_lo[5071:5056]},
     {storeUnit_maskInput_lo[5055:5040]},
     {storeUnit_maskInput_lo[5039:5024]},
     {storeUnit_maskInput_lo[5023:5008]},
     {storeUnit_maskInput_lo[5007:4992]},
     {storeUnit_maskInput_lo[4991:4976]},
     {storeUnit_maskInput_lo[4975:4960]},
     {storeUnit_maskInput_lo[4959:4944]},
     {storeUnit_maskInput_lo[4943:4928]},
     {storeUnit_maskInput_lo[4927:4912]},
     {storeUnit_maskInput_lo[4911:4896]},
     {storeUnit_maskInput_lo[4895:4880]},
     {storeUnit_maskInput_lo[4879:4864]},
     {storeUnit_maskInput_lo[4863:4848]},
     {storeUnit_maskInput_lo[4847:4832]},
     {storeUnit_maskInput_lo[4831:4816]},
     {storeUnit_maskInput_lo[4815:4800]},
     {storeUnit_maskInput_lo[4799:4784]},
     {storeUnit_maskInput_lo[4783:4768]},
     {storeUnit_maskInput_lo[4767:4752]},
     {storeUnit_maskInput_lo[4751:4736]},
     {storeUnit_maskInput_lo[4735:4720]},
     {storeUnit_maskInput_lo[4719:4704]},
     {storeUnit_maskInput_lo[4703:4688]},
     {storeUnit_maskInput_lo[4687:4672]},
     {storeUnit_maskInput_lo[4671:4656]},
     {storeUnit_maskInput_lo[4655:4640]},
     {storeUnit_maskInput_lo[4639:4624]},
     {storeUnit_maskInput_lo[4623:4608]},
     {storeUnit_maskInput_lo[4607:4592]},
     {storeUnit_maskInput_lo[4591:4576]},
     {storeUnit_maskInput_lo[4575:4560]},
     {storeUnit_maskInput_lo[4559:4544]},
     {storeUnit_maskInput_lo[4543:4528]},
     {storeUnit_maskInput_lo[4527:4512]},
     {storeUnit_maskInput_lo[4511:4496]},
     {storeUnit_maskInput_lo[4495:4480]},
     {storeUnit_maskInput_lo[4479:4464]},
     {storeUnit_maskInput_lo[4463:4448]},
     {storeUnit_maskInput_lo[4447:4432]},
     {storeUnit_maskInput_lo[4431:4416]},
     {storeUnit_maskInput_lo[4415:4400]},
     {storeUnit_maskInput_lo[4399:4384]},
     {storeUnit_maskInput_lo[4383:4368]},
     {storeUnit_maskInput_lo[4367:4352]},
     {storeUnit_maskInput_lo[4351:4336]},
     {storeUnit_maskInput_lo[4335:4320]},
     {storeUnit_maskInput_lo[4319:4304]},
     {storeUnit_maskInput_lo[4303:4288]},
     {storeUnit_maskInput_lo[4287:4272]},
     {storeUnit_maskInput_lo[4271:4256]},
     {storeUnit_maskInput_lo[4255:4240]},
     {storeUnit_maskInput_lo[4239:4224]},
     {storeUnit_maskInput_lo[4223:4208]},
     {storeUnit_maskInput_lo[4207:4192]},
     {storeUnit_maskInput_lo[4191:4176]},
     {storeUnit_maskInput_lo[4175:4160]},
     {storeUnit_maskInput_lo[4159:4144]},
     {storeUnit_maskInput_lo[4143:4128]},
     {storeUnit_maskInput_lo[4127:4112]},
     {storeUnit_maskInput_lo[4111:4096]},
     {storeUnit_maskInput_lo[4095:4080]},
     {storeUnit_maskInput_lo[4079:4064]},
     {storeUnit_maskInput_lo[4063:4048]},
     {storeUnit_maskInput_lo[4047:4032]},
     {storeUnit_maskInput_lo[4031:4016]},
     {storeUnit_maskInput_lo[4015:4000]},
     {storeUnit_maskInput_lo[3999:3984]},
     {storeUnit_maskInput_lo[3983:3968]},
     {storeUnit_maskInput_lo[3967:3952]},
     {storeUnit_maskInput_lo[3951:3936]},
     {storeUnit_maskInput_lo[3935:3920]},
     {storeUnit_maskInput_lo[3919:3904]},
     {storeUnit_maskInput_lo[3903:3888]},
     {storeUnit_maskInput_lo[3887:3872]},
     {storeUnit_maskInput_lo[3871:3856]},
     {storeUnit_maskInput_lo[3855:3840]},
     {storeUnit_maskInput_lo[3839:3824]},
     {storeUnit_maskInput_lo[3823:3808]},
     {storeUnit_maskInput_lo[3807:3792]},
     {storeUnit_maskInput_lo[3791:3776]},
     {storeUnit_maskInput_lo[3775:3760]},
     {storeUnit_maskInput_lo[3759:3744]},
     {storeUnit_maskInput_lo[3743:3728]},
     {storeUnit_maskInput_lo[3727:3712]},
     {storeUnit_maskInput_lo[3711:3696]},
     {storeUnit_maskInput_lo[3695:3680]},
     {storeUnit_maskInput_lo[3679:3664]},
     {storeUnit_maskInput_lo[3663:3648]},
     {storeUnit_maskInput_lo[3647:3632]},
     {storeUnit_maskInput_lo[3631:3616]},
     {storeUnit_maskInput_lo[3615:3600]},
     {storeUnit_maskInput_lo[3599:3584]},
     {storeUnit_maskInput_lo[3583:3568]},
     {storeUnit_maskInput_lo[3567:3552]},
     {storeUnit_maskInput_lo[3551:3536]},
     {storeUnit_maskInput_lo[3535:3520]},
     {storeUnit_maskInput_lo[3519:3504]},
     {storeUnit_maskInput_lo[3503:3488]},
     {storeUnit_maskInput_lo[3487:3472]},
     {storeUnit_maskInput_lo[3471:3456]},
     {storeUnit_maskInput_lo[3455:3440]},
     {storeUnit_maskInput_lo[3439:3424]},
     {storeUnit_maskInput_lo[3423:3408]},
     {storeUnit_maskInput_lo[3407:3392]},
     {storeUnit_maskInput_lo[3391:3376]},
     {storeUnit_maskInput_lo[3375:3360]},
     {storeUnit_maskInput_lo[3359:3344]},
     {storeUnit_maskInput_lo[3343:3328]},
     {storeUnit_maskInput_lo[3327:3312]},
     {storeUnit_maskInput_lo[3311:3296]},
     {storeUnit_maskInput_lo[3295:3280]},
     {storeUnit_maskInput_lo[3279:3264]},
     {storeUnit_maskInput_lo[3263:3248]},
     {storeUnit_maskInput_lo[3247:3232]},
     {storeUnit_maskInput_lo[3231:3216]},
     {storeUnit_maskInput_lo[3215:3200]},
     {storeUnit_maskInput_lo[3199:3184]},
     {storeUnit_maskInput_lo[3183:3168]},
     {storeUnit_maskInput_lo[3167:3152]},
     {storeUnit_maskInput_lo[3151:3136]},
     {storeUnit_maskInput_lo[3135:3120]},
     {storeUnit_maskInput_lo[3119:3104]},
     {storeUnit_maskInput_lo[3103:3088]},
     {storeUnit_maskInput_lo[3087:3072]},
     {storeUnit_maskInput_lo[3071:3056]},
     {storeUnit_maskInput_lo[3055:3040]},
     {storeUnit_maskInput_lo[3039:3024]},
     {storeUnit_maskInput_lo[3023:3008]},
     {storeUnit_maskInput_lo[3007:2992]},
     {storeUnit_maskInput_lo[2991:2976]},
     {storeUnit_maskInput_lo[2975:2960]},
     {storeUnit_maskInput_lo[2959:2944]},
     {storeUnit_maskInput_lo[2943:2928]},
     {storeUnit_maskInput_lo[2927:2912]},
     {storeUnit_maskInput_lo[2911:2896]},
     {storeUnit_maskInput_lo[2895:2880]},
     {storeUnit_maskInput_lo[2879:2864]},
     {storeUnit_maskInput_lo[2863:2848]},
     {storeUnit_maskInput_lo[2847:2832]},
     {storeUnit_maskInput_lo[2831:2816]},
     {storeUnit_maskInput_lo[2815:2800]},
     {storeUnit_maskInput_lo[2799:2784]},
     {storeUnit_maskInput_lo[2783:2768]},
     {storeUnit_maskInput_lo[2767:2752]},
     {storeUnit_maskInput_lo[2751:2736]},
     {storeUnit_maskInput_lo[2735:2720]},
     {storeUnit_maskInput_lo[2719:2704]},
     {storeUnit_maskInput_lo[2703:2688]},
     {storeUnit_maskInput_lo[2687:2672]},
     {storeUnit_maskInput_lo[2671:2656]},
     {storeUnit_maskInput_lo[2655:2640]},
     {storeUnit_maskInput_lo[2639:2624]},
     {storeUnit_maskInput_lo[2623:2608]},
     {storeUnit_maskInput_lo[2607:2592]},
     {storeUnit_maskInput_lo[2591:2576]},
     {storeUnit_maskInput_lo[2575:2560]},
     {storeUnit_maskInput_lo[2559:2544]},
     {storeUnit_maskInput_lo[2543:2528]},
     {storeUnit_maskInput_lo[2527:2512]},
     {storeUnit_maskInput_lo[2511:2496]},
     {storeUnit_maskInput_lo[2495:2480]},
     {storeUnit_maskInput_lo[2479:2464]},
     {storeUnit_maskInput_lo[2463:2448]},
     {storeUnit_maskInput_lo[2447:2432]},
     {storeUnit_maskInput_lo[2431:2416]},
     {storeUnit_maskInput_lo[2415:2400]},
     {storeUnit_maskInput_lo[2399:2384]},
     {storeUnit_maskInput_lo[2383:2368]},
     {storeUnit_maskInput_lo[2367:2352]},
     {storeUnit_maskInput_lo[2351:2336]},
     {storeUnit_maskInput_lo[2335:2320]},
     {storeUnit_maskInput_lo[2319:2304]},
     {storeUnit_maskInput_lo[2303:2288]},
     {storeUnit_maskInput_lo[2287:2272]},
     {storeUnit_maskInput_lo[2271:2256]},
     {storeUnit_maskInput_lo[2255:2240]},
     {storeUnit_maskInput_lo[2239:2224]},
     {storeUnit_maskInput_lo[2223:2208]},
     {storeUnit_maskInput_lo[2207:2192]},
     {storeUnit_maskInput_lo[2191:2176]},
     {storeUnit_maskInput_lo[2175:2160]},
     {storeUnit_maskInput_lo[2159:2144]},
     {storeUnit_maskInput_lo[2143:2128]},
     {storeUnit_maskInput_lo[2127:2112]},
     {storeUnit_maskInput_lo[2111:2096]},
     {storeUnit_maskInput_lo[2095:2080]},
     {storeUnit_maskInput_lo[2079:2064]},
     {storeUnit_maskInput_lo[2063:2048]},
     {storeUnit_maskInput_lo[2047:2032]},
     {storeUnit_maskInput_lo[2031:2016]},
     {storeUnit_maskInput_lo[2015:2000]},
     {storeUnit_maskInput_lo[1999:1984]},
     {storeUnit_maskInput_lo[1983:1968]},
     {storeUnit_maskInput_lo[1967:1952]},
     {storeUnit_maskInput_lo[1951:1936]},
     {storeUnit_maskInput_lo[1935:1920]},
     {storeUnit_maskInput_lo[1919:1904]},
     {storeUnit_maskInput_lo[1903:1888]},
     {storeUnit_maskInput_lo[1887:1872]},
     {storeUnit_maskInput_lo[1871:1856]},
     {storeUnit_maskInput_lo[1855:1840]},
     {storeUnit_maskInput_lo[1839:1824]},
     {storeUnit_maskInput_lo[1823:1808]},
     {storeUnit_maskInput_lo[1807:1792]},
     {storeUnit_maskInput_lo[1791:1776]},
     {storeUnit_maskInput_lo[1775:1760]},
     {storeUnit_maskInput_lo[1759:1744]},
     {storeUnit_maskInput_lo[1743:1728]},
     {storeUnit_maskInput_lo[1727:1712]},
     {storeUnit_maskInput_lo[1711:1696]},
     {storeUnit_maskInput_lo[1695:1680]},
     {storeUnit_maskInput_lo[1679:1664]},
     {storeUnit_maskInput_lo[1663:1648]},
     {storeUnit_maskInput_lo[1647:1632]},
     {storeUnit_maskInput_lo[1631:1616]},
     {storeUnit_maskInput_lo[1615:1600]},
     {storeUnit_maskInput_lo[1599:1584]},
     {storeUnit_maskInput_lo[1583:1568]},
     {storeUnit_maskInput_lo[1567:1552]},
     {storeUnit_maskInput_lo[1551:1536]},
     {storeUnit_maskInput_lo[1535:1520]},
     {storeUnit_maskInput_lo[1519:1504]},
     {storeUnit_maskInput_lo[1503:1488]},
     {storeUnit_maskInput_lo[1487:1472]},
     {storeUnit_maskInput_lo[1471:1456]},
     {storeUnit_maskInput_lo[1455:1440]},
     {storeUnit_maskInput_lo[1439:1424]},
     {storeUnit_maskInput_lo[1423:1408]},
     {storeUnit_maskInput_lo[1407:1392]},
     {storeUnit_maskInput_lo[1391:1376]},
     {storeUnit_maskInput_lo[1375:1360]},
     {storeUnit_maskInput_lo[1359:1344]},
     {storeUnit_maskInput_lo[1343:1328]},
     {storeUnit_maskInput_lo[1327:1312]},
     {storeUnit_maskInput_lo[1311:1296]},
     {storeUnit_maskInput_lo[1295:1280]},
     {storeUnit_maskInput_lo[1279:1264]},
     {storeUnit_maskInput_lo[1263:1248]},
     {storeUnit_maskInput_lo[1247:1232]},
     {storeUnit_maskInput_lo[1231:1216]},
     {storeUnit_maskInput_lo[1215:1200]},
     {storeUnit_maskInput_lo[1199:1184]},
     {storeUnit_maskInput_lo[1183:1168]},
     {storeUnit_maskInput_lo[1167:1152]},
     {storeUnit_maskInput_lo[1151:1136]},
     {storeUnit_maskInput_lo[1135:1120]},
     {storeUnit_maskInput_lo[1119:1104]},
     {storeUnit_maskInput_lo[1103:1088]},
     {storeUnit_maskInput_lo[1087:1072]},
     {storeUnit_maskInput_lo[1071:1056]},
     {storeUnit_maskInput_lo[1055:1040]},
     {storeUnit_maskInput_lo[1039:1024]},
     {storeUnit_maskInput_lo[1023:1008]},
     {storeUnit_maskInput_lo[1007:992]},
     {storeUnit_maskInput_lo[991:976]},
     {storeUnit_maskInput_lo[975:960]},
     {storeUnit_maskInput_lo[959:944]},
     {storeUnit_maskInput_lo[943:928]},
     {storeUnit_maskInput_lo[927:912]},
     {storeUnit_maskInput_lo[911:896]},
     {storeUnit_maskInput_lo[895:880]},
     {storeUnit_maskInput_lo[879:864]},
     {storeUnit_maskInput_lo[863:848]},
     {storeUnit_maskInput_lo[847:832]},
     {storeUnit_maskInput_lo[831:816]},
     {storeUnit_maskInput_lo[815:800]},
     {storeUnit_maskInput_lo[799:784]},
     {storeUnit_maskInput_lo[783:768]},
     {storeUnit_maskInput_lo[767:752]},
     {storeUnit_maskInput_lo[751:736]},
     {storeUnit_maskInput_lo[735:720]},
     {storeUnit_maskInput_lo[719:704]},
     {storeUnit_maskInput_lo[703:688]},
     {storeUnit_maskInput_lo[687:672]},
     {storeUnit_maskInput_lo[671:656]},
     {storeUnit_maskInput_lo[655:640]},
     {storeUnit_maskInput_lo[639:624]},
     {storeUnit_maskInput_lo[623:608]},
     {storeUnit_maskInput_lo[607:592]},
     {storeUnit_maskInput_lo[591:576]},
     {storeUnit_maskInput_lo[575:560]},
     {storeUnit_maskInput_lo[559:544]},
     {storeUnit_maskInput_lo[543:528]},
     {storeUnit_maskInput_lo[527:512]},
     {storeUnit_maskInput_lo[511:496]},
     {storeUnit_maskInput_lo[495:480]},
     {storeUnit_maskInput_lo[479:464]},
     {storeUnit_maskInput_lo[463:448]},
     {storeUnit_maskInput_lo[447:432]},
     {storeUnit_maskInput_lo[431:416]},
     {storeUnit_maskInput_lo[415:400]},
     {storeUnit_maskInput_lo[399:384]},
     {storeUnit_maskInput_lo[383:368]},
     {storeUnit_maskInput_lo[367:352]},
     {storeUnit_maskInput_lo[351:336]},
     {storeUnit_maskInput_lo[335:320]},
     {storeUnit_maskInput_lo[319:304]},
     {storeUnit_maskInput_lo[303:288]},
     {storeUnit_maskInput_lo[287:272]},
     {storeUnit_maskInput_lo[271:256]},
     {storeUnit_maskInput_lo[255:240]},
     {storeUnit_maskInput_lo[239:224]},
     {storeUnit_maskInput_lo[223:208]},
     {storeUnit_maskInput_lo[207:192]},
     {storeUnit_maskInput_lo[191:176]},
     {storeUnit_maskInput_lo[175:160]},
     {storeUnit_maskInput_lo[159:144]},
     {storeUnit_maskInput_lo[143:128]},
     {storeUnit_maskInput_lo[127:112]},
     {storeUnit_maskInput_lo[111:96]},
     {storeUnit_maskInput_lo[95:80]},
     {storeUnit_maskInput_lo[79:64]},
     {storeUnit_maskInput_lo[63:48]},
     {storeUnit_maskInput_lo[47:32]},
     {storeUnit_maskInput_lo[31:16]},
     {storeUnit_maskInput_lo[15:0]}};
  wire [10:0]         maskSelect_2 = _otherUnit_maskSelect_valid ? _otherUnit_maskSelect_bits : 11'h0;
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_lo_lo = {otherUnit_maskInput_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_lo_hi_hi = {otherUnit_maskInput_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_lo_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_lo_hi = {otherUnit_maskInput_lo_lo_hi_hi, otherUnit_maskInput_lo_lo_hi_lo};
  wire [8191:0]       otherUnit_maskInput_lo_lo = {otherUnit_maskInput_lo_lo_hi, otherUnit_maskInput_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_hi_lo = {otherUnit_maskInput_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_lo_hi_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_lo_hi_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_lo_hi_hi = {otherUnit_maskInput_lo_hi_hi_hi, otherUnit_maskInput_lo_hi_hi_lo};
  wire [8191:0]       otherUnit_maskInput_lo_hi = {otherUnit_maskInput_lo_hi_hi, otherUnit_maskInput_lo_hi_lo};
  wire [16383:0]      otherUnit_maskInput_lo = {otherUnit_maskInput_lo_hi, otherUnit_maskInput_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_lo_lo = {otherUnit_maskInput_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_lo_hi_hi = {otherUnit_maskInput_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_lo_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_lo_hi = {otherUnit_maskInput_hi_lo_hi_hi, otherUnit_maskInput_hi_lo_hi_lo};
  wire [8191:0]       otherUnit_maskInput_hi_lo = {otherUnit_maskInput_hi_lo_hi, otherUnit_maskInput_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_lo_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_hi_lo = {otherUnit_maskInput_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_lo_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [127:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [255:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [511:0]        otherUnit_maskInput_hi_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_hi_lo};
  wire [1023:0]       otherUnit_maskInput_hi_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_hi_lo};
  wire [2047:0]       otherUnit_maskInput_hi_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_hi_lo};
  wire [4095:0]       otherUnit_maskInput_hi_hi_hi = {otherUnit_maskInput_hi_hi_hi_hi, otherUnit_maskInput_hi_hi_hi_lo};
  wire [8191:0]       otherUnit_maskInput_hi_hi = {otherUnit_maskInput_hi_hi_hi, otherUnit_maskInput_hi_hi_lo};
  wire [16383:0]      otherUnit_maskInput_hi = {otherUnit_maskInput_hi_hi, otherUnit_maskInput_hi_lo};
  wire [2047:0][15:0] _GEN_513 =
    {{otherUnit_maskInput_hi[16383:16368]},
     {otherUnit_maskInput_hi[16367:16352]},
     {otherUnit_maskInput_hi[16351:16336]},
     {otherUnit_maskInput_hi[16335:16320]},
     {otherUnit_maskInput_hi[16319:16304]},
     {otherUnit_maskInput_hi[16303:16288]},
     {otherUnit_maskInput_hi[16287:16272]},
     {otherUnit_maskInput_hi[16271:16256]},
     {otherUnit_maskInput_hi[16255:16240]},
     {otherUnit_maskInput_hi[16239:16224]},
     {otherUnit_maskInput_hi[16223:16208]},
     {otherUnit_maskInput_hi[16207:16192]},
     {otherUnit_maskInput_hi[16191:16176]},
     {otherUnit_maskInput_hi[16175:16160]},
     {otherUnit_maskInput_hi[16159:16144]},
     {otherUnit_maskInput_hi[16143:16128]},
     {otherUnit_maskInput_hi[16127:16112]},
     {otherUnit_maskInput_hi[16111:16096]},
     {otherUnit_maskInput_hi[16095:16080]},
     {otherUnit_maskInput_hi[16079:16064]},
     {otherUnit_maskInput_hi[16063:16048]},
     {otherUnit_maskInput_hi[16047:16032]},
     {otherUnit_maskInput_hi[16031:16016]},
     {otherUnit_maskInput_hi[16015:16000]},
     {otherUnit_maskInput_hi[15999:15984]},
     {otherUnit_maskInput_hi[15983:15968]},
     {otherUnit_maskInput_hi[15967:15952]},
     {otherUnit_maskInput_hi[15951:15936]},
     {otherUnit_maskInput_hi[15935:15920]},
     {otherUnit_maskInput_hi[15919:15904]},
     {otherUnit_maskInput_hi[15903:15888]},
     {otherUnit_maskInput_hi[15887:15872]},
     {otherUnit_maskInput_hi[15871:15856]},
     {otherUnit_maskInput_hi[15855:15840]},
     {otherUnit_maskInput_hi[15839:15824]},
     {otherUnit_maskInput_hi[15823:15808]},
     {otherUnit_maskInput_hi[15807:15792]},
     {otherUnit_maskInput_hi[15791:15776]},
     {otherUnit_maskInput_hi[15775:15760]},
     {otherUnit_maskInput_hi[15759:15744]},
     {otherUnit_maskInput_hi[15743:15728]},
     {otherUnit_maskInput_hi[15727:15712]},
     {otherUnit_maskInput_hi[15711:15696]},
     {otherUnit_maskInput_hi[15695:15680]},
     {otherUnit_maskInput_hi[15679:15664]},
     {otherUnit_maskInput_hi[15663:15648]},
     {otherUnit_maskInput_hi[15647:15632]},
     {otherUnit_maskInput_hi[15631:15616]},
     {otherUnit_maskInput_hi[15615:15600]},
     {otherUnit_maskInput_hi[15599:15584]},
     {otherUnit_maskInput_hi[15583:15568]},
     {otherUnit_maskInput_hi[15567:15552]},
     {otherUnit_maskInput_hi[15551:15536]},
     {otherUnit_maskInput_hi[15535:15520]},
     {otherUnit_maskInput_hi[15519:15504]},
     {otherUnit_maskInput_hi[15503:15488]},
     {otherUnit_maskInput_hi[15487:15472]},
     {otherUnit_maskInput_hi[15471:15456]},
     {otherUnit_maskInput_hi[15455:15440]},
     {otherUnit_maskInput_hi[15439:15424]},
     {otherUnit_maskInput_hi[15423:15408]},
     {otherUnit_maskInput_hi[15407:15392]},
     {otherUnit_maskInput_hi[15391:15376]},
     {otherUnit_maskInput_hi[15375:15360]},
     {otherUnit_maskInput_hi[15359:15344]},
     {otherUnit_maskInput_hi[15343:15328]},
     {otherUnit_maskInput_hi[15327:15312]},
     {otherUnit_maskInput_hi[15311:15296]},
     {otherUnit_maskInput_hi[15295:15280]},
     {otherUnit_maskInput_hi[15279:15264]},
     {otherUnit_maskInput_hi[15263:15248]},
     {otherUnit_maskInput_hi[15247:15232]},
     {otherUnit_maskInput_hi[15231:15216]},
     {otherUnit_maskInput_hi[15215:15200]},
     {otherUnit_maskInput_hi[15199:15184]},
     {otherUnit_maskInput_hi[15183:15168]},
     {otherUnit_maskInput_hi[15167:15152]},
     {otherUnit_maskInput_hi[15151:15136]},
     {otherUnit_maskInput_hi[15135:15120]},
     {otherUnit_maskInput_hi[15119:15104]},
     {otherUnit_maskInput_hi[15103:15088]},
     {otherUnit_maskInput_hi[15087:15072]},
     {otherUnit_maskInput_hi[15071:15056]},
     {otherUnit_maskInput_hi[15055:15040]},
     {otherUnit_maskInput_hi[15039:15024]},
     {otherUnit_maskInput_hi[15023:15008]},
     {otherUnit_maskInput_hi[15007:14992]},
     {otherUnit_maskInput_hi[14991:14976]},
     {otherUnit_maskInput_hi[14975:14960]},
     {otherUnit_maskInput_hi[14959:14944]},
     {otherUnit_maskInput_hi[14943:14928]},
     {otherUnit_maskInput_hi[14927:14912]},
     {otherUnit_maskInput_hi[14911:14896]},
     {otherUnit_maskInput_hi[14895:14880]},
     {otherUnit_maskInput_hi[14879:14864]},
     {otherUnit_maskInput_hi[14863:14848]},
     {otherUnit_maskInput_hi[14847:14832]},
     {otherUnit_maskInput_hi[14831:14816]},
     {otherUnit_maskInput_hi[14815:14800]},
     {otherUnit_maskInput_hi[14799:14784]},
     {otherUnit_maskInput_hi[14783:14768]},
     {otherUnit_maskInput_hi[14767:14752]},
     {otherUnit_maskInput_hi[14751:14736]},
     {otherUnit_maskInput_hi[14735:14720]},
     {otherUnit_maskInput_hi[14719:14704]},
     {otherUnit_maskInput_hi[14703:14688]},
     {otherUnit_maskInput_hi[14687:14672]},
     {otherUnit_maskInput_hi[14671:14656]},
     {otherUnit_maskInput_hi[14655:14640]},
     {otherUnit_maskInput_hi[14639:14624]},
     {otherUnit_maskInput_hi[14623:14608]},
     {otherUnit_maskInput_hi[14607:14592]},
     {otherUnit_maskInput_hi[14591:14576]},
     {otherUnit_maskInput_hi[14575:14560]},
     {otherUnit_maskInput_hi[14559:14544]},
     {otherUnit_maskInput_hi[14543:14528]},
     {otherUnit_maskInput_hi[14527:14512]},
     {otherUnit_maskInput_hi[14511:14496]},
     {otherUnit_maskInput_hi[14495:14480]},
     {otherUnit_maskInput_hi[14479:14464]},
     {otherUnit_maskInput_hi[14463:14448]},
     {otherUnit_maskInput_hi[14447:14432]},
     {otherUnit_maskInput_hi[14431:14416]},
     {otherUnit_maskInput_hi[14415:14400]},
     {otherUnit_maskInput_hi[14399:14384]},
     {otherUnit_maskInput_hi[14383:14368]},
     {otherUnit_maskInput_hi[14367:14352]},
     {otherUnit_maskInput_hi[14351:14336]},
     {otherUnit_maskInput_hi[14335:14320]},
     {otherUnit_maskInput_hi[14319:14304]},
     {otherUnit_maskInput_hi[14303:14288]},
     {otherUnit_maskInput_hi[14287:14272]},
     {otherUnit_maskInput_hi[14271:14256]},
     {otherUnit_maskInput_hi[14255:14240]},
     {otherUnit_maskInput_hi[14239:14224]},
     {otherUnit_maskInput_hi[14223:14208]},
     {otherUnit_maskInput_hi[14207:14192]},
     {otherUnit_maskInput_hi[14191:14176]},
     {otherUnit_maskInput_hi[14175:14160]},
     {otherUnit_maskInput_hi[14159:14144]},
     {otherUnit_maskInput_hi[14143:14128]},
     {otherUnit_maskInput_hi[14127:14112]},
     {otherUnit_maskInput_hi[14111:14096]},
     {otherUnit_maskInput_hi[14095:14080]},
     {otherUnit_maskInput_hi[14079:14064]},
     {otherUnit_maskInput_hi[14063:14048]},
     {otherUnit_maskInput_hi[14047:14032]},
     {otherUnit_maskInput_hi[14031:14016]},
     {otherUnit_maskInput_hi[14015:14000]},
     {otherUnit_maskInput_hi[13999:13984]},
     {otherUnit_maskInput_hi[13983:13968]},
     {otherUnit_maskInput_hi[13967:13952]},
     {otherUnit_maskInput_hi[13951:13936]},
     {otherUnit_maskInput_hi[13935:13920]},
     {otherUnit_maskInput_hi[13919:13904]},
     {otherUnit_maskInput_hi[13903:13888]},
     {otherUnit_maskInput_hi[13887:13872]},
     {otherUnit_maskInput_hi[13871:13856]},
     {otherUnit_maskInput_hi[13855:13840]},
     {otherUnit_maskInput_hi[13839:13824]},
     {otherUnit_maskInput_hi[13823:13808]},
     {otherUnit_maskInput_hi[13807:13792]},
     {otherUnit_maskInput_hi[13791:13776]},
     {otherUnit_maskInput_hi[13775:13760]},
     {otherUnit_maskInput_hi[13759:13744]},
     {otherUnit_maskInput_hi[13743:13728]},
     {otherUnit_maskInput_hi[13727:13712]},
     {otherUnit_maskInput_hi[13711:13696]},
     {otherUnit_maskInput_hi[13695:13680]},
     {otherUnit_maskInput_hi[13679:13664]},
     {otherUnit_maskInput_hi[13663:13648]},
     {otherUnit_maskInput_hi[13647:13632]},
     {otherUnit_maskInput_hi[13631:13616]},
     {otherUnit_maskInput_hi[13615:13600]},
     {otherUnit_maskInput_hi[13599:13584]},
     {otherUnit_maskInput_hi[13583:13568]},
     {otherUnit_maskInput_hi[13567:13552]},
     {otherUnit_maskInput_hi[13551:13536]},
     {otherUnit_maskInput_hi[13535:13520]},
     {otherUnit_maskInput_hi[13519:13504]},
     {otherUnit_maskInput_hi[13503:13488]},
     {otherUnit_maskInput_hi[13487:13472]},
     {otherUnit_maskInput_hi[13471:13456]},
     {otherUnit_maskInput_hi[13455:13440]},
     {otherUnit_maskInput_hi[13439:13424]},
     {otherUnit_maskInput_hi[13423:13408]},
     {otherUnit_maskInput_hi[13407:13392]},
     {otherUnit_maskInput_hi[13391:13376]},
     {otherUnit_maskInput_hi[13375:13360]},
     {otherUnit_maskInput_hi[13359:13344]},
     {otherUnit_maskInput_hi[13343:13328]},
     {otherUnit_maskInput_hi[13327:13312]},
     {otherUnit_maskInput_hi[13311:13296]},
     {otherUnit_maskInput_hi[13295:13280]},
     {otherUnit_maskInput_hi[13279:13264]},
     {otherUnit_maskInput_hi[13263:13248]},
     {otherUnit_maskInput_hi[13247:13232]},
     {otherUnit_maskInput_hi[13231:13216]},
     {otherUnit_maskInput_hi[13215:13200]},
     {otherUnit_maskInput_hi[13199:13184]},
     {otherUnit_maskInput_hi[13183:13168]},
     {otherUnit_maskInput_hi[13167:13152]},
     {otherUnit_maskInput_hi[13151:13136]},
     {otherUnit_maskInput_hi[13135:13120]},
     {otherUnit_maskInput_hi[13119:13104]},
     {otherUnit_maskInput_hi[13103:13088]},
     {otherUnit_maskInput_hi[13087:13072]},
     {otherUnit_maskInput_hi[13071:13056]},
     {otherUnit_maskInput_hi[13055:13040]},
     {otherUnit_maskInput_hi[13039:13024]},
     {otherUnit_maskInput_hi[13023:13008]},
     {otherUnit_maskInput_hi[13007:12992]},
     {otherUnit_maskInput_hi[12991:12976]},
     {otherUnit_maskInput_hi[12975:12960]},
     {otherUnit_maskInput_hi[12959:12944]},
     {otherUnit_maskInput_hi[12943:12928]},
     {otherUnit_maskInput_hi[12927:12912]},
     {otherUnit_maskInput_hi[12911:12896]},
     {otherUnit_maskInput_hi[12895:12880]},
     {otherUnit_maskInput_hi[12879:12864]},
     {otherUnit_maskInput_hi[12863:12848]},
     {otherUnit_maskInput_hi[12847:12832]},
     {otherUnit_maskInput_hi[12831:12816]},
     {otherUnit_maskInput_hi[12815:12800]},
     {otherUnit_maskInput_hi[12799:12784]},
     {otherUnit_maskInput_hi[12783:12768]},
     {otherUnit_maskInput_hi[12767:12752]},
     {otherUnit_maskInput_hi[12751:12736]},
     {otherUnit_maskInput_hi[12735:12720]},
     {otherUnit_maskInput_hi[12719:12704]},
     {otherUnit_maskInput_hi[12703:12688]},
     {otherUnit_maskInput_hi[12687:12672]},
     {otherUnit_maskInput_hi[12671:12656]},
     {otherUnit_maskInput_hi[12655:12640]},
     {otherUnit_maskInput_hi[12639:12624]},
     {otherUnit_maskInput_hi[12623:12608]},
     {otherUnit_maskInput_hi[12607:12592]},
     {otherUnit_maskInput_hi[12591:12576]},
     {otherUnit_maskInput_hi[12575:12560]},
     {otherUnit_maskInput_hi[12559:12544]},
     {otherUnit_maskInput_hi[12543:12528]},
     {otherUnit_maskInput_hi[12527:12512]},
     {otherUnit_maskInput_hi[12511:12496]},
     {otherUnit_maskInput_hi[12495:12480]},
     {otherUnit_maskInput_hi[12479:12464]},
     {otherUnit_maskInput_hi[12463:12448]},
     {otherUnit_maskInput_hi[12447:12432]},
     {otherUnit_maskInput_hi[12431:12416]},
     {otherUnit_maskInput_hi[12415:12400]},
     {otherUnit_maskInput_hi[12399:12384]},
     {otherUnit_maskInput_hi[12383:12368]},
     {otherUnit_maskInput_hi[12367:12352]},
     {otherUnit_maskInput_hi[12351:12336]},
     {otherUnit_maskInput_hi[12335:12320]},
     {otherUnit_maskInput_hi[12319:12304]},
     {otherUnit_maskInput_hi[12303:12288]},
     {otherUnit_maskInput_hi[12287:12272]},
     {otherUnit_maskInput_hi[12271:12256]},
     {otherUnit_maskInput_hi[12255:12240]},
     {otherUnit_maskInput_hi[12239:12224]},
     {otherUnit_maskInput_hi[12223:12208]},
     {otherUnit_maskInput_hi[12207:12192]},
     {otherUnit_maskInput_hi[12191:12176]},
     {otherUnit_maskInput_hi[12175:12160]},
     {otherUnit_maskInput_hi[12159:12144]},
     {otherUnit_maskInput_hi[12143:12128]},
     {otherUnit_maskInput_hi[12127:12112]},
     {otherUnit_maskInput_hi[12111:12096]},
     {otherUnit_maskInput_hi[12095:12080]},
     {otherUnit_maskInput_hi[12079:12064]},
     {otherUnit_maskInput_hi[12063:12048]},
     {otherUnit_maskInput_hi[12047:12032]},
     {otherUnit_maskInput_hi[12031:12016]},
     {otherUnit_maskInput_hi[12015:12000]},
     {otherUnit_maskInput_hi[11999:11984]},
     {otherUnit_maskInput_hi[11983:11968]},
     {otherUnit_maskInput_hi[11967:11952]},
     {otherUnit_maskInput_hi[11951:11936]},
     {otherUnit_maskInput_hi[11935:11920]},
     {otherUnit_maskInput_hi[11919:11904]},
     {otherUnit_maskInput_hi[11903:11888]},
     {otherUnit_maskInput_hi[11887:11872]},
     {otherUnit_maskInput_hi[11871:11856]},
     {otherUnit_maskInput_hi[11855:11840]},
     {otherUnit_maskInput_hi[11839:11824]},
     {otherUnit_maskInput_hi[11823:11808]},
     {otherUnit_maskInput_hi[11807:11792]},
     {otherUnit_maskInput_hi[11791:11776]},
     {otherUnit_maskInput_hi[11775:11760]},
     {otherUnit_maskInput_hi[11759:11744]},
     {otherUnit_maskInput_hi[11743:11728]},
     {otherUnit_maskInput_hi[11727:11712]},
     {otherUnit_maskInput_hi[11711:11696]},
     {otherUnit_maskInput_hi[11695:11680]},
     {otherUnit_maskInput_hi[11679:11664]},
     {otherUnit_maskInput_hi[11663:11648]},
     {otherUnit_maskInput_hi[11647:11632]},
     {otherUnit_maskInput_hi[11631:11616]},
     {otherUnit_maskInput_hi[11615:11600]},
     {otherUnit_maskInput_hi[11599:11584]},
     {otherUnit_maskInput_hi[11583:11568]},
     {otherUnit_maskInput_hi[11567:11552]},
     {otherUnit_maskInput_hi[11551:11536]},
     {otherUnit_maskInput_hi[11535:11520]},
     {otherUnit_maskInput_hi[11519:11504]},
     {otherUnit_maskInput_hi[11503:11488]},
     {otherUnit_maskInput_hi[11487:11472]},
     {otherUnit_maskInput_hi[11471:11456]},
     {otherUnit_maskInput_hi[11455:11440]},
     {otherUnit_maskInput_hi[11439:11424]},
     {otherUnit_maskInput_hi[11423:11408]},
     {otherUnit_maskInput_hi[11407:11392]},
     {otherUnit_maskInput_hi[11391:11376]},
     {otherUnit_maskInput_hi[11375:11360]},
     {otherUnit_maskInput_hi[11359:11344]},
     {otherUnit_maskInput_hi[11343:11328]},
     {otherUnit_maskInput_hi[11327:11312]},
     {otherUnit_maskInput_hi[11311:11296]},
     {otherUnit_maskInput_hi[11295:11280]},
     {otherUnit_maskInput_hi[11279:11264]},
     {otherUnit_maskInput_hi[11263:11248]},
     {otherUnit_maskInput_hi[11247:11232]},
     {otherUnit_maskInput_hi[11231:11216]},
     {otherUnit_maskInput_hi[11215:11200]},
     {otherUnit_maskInput_hi[11199:11184]},
     {otherUnit_maskInput_hi[11183:11168]},
     {otherUnit_maskInput_hi[11167:11152]},
     {otherUnit_maskInput_hi[11151:11136]},
     {otherUnit_maskInput_hi[11135:11120]},
     {otherUnit_maskInput_hi[11119:11104]},
     {otherUnit_maskInput_hi[11103:11088]},
     {otherUnit_maskInput_hi[11087:11072]},
     {otherUnit_maskInput_hi[11071:11056]},
     {otherUnit_maskInput_hi[11055:11040]},
     {otherUnit_maskInput_hi[11039:11024]},
     {otherUnit_maskInput_hi[11023:11008]},
     {otherUnit_maskInput_hi[11007:10992]},
     {otherUnit_maskInput_hi[10991:10976]},
     {otherUnit_maskInput_hi[10975:10960]},
     {otherUnit_maskInput_hi[10959:10944]},
     {otherUnit_maskInput_hi[10943:10928]},
     {otherUnit_maskInput_hi[10927:10912]},
     {otherUnit_maskInput_hi[10911:10896]},
     {otherUnit_maskInput_hi[10895:10880]},
     {otherUnit_maskInput_hi[10879:10864]},
     {otherUnit_maskInput_hi[10863:10848]},
     {otherUnit_maskInput_hi[10847:10832]},
     {otherUnit_maskInput_hi[10831:10816]},
     {otherUnit_maskInput_hi[10815:10800]},
     {otherUnit_maskInput_hi[10799:10784]},
     {otherUnit_maskInput_hi[10783:10768]},
     {otherUnit_maskInput_hi[10767:10752]},
     {otherUnit_maskInput_hi[10751:10736]},
     {otherUnit_maskInput_hi[10735:10720]},
     {otherUnit_maskInput_hi[10719:10704]},
     {otherUnit_maskInput_hi[10703:10688]},
     {otherUnit_maskInput_hi[10687:10672]},
     {otherUnit_maskInput_hi[10671:10656]},
     {otherUnit_maskInput_hi[10655:10640]},
     {otherUnit_maskInput_hi[10639:10624]},
     {otherUnit_maskInput_hi[10623:10608]},
     {otherUnit_maskInput_hi[10607:10592]},
     {otherUnit_maskInput_hi[10591:10576]},
     {otherUnit_maskInput_hi[10575:10560]},
     {otherUnit_maskInput_hi[10559:10544]},
     {otherUnit_maskInput_hi[10543:10528]},
     {otherUnit_maskInput_hi[10527:10512]},
     {otherUnit_maskInput_hi[10511:10496]},
     {otherUnit_maskInput_hi[10495:10480]},
     {otherUnit_maskInput_hi[10479:10464]},
     {otherUnit_maskInput_hi[10463:10448]},
     {otherUnit_maskInput_hi[10447:10432]},
     {otherUnit_maskInput_hi[10431:10416]},
     {otherUnit_maskInput_hi[10415:10400]},
     {otherUnit_maskInput_hi[10399:10384]},
     {otherUnit_maskInput_hi[10383:10368]},
     {otherUnit_maskInput_hi[10367:10352]},
     {otherUnit_maskInput_hi[10351:10336]},
     {otherUnit_maskInput_hi[10335:10320]},
     {otherUnit_maskInput_hi[10319:10304]},
     {otherUnit_maskInput_hi[10303:10288]},
     {otherUnit_maskInput_hi[10287:10272]},
     {otherUnit_maskInput_hi[10271:10256]},
     {otherUnit_maskInput_hi[10255:10240]},
     {otherUnit_maskInput_hi[10239:10224]},
     {otherUnit_maskInput_hi[10223:10208]},
     {otherUnit_maskInput_hi[10207:10192]},
     {otherUnit_maskInput_hi[10191:10176]},
     {otherUnit_maskInput_hi[10175:10160]},
     {otherUnit_maskInput_hi[10159:10144]},
     {otherUnit_maskInput_hi[10143:10128]},
     {otherUnit_maskInput_hi[10127:10112]},
     {otherUnit_maskInput_hi[10111:10096]},
     {otherUnit_maskInput_hi[10095:10080]},
     {otherUnit_maskInput_hi[10079:10064]},
     {otherUnit_maskInput_hi[10063:10048]},
     {otherUnit_maskInput_hi[10047:10032]},
     {otherUnit_maskInput_hi[10031:10016]},
     {otherUnit_maskInput_hi[10015:10000]},
     {otherUnit_maskInput_hi[9999:9984]},
     {otherUnit_maskInput_hi[9983:9968]},
     {otherUnit_maskInput_hi[9967:9952]},
     {otherUnit_maskInput_hi[9951:9936]},
     {otherUnit_maskInput_hi[9935:9920]},
     {otherUnit_maskInput_hi[9919:9904]},
     {otherUnit_maskInput_hi[9903:9888]},
     {otherUnit_maskInput_hi[9887:9872]},
     {otherUnit_maskInput_hi[9871:9856]},
     {otherUnit_maskInput_hi[9855:9840]},
     {otherUnit_maskInput_hi[9839:9824]},
     {otherUnit_maskInput_hi[9823:9808]},
     {otherUnit_maskInput_hi[9807:9792]},
     {otherUnit_maskInput_hi[9791:9776]},
     {otherUnit_maskInput_hi[9775:9760]},
     {otherUnit_maskInput_hi[9759:9744]},
     {otherUnit_maskInput_hi[9743:9728]},
     {otherUnit_maskInput_hi[9727:9712]},
     {otherUnit_maskInput_hi[9711:9696]},
     {otherUnit_maskInput_hi[9695:9680]},
     {otherUnit_maskInput_hi[9679:9664]},
     {otherUnit_maskInput_hi[9663:9648]},
     {otherUnit_maskInput_hi[9647:9632]},
     {otherUnit_maskInput_hi[9631:9616]},
     {otherUnit_maskInput_hi[9615:9600]},
     {otherUnit_maskInput_hi[9599:9584]},
     {otherUnit_maskInput_hi[9583:9568]},
     {otherUnit_maskInput_hi[9567:9552]},
     {otherUnit_maskInput_hi[9551:9536]},
     {otherUnit_maskInput_hi[9535:9520]},
     {otherUnit_maskInput_hi[9519:9504]},
     {otherUnit_maskInput_hi[9503:9488]},
     {otherUnit_maskInput_hi[9487:9472]},
     {otherUnit_maskInput_hi[9471:9456]},
     {otherUnit_maskInput_hi[9455:9440]},
     {otherUnit_maskInput_hi[9439:9424]},
     {otherUnit_maskInput_hi[9423:9408]},
     {otherUnit_maskInput_hi[9407:9392]},
     {otherUnit_maskInput_hi[9391:9376]},
     {otherUnit_maskInput_hi[9375:9360]},
     {otherUnit_maskInput_hi[9359:9344]},
     {otherUnit_maskInput_hi[9343:9328]},
     {otherUnit_maskInput_hi[9327:9312]},
     {otherUnit_maskInput_hi[9311:9296]},
     {otherUnit_maskInput_hi[9295:9280]},
     {otherUnit_maskInput_hi[9279:9264]},
     {otherUnit_maskInput_hi[9263:9248]},
     {otherUnit_maskInput_hi[9247:9232]},
     {otherUnit_maskInput_hi[9231:9216]},
     {otherUnit_maskInput_hi[9215:9200]},
     {otherUnit_maskInput_hi[9199:9184]},
     {otherUnit_maskInput_hi[9183:9168]},
     {otherUnit_maskInput_hi[9167:9152]},
     {otherUnit_maskInput_hi[9151:9136]},
     {otherUnit_maskInput_hi[9135:9120]},
     {otherUnit_maskInput_hi[9119:9104]},
     {otherUnit_maskInput_hi[9103:9088]},
     {otherUnit_maskInput_hi[9087:9072]},
     {otherUnit_maskInput_hi[9071:9056]},
     {otherUnit_maskInput_hi[9055:9040]},
     {otherUnit_maskInput_hi[9039:9024]},
     {otherUnit_maskInput_hi[9023:9008]},
     {otherUnit_maskInput_hi[9007:8992]},
     {otherUnit_maskInput_hi[8991:8976]},
     {otherUnit_maskInput_hi[8975:8960]},
     {otherUnit_maskInput_hi[8959:8944]},
     {otherUnit_maskInput_hi[8943:8928]},
     {otherUnit_maskInput_hi[8927:8912]},
     {otherUnit_maskInput_hi[8911:8896]},
     {otherUnit_maskInput_hi[8895:8880]},
     {otherUnit_maskInput_hi[8879:8864]},
     {otherUnit_maskInput_hi[8863:8848]},
     {otherUnit_maskInput_hi[8847:8832]},
     {otherUnit_maskInput_hi[8831:8816]},
     {otherUnit_maskInput_hi[8815:8800]},
     {otherUnit_maskInput_hi[8799:8784]},
     {otherUnit_maskInput_hi[8783:8768]},
     {otherUnit_maskInput_hi[8767:8752]},
     {otherUnit_maskInput_hi[8751:8736]},
     {otherUnit_maskInput_hi[8735:8720]},
     {otherUnit_maskInput_hi[8719:8704]},
     {otherUnit_maskInput_hi[8703:8688]},
     {otherUnit_maskInput_hi[8687:8672]},
     {otherUnit_maskInput_hi[8671:8656]},
     {otherUnit_maskInput_hi[8655:8640]},
     {otherUnit_maskInput_hi[8639:8624]},
     {otherUnit_maskInput_hi[8623:8608]},
     {otherUnit_maskInput_hi[8607:8592]},
     {otherUnit_maskInput_hi[8591:8576]},
     {otherUnit_maskInput_hi[8575:8560]},
     {otherUnit_maskInput_hi[8559:8544]},
     {otherUnit_maskInput_hi[8543:8528]},
     {otherUnit_maskInput_hi[8527:8512]},
     {otherUnit_maskInput_hi[8511:8496]},
     {otherUnit_maskInput_hi[8495:8480]},
     {otherUnit_maskInput_hi[8479:8464]},
     {otherUnit_maskInput_hi[8463:8448]},
     {otherUnit_maskInput_hi[8447:8432]},
     {otherUnit_maskInput_hi[8431:8416]},
     {otherUnit_maskInput_hi[8415:8400]},
     {otherUnit_maskInput_hi[8399:8384]},
     {otherUnit_maskInput_hi[8383:8368]},
     {otherUnit_maskInput_hi[8367:8352]},
     {otherUnit_maskInput_hi[8351:8336]},
     {otherUnit_maskInput_hi[8335:8320]},
     {otherUnit_maskInput_hi[8319:8304]},
     {otherUnit_maskInput_hi[8303:8288]},
     {otherUnit_maskInput_hi[8287:8272]},
     {otherUnit_maskInput_hi[8271:8256]},
     {otherUnit_maskInput_hi[8255:8240]},
     {otherUnit_maskInput_hi[8239:8224]},
     {otherUnit_maskInput_hi[8223:8208]},
     {otherUnit_maskInput_hi[8207:8192]},
     {otherUnit_maskInput_hi[8191:8176]},
     {otherUnit_maskInput_hi[8175:8160]},
     {otherUnit_maskInput_hi[8159:8144]},
     {otherUnit_maskInput_hi[8143:8128]},
     {otherUnit_maskInput_hi[8127:8112]},
     {otherUnit_maskInput_hi[8111:8096]},
     {otherUnit_maskInput_hi[8095:8080]},
     {otherUnit_maskInput_hi[8079:8064]},
     {otherUnit_maskInput_hi[8063:8048]},
     {otherUnit_maskInput_hi[8047:8032]},
     {otherUnit_maskInput_hi[8031:8016]},
     {otherUnit_maskInput_hi[8015:8000]},
     {otherUnit_maskInput_hi[7999:7984]},
     {otherUnit_maskInput_hi[7983:7968]},
     {otherUnit_maskInput_hi[7967:7952]},
     {otherUnit_maskInput_hi[7951:7936]},
     {otherUnit_maskInput_hi[7935:7920]},
     {otherUnit_maskInput_hi[7919:7904]},
     {otherUnit_maskInput_hi[7903:7888]},
     {otherUnit_maskInput_hi[7887:7872]},
     {otherUnit_maskInput_hi[7871:7856]},
     {otherUnit_maskInput_hi[7855:7840]},
     {otherUnit_maskInput_hi[7839:7824]},
     {otherUnit_maskInput_hi[7823:7808]},
     {otherUnit_maskInput_hi[7807:7792]},
     {otherUnit_maskInput_hi[7791:7776]},
     {otherUnit_maskInput_hi[7775:7760]},
     {otherUnit_maskInput_hi[7759:7744]},
     {otherUnit_maskInput_hi[7743:7728]},
     {otherUnit_maskInput_hi[7727:7712]},
     {otherUnit_maskInput_hi[7711:7696]},
     {otherUnit_maskInput_hi[7695:7680]},
     {otherUnit_maskInput_hi[7679:7664]},
     {otherUnit_maskInput_hi[7663:7648]},
     {otherUnit_maskInput_hi[7647:7632]},
     {otherUnit_maskInput_hi[7631:7616]},
     {otherUnit_maskInput_hi[7615:7600]},
     {otherUnit_maskInput_hi[7599:7584]},
     {otherUnit_maskInput_hi[7583:7568]},
     {otherUnit_maskInput_hi[7567:7552]},
     {otherUnit_maskInput_hi[7551:7536]},
     {otherUnit_maskInput_hi[7535:7520]},
     {otherUnit_maskInput_hi[7519:7504]},
     {otherUnit_maskInput_hi[7503:7488]},
     {otherUnit_maskInput_hi[7487:7472]},
     {otherUnit_maskInput_hi[7471:7456]},
     {otherUnit_maskInput_hi[7455:7440]},
     {otherUnit_maskInput_hi[7439:7424]},
     {otherUnit_maskInput_hi[7423:7408]},
     {otherUnit_maskInput_hi[7407:7392]},
     {otherUnit_maskInput_hi[7391:7376]},
     {otherUnit_maskInput_hi[7375:7360]},
     {otherUnit_maskInput_hi[7359:7344]},
     {otherUnit_maskInput_hi[7343:7328]},
     {otherUnit_maskInput_hi[7327:7312]},
     {otherUnit_maskInput_hi[7311:7296]},
     {otherUnit_maskInput_hi[7295:7280]},
     {otherUnit_maskInput_hi[7279:7264]},
     {otherUnit_maskInput_hi[7263:7248]},
     {otherUnit_maskInput_hi[7247:7232]},
     {otherUnit_maskInput_hi[7231:7216]},
     {otherUnit_maskInput_hi[7215:7200]},
     {otherUnit_maskInput_hi[7199:7184]},
     {otherUnit_maskInput_hi[7183:7168]},
     {otherUnit_maskInput_hi[7167:7152]},
     {otherUnit_maskInput_hi[7151:7136]},
     {otherUnit_maskInput_hi[7135:7120]},
     {otherUnit_maskInput_hi[7119:7104]},
     {otherUnit_maskInput_hi[7103:7088]},
     {otherUnit_maskInput_hi[7087:7072]},
     {otherUnit_maskInput_hi[7071:7056]},
     {otherUnit_maskInput_hi[7055:7040]},
     {otherUnit_maskInput_hi[7039:7024]},
     {otherUnit_maskInput_hi[7023:7008]},
     {otherUnit_maskInput_hi[7007:6992]},
     {otherUnit_maskInput_hi[6991:6976]},
     {otherUnit_maskInput_hi[6975:6960]},
     {otherUnit_maskInput_hi[6959:6944]},
     {otherUnit_maskInput_hi[6943:6928]},
     {otherUnit_maskInput_hi[6927:6912]},
     {otherUnit_maskInput_hi[6911:6896]},
     {otherUnit_maskInput_hi[6895:6880]},
     {otherUnit_maskInput_hi[6879:6864]},
     {otherUnit_maskInput_hi[6863:6848]},
     {otherUnit_maskInput_hi[6847:6832]},
     {otherUnit_maskInput_hi[6831:6816]},
     {otherUnit_maskInput_hi[6815:6800]},
     {otherUnit_maskInput_hi[6799:6784]},
     {otherUnit_maskInput_hi[6783:6768]},
     {otherUnit_maskInput_hi[6767:6752]},
     {otherUnit_maskInput_hi[6751:6736]},
     {otherUnit_maskInput_hi[6735:6720]},
     {otherUnit_maskInput_hi[6719:6704]},
     {otherUnit_maskInput_hi[6703:6688]},
     {otherUnit_maskInput_hi[6687:6672]},
     {otherUnit_maskInput_hi[6671:6656]},
     {otherUnit_maskInput_hi[6655:6640]},
     {otherUnit_maskInput_hi[6639:6624]},
     {otherUnit_maskInput_hi[6623:6608]},
     {otherUnit_maskInput_hi[6607:6592]},
     {otherUnit_maskInput_hi[6591:6576]},
     {otherUnit_maskInput_hi[6575:6560]},
     {otherUnit_maskInput_hi[6559:6544]},
     {otherUnit_maskInput_hi[6543:6528]},
     {otherUnit_maskInput_hi[6527:6512]},
     {otherUnit_maskInput_hi[6511:6496]},
     {otherUnit_maskInput_hi[6495:6480]},
     {otherUnit_maskInput_hi[6479:6464]},
     {otherUnit_maskInput_hi[6463:6448]},
     {otherUnit_maskInput_hi[6447:6432]},
     {otherUnit_maskInput_hi[6431:6416]},
     {otherUnit_maskInput_hi[6415:6400]},
     {otherUnit_maskInput_hi[6399:6384]},
     {otherUnit_maskInput_hi[6383:6368]},
     {otherUnit_maskInput_hi[6367:6352]},
     {otherUnit_maskInput_hi[6351:6336]},
     {otherUnit_maskInput_hi[6335:6320]},
     {otherUnit_maskInput_hi[6319:6304]},
     {otherUnit_maskInput_hi[6303:6288]},
     {otherUnit_maskInput_hi[6287:6272]},
     {otherUnit_maskInput_hi[6271:6256]},
     {otherUnit_maskInput_hi[6255:6240]},
     {otherUnit_maskInput_hi[6239:6224]},
     {otherUnit_maskInput_hi[6223:6208]},
     {otherUnit_maskInput_hi[6207:6192]},
     {otherUnit_maskInput_hi[6191:6176]},
     {otherUnit_maskInput_hi[6175:6160]},
     {otherUnit_maskInput_hi[6159:6144]},
     {otherUnit_maskInput_hi[6143:6128]},
     {otherUnit_maskInput_hi[6127:6112]},
     {otherUnit_maskInput_hi[6111:6096]},
     {otherUnit_maskInput_hi[6095:6080]},
     {otherUnit_maskInput_hi[6079:6064]},
     {otherUnit_maskInput_hi[6063:6048]},
     {otherUnit_maskInput_hi[6047:6032]},
     {otherUnit_maskInput_hi[6031:6016]},
     {otherUnit_maskInput_hi[6015:6000]},
     {otherUnit_maskInput_hi[5999:5984]},
     {otherUnit_maskInput_hi[5983:5968]},
     {otherUnit_maskInput_hi[5967:5952]},
     {otherUnit_maskInput_hi[5951:5936]},
     {otherUnit_maskInput_hi[5935:5920]},
     {otherUnit_maskInput_hi[5919:5904]},
     {otherUnit_maskInput_hi[5903:5888]},
     {otherUnit_maskInput_hi[5887:5872]},
     {otherUnit_maskInput_hi[5871:5856]},
     {otherUnit_maskInput_hi[5855:5840]},
     {otherUnit_maskInput_hi[5839:5824]},
     {otherUnit_maskInput_hi[5823:5808]},
     {otherUnit_maskInput_hi[5807:5792]},
     {otherUnit_maskInput_hi[5791:5776]},
     {otherUnit_maskInput_hi[5775:5760]},
     {otherUnit_maskInput_hi[5759:5744]},
     {otherUnit_maskInput_hi[5743:5728]},
     {otherUnit_maskInput_hi[5727:5712]},
     {otherUnit_maskInput_hi[5711:5696]},
     {otherUnit_maskInput_hi[5695:5680]},
     {otherUnit_maskInput_hi[5679:5664]},
     {otherUnit_maskInput_hi[5663:5648]},
     {otherUnit_maskInput_hi[5647:5632]},
     {otherUnit_maskInput_hi[5631:5616]},
     {otherUnit_maskInput_hi[5615:5600]},
     {otherUnit_maskInput_hi[5599:5584]},
     {otherUnit_maskInput_hi[5583:5568]},
     {otherUnit_maskInput_hi[5567:5552]},
     {otherUnit_maskInput_hi[5551:5536]},
     {otherUnit_maskInput_hi[5535:5520]},
     {otherUnit_maskInput_hi[5519:5504]},
     {otherUnit_maskInput_hi[5503:5488]},
     {otherUnit_maskInput_hi[5487:5472]},
     {otherUnit_maskInput_hi[5471:5456]},
     {otherUnit_maskInput_hi[5455:5440]},
     {otherUnit_maskInput_hi[5439:5424]},
     {otherUnit_maskInput_hi[5423:5408]},
     {otherUnit_maskInput_hi[5407:5392]},
     {otherUnit_maskInput_hi[5391:5376]},
     {otherUnit_maskInput_hi[5375:5360]},
     {otherUnit_maskInput_hi[5359:5344]},
     {otherUnit_maskInput_hi[5343:5328]},
     {otherUnit_maskInput_hi[5327:5312]},
     {otherUnit_maskInput_hi[5311:5296]},
     {otherUnit_maskInput_hi[5295:5280]},
     {otherUnit_maskInput_hi[5279:5264]},
     {otherUnit_maskInput_hi[5263:5248]},
     {otherUnit_maskInput_hi[5247:5232]},
     {otherUnit_maskInput_hi[5231:5216]},
     {otherUnit_maskInput_hi[5215:5200]},
     {otherUnit_maskInput_hi[5199:5184]},
     {otherUnit_maskInput_hi[5183:5168]},
     {otherUnit_maskInput_hi[5167:5152]},
     {otherUnit_maskInput_hi[5151:5136]},
     {otherUnit_maskInput_hi[5135:5120]},
     {otherUnit_maskInput_hi[5119:5104]},
     {otherUnit_maskInput_hi[5103:5088]},
     {otherUnit_maskInput_hi[5087:5072]},
     {otherUnit_maskInput_hi[5071:5056]},
     {otherUnit_maskInput_hi[5055:5040]},
     {otherUnit_maskInput_hi[5039:5024]},
     {otherUnit_maskInput_hi[5023:5008]},
     {otherUnit_maskInput_hi[5007:4992]},
     {otherUnit_maskInput_hi[4991:4976]},
     {otherUnit_maskInput_hi[4975:4960]},
     {otherUnit_maskInput_hi[4959:4944]},
     {otherUnit_maskInput_hi[4943:4928]},
     {otherUnit_maskInput_hi[4927:4912]},
     {otherUnit_maskInput_hi[4911:4896]},
     {otherUnit_maskInput_hi[4895:4880]},
     {otherUnit_maskInput_hi[4879:4864]},
     {otherUnit_maskInput_hi[4863:4848]},
     {otherUnit_maskInput_hi[4847:4832]},
     {otherUnit_maskInput_hi[4831:4816]},
     {otherUnit_maskInput_hi[4815:4800]},
     {otherUnit_maskInput_hi[4799:4784]},
     {otherUnit_maskInput_hi[4783:4768]},
     {otherUnit_maskInput_hi[4767:4752]},
     {otherUnit_maskInput_hi[4751:4736]},
     {otherUnit_maskInput_hi[4735:4720]},
     {otherUnit_maskInput_hi[4719:4704]},
     {otherUnit_maskInput_hi[4703:4688]},
     {otherUnit_maskInput_hi[4687:4672]},
     {otherUnit_maskInput_hi[4671:4656]},
     {otherUnit_maskInput_hi[4655:4640]},
     {otherUnit_maskInput_hi[4639:4624]},
     {otherUnit_maskInput_hi[4623:4608]},
     {otherUnit_maskInput_hi[4607:4592]},
     {otherUnit_maskInput_hi[4591:4576]},
     {otherUnit_maskInput_hi[4575:4560]},
     {otherUnit_maskInput_hi[4559:4544]},
     {otherUnit_maskInput_hi[4543:4528]},
     {otherUnit_maskInput_hi[4527:4512]},
     {otherUnit_maskInput_hi[4511:4496]},
     {otherUnit_maskInput_hi[4495:4480]},
     {otherUnit_maskInput_hi[4479:4464]},
     {otherUnit_maskInput_hi[4463:4448]},
     {otherUnit_maskInput_hi[4447:4432]},
     {otherUnit_maskInput_hi[4431:4416]},
     {otherUnit_maskInput_hi[4415:4400]},
     {otherUnit_maskInput_hi[4399:4384]},
     {otherUnit_maskInput_hi[4383:4368]},
     {otherUnit_maskInput_hi[4367:4352]},
     {otherUnit_maskInput_hi[4351:4336]},
     {otherUnit_maskInput_hi[4335:4320]},
     {otherUnit_maskInput_hi[4319:4304]},
     {otherUnit_maskInput_hi[4303:4288]},
     {otherUnit_maskInput_hi[4287:4272]},
     {otherUnit_maskInput_hi[4271:4256]},
     {otherUnit_maskInput_hi[4255:4240]},
     {otherUnit_maskInput_hi[4239:4224]},
     {otherUnit_maskInput_hi[4223:4208]},
     {otherUnit_maskInput_hi[4207:4192]},
     {otherUnit_maskInput_hi[4191:4176]},
     {otherUnit_maskInput_hi[4175:4160]},
     {otherUnit_maskInput_hi[4159:4144]},
     {otherUnit_maskInput_hi[4143:4128]},
     {otherUnit_maskInput_hi[4127:4112]},
     {otherUnit_maskInput_hi[4111:4096]},
     {otherUnit_maskInput_hi[4095:4080]},
     {otherUnit_maskInput_hi[4079:4064]},
     {otherUnit_maskInput_hi[4063:4048]},
     {otherUnit_maskInput_hi[4047:4032]},
     {otherUnit_maskInput_hi[4031:4016]},
     {otherUnit_maskInput_hi[4015:4000]},
     {otherUnit_maskInput_hi[3999:3984]},
     {otherUnit_maskInput_hi[3983:3968]},
     {otherUnit_maskInput_hi[3967:3952]},
     {otherUnit_maskInput_hi[3951:3936]},
     {otherUnit_maskInput_hi[3935:3920]},
     {otherUnit_maskInput_hi[3919:3904]},
     {otherUnit_maskInput_hi[3903:3888]},
     {otherUnit_maskInput_hi[3887:3872]},
     {otherUnit_maskInput_hi[3871:3856]},
     {otherUnit_maskInput_hi[3855:3840]},
     {otherUnit_maskInput_hi[3839:3824]},
     {otherUnit_maskInput_hi[3823:3808]},
     {otherUnit_maskInput_hi[3807:3792]},
     {otherUnit_maskInput_hi[3791:3776]},
     {otherUnit_maskInput_hi[3775:3760]},
     {otherUnit_maskInput_hi[3759:3744]},
     {otherUnit_maskInput_hi[3743:3728]},
     {otherUnit_maskInput_hi[3727:3712]},
     {otherUnit_maskInput_hi[3711:3696]},
     {otherUnit_maskInput_hi[3695:3680]},
     {otherUnit_maskInput_hi[3679:3664]},
     {otherUnit_maskInput_hi[3663:3648]},
     {otherUnit_maskInput_hi[3647:3632]},
     {otherUnit_maskInput_hi[3631:3616]},
     {otherUnit_maskInput_hi[3615:3600]},
     {otherUnit_maskInput_hi[3599:3584]},
     {otherUnit_maskInput_hi[3583:3568]},
     {otherUnit_maskInput_hi[3567:3552]},
     {otherUnit_maskInput_hi[3551:3536]},
     {otherUnit_maskInput_hi[3535:3520]},
     {otherUnit_maskInput_hi[3519:3504]},
     {otherUnit_maskInput_hi[3503:3488]},
     {otherUnit_maskInput_hi[3487:3472]},
     {otherUnit_maskInput_hi[3471:3456]},
     {otherUnit_maskInput_hi[3455:3440]},
     {otherUnit_maskInput_hi[3439:3424]},
     {otherUnit_maskInput_hi[3423:3408]},
     {otherUnit_maskInput_hi[3407:3392]},
     {otherUnit_maskInput_hi[3391:3376]},
     {otherUnit_maskInput_hi[3375:3360]},
     {otherUnit_maskInput_hi[3359:3344]},
     {otherUnit_maskInput_hi[3343:3328]},
     {otherUnit_maskInput_hi[3327:3312]},
     {otherUnit_maskInput_hi[3311:3296]},
     {otherUnit_maskInput_hi[3295:3280]},
     {otherUnit_maskInput_hi[3279:3264]},
     {otherUnit_maskInput_hi[3263:3248]},
     {otherUnit_maskInput_hi[3247:3232]},
     {otherUnit_maskInput_hi[3231:3216]},
     {otherUnit_maskInput_hi[3215:3200]},
     {otherUnit_maskInput_hi[3199:3184]},
     {otherUnit_maskInput_hi[3183:3168]},
     {otherUnit_maskInput_hi[3167:3152]},
     {otherUnit_maskInput_hi[3151:3136]},
     {otherUnit_maskInput_hi[3135:3120]},
     {otherUnit_maskInput_hi[3119:3104]},
     {otherUnit_maskInput_hi[3103:3088]},
     {otherUnit_maskInput_hi[3087:3072]},
     {otherUnit_maskInput_hi[3071:3056]},
     {otherUnit_maskInput_hi[3055:3040]},
     {otherUnit_maskInput_hi[3039:3024]},
     {otherUnit_maskInput_hi[3023:3008]},
     {otherUnit_maskInput_hi[3007:2992]},
     {otherUnit_maskInput_hi[2991:2976]},
     {otherUnit_maskInput_hi[2975:2960]},
     {otherUnit_maskInput_hi[2959:2944]},
     {otherUnit_maskInput_hi[2943:2928]},
     {otherUnit_maskInput_hi[2927:2912]},
     {otherUnit_maskInput_hi[2911:2896]},
     {otherUnit_maskInput_hi[2895:2880]},
     {otherUnit_maskInput_hi[2879:2864]},
     {otherUnit_maskInput_hi[2863:2848]},
     {otherUnit_maskInput_hi[2847:2832]},
     {otherUnit_maskInput_hi[2831:2816]},
     {otherUnit_maskInput_hi[2815:2800]},
     {otherUnit_maskInput_hi[2799:2784]},
     {otherUnit_maskInput_hi[2783:2768]},
     {otherUnit_maskInput_hi[2767:2752]},
     {otherUnit_maskInput_hi[2751:2736]},
     {otherUnit_maskInput_hi[2735:2720]},
     {otherUnit_maskInput_hi[2719:2704]},
     {otherUnit_maskInput_hi[2703:2688]},
     {otherUnit_maskInput_hi[2687:2672]},
     {otherUnit_maskInput_hi[2671:2656]},
     {otherUnit_maskInput_hi[2655:2640]},
     {otherUnit_maskInput_hi[2639:2624]},
     {otherUnit_maskInput_hi[2623:2608]},
     {otherUnit_maskInput_hi[2607:2592]},
     {otherUnit_maskInput_hi[2591:2576]},
     {otherUnit_maskInput_hi[2575:2560]},
     {otherUnit_maskInput_hi[2559:2544]},
     {otherUnit_maskInput_hi[2543:2528]},
     {otherUnit_maskInput_hi[2527:2512]},
     {otherUnit_maskInput_hi[2511:2496]},
     {otherUnit_maskInput_hi[2495:2480]},
     {otherUnit_maskInput_hi[2479:2464]},
     {otherUnit_maskInput_hi[2463:2448]},
     {otherUnit_maskInput_hi[2447:2432]},
     {otherUnit_maskInput_hi[2431:2416]},
     {otherUnit_maskInput_hi[2415:2400]},
     {otherUnit_maskInput_hi[2399:2384]},
     {otherUnit_maskInput_hi[2383:2368]},
     {otherUnit_maskInput_hi[2367:2352]},
     {otherUnit_maskInput_hi[2351:2336]},
     {otherUnit_maskInput_hi[2335:2320]},
     {otherUnit_maskInput_hi[2319:2304]},
     {otherUnit_maskInput_hi[2303:2288]},
     {otherUnit_maskInput_hi[2287:2272]},
     {otherUnit_maskInput_hi[2271:2256]},
     {otherUnit_maskInput_hi[2255:2240]},
     {otherUnit_maskInput_hi[2239:2224]},
     {otherUnit_maskInput_hi[2223:2208]},
     {otherUnit_maskInput_hi[2207:2192]},
     {otherUnit_maskInput_hi[2191:2176]},
     {otherUnit_maskInput_hi[2175:2160]},
     {otherUnit_maskInput_hi[2159:2144]},
     {otherUnit_maskInput_hi[2143:2128]},
     {otherUnit_maskInput_hi[2127:2112]},
     {otherUnit_maskInput_hi[2111:2096]},
     {otherUnit_maskInput_hi[2095:2080]},
     {otherUnit_maskInput_hi[2079:2064]},
     {otherUnit_maskInput_hi[2063:2048]},
     {otherUnit_maskInput_hi[2047:2032]},
     {otherUnit_maskInput_hi[2031:2016]},
     {otherUnit_maskInput_hi[2015:2000]},
     {otherUnit_maskInput_hi[1999:1984]},
     {otherUnit_maskInput_hi[1983:1968]},
     {otherUnit_maskInput_hi[1967:1952]},
     {otherUnit_maskInput_hi[1951:1936]},
     {otherUnit_maskInput_hi[1935:1920]},
     {otherUnit_maskInput_hi[1919:1904]},
     {otherUnit_maskInput_hi[1903:1888]},
     {otherUnit_maskInput_hi[1887:1872]},
     {otherUnit_maskInput_hi[1871:1856]},
     {otherUnit_maskInput_hi[1855:1840]},
     {otherUnit_maskInput_hi[1839:1824]},
     {otherUnit_maskInput_hi[1823:1808]},
     {otherUnit_maskInput_hi[1807:1792]},
     {otherUnit_maskInput_hi[1791:1776]},
     {otherUnit_maskInput_hi[1775:1760]},
     {otherUnit_maskInput_hi[1759:1744]},
     {otherUnit_maskInput_hi[1743:1728]},
     {otherUnit_maskInput_hi[1727:1712]},
     {otherUnit_maskInput_hi[1711:1696]},
     {otherUnit_maskInput_hi[1695:1680]},
     {otherUnit_maskInput_hi[1679:1664]},
     {otherUnit_maskInput_hi[1663:1648]},
     {otherUnit_maskInput_hi[1647:1632]},
     {otherUnit_maskInput_hi[1631:1616]},
     {otherUnit_maskInput_hi[1615:1600]},
     {otherUnit_maskInput_hi[1599:1584]},
     {otherUnit_maskInput_hi[1583:1568]},
     {otherUnit_maskInput_hi[1567:1552]},
     {otherUnit_maskInput_hi[1551:1536]},
     {otherUnit_maskInput_hi[1535:1520]},
     {otherUnit_maskInput_hi[1519:1504]},
     {otherUnit_maskInput_hi[1503:1488]},
     {otherUnit_maskInput_hi[1487:1472]},
     {otherUnit_maskInput_hi[1471:1456]},
     {otherUnit_maskInput_hi[1455:1440]},
     {otherUnit_maskInput_hi[1439:1424]},
     {otherUnit_maskInput_hi[1423:1408]},
     {otherUnit_maskInput_hi[1407:1392]},
     {otherUnit_maskInput_hi[1391:1376]},
     {otherUnit_maskInput_hi[1375:1360]},
     {otherUnit_maskInput_hi[1359:1344]},
     {otherUnit_maskInput_hi[1343:1328]},
     {otherUnit_maskInput_hi[1327:1312]},
     {otherUnit_maskInput_hi[1311:1296]},
     {otherUnit_maskInput_hi[1295:1280]},
     {otherUnit_maskInput_hi[1279:1264]},
     {otherUnit_maskInput_hi[1263:1248]},
     {otherUnit_maskInput_hi[1247:1232]},
     {otherUnit_maskInput_hi[1231:1216]},
     {otherUnit_maskInput_hi[1215:1200]},
     {otherUnit_maskInput_hi[1199:1184]},
     {otherUnit_maskInput_hi[1183:1168]},
     {otherUnit_maskInput_hi[1167:1152]},
     {otherUnit_maskInput_hi[1151:1136]},
     {otherUnit_maskInput_hi[1135:1120]},
     {otherUnit_maskInput_hi[1119:1104]},
     {otherUnit_maskInput_hi[1103:1088]},
     {otherUnit_maskInput_hi[1087:1072]},
     {otherUnit_maskInput_hi[1071:1056]},
     {otherUnit_maskInput_hi[1055:1040]},
     {otherUnit_maskInput_hi[1039:1024]},
     {otherUnit_maskInput_hi[1023:1008]},
     {otherUnit_maskInput_hi[1007:992]},
     {otherUnit_maskInput_hi[991:976]},
     {otherUnit_maskInput_hi[975:960]},
     {otherUnit_maskInput_hi[959:944]},
     {otherUnit_maskInput_hi[943:928]},
     {otherUnit_maskInput_hi[927:912]},
     {otherUnit_maskInput_hi[911:896]},
     {otherUnit_maskInput_hi[895:880]},
     {otherUnit_maskInput_hi[879:864]},
     {otherUnit_maskInput_hi[863:848]},
     {otherUnit_maskInput_hi[847:832]},
     {otherUnit_maskInput_hi[831:816]},
     {otherUnit_maskInput_hi[815:800]},
     {otherUnit_maskInput_hi[799:784]},
     {otherUnit_maskInput_hi[783:768]},
     {otherUnit_maskInput_hi[767:752]},
     {otherUnit_maskInput_hi[751:736]},
     {otherUnit_maskInput_hi[735:720]},
     {otherUnit_maskInput_hi[719:704]},
     {otherUnit_maskInput_hi[703:688]},
     {otherUnit_maskInput_hi[687:672]},
     {otherUnit_maskInput_hi[671:656]},
     {otherUnit_maskInput_hi[655:640]},
     {otherUnit_maskInput_hi[639:624]},
     {otherUnit_maskInput_hi[623:608]},
     {otherUnit_maskInput_hi[607:592]},
     {otherUnit_maskInput_hi[591:576]},
     {otherUnit_maskInput_hi[575:560]},
     {otherUnit_maskInput_hi[559:544]},
     {otherUnit_maskInput_hi[543:528]},
     {otherUnit_maskInput_hi[527:512]},
     {otherUnit_maskInput_hi[511:496]},
     {otherUnit_maskInput_hi[495:480]},
     {otherUnit_maskInput_hi[479:464]},
     {otherUnit_maskInput_hi[463:448]},
     {otherUnit_maskInput_hi[447:432]},
     {otherUnit_maskInput_hi[431:416]},
     {otherUnit_maskInput_hi[415:400]},
     {otherUnit_maskInput_hi[399:384]},
     {otherUnit_maskInput_hi[383:368]},
     {otherUnit_maskInput_hi[367:352]},
     {otherUnit_maskInput_hi[351:336]},
     {otherUnit_maskInput_hi[335:320]},
     {otherUnit_maskInput_hi[319:304]},
     {otherUnit_maskInput_hi[303:288]},
     {otherUnit_maskInput_hi[287:272]},
     {otherUnit_maskInput_hi[271:256]},
     {otherUnit_maskInput_hi[255:240]},
     {otherUnit_maskInput_hi[239:224]},
     {otherUnit_maskInput_hi[223:208]},
     {otherUnit_maskInput_hi[207:192]},
     {otherUnit_maskInput_hi[191:176]},
     {otherUnit_maskInput_hi[175:160]},
     {otherUnit_maskInput_hi[159:144]},
     {otherUnit_maskInput_hi[143:128]},
     {otherUnit_maskInput_hi[127:112]},
     {otherUnit_maskInput_hi[111:96]},
     {otherUnit_maskInput_hi[95:80]},
     {otherUnit_maskInput_hi[79:64]},
     {otherUnit_maskInput_hi[63:48]},
     {otherUnit_maskInput_hi[47:32]},
     {otherUnit_maskInput_hi[31:16]},
     {otherUnit_maskInput_hi[15:0]},
     {otherUnit_maskInput_lo[16383:16368]},
     {otherUnit_maskInput_lo[16367:16352]},
     {otherUnit_maskInput_lo[16351:16336]},
     {otherUnit_maskInput_lo[16335:16320]},
     {otherUnit_maskInput_lo[16319:16304]},
     {otherUnit_maskInput_lo[16303:16288]},
     {otherUnit_maskInput_lo[16287:16272]},
     {otherUnit_maskInput_lo[16271:16256]},
     {otherUnit_maskInput_lo[16255:16240]},
     {otherUnit_maskInput_lo[16239:16224]},
     {otherUnit_maskInput_lo[16223:16208]},
     {otherUnit_maskInput_lo[16207:16192]},
     {otherUnit_maskInput_lo[16191:16176]},
     {otherUnit_maskInput_lo[16175:16160]},
     {otherUnit_maskInput_lo[16159:16144]},
     {otherUnit_maskInput_lo[16143:16128]},
     {otherUnit_maskInput_lo[16127:16112]},
     {otherUnit_maskInput_lo[16111:16096]},
     {otherUnit_maskInput_lo[16095:16080]},
     {otherUnit_maskInput_lo[16079:16064]},
     {otherUnit_maskInput_lo[16063:16048]},
     {otherUnit_maskInput_lo[16047:16032]},
     {otherUnit_maskInput_lo[16031:16016]},
     {otherUnit_maskInput_lo[16015:16000]},
     {otherUnit_maskInput_lo[15999:15984]},
     {otherUnit_maskInput_lo[15983:15968]},
     {otherUnit_maskInput_lo[15967:15952]},
     {otherUnit_maskInput_lo[15951:15936]},
     {otherUnit_maskInput_lo[15935:15920]},
     {otherUnit_maskInput_lo[15919:15904]},
     {otherUnit_maskInput_lo[15903:15888]},
     {otherUnit_maskInput_lo[15887:15872]},
     {otherUnit_maskInput_lo[15871:15856]},
     {otherUnit_maskInput_lo[15855:15840]},
     {otherUnit_maskInput_lo[15839:15824]},
     {otherUnit_maskInput_lo[15823:15808]},
     {otherUnit_maskInput_lo[15807:15792]},
     {otherUnit_maskInput_lo[15791:15776]},
     {otherUnit_maskInput_lo[15775:15760]},
     {otherUnit_maskInput_lo[15759:15744]},
     {otherUnit_maskInput_lo[15743:15728]},
     {otherUnit_maskInput_lo[15727:15712]},
     {otherUnit_maskInput_lo[15711:15696]},
     {otherUnit_maskInput_lo[15695:15680]},
     {otherUnit_maskInput_lo[15679:15664]},
     {otherUnit_maskInput_lo[15663:15648]},
     {otherUnit_maskInput_lo[15647:15632]},
     {otherUnit_maskInput_lo[15631:15616]},
     {otherUnit_maskInput_lo[15615:15600]},
     {otherUnit_maskInput_lo[15599:15584]},
     {otherUnit_maskInput_lo[15583:15568]},
     {otherUnit_maskInput_lo[15567:15552]},
     {otherUnit_maskInput_lo[15551:15536]},
     {otherUnit_maskInput_lo[15535:15520]},
     {otherUnit_maskInput_lo[15519:15504]},
     {otherUnit_maskInput_lo[15503:15488]},
     {otherUnit_maskInput_lo[15487:15472]},
     {otherUnit_maskInput_lo[15471:15456]},
     {otherUnit_maskInput_lo[15455:15440]},
     {otherUnit_maskInput_lo[15439:15424]},
     {otherUnit_maskInput_lo[15423:15408]},
     {otherUnit_maskInput_lo[15407:15392]},
     {otherUnit_maskInput_lo[15391:15376]},
     {otherUnit_maskInput_lo[15375:15360]},
     {otherUnit_maskInput_lo[15359:15344]},
     {otherUnit_maskInput_lo[15343:15328]},
     {otherUnit_maskInput_lo[15327:15312]},
     {otherUnit_maskInput_lo[15311:15296]},
     {otherUnit_maskInput_lo[15295:15280]},
     {otherUnit_maskInput_lo[15279:15264]},
     {otherUnit_maskInput_lo[15263:15248]},
     {otherUnit_maskInput_lo[15247:15232]},
     {otherUnit_maskInput_lo[15231:15216]},
     {otherUnit_maskInput_lo[15215:15200]},
     {otherUnit_maskInput_lo[15199:15184]},
     {otherUnit_maskInput_lo[15183:15168]},
     {otherUnit_maskInput_lo[15167:15152]},
     {otherUnit_maskInput_lo[15151:15136]},
     {otherUnit_maskInput_lo[15135:15120]},
     {otherUnit_maskInput_lo[15119:15104]},
     {otherUnit_maskInput_lo[15103:15088]},
     {otherUnit_maskInput_lo[15087:15072]},
     {otherUnit_maskInput_lo[15071:15056]},
     {otherUnit_maskInput_lo[15055:15040]},
     {otherUnit_maskInput_lo[15039:15024]},
     {otherUnit_maskInput_lo[15023:15008]},
     {otherUnit_maskInput_lo[15007:14992]},
     {otherUnit_maskInput_lo[14991:14976]},
     {otherUnit_maskInput_lo[14975:14960]},
     {otherUnit_maskInput_lo[14959:14944]},
     {otherUnit_maskInput_lo[14943:14928]},
     {otherUnit_maskInput_lo[14927:14912]},
     {otherUnit_maskInput_lo[14911:14896]},
     {otherUnit_maskInput_lo[14895:14880]},
     {otherUnit_maskInput_lo[14879:14864]},
     {otherUnit_maskInput_lo[14863:14848]},
     {otherUnit_maskInput_lo[14847:14832]},
     {otherUnit_maskInput_lo[14831:14816]},
     {otherUnit_maskInput_lo[14815:14800]},
     {otherUnit_maskInput_lo[14799:14784]},
     {otherUnit_maskInput_lo[14783:14768]},
     {otherUnit_maskInput_lo[14767:14752]},
     {otherUnit_maskInput_lo[14751:14736]},
     {otherUnit_maskInput_lo[14735:14720]},
     {otherUnit_maskInput_lo[14719:14704]},
     {otherUnit_maskInput_lo[14703:14688]},
     {otherUnit_maskInput_lo[14687:14672]},
     {otherUnit_maskInput_lo[14671:14656]},
     {otherUnit_maskInput_lo[14655:14640]},
     {otherUnit_maskInput_lo[14639:14624]},
     {otherUnit_maskInput_lo[14623:14608]},
     {otherUnit_maskInput_lo[14607:14592]},
     {otherUnit_maskInput_lo[14591:14576]},
     {otherUnit_maskInput_lo[14575:14560]},
     {otherUnit_maskInput_lo[14559:14544]},
     {otherUnit_maskInput_lo[14543:14528]},
     {otherUnit_maskInput_lo[14527:14512]},
     {otherUnit_maskInput_lo[14511:14496]},
     {otherUnit_maskInput_lo[14495:14480]},
     {otherUnit_maskInput_lo[14479:14464]},
     {otherUnit_maskInput_lo[14463:14448]},
     {otherUnit_maskInput_lo[14447:14432]},
     {otherUnit_maskInput_lo[14431:14416]},
     {otherUnit_maskInput_lo[14415:14400]},
     {otherUnit_maskInput_lo[14399:14384]},
     {otherUnit_maskInput_lo[14383:14368]},
     {otherUnit_maskInput_lo[14367:14352]},
     {otherUnit_maskInput_lo[14351:14336]},
     {otherUnit_maskInput_lo[14335:14320]},
     {otherUnit_maskInput_lo[14319:14304]},
     {otherUnit_maskInput_lo[14303:14288]},
     {otherUnit_maskInput_lo[14287:14272]},
     {otherUnit_maskInput_lo[14271:14256]},
     {otherUnit_maskInput_lo[14255:14240]},
     {otherUnit_maskInput_lo[14239:14224]},
     {otherUnit_maskInput_lo[14223:14208]},
     {otherUnit_maskInput_lo[14207:14192]},
     {otherUnit_maskInput_lo[14191:14176]},
     {otherUnit_maskInput_lo[14175:14160]},
     {otherUnit_maskInput_lo[14159:14144]},
     {otherUnit_maskInput_lo[14143:14128]},
     {otherUnit_maskInput_lo[14127:14112]},
     {otherUnit_maskInput_lo[14111:14096]},
     {otherUnit_maskInput_lo[14095:14080]},
     {otherUnit_maskInput_lo[14079:14064]},
     {otherUnit_maskInput_lo[14063:14048]},
     {otherUnit_maskInput_lo[14047:14032]},
     {otherUnit_maskInput_lo[14031:14016]},
     {otherUnit_maskInput_lo[14015:14000]},
     {otherUnit_maskInput_lo[13999:13984]},
     {otherUnit_maskInput_lo[13983:13968]},
     {otherUnit_maskInput_lo[13967:13952]},
     {otherUnit_maskInput_lo[13951:13936]},
     {otherUnit_maskInput_lo[13935:13920]},
     {otherUnit_maskInput_lo[13919:13904]},
     {otherUnit_maskInput_lo[13903:13888]},
     {otherUnit_maskInput_lo[13887:13872]},
     {otherUnit_maskInput_lo[13871:13856]},
     {otherUnit_maskInput_lo[13855:13840]},
     {otherUnit_maskInput_lo[13839:13824]},
     {otherUnit_maskInput_lo[13823:13808]},
     {otherUnit_maskInput_lo[13807:13792]},
     {otherUnit_maskInput_lo[13791:13776]},
     {otherUnit_maskInput_lo[13775:13760]},
     {otherUnit_maskInput_lo[13759:13744]},
     {otherUnit_maskInput_lo[13743:13728]},
     {otherUnit_maskInput_lo[13727:13712]},
     {otherUnit_maskInput_lo[13711:13696]},
     {otherUnit_maskInput_lo[13695:13680]},
     {otherUnit_maskInput_lo[13679:13664]},
     {otherUnit_maskInput_lo[13663:13648]},
     {otherUnit_maskInput_lo[13647:13632]},
     {otherUnit_maskInput_lo[13631:13616]},
     {otherUnit_maskInput_lo[13615:13600]},
     {otherUnit_maskInput_lo[13599:13584]},
     {otherUnit_maskInput_lo[13583:13568]},
     {otherUnit_maskInput_lo[13567:13552]},
     {otherUnit_maskInput_lo[13551:13536]},
     {otherUnit_maskInput_lo[13535:13520]},
     {otherUnit_maskInput_lo[13519:13504]},
     {otherUnit_maskInput_lo[13503:13488]},
     {otherUnit_maskInput_lo[13487:13472]},
     {otherUnit_maskInput_lo[13471:13456]},
     {otherUnit_maskInput_lo[13455:13440]},
     {otherUnit_maskInput_lo[13439:13424]},
     {otherUnit_maskInput_lo[13423:13408]},
     {otherUnit_maskInput_lo[13407:13392]},
     {otherUnit_maskInput_lo[13391:13376]},
     {otherUnit_maskInput_lo[13375:13360]},
     {otherUnit_maskInput_lo[13359:13344]},
     {otherUnit_maskInput_lo[13343:13328]},
     {otherUnit_maskInput_lo[13327:13312]},
     {otherUnit_maskInput_lo[13311:13296]},
     {otherUnit_maskInput_lo[13295:13280]},
     {otherUnit_maskInput_lo[13279:13264]},
     {otherUnit_maskInput_lo[13263:13248]},
     {otherUnit_maskInput_lo[13247:13232]},
     {otherUnit_maskInput_lo[13231:13216]},
     {otherUnit_maskInput_lo[13215:13200]},
     {otherUnit_maskInput_lo[13199:13184]},
     {otherUnit_maskInput_lo[13183:13168]},
     {otherUnit_maskInput_lo[13167:13152]},
     {otherUnit_maskInput_lo[13151:13136]},
     {otherUnit_maskInput_lo[13135:13120]},
     {otherUnit_maskInput_lo[13119:13104]},
     {otherUnit_maskInput_lo[13103:13088]},
     {otherUnit_maskInput_lo[13087:13072]},
     {otherUnit_maskInput_lo[13071:13056]},
     {otherUnit_maskInput_lo[13055:13040]},
     {otherUnit_maskInput_lo[13039:13024]},
     {otherUnit_maskInput_lo[13023:13008]},
     {otherUnit_maskInput_lo[13007:12992]},
     {otherUnit_maskInput_lo[12991:12976]},
     {otherUnit_maskInput_lo[12975:12960]},
     {otherUnit_maskInput_lo[12959:12944]},
     {otherUnit_maskInput_lo[12943:12928]},
     {otherUnit_maskInput_lo[12927:12912]},
     {otherUnit_maskInput_lo[12911:12896]},
     {otherUnit_maskInput_lo[12895:12880]},
     {otherUnit_maskInput_lo[12879:12864]},
     {otherUnit_maskInput_lo[12863:12848]},
     {otherUnit_maskInput_lo[12847:12832]},
     {otherUnit_maskInput_lo[12831:12816]},
     {otherUnit_maskInput_lo[12815:12800]},
     {otherUnit_maskInput_lo[12799:12784]},
     {otherUnit_maskInput_lo[12783:12768]},
     {otherUnit_maskInput_lo[12767:12752]},
     {otherUnit_maskInput_lo[12751:12736]},
     {otherUnit_maskInput_lo[12735:12720]},
     {otherUnit_maskInput_lo[12719:12704]},
     {otherUnit_maskInput_lo[12703:12688]},
     {otherUnit_maskInput_lo[12687:12672]},
     {otherUnit_maskInput_lo[12671:12656]},
     {otherUnit_maskInput_lo[12655:12640]},
     {otherUnit_maskInput_lo[12639:12624]},
     {otherUnit_maskInput_lo[12623:12608]},
     {otherUnit_maskInput_lo[12607:12592]},
     {otherUnit_maskInput_lo[12591:12576]},
     {otherUnit_maskInput_lo[12575:12560]},
     {otherUnit_maskInput_lo[12559:12544]},
     {otherUnit_maskInput_lo[12543:12528]},
     {otherUnit_maskInput_lo[12527:12512]},
     {otherUnit_maskInput_lo[12511:12496]},
     {otherUnit_maskInput_lo[12495:12480]},
     {otherUnit_maskInput_lo[12479:12464]},
     {otherUnit_maskInput_lo[12463:12448]},
     {otherUnit_maskInput_lo[12447:12432]},
     {otherUnit_maskInput_lo[12431:12416]},
     {otherUnit_maskInput_lo[12415:12400]},
     {otherUnit_maskInput_lo[12399:12384]},
     {otherUnit_maskInput_lo[12383:12368]},
     {otherUnit_maskInput_lo[12367:12352]},
     {otherUnit_maskInput_lo[12351:12336]},
     {otherUnit_maskInput_lo[12335:12320]},
     {otherUnit_maskInput_lo[12319:12304]},
     {otherUnit_maskInput_lo[12303:12288]},
     {otherUnit_maskInput_lo[12287:12272]},
     {otherUnit_maskInput_lo[12271:12256]},
     {otherUnit_maskInput_lo[12255:12240]},
     {otherUnit_maskInput_lo[12239:12224]},
     {otherUnit_maskInput_lo[12223:12208]},
     {otherUnit_maskInput_lo[12207:12192]},
     {otherUnit_maskInput_lo[12191:12176]},
     {otherUnit_maskInput_lo[12175:12160]},
     {otherUnit_maskInput_lo[12159:12144]},
     {otherUnit_maskInput_lo[12143:12128]},
     {otherUnit_maskInput_lo[12127:12112]},
     {otherUnit_maskInput_lo[12111:12096]},
     {otherUnit_maskInput_lo[12095:12080]},
     {otherUnit_maskInput_lo[12079:12064]},
     {otherUnit_maskInput_lo[12063:12048]},
     {otherUnit_maskInput_lo[12047:12032]},
     {otherUnit_maskInput_lo[12031:12016]},
     {otherUnit_maskInput_lo[12015:12000]},
     {otherUnit_maskInput_lo[11999:11984]},
     {otherUnit_maskInput_lo[11983:11968]},
     {otherUnit_maskInput_lo[11967:11952]},
     {otherUnit_maskInput_lo[11951:11936]},
     {otherUnit_maskInput_lo[11935:11920]},
     {otherUnit_maskInput_lo[11919:11904]},
     {otherUnit_maskInput_lo[11903:11888]},
     {otherUnit_maskInput_lo[11887:11872]},
     {otherUnit_maskInput_lo[11871:11856]},
     {otherUnit_maskInput_lo[11855:11840]},
     {otherUnit_maskInput_lo[11839:11824]},
     {otherUnit_maskInput_lo[11823:11808]},
     {otherUnit_maskInput_lo[11807:11792]},
     {otherUnit_maskInput_lo[11791:11776]},
     {otherUnit_maskInput_lo[11775:11760]},
     {otherUnit_maskInput_lo[11759:11744]},
     {otherUnit_maskInput_lo[11743:11728]},
     {otherUnit_maskInput_lo[11727:11712]},
     {otherUnit_maskInput_lo[11711:11696]},
     {otherUnit_maskInput_lo[11695:11680]},
     {otherUnit_maskInput_lo[11679:11664]},
     {otherUnit_maskInput_lo[11663:11648]},
     {otherUnit_maskInput_lo[11647:11632]},
     {otherUnit_maskInput_lo[11631:11616]},
     {otherUnit_maskInput_lo[11615:11600]},
     {otherUnit_maskInput_lo[11599:11584]},
     {otherUnit_maskInput_lo[11583:11568]},
     {otherUnit_maskInput_lo[11567:11552]},
     {otherUnit_maskInput_lo[11551:11536]},
     {otherUnit_maskInput_lo[11535:11520]},
     {otherUnit_maskInput_lo[11519:11504]},
     {otherUnit_maskInput_lo[11503:11488]},
     {otherUnit_maskInput_lo[11487:11472]},
     {otherUnit_maskInput_lo[11471:11456]},
     {otherUnit_maskInput_lo[11455:11440]},
     {otherUnit_maskInput_lo[11439:11424]},
     {otherUnit_maskInput_lo[11423:11408]},
     {otherUnit_maskInput_lo[11407:11392]},
     {otherUnit_maskInput_lo[11391:11376]},
     {otherUnit_maskInput_lo[11375:11360]},
     {otherUnit_maskInput_lo[11359:11344]},
     {otherUnit_maskInput_lo[11343:11328]},
     {otherUnit_maskInput_lo[11327:11312]},
     {otherUnit_maskInput_lo[11311:11296]},
     {otherUnit_maskInput_lo[11295:11280]},
     {otherUnit_maskInput_lo[11279:11264]},
     {otherUnit_maskInput_lo[11263:11248]},
     {otherUnit_maskInput_lo[11247:11232]},
     {otherUnit_maskInput_lo[11231:11216]},
     {otherUnit_maskInput_lo[11215:11200]},
     {otherUnit_maskInput_lo[11199:11184]},
     {otherUnit_maskInput_lo[11183:11168]},
     {otherUnit_maskInput_lo[11167:11152]},
     {otherUnit_maskInput_lo[11151:11136]},
     {otherUnit_maskInput_lo[11135:11120]},
     {otherUnit_maskInput_lo[11119:11104]},
     {otherUnit_maskInput_lo[11103:11088]},
     {otherUnit_maskInput_lo[11087:11072]},
     {otherUnit_maskInput_lo[11071:11056]},
     {otherUnit_maskInput_lo[11055:11040]},
     {otherUnit_maskInput_lo[11039:11024]},
     {otherUnit_maskInput_lo[11023:11008]},
     {otherUnit_maskInput_lo[11007:10992]},
     {otherUnit_maskInput_lo[10991:10976]},
     {otherUnit_maskInput_lo[10975:10960]},
     {otherUnit_maskInput_lo[10959:10944]},
     {otherUnit_maskInput_lo[10943:10928]},
     {otherUnit_maskInput_lo[10927:10912]},
     {otherUnit_maskInput_lo[10911:10896]},
     {otherUnit_maskInput_lo[10895:10880]},
     {otherUnit_maskInput_lo[10879:10864]},
     {otherUnit_maskInput_lo[10863:10848]},
     {otherUnit_maskInput_lo[10847:10832]},
     {otherUnit_maskInput_lo[10831:10816]},
     {otherUnit_maskInput_lo[10815:10800]},
     {otherUnit_maskInput_lo[10799:10784]},
     {otherUnit_maskInput_lo[10783:10768]},
     {otherUnit_maskInput_lo[10767:10752]},
     {otherUnit_maskInput_lo[10751:10736]},
     {otherUnit_maskInput_lo[10735:10720]},
     {otherUnit_maskInput_lo[10719:10704]},
     {otherUnit_maskInput_lo[10703:10688]},
     {otherUnit_maskInput_lo[10687:10672]},
     {otherUnit_maskInput_lo[10671:10656]},
     {otherUnit_maskInput_lo[10655:10640]},
     {otherUnit_maskInput_lo[10639:10624]},
     {otherUnit_maskInput_lo[10623:10608]},
     {otherUnit_maskInput_lo[10607:10592]},
     {otherUnit_maskInput_lo[10591:10576]},
     {otherUnit_maskInput_lo[10575:10560]},
     {otherUnit_maskInput_lo[10559:10544]},
     {otherUnit_maskInput_lo[10543:10528]},
     {otherUnit_maskInput_lo[10527:10512]},
     {otherUnit_maskInput_lo[10511:10496]},
     {otherUnit_maskInput_lo[10495:10480]},
     {otherUnit_maskInput_lo[10479:10464]},
     {otherUnit_maskInput_lo[10463:10448]},
     {otherUnit_maskInput_lo[10447:10432]},
     {otherUnit_maskInput_lo[10431:10416]},
     {otherUnit_maskInput_lo[10415:10400]},
     {otherUnit_maskInput_lo[10399:10384]},
     {otherUnit_maskInput_lo[10383:10368]},
     {otherUnit_maskInput_lo[10367:10352]},
     {otherUnit_maskInput_lo[10351:10336]},
     {otherUnit_maskInput_lo[10335:10320]},
     {otherUnit_maskInput_lo[10319:10304]},
     {otherUnit_maskInput_lo[10303:10288]},
     {otherUnit_maskInput_lo[10287:10272]},
     {otherUnit_maskInput_lo[10271:10256]},
     {otherUnit_maskInput_lo[10255:10240]},
     {otherUnit_maskInput_lo[10239:10224]},
     {otherUnit_maskInput_lo[10223:10208]},
     {otherUnit_maskInput_lo[10207:10192]},
     {otherUnit_maskInput_lo[10191:10176]},
     {otherUnit_maskInput_lo[10175:10160]},
     {otherUnit_maskInput_lo[10159:10144]},
     {otherUnit_maskInput_lo[10143:10128]},
     {otherUnit_maskInput_lo[10127:10112]},
     {otherUnit_maskInput_lo[10111:10096]},
     {otherUnit_maskInput_lo[10095:10080]},
     {otherUnit_maskInput_lo[10079:10064]},
     {otherUnit_maskInput_lo[10063:10048]},
     {otherUnit_maskInput_lo[10047:10032]},
     {otherUnit_maskInput_lo[10031:10016]},
     {otherUnit_maskInput_lo[10015:10000]},
     {otherUnit_maskInput_lo[9999:9984]},
     {otherUnit_maskInput_lo[9983:9968]},
     {otherUnit_maskInput_lo[9967:9952]},
     {otherUnit_maskInput_lo[9951:9936]},
     {otherUnit_maskInput_lo[9935:9920]},
     {otherUnit_maskInput_lo[9919:9904]},
     {otherUnit_maskInput_lo[9903:9888]},
     {otherUnit_maskInput_lo[9887:9872]},
     {otherUnit_maskInput_lo[9871:9856]},
     {otherUnit_maskInput_lo[9855:9840]},
     {otherUnit_maskInput_lo[9839:9824]},
     {otherUnit_maskInput_lo[9823:9808]},
     {otherUnit_maskInput_lo[9807:9792]},
     {otherUnit_maskInput_lo[9791:9776]},
     {otherUnit_maskInput_lo[9775:9760]},
     {otherUnit_maskInput_lo[9759:9744]},
     {otherUnit_maskInput_lo[9743:9728]},
     {otherUnit_maskInput_lo[9727:9712]},
     {otherUnit_maskInput_lo[9711:9696]},
     {otherUnit_maskInput_lo[9695:9680]},
     {otherUnit_maskInput_lo[9679:9664]},
     {otherUnit_maskInput_lo[9663:9648]},
     {otherUnit_maskInput_lo[9647:9632]},
     {otherUnit_maskInput_lo[9631:9616]},
     {otherUnit_maskInput_lo[9615:9600]},
     {otherUnit_maskInput_lo[9599:9584]},
     {otherUnit_maskInput_lo[9583:9568]},
     {otherUnit_maskInput_lo[9567:9552]},
     {otherUnit_maskInput_lo[9551:9536]},
     {otherUnit_maskInput_lo[9535:9520]},
     {otherUnit_maskInput_lo[9519:9504]},
     {otherUnit_maskInput_lo[9503:9488]},
     {otherUnit_maskInput_lo[9487:9472]},
     {otherUnit_maskInput_lo[9471:9456]},
     {otherUnit_maskInput_lo[9455:9440]},
     {otherUnit_maskInput_lo[9439:9424]},
     {otherUnit_maskInput_lo[9423:9408]},
     {otherUnit_maskInput_lo[9407:9392]},
     {otherUnit_maskInput_lo[9391:9376]},
     {otherUnit_maskInput_lo[9375:9360]},
     {otherUnit_maskInput_lo[9359:9344]},
     {otherUnit_maskInput_lo[9343:9328]},
     {otherUnit_maskInput_lo[9327:9312]},
     {otherUnit_maskInput_lo[9311:9296]},
     {otherUnit_maskInput_lo[9295:9280]},
     {otherUnit_maskInput_lo[9279:9264]},
     {otherUnit_maskInput_lo[9263:9248]},
     {otherUnit_maskInput_lo[9247:9232]},
     {otherUnit_maskInput_lo[9231:9216]},
     {otherUnit_maskInput_lo[9215:9200]},
     {otherUnit_maskInput_lo[9199:9184]},
     {otherUnit_maskInput_lo[9183:9168]},
     {otherUnit_maskInput_lo[9167:9152]},
     {otherUnit_maskInput_lo[9151:9136]},
     {otherUnit_maskInput_lo[9135:9120]},
     {otherUnit_maskInput_lo[9119:9104]},
     {otherUnit_maskInput_lo[9103:9088]},
     {otherUnit_maskInput_lo[9087:9072]},
     {otherUnit_maskInput_lo[9071:9056]},
     {otherUnit_maskInput_lo[9055:9040]},
     {otherUnit_maskInput_lo[9039:9024]},
     {otherUnit_maskInput_lo[9023:9008]},
     {otherUnit_maskInput_lo[9007:8992]},
     {otherUnit_maskInput_lo[8991:8976]},
     {otherUnit_maskInput_lo[8975:8960]},
     {otherUnit_maskInput_lo[8959:8944]},
     {otherUnit_maskInput_lo[8943:8928]},
     {otherUnit_maskInput_lo[8927:8912]},
     {otherUnit_maskInput_lo[8911:8896]},
     {otherUnit_maskInput_lo[8895:8880]},
     {otherUnit_maskInput_lo[8879:8864]},
     {otherUnit_maskInput_lo[8863:8848]},
     {otherUnit_maskInput_lo[8847:8832]},
     {otherUnit_maskInput_lo[8831:8816]},
     {otherUnit_maskInput_lo[8815:8800]},
     {otherUnit_maskInput_lo[8799:8784]},
     {otherUnit_maskInput_lo[8783:8768]},
     {otherUnit_maskInput_lo[8767:8752]},
     {otherUnit_maskInput_lo[8751:8736]},
     {otherUnit_maskInput_lo[8735:8720]},
     {otherUnit_maskInput_lo[8719:8704]},
     {otherUnit_maskInput_lo[8703:8688]},
     {otherUnit_maskInput_lo[8687:8672]},
     {otherUnit_maskInput_lo[8671:8656]},
     {otherUnit_maskInput_lo[8655:8640]},
     {otherUnit_maskInput_lo[8639:8624]},
     {otherUnit_maskInput_lo[8623:8608]},
     {otherUnit_maskInput_lo[8607:8592]},
     {otherUnit_maskInput_lo[8591:8576]},
     {otherUnit_maskInput_lo[8575:8560]},
     {otherUnit_maskInput_lo[8559:8544]},
     {otherUnit_maskInput_lo[8543:8528]},
     {otherUnit_maskInput_lo[8527:8512]},
     {otherUnit_maskInput_lo[8511:8496]},
     {otherUnit_maskInput_lo[8495:8480]},
     {otherUnit_maskInput_lo[8479:8464]},
     {otherUnit_maskInput_lo[8463:8448]},
     {otherUnit_maskInput_lo[8447:8432]},
     {otherUnit_maskInput_lo[8431:8416]},
     {otherUnit_maskInput_lo[8415:8400]},
     {otherUnit_maskInput_lo[8399:8384]},
     {otherUnit_maskInput_lo[8383:8368]},
     {otherUnit_maskInput_lo[8367:8352]},
     {otherUnit_maskInput_lo[8351:8336]},
     {otherUnit_maskInput_lo[8335:8320]},
     {otherUnit_maskInput_lo[8319:8304]},
     {otherUnit_maskInput_lo[8303:8288]},
     {otherUnit_maskInput_lo[8287:8272]},
     {otherUnit_maskInput_lo[8271:8256]},
     {otherUnit_maskInput_lo[8255:8240]},
     {otherUnit_maskInput_lo[8239:8224]},
     {otherUnit_maskInput_lo[8223:8208]},
     {otherUnit_maskInput_lo[8207:8192]},
     {otherUnit_maskInput_lo[8191:8176]},
     {otherUnit_maskInput_lo[8175:8160]},
     {otherUnit_maskInput_lo[8159:8144]},
     {otherUnit_maskInput_lo[8143:8128]},
     {otherUnit_maskInput_lo[8127:8112]},
     {otherUnit_maskInput_lo[8111:8096]},
     {otherUnit_maskInput_lo[8095:8080]},
     {otherUnit_maskInput_lo[8079:8064]},
     {otherUnit_maskInput_lo[8063:8048]},
     {otherUnit_maskInput_lo[8047:8032]},
     {otherUnit_maskInput_lo[8031:8016]},
     {otherUnit_maskInput_lo[8015:8000]},
     {otherUnit_maskInput_lo[7999:7984]},
     {otherUnit_maskInput_lo[7983:7968]},
     {otherUnit_maskInput_lo[7967:7952]},
     {otherUnit_maskInput_lo[7951:7936]},
     {otherUnit_maskInput_lo[7935:7920]},
     {otherUnit_maskInput_lo[7919:7904]},
     {otherUnit_maskInput_lo[7903:7888]},
     {otherUnit_maskInput_lo[7887:7872]},
     {otherUnit_maskInput_lo[7871:7856]},
     {otherUnit_maskInput_lo[7855:7840]},
     {otherUnit_maskInput_lo[7839:7824]},
     {otherUnit_maskInput_lo[7823:7808]},
     {otherUnit_maskInput_lo[7807:7792]},
     {otherUnit_maskInput_lo[7791:7776]},
     {otherUnit_maskInput_lo[7775:7760]},
     {otherUnit_maskInput_lo[7759:7744]},
     {otherUnit_maskInput_lo[7743:7728]},
     {otherUnit_maskInput_lo[7727:7712]},
     {otherUnit_maskInput_lo[7711:7696]},
     {otherUnit_maskInput_lo[7695:7680]},
     {otherUnit_maskInput_lo[7679:7664]},
     {otherUnit_maskInput_lo[7663:7648]},
     {otherUnit_maskInput_lo[7647:7632]},
     {otherUnit_maskInput_lo[7631:7616]},
     {otherUnit_maskInput_lo[7615:7600]},
     {otherUnit_maskInput_lo[7599:7584]},
     {otherUnit_maskInput_lo[7583:7568]},
     {otherUnit_maskInput_lo[7567:7552]},
     {otherUnit_maskInput_lo[7551:7536]},
     {otherUnit_maskInput_lo[7535:7520]},
     {otherUnit_maskInput_lo[7519:7504]},
     {otherUnit_maskInput_lo[7503:7488]},
     {otherUnit_maskInput_lo[7487:7472]},
     {otherUnit_maskInput_lo[7471:7456]},
     {otherUnit_maskInput_lo[7455:7440]},
     {otherUnit_maskInput_lo[7439:7424]},
     {otherUnit_maskInput_lo[7423:7408]},
     {otherUnit_maskInput_lo[7407:7392]},
     {otherUnit_maskInput_lo[7391:7376]},
     {otherUnit_maskInput_lo[7375:7360]},
     {otherUnit_maskInput_lo[7359:7344]},
     {otherUnit_maskInput_lo[7343:7328]},
     {otherUnit_maskInput_lo[7327:7312]},
     {otherUnit_maskInput_lo[7311:7296]},
     {otherUnit_maskInput_lo[7295:7280]},
     {otherUnit_maskInput_lo[7279:7264]},
     {otherUnit_maskInput_lo[7263:7248]},
     {otherUnit_maskInput_lo[7247:7232]},
     {otherUnit_maskInput_lo[7231:7216]},
     {otherUnit_maskInput_lo[7215:7200]},
     {otherUnit_maskInput_lo[7199:7184]},
     {otherUnit_maskInput_lo[7183:7168]},
     {otherUnit_maskInput_lo[7167:7152]},
     {otherUnit_maskInput_lo[7151:7136]},
     {otherUnit_maskInput_lo[7135:7120]},
     {otherUnit_maskInput_lo[7119:7104]},
     {otherUnit_maskInput_lo[7103:7088]},
     {otherUnit_maskInput_lo[7087:7072]},
     {otherUnit_maskInput_lo[7071:7056]},
     {otherUnit_maskInput_lo[7055:7040]},
     {otherUnit_maskInput_lo[7039:7024]},
     {otherUnit_maskInput_lo[7023:7008]},
     {otherUnit_maskInput_lo[7007:6992]},
     {otherUnit_maskInput_lo[6991:6976]},
     {otherUnit_maskInput_lo[6975:6960]},
     {otherUnit_maskInput_lo[6959:6944]},
     {otherUnit_maskInput_lo[6943:6928]},
     {otherUnit_maskInput_lo[6927:6912]},
     {otherUnit_maskInput_lo[6911:6896]},
     {otherUnit_maskInput_lo[6895:6880]},
     {otherUnit_maskInput_lo[6879:6864]},
     {otherUnit_maskInput_lo[6863:6848]},
     {otherUnit_maskInput_lo[6847:6832]},
     {otherUnit_maskInput_lo[6831:6816]},
     {otherUnit_maskInput_lo[6815:6800]},
     {otherUnit_maskInput_lo[6799:6784]},
     {otherUnit_maskInput_lo[6783:6768]},
     {otherUnit_maskInput_lo[6767:6752]},
     {otherUnit_maskInput_lo[6751:6736]},
     {otherUnit_maskInput_lo[6735:6720]},
     {otherUnit_maskInput_lo[6719:6704]},
     {otherUnit_maskInput_lo[6703:6688]},
     {otherUnit_maskInput_lo[6687:6672]},
     {otherUnit_maskInput_lo[6671:6656]},
     {otherUnit_maskInput_lo[6655:6640]},
     {otherUnit_maskInput_lo[6639:6624]},
     {otherUnit_maskInput_lo[6623:6608]},
     {otherUnit_maskInput_lo[6607:6592]},
     {otherUnit_maskInput_lo[6591:6576]},
     {otherUnit_maskInput_lo[6575:6560]},
     {otherUnit_maskInput_lo[6559:6544]},
     {otherUnit_maskInput_lo[6543:6528]},
     {otherUnit_maskInput_lo[6527:6512]},
     {otherUnit_maskInput_lo[6511:6496]},
     {otherUnit_maskInput_lo[6495:6480]},
     {otherUnit_maskInput_lo[6479:6464]},
     {otherUnit_maskInput_lo[6463:6448]},
     {otherUnit_maskInput_lo[6447:6432]},
     {otherUnit_maskInput_lo[6431:6416]},
     {otherUnit_maskInput_lo[6415:6400]},
     {otherUnit_maskInput_lo[6399:6384]},
     {otherUnit_maskInput_lo[6383:6368]},
     {otherUnit_maskInput_lo[6367:6352]},
     {otherUnit_maskInput_lo[6351:6336]},
     {otherUnit_maskInput_lo[6335:6320]},
     {otherUnit_maskInput_lo[6319:6304]},
     {otherUnit_maskInput_lo[6303:6288]},
     {otherUnit_maskInput_lo[6287:6272]},
     {otherUnit_maskInput_lo[6271:6256]},
     {otherUnit_maskInput_lo[6255:6240]},
     {otherUnit_maskInput_lo[6239:6224]},
     {otherUnit_maskInput_lo[6223:6208]},
     {otherUnit_maskInput_lo[6207:6192]},
     {otherUnit_maskInput_lo[6191:6176]},
     {otherUnit_maskInput_lo[6175:6160]},
     {otherUnit_maskInput_lo[6159:6144]},
     {otherUnit_maskInput_lo[6143:6128]},
     {otherUnit_maskInput_lo[6127:6112]},
     {otherUnit_maskInput_lo[6111:6096]},
     {otherUnit_maskInput_lo[6095:6080]},
     {otherUnit_maskInput_lo[6079:6064]},
     {otherUnit_maskInput_lo[6063:6048]},
     {otherUnit_maskInput_lo[6047:6032]},
     {otherUnit_maskInput_lo[6031:6016]},
     {otherUnit_maskInput_lo[6015:6000]},
     {otherUnit_maskInput_lo[5999:5984]},
     {otherUnit_maskInput_lo[5983:5968]},
     {otherUnit_maskInput_lo[5967:5952]},
     {otherUnit_maskInput_lo[5951:5936]},
     {otherUnit_maskInput_lo[5935:5920]},
     {otherUnit_maskInput_lo[5919:5904]},
     {otherUnit_maskInput_lo[5903:5888]},
     {otherUnit_maskInput_lo[5887:5872]},
     {otherUnit_maskInput_lo[5871:5856]},
     {otherUnit_maskInput_lo[5855:5840]},
     {otherUnit_maskInput_lo[5839:5824]},
     {otherUnit_maskInput_lo[5823:5808]},
     {otherUnit_maskInput_lo[5807:5792]},
     {otherUnit_maskInput_lo[5791:5776]},
     {otherUnit_maskInput_lo[5775:5760]},
     {otherUnit_maskInput_lo[5759:5744]},
     {otherUnit_maskInput_lo[5743:5728]},
     {otherUnit_maskInput_lo[5727:5712]},
     {otherUnit_maskInput_lo[5711:5696]},
     {otherUnit_maskInput_lo[5695:5680]},
     {otherUnit_maskInput_lo[5679:5664]},
     {otherUnit_maskInput_lo[5663:5648]},
     {otherUnit_maskInput_lo[5647:5632]},
     {otherUnit_maskInput_lo[5631:5616]},
     {otherUnit_maskInput_lo[5615:5600]},
     {otherUnit_maskInput_lo[5599:5584]},
     {otherUnit_maskInput_lo[5583:5568]},
     {otherUnit_maskInput_lo[5567:5552]},
     {otherUnit_maskInput_lo[5551:5536]},
     {otherUnit_maskInput_lo[5535:5520]},
     {otherUnit_maskInput_lo[5519:5504]},
     {otherUnit_maskInput_lo[5503:5488]},
     {otherUnit_maskInput_lo[5487:5472]},
     {otherUnit_maskInput_lo[5471:5456]},
     {otherUnit_maskInput_lo[5455:5440]},
     {otherUnit_maskInput_lo[5439:5424]},
     {otherUnit_maskInput_lo[5423:5408]},
     {otherUnit_maskInput_lo[5407:5392]},
     {otherUnit_maskInput_lo[5391:5376]},
     {otherUnit_maskInput_lo[5375:5360]},
     {otherUnit_maskInput_lo[5359:5344]},
     {otherUnit_maskInput_lo[5343:5328]},
     {otherUnit_maskInput_lo[5327:5312]},
     {otherUnit_maskInput_lo[5311:5296]},
     {otherUnit_maskInput_lo[5295:5280]},
     {otherUnit_maskInput_lo[5279:5264]},
     {otherUnit_maskInput_lo[5263:5248]},
     {otherUnit_maskInput_lo[5247:5232]},
     {otherUnit_maskInput_lo[5231:5216]},
     {otherUnit_maskInput_lo[5215:5200]},
     {otherUnit_maskInput_lo[5199:5184]},
     {otherUnit_maskInput_lo[5183:5168]},
     {otherUnit_maskInput_lo[5167:5152]},
     {otherUnit_maskInput_lo[5151:5136]},
     {otherUnit_maskInput_lo[5135:5120]},
     {otherUnit_maskInput_lo[5119:5104]},
     {otherUnit_maskInput_lo[5103:5088]},
     {otherUnit_maskInput_lo[5087:5072]},
     {otherUnit_maskInput_lo[5071:5056]},
     {otherUnit_maskInput_lo[5055:5040]},
     {otherUnit_maskInput_lo[5039:5024]},
     {otherUnit_maskInput_lo[5023:5008]},
     {otherUnit_maskInput_lo[5007:4992]},
     {otherUnit_maskInput_lo[4991:4976]},
     {otherUnit_maskInput_lo[4975:4960]},
     {otherUnit_maskInput_lo[4959:4944]},
     {otherUnit_maskInput_lo[4943:4928]},
     {otherUnit_maskInput_lo[4927:4912]},
     {otherUnit_maskInput_lo[4911:4896]},
     {otherUnit_maskInput_lo[4895:4880]},
     {otherUnit_maskInput_lo[4879:4864]},
     {otherUnit_maskInput_lo[4863:4848]},
     {otherUnit_maskInput_lo[4847:4832]},
     {otherUnit_maskInput_lo[4831:4816]},
     {otherUnit_maskInput_lo[4815:4800]},
     {otherUnit_maskInput_lo[4799:4784]},
     {otherUnit_maskInput_lo[4783:4768]},
     {otherUnit_maskInput_lo[4767:4752]},
     {otherUnit_maskInput_lo[4751:4736]},
     {otherUnit_maskInput_lo[4735:4720]},
     {otherUnit_maskInput_lo[4719:4704]},
     {otherUnit_maskInput_lo[4703:4688]},
     {otherUnit_maskInput_lo[4687:4672]},
     {otherUnit_maskInput_lo[4671:4656]},
     {otherUnit_maskInput_lo[4655:4640]},
     {otherUnit_maskInput_lo[4639:4624]},
     {otherUnit_maskInput_lo[4623:4608]},
     {otherUnit_maskInput_lo[4607:4592]},
     {otherUnit_maskInput_lo[4591:4576]},
     {otherUnit_maskInput_lo[4575:4560]},
     {otherUnit_maskInput_lo[4559:4544]},
     {otherUnit_maskInput_lo[4543:4528]},
     {otherUnit_maskInput_lo[4527:4512]},
     {otherUnit_maskInput_lo[4511:4496]},
     {otherUnit_maskInput_lo[4495:4480]},
     {otherUnit_maskInput_lo[4479:4464]},
     {otherUnit_maskInput_lo[4463:4448]},
     {otherUnit_maskInput_lo[4447:4432]},
     {otherUnit_maskInput_lo[4431:4416]},
     {otherUnit_maskInput_lo[4415:4400]},
     {otherUnit_maskInput_lo[4399:4384]},
     {otherUnit_maskInput_lo[4383:4368]},
     {otherUnit_maskInput_lo[4367:4352]},
     {otherUnit_maskInput_lo[4351:4336]},
     {otherUnit_maskInput_lo[4335:4320]},
     {otherUnit_maskInput_lo[4319:4304]},
     {otherUnit_maskInput_lo[4303:4288]},
     {otherUnit_maskInput_lo[4287:4272]},
     {otherUnit_maskInput_lo[4271:4256]},
     {otherUnit_maskInput_lo[4255:4240]},
     {otherUnit_maskInput_lo[4239:4224]},
     {otherUnit_maskInput_lo[4223:4208]},
     {otherUnit_maskInput_lo[4207:4192]},
     {otherUnit_maskInput_lo[4191:4176]},
     {otherUnit_maskInput_lo[4175:4160]},
     {otherUnit_maskInput_lo[4159:4144]},
     {otherUnit_maskInput_lo[4143:4128]},
     {otherUnit_maskInput_lo[4127:4112]},
     {otherUnit_maskInput_lo[4111:4096]},
     {otherUnit_maskInput_lo[4095:4080]},
     {otherUnit_maskInput_lo[4079:4064]},
     {otherUnit_maskInput_lo[4063:4048]},
     {otherUnit_maskInput_lo[4047:4032]},
     {otherUnit_maskInput_lo[4031:4016]},
     {otherUnit_maskInput_lo[4015:4000]},
     {otherUnit_maskInput_lo[3999:3984]},
     {otherUnit_maskInput_lo[3983:3968]},
     {otherUnit_maskInput_lo[3967:3952]},
     {otherUnit_maskInput_lo[3951:3936]},
     {otherUnit_maskInput_lo[3935:3920]},
     {otherUnit_maskInput_lo[3919:3904]},
     {otherUnit_maskInput_lo[3903:3888]},
     {otherUnit_maskInput_lo[3887:3872]},
     {otherUnit_maskInput_lo[3871:3856]},
     {otherUnit_maskInput_lo[3855:3840]},
     {otherUnit_maskInput_lo[3839:3824]},
     {otherUnit_maskInput_lo[3823:3808]},
     {otherUnit_maskInput_lo[3807:3792]},
     {otherUnit_maskInput_lo[3791:3776]},
     {otherUnit_maskInput_lo[3775:3760]},
     {otherUnit_maskInput_lo[3759:3744]},
     {otherUnit_maskInput_lo[3743:3728]},
     {otherUnit_maskInput_lo[3727:3712]},
     {otherUnit_maskInput_lo[3711:3696]},
     {otherUnit_maskInput_lo[3695:3680]},
     {otherUnit_maskInput_lo[3679:3664]},
     {otherUnit_maskInput_lo[3663:3648]},
     {otherUnit_maskInput_lo[3647:3632]},
     {otherUnit_maskInput_lo[3631:3616]},
     {otherUnit_maskInput_lo[3615:3600]},
     {otherUnit_maskInput_lo[3599:3584]},
     {otherUnit_maskInput_lo[3583:3568]},
     {otherUnit_maskInput_lo[3567:3552]},
     {otherUnit_maskInput_lo[3551:3536]},
     {otherUnit_maskInput_lo[3535:3520]},
     {otherUnit_maskInput_lo[3519:3504]},
     {otherUnit_maskInput_lo[3503:3488]},
     {otherUnit_maskInput_lo[3487:3472]},
     {otherUnit_maskInput_lo[3471:3456]},
     {otherUnit_maskInput_lo[3455:3440]},
     {otherUnit_maskInput_lo[3439:3424]},
     {otherUnit_maskInput_lo[3423:3408]},
     {otherUnit_maskInput_lo[3407:3392]},
     {otherUnit_maskInput_lo[3391:3376]},
     {otherUnit_maskInput_lo[3375:3360]},
     {otherUnit_maskInput_lo[3359:3344]},
     {otherUnit_maskInput_lo[3343:3328]},
     {otherUnit_maskInput_lo[3327:3312]},
     {otherUnit_maskInput_lo[3311:3296]},
     {otherUnit_maskInput_lo[3295:3280]},
     {otherUnit_maskInput_lo[3279:3264]},
     {otherUnit_maskInput_lo[3263:3248]},
     {otherUnit_maskInput_lo[3247:3232]},
     {otherUnit_maskInput_lo[3231:3216]},
     {otherUnit_maskInput_lo[3215:3200]},
     {otherUnit_maskInput_lo[3199:3184]},
     {otherUnit_maskInput_lo[3183:3168]},
     {otherUnit_maskInput_lo[3167:3152]},
     {otherUnit_maskInput_lo[3151:3136]},
     {otherUnit_maskInput_lo[3135:3120]},
     {otherUnit_maskInput_lo[3119:3104]},
     {otherUnit_maskInput_lo[3103:3088]},
     {otherUnit_maskInput_lo[3087:3072]},
     {otherUnit_maskInput_lo[3071:3056]},
     {otherUnit_maskInput_lo[3055:3040]},
     {otherUnit_maskInput_lo[3039:3024]},
     {otherUnit_maskInput_lo[3023:3008]},
     {otherUnit_maskInput_lo[3007:2992]},
     {otherUnit_maskInput_lo[2991:2976]},
     {otherUnit_maskInput_lo[2975:2960]},
     {otherUnit_maskInput_lo[2959:2944]},
     {otherUnit_maskInput_lo[2943:2928]},
     {otherUnit_maskInput_lo[2927:2912]},
     {otherUnit_maskInput_lo[2911:2896]},
     {otherUnit_maskInput_lo[2895:2880]},
     {otherUnit_maskInput_lo[2879:2864]},
     {otherUnit_maskInput_lo[2863:2848]},
     {otherUnit_maskInput_lo[2847:2832]},
     {otherUnit_maskInput_lo[2831:2816]},
     {otherUnit_maskInput_lo[2815:2800]},
     {otherUnit_maskInput_lo[2799:2784]},
     {otherUnit_maskInput_lo[2783:2768]},
     {otherUnit_maskInput_lo[2767:2752]},
     {otherUnit_maskInput_lo[2751:2736]},
     {otherUnit_maskInput_lo[2735:2720]},
     {otherUnit_maskInput_lo[2719:2704]},
     {otherUnit_maskInput_lo[2703:2688]},
     {otherUnit_maskInput_lo[2687:2672]},
     {otherUnit_maskInput_lo[2671:2656]},
     {otherUnit_maskInput_lo[2655:2640]},
     {otherUnit_maskInput_lo[2639:2624]},
     {otherUnit_maskInput_lo[2623:2608]},
     {otherUnit_maskInput_lo[2607:2592]},
     {otherUnit_maskInput_lo[2591:2576]},
     {otherUnit_maskInput_lo[2575:2560]},
     {otherUnit_maskInput_lo[2559:2544]},
     {otherUnit_maskInput_lo[2543:2528]},
     {otherUnit_maskInput_lo[2527:2512]},
     {otherUnit_maskInput_lo[2511:2496]},
     {otherUnit_maskInput_lo[2495:2480]},
     {otherUnit_maskInput_lo[2479:2464]},
     {otherUnit_maskInput_lo[2463:2448]},
     {otherUnit_maskInput_lo[2447:2432]},
     {otherUnit_maskInput_lo[2431:2416]},
     {otherUnit_maskInput_lo[2415:2400]},
     {otherUnit_maskInput_lo[2399:2384]},
     {otherUnit_maskInput_lo[2383:2368]},
     {otherUnit_maskInput_lo[2367:2352]},
     {otherUnit_maskInput_lo[2351:2336]},
     {otherUnit_maskInput_lo[2335:2320]},
     {otherUnit_maskInput_lo[2319:2304]},
     {otherUnit_maskInput_lo[2303:2288]},
     {otherUnit_maskInput_lo[2287:2272]},
     {otherUnit_maskInput_lo[2271:2256]},
     {otherUnit_maskInput_lo[2255:2240]},
     {otherUnit_maskInput_lo[2239:2224]},
     {otherUnit_maskInput_lo[2223:2208]},
     {otherUnit_maskInput_lo[2207:2192]},
     {otherUnit_maskInput_lo[2191:2176]},
     {otherUnit_maskInput_lo[2175:2160]},
     {otherUnit_maskInput_lo[2159:2144]},
     {otherUnit_maskInput_lo[2143:2128]},
     {otherUnit_maskInput_lo[2127:2112]},
     {otherUnit_maskInput_lo[2111:2096]},
     {otherUnit_maskInput_lo[2095:2080]},
     {otherUnit_maskInput_lo[2079:2064]},
     {otherUnit_maskInput_lo[2063:2048]},
     {otherUnit_maskInput_lo[2047:2032]},
     {otherUnit_maskInput_lo[2031:2016]},
     {otherUnit_maskInput_lo[2015:2000]},
     {otherUnit_maskInput_lo[1999:1984]},
     {otherUnit_maskInput_lo[1983:1968]},
     {otherUnit_maskInput_lo[1967:1952]},
     {otherUnit_maskInput_lo[1951:1936]},
     {otherUnit_maskInput_lo[1935:1920]},
     {otherUnit_maskInput_lo[1919:1904]},
     {otherUnit_maskInput_lo[1903:1888]},
     {otherUnit_maskInput_lo[1887:1872]},
     {otherUnit_maskInput_lo[1871:1856]},
     {otherUnit_maskInput_lo[1855:1840]},
     {otherUnit_maskInput_lo[1839:1824]},
     {otherUnit_maskInput_lo[1823:1808]},
     {otherUnit_maskInput_lo[1807:1792]},
     {otherUnit_maskInput_lo[1791:1776]},
     {otherUnit_maskInput_lo[1775:1760]},
     {otherUnit_maskInput_lo[1759:1744]},
     {otherUnit_maskInput_lo[1743:1728]},
     {otherUnit_maskInput_lo[1727:1712]},
     {otherUnit_maskInput_lo[1711:1696]},
     {otherUnit_maskInput_lo[1695:1680]},
     {otherUnit_maskInput_lo[1679:1664]},
     {otherUnit_maskInput_lo[1663:1648]},
     {otherUnit_maskInput_lo[1647:1632]},
     {otherUnit_maskInput_lo[1631:1616]},
     {otherUnit_maskInput_lo[1615:1600]},
     {otherUnit_maskInput_lo[1599:1584]},
     {otherUnit_maskInput_lo[1583:1568]},
     {otherUnit_maskInput_lo[1567:1552]},
     {otherUnit_maskInput_lo[1551:1536]},
     {otherUnit_maskInput_lo[1535:1520]},
     {otherUnit_maskInput_lo[1519:1504]},
     {otherUnit_maskInput_lo[1503:1488]},
     {otherUnit_maskInput_lo[1487:1472]},
     {otherUnit_maskInput_lo[1471:1456]},
     {otherUnit_maskInput_lo[1455:1440]},
     {otherUnit_maskInput_lo[1439:1424]},
     {otherUnit_maskInput_lo[1423:1408]},
     {otherUnit_maskInput_lo[1407:1392]},
     {otherUnit_maskInput_lo[1391:1376]},
     {otherUnit_maskInput_lo[1375:1360]},
     {otherUnit_maskInput_lo[1359:1344]},
     {otherUnit_maskInput_lo[1343:1328]},
     {otherUnit_maskInput_lo[1327:1312]},
     {otherUnit_maskInput_lo[1311:1296]},
     {otherUnit_maskInput_lo[1295:1280]},
     {otherUnit_maskInput_lo[1279:1264]},
     {otherUnit_maskInput_lo[1263:1248]},
     {otherUnit_maskInput_lo[1247:1232]},
     {otherUnit_maskInput_lo[1231:1216]},
     {otherUnit_maskInput_lo[1215:1200]},
     {otherUnit_maskInput_lo[1199:1184]},
     {otherUnit_maskInput_lo[1183:1168]},
     {otherUnit_maskInput_lo[1167:1152]},
     {otherUnit_maskInput_lo[1151:1136]},
     {otherUnit_maskInput_lo[1135:1120]},
     {otherUnit_maskInput_lo[1119:1104]},
     {otherUnit_maskInput_lo[1103:1088]},
     {otherUnit_maskInput_lo[1087:1072]},
     {otherUnit_maskInput_lo[1071:1056]},
     {otherUnit_maskInput_lo[1055:1040]},
     {otherUnit_maskInput_lo[1039:1024]},
     {otherUnit_maskInput_lo[1023:1008]},
     {otherUnit_maskInput_lo[1007:992]},
     {otherUnit_maskInput_lo[991:976]},
     {otherUnit_maskInput_lo[975:960]},
     {otherUnit_maskInput_lo[959:944]},
     {otherUnit_maskInput_lo[943:928]},
     {otherUnit_maskInput_lo[927:912]},
     {otherUnit_maskInput_lo[911:896]},
     {otherUnit_maskInput_lo[895:880]},
     {otherUnit_maskInput_lo[879:864]},
     {otherUnit_maskInput_lo[863:848]},
     {otherUnit_maskInput_lo[847:832]},
     {otherUnit_maskInput_lo[831:816]},
     {otherUnit_maskInput_lo[815:800]},
     {otherUnit_maskInput_lo[799:784]},
     {otherUnit_maskInput_lo[783:768]},
     {otherUnit_maskInput_lo[767:752]},
     {otherUnit_maskInput_lo[751:736]},
     {otherUnit_maskInput_lo[735:720]},
     {otherUnit_maskInput_lo[719:704]},
     {otherUnit_maskInput_lo[703:688]},
     {otherUnit_maskInput_lo[687:672]},
     {otherUnit_maskInput_lo[671:656]},
     {otherUnit_maskInput_lo[655:640]},
     {otherUnit_maskInput_lo[639:624]},
     {otherUnit_maskInput_lo[623:608]},
     {otherUnit_maskInput_lo[607:592]},
     {otherUnit_maskInput_lo[591:576]},
     {otherUnit_maskInput_lo[575:560]},
     {otherUnit_maskInput_lo[559:544]},
     {otherUnit_maskInput_lo[543:528]},
     {otherUnit_maskInput_lo[527:512]},
     {otherUnit_maskInput_lo[511:496]},
     {otherUnit_maskInput_lo[495:480]},
     {otherUnit_maskInput_lo[479:464]},
     {otherUnit_maskInput_lo[463:448]},
     {otherUnit_maskInput_lo[447:432]},
     {otherUnit_maskInput_lo[431:416]},
     {otherUnit_maskInput_lo[415:400]},
     {otherUnit_maskInput_lo[399:384]},
     {otherUnit_maskInput_lo[383:368]},
     {otherUnit_maskInput_lo[367:352]},
     {otherUnit_maskInput_lo[351:336]},
     {otherUnit_maskInput_lo[335:320]},
     {otherUnit_maskInput_lo[319:304]},
     {otherUnit_maskInput_lo[303:288]},
     {otherUnit_maskInput_lo[287:272]},
     {otherUnit_maskInput_lo[271:256]},
     {otherUnit_maskInput_lo[255:240]},
     {otherUnit_maskInput_lo[239:224]},
     {otherUnit_maskInput_lo[223:208]},
     {otherUnit_maskInput_lo[207:192]},
     {otherUnit_maskInput_lo[191:176]},
     {otherUnit_maskInput_lo[175:160]},
     {otherUnit_maskInput_lo[159:144]},
     {otherUnit_maskInput_lo[143:128]},
     {otherUnit_maskInput_lo[127:112]},
     {otherUnit_maskInput_lo[111:96]},
     {otherUnit_maskInput_lo[95:80]},
     {otherUnit_maskInput_lo[79:64]},
     {otherUnit_maskInput_lo[63:48]},
     {otherUnit_maskInput_lo[47:32]},
     {otherUnit_maskInput_lo[31:16]},
     {otherUnit_maskInput_lo[15:0]}};
  wire                vrfWritePort_0_valid_0 = writeQueueVec_0_deq_valid;
  wire [4:0]          vrfWritePort_0_bits_vd_0 = writeQueueVec_0_deq_bits_data_vd;
  wire [7:0]          vrfWritePort_0_bits_offset_0 = writeQueueVec_0_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_0_bits_mask_0 = writeQueueVec_0_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_0_bits_data_0 = writeQueueVec_0_deq_bits_data_data;
  wire                vrfWritePort_0_bits_last_0 = writeQueueVec_0_deq_bits_data_last;
  wire [2:0]          vrfWritePort_0_bits_instructionIndex_0 = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_enq_bits = writeQueueVec_0_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_0_enq_bits_data_data;
  wire                writeQueueVec_0_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi = {writeQueueVec_0_enq_bits_data_data, writeQueueVec_0_enq_bits_data_last};
  wire [2:0]          writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo = {writeQueueVec_dataIn_lo_hi, writeQueueVec_0_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_0_enq_bits_data_vd;
  wire [7:0]          writeQueueVec_0_enq_bits_data_offset;
  wire [12:0]         writeQueueVec_dataIn_hi_hi = {writeQueueVec_0_enq_bits_data_vd, writeQueueVec_0_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_0_enq_bits_data_mask;
  wire [16:0]         writeQueueVec_dataIn_hi = {writeQueueVec_dataIn_hi_hi, writeQueueVec_0_enq_bits_data_mask};
  wire [56:0]         writeQueueVec_dataIn = {writeQueueVec_dataIn_hi, writeQueueVec_dataIn_lo, 4'h1};
  wire [3:0]          writeQueueVec_dataOut_targetLane = _writeQueueVec_fifo_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_data_instructionIndex = _writeQueueVec_fifo_data_out[6:4];
  wire                writeQueueVec_dataOut_data_last = _writeQueueVec_fifo_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_data_data = _writeQueueVec_fifo_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_data_mask = _writeQueueVec_fifo_data_out[43:40];
  wire [7:0]          writeQueueVec_dataOut_data_offset = _writeQueueVec_fifo_data_out[51:44];
  wire [4:0]          writeQueueVec_dataOut_data_vd = _writeQueueVec_fifo_data_out[56:52];
  wire                writeQueueVec_0_enq_ready = ~_writeQueueVec_fifo_full;
  wire                writeQueueVec_0_enq_valid;
  wire                _probeWire_slots_0_writeValid_T = writeQueueVec_0_enq_ready & writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_valid = ~_writeQueueVec_fifo_empty | writeQueueVec_0_enq_valid;
  assign writeQueueVec_0_deq_bits_data_vd = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_vd : writeQueueVec_dataOut_data_vd;
  assign writeQueueVec_0_deq_bits_data_offset = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_offset : writeQueueVec_dataOut_data_offset;
  assign writeQueueVec_0_deq_bits_data_mask = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_mask : writeQueueVec_dataOut_data_mask;
  assign writeQueueVec_0_deq_bits_data_data = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_data : writeQueueVec_dataOut_data_data;
  assign writeQueueVec_0_deq_bits_data_last = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_last : writeQueueVec_dataOut_data_last;
  assign writeQueueVec_0_deq_bits_data_instructionIndex = _writeQueueVec_fifo_empty ? writeQueueVec_0_enq_bits_data_instructionIndex : writeQueueVec_dataOut_data_instructionIndex;
  wire [3:0]          writeQueueVec_0_deq_bits_targetLane = _writeQueueVec_fifo_empty ? 4'h1 : writeQueueVec_dataOut_targetLane;
  wire                vrfWritePort_1_valid_0 = writeQueueVec_1_deq_valid;
  wire [4:0]          vrfWritePort_1_bits_vd_0 = writeQueueVec_1_deq_bits_data_vd;
  wire [7:0]          vrfWritePort_1_bits_offset_0 = writeQueueVec_1_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_1_bits_mask_0 = writeQueueVec_1_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_1_bits_data_0 = writeQueueVec_1_deq_bits_data_data;
  wire                vrfWritePort_1_bits_last_0 = writeQueueVec_1_deq_bits_data_last;
  wire [2:0]          vrfWritePort_1_bits_instructionIndex_0 = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_1_enq_bits = writeQueueVec_1_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_1_enq_bits_data_data;
  wire                writeQueueVec_1_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi_1 = {writeQueueVec_1_enq_bits_data_data, writeQueueVec_1_enq_bits_data_last};
  wire [2:0]          writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo_1 = {writeQueueVec_dataIn_lo_hi_1, writeQueueVec_1_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_1_enq_bits_data_vd;
  wire [7:0]          writeQueueVec_1_enq_bits_data_offset;
  wire [12:0]         writeQueueVec_dataIn_hi_hi_1 = {writeQueueVec_1_enq_bits_data_vd, writeQueueVec_1_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_1_enq_bits_data_mask;
  wire [16:0]         writeQueueVec_dataIn_hi_1 = {writeQueueVec_dataIn_hi_hi_1, writeQueueVec_1_enq_bits_data_mask};
  wire [56:0]         writeQueueVec_dataIn_1 = {writeQueueVec_dataIn_hi_1, writeQueueVec_dataIn_lo_1, 4'h2};
  wire [3:0]          writeQueueVec_dataOut_1_targetLane = _writeQueueVec_fifo_1_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_1_data_instructionIndex = _writeQueueVec_fifo_1_data_out[6:4];
  wire                writeQueueVec_dataOut_1_data_last = _writeQueueVec_fifo_1_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_1_data_data = _writeQueueVec_fifo_1_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_1_data_mask = _writeQueueVec_fifo_1_data_out[43:40];
  wire [7:0]          writeQueueVec_dataOut_1_data_offset = _writeQueueVec_fifo_1_data_out[51:44];
  wire [4:0]          writeQueueVec_dataOut_1_data_vd = _writeQueueVec_fifo_1_data_out[56:52];
  wire                writeQueueVec_1_enq_ready = ~_writeQueueVec_fifo_1_full;
  wire                writeQueueVec_1_enq_valid;
  wire                _probeWire_slots_1_writeValid_T = writeQueueVec_1_enq_ready & writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_valid = ~_writeQueueVec_fifo_1_empty | writeQueueVec_1_enq_valid;
  assign writeQueueVec_1_deq_bits_data_vd = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_vd : writeQueueVec_dataOut_1_data_vd;
  assign writeQueueVec_1_deq_bits_data_offset = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_offset : writeQueueVec_dataOut_1_data_offset;
  assign writeQueueVec_1_deq_bits_data_mask = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_mask : writeQueueVec_dataOut_1_data_mask;
  assign writeQueueVec_1_deq_bits_data_data = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_data : writeQueueVec_dataOut_1_data_data;
  assign writeQueueVec_1_deq_bits_data_last = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_last : writeQueueVec_dataOut_1_data_last;
  assign writeQueueVec_1_deq_bits_data_instructionIndex = _writeQueueVec_fifo_1_empty ? writeQueueVec_1_enq_bits_data_instructionIndex : writeQueueVec_dataOut_1_data_instructionIndex;
  wire [3:0]          writeQueueVec_1_deq_bits_targetLane = _writeQueueVec_fifo_1_empty ? 4'h2 : writeQueueVec_dataOut_1_targetLane;
  wire                vrfWritePort_2_valid_0 = writeQueueVec_2_deq_valid;
  wire [4:0]          vrfWritePort_2_bits_vd_0 = writeQueueVec_2_deq_bits_data_vd;
  wire [7:0]          vrfWritePort_2_bits_offset_0 = writeQueueVec_2_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_2_bits_mask_0 = writeQueueVec_2_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_2_bits_data_0 = writeQueueVec_2_deq_bits_data_data;
  wire                vrfWritePort_2_bits_last_0 = writeQueueVec_2_deq_bits_data_last;
  wire [2:0]          vrfWritePort_2_bits_instructionIndex_0 = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_2_enq_bits = writeQueueVec_2_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_2_enq_bits_data_data;
  wire                writeQueueVec_2_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi_2 = {writeQueueVec_2_enq_bits_data_data, writeQueueVec_2_enq_bits_data_last};
  wire [2:0]          writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo_2 = {writeQueueVec_dataIn_lo_hi_2, writeQueueVec_2_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_2_enq_bits_data_vd;
  wire [7:0]          writeQueueVec_2_enq_bits_data_offset;
  wire [12:0]         writeQueueVec_dataIn_hi_hi_2 = {writeQueueVec_2_enq_bits_data_vd, writeQueueVec_2_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_2_enq_bits_data_mask;
  wire [16:0]         writeQueueVec_dataIn_hi_2 = {writeQueueVec_dataIn_hi_hi_2, writeQueueVec_2_enq_bits_data_mask};
  wire [56:0]         writeQueueVec_dataIn_2 = {writeQueueVec_dataIn_hi_2, writeQueueVec_dataIn_lo_2, 4'h4};
  wire [3:0]          writeQueueVec_dataOut_2_targetLane = _writeQueueVec_fifo_2_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_2_data_instructionIndex = _writeQueueVec_fifo_2_data_out[6:4];
  wire                writeQueueVec_dataOut_2_data_last = _writeQueueVec_fifo_2_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_2_data_data = _writeQueueVec_fifo_2_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_2_data_mask = _writeQueueVec_fifo_2_data_out[43:40];
  wire [7:0]          writeQueueVec_dataOut_2_data_offset = _writeQueueVec_fifo_2_data_out[51:44];
  wire [4:0]          writeQueueVec_dataOut_2_data_vd = _writeQueueVec_fifo_2_data_out[56:52];
  wire                writeQueueVec_2_enq_ready = ~_writeQueueVec_fifo_2_full;
  wire                writeQueueVec_2_enq_valid;
  wire                _probeWire_slots_2_writeValid_T = writeQueueVec_2_enq_ready & writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_valid = ~_writeQueueVec_fifo_2_empty | writeQueueVec_2_enq_valid;
  assign writeQueueVec_2_deq_bits_data_vd = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_vd : writeQueueVec_dataOut_2_data_vd;
  assign writeQueueVec_2_deq_bits_data_offset = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_offset : writeQueueVec_dataOut_2_data_offset;
  assign writeQueueVec_2_deq_bits_data_mask = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_mask : writeQueueVec_dataOut_2_data_mask;
  assign writeQueueVec_2_deq_bits_data_data = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_data : writeQueueVec_dataOut_2_data_data;
  assign writeQueueVec_2_deq_bits_data_last = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_last : writeQueueVec_dataOut_2_data_last;
  assign writeQueueVec_2_deq_bits_data_instructionIndex = _writeQueueVec_fifo_2_empty ? writeQueueVec_2_enq_bits_data_instructionIndex : writeQueueVec_dataOut_2_data_instructionIndex;
  wire [3:0]          writeQueueVec_2_deq_bits_targetLane = _writeQueueVec_fifo_2_empty ? 4'h4 : writeQueueVec_dataOut_2_targetLane;
  wire                vrfWritePort_3_valid_0 = writeQueueVec_3_deq_valid;
  wire [4:0]          vrfWritePort_3_bits_vd_0 = writeQueueVec_3_deq_bits_data_vd;
  wire [7:0]          vrfWritePort_3_bits_offset_0 = writeQueueVec_3_deq_bits_data_offset;
  wire [3:0]          vrfWritePort_3_bits_mask_0 = writeQueueVec_3_deq_bits_data_mask;
  wire [31:0]         vrfWritePort_3_bits_data_0 = writeQueueVec_3_deq_bits_data_data;
  wire                vrfWritePort_3_bits_last_0 = writeQueueVec_3_deq_bits_data_last;
  wire [2:0]          vrfWritePort_3_bits_instructionIndex_0 = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [2:0]          writeIndexQueue_3_enq_bits = writeQueueVec_3_deq_bits_data_instructionIndex;
  wire [31:0]         writeQueueVec_3_enq_bits_data_data;
  wire                writeQueueVec_3_enq_bits_data_last;
  wire [32:0]         writeQueueVec_dataIn_lo_hi_3 = {writeQueueVec_3_enq_bits_data_data, writeQueueVec_3_enq_bits_data_last};
  wire [2:0]          writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [35:0]         writeQueueVec_dataIn_lo_3 = {writeQueueVec_dataIn_lo_hi_3, writeQueueVec_3_enq_bits_data_instructionIndex};
  wire [4:0]          writeQueueVec_3_enq_bits_data_vd;
  wire [7:0]          writeQueueVec_3_enq_bits_data_offset;
  wire [12:0]         writeQueueVec_dataIn_hi_hi_3 = {writeQueueVec_3_enq_bits_data_vd, writeQueueVec_3_enq_bits_data_offset};
  wire [3:0]          writeQueueVec_3_enq_bits_data_mask;
  wire [16:0]         writeQueueVec_dataIn_hi_3 = {writeQueueVec_dataIn_hi_hi_3, writeQueueVec_3_enq_bits_data_mask};
  wire [56:0]         writeQueueVec_dataIn_3 = {writeQueueVec_dataIn_hi_3, writeQueueVec_dataIn_lo_3, 4'h8};
  wire [3:0]          writeQueueVec_dataOut_3_targetLane = _writeQueueVec_fifo_3_data_out[3:0];
  wire [2:0]          writeQueueVec_dataOut_3_data_instructionIndex = _writeQueueVec_fifo_3_data_out[6:4];
  wire                writeQueueVec_dataOut_3_data_last = _writeQueueVec_fifo_3_data_out[7];
  wire [31:0]         writeQueueVec_dataOut_3_data_data = _writeQueueVec_fifo_3_data_out[39:8];
  wire [3:0]          writeQueueVec_dataOut_3_data_mask = _writeQueueVec_fifo_3_data_out[43:40];
  wire [7:0]          writeQueueVec_dataOut_3_data_offset = _writeQueueVec_fifo_3_data_out[51:44];
  wire [4:0]          writeQueueVec_dataOut_3_data_vd = _writeQueueVec_fifo_3_data_out[56:52];
  wire                writeQueueVec_3_enq_ready = ~_writeQueueVec_fifo_3_full;
  wire                writeQueueVec_3_enq_valid;
  wire                _probeWire_slots_3_writeValid_T = writeQueueVec_3_enq_ready & writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_valid = ~_writeQueueVec_fifo_3_empty | writeQueueVec_3_enq_valid;
  assign writeQueueVec_3_deq_bits_data_vd = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_vd : writeQueueVec_dataOut_3_data_vd;
  assign writeQueueVec_3_deq_bits_data_offset = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_offset : writeQueueVec_dataOut_3_data_offset;
  assign writeQueueVec_3_deq_bits_data_mask = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_mask : writeQueueVec_dataOut_3_data_mask;
  assign writeQueueVec_3_deq_bits_data_data = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_data : writeQueueVec_dataOut_3_data_data;
  assign writeQueueVec_3_deq_bits_data_last = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_last : writeQueueVec_dataOut_3_data_last;
  assign writeQueueVec_3_deq_bits_data_instructionIndex = _writeQueueVec_fifo_3_empty ? writeQueueVec_3_enq_bits_data_instructionIndex : writeQueueVec_dataOut_3_data_instructionIndex;
  wire [3:0]          writeQueueVec_3_deq_bits_targetLane = _writeQueueVec_fifo_3_empty ? 4'h8 : writeQueueVec_dataOut_3_targetLane;
  wire                otherUnitTargetQueue_deq_valid;
  assign otherUnitTargetQueue_deq_valid = ~_otherUnitTargetQueue_fifo_empty;
  wire                otherUnitTargetQueue_deq_ready;
  wire                otherUnitTargetQueue_enq_ready = ~_otherUnitTargetQueue_fifo_full | otherUnitTargetQueue_deq_ready;
  wire                otherUnitTargetQueue_enq_valid;
  wire                otherUnitDataQueueVec_0_enq_ready = ~_otherUnitDataQueueVec_fifo_full;
  wire                otherUnitDataQueueVec_0_deq_ready;
  wire                otherUnitDataQueueVec_0_enq_valid;
  wire                otherUnitDataQueueVec_0_deq_valid = ~_otherUnitDataQueueVec_fifo_empty | otherUnitDataQueueVec_0_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_0_deq_bits = _otherUnitDataQueueVec_fifo_empty ? otherUnitDataQueueVec_0_enq_bits : _otherUnitDataQueueVec_fifo_data_out;
  wire                otherUnitDataQueueVec_1_enq_ready = ~_otherUnitDataQueueVec_fifo_1_full;
  wire                otherUnitDataQueueVec_1_deq_ready;
  wire                otherUnitDataQueueVec_1_enq_valid;
  wire                otherUnitDataQueueVec_1_deq_valid = ~_otherUnitDataQueueVec_fifo_1_empty | otherUnitDataQueueVec_1_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_1_deq_bits = _otherUnitDataQueueVec_fifo_1_empty ? otherUnitDataQueueVec_1_enq_bits : _otherUnitDataQueueVec_fifo_1_data_out;
  wire                otherUnitDataQueueVec_2_enq_ready = ~_otherUnitDataQueueVec_fifo_2_full;
  wire                otherUnitDataQueueVec_2_deq_ready;
  wire                otherUnitDataQueueVec_2_enq_valid;
  wire                otherUnitDataQueueVec_2_deq_valid = ~_otherUnitDataQueueVec_fifo_2_empty | otherUnitDataQueueVec_2_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_2_deq_bits = _otherUnitDataQueueVec_fifo_2_empty ? otherUnitDataQueueVec_2_enq_bits : _otherUnitDataQueueVec_fifo_2_data_out;
  wire                otherUnitDataQueueVec_3_enq_ready = ~_otherUnitDataQueueVec_fifo_3_full;
  wire                otherUnitDataQueueVec_3_deq_ready;
  wire                otherUnitDataQueueVec_3_enq_valid;
  wire                otherUnitDataQueueVec_3_deq_valid = ~_otherUnitDataQueueVec_fifo_3_empty | otherUnitDataQueueVec_3_enq_valid;
  wire [31:0]         otherUnitDataQueueVec_3_deq_bits = _otherUnitDataQueueVec_fifo_3_empty ? otherUnitDataQueueVec_3_enq_bits : _otherUnitDataQueueVec_fifo_3_data_out;
  wire [3:0]          otherTryReadVrf = _otherUnit_vrfReadDataPorts_valid ? _otherUnit_status_targetLane : 4'h0;
  wire                vrfReadDataPorts_0_valid_0 = otherTryReadVrf[0] | _storeUnit_vrfReadDataPorts_0_valid;
  wire [4:0]          vrfReadDataPorts_0_bits_vs_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_0_bits_vs;
  wire [7:0]          vrfReadDataPorts_0_bits_offset_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_0_bits_offset;
  wire [2:0]          vrfReadDataPorts_0_bits_instructionIndex_0 = otherTryReadVrf[0] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_0_bits_instructionIndex;
  wire                otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_0_enq_valid = vrfReadResults_0_valid & ~otherUnitTargetQueue_empty;
  wire [3:0]          dataDeqFire;
  assign otherUnitDataQueueVec_0_deq_ready = dataDeqFire[0];
  wire                vrfReadDataPorts_1_valid_0 = otherTryReadVrf[1] | _storeUnit_vrfReadDataPorts_1_valid;
  wire [4:0]          vrfReadDataPorts_1_bits_vs_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_1_bits_vs;
  wire [7:0]          vrfReadDataPorts_1_bits_offset_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_1_bits_offset;
  wire [2:0]          vrfReadDataPorts_1_bits_instructionIndex_0 = otherTryReadVrf[1] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_1_bits_instructionIndex;
  assign otherUnitDataQueueVec_1_enq_valid = vrfReadResults_1_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_1_deq_ready = dataDeqFire[1];
  wire                vrfReadDataPorts_2_valid_0 = otherTryReadVrf[2] | _storeUnit_vrfReadDataPorts_2_valid;
  wire [4:0]          vrfReadDataPorts_2_bits_vs_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_2_bits_vs;
  wire [7:0]          vrfReadDataPorts_2_bits_offset_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_2_bits_offset;
  wire [2:0]          vrfReadDataPorts_2_bits_instructionIndex_0 = otherTryReadVrf[2] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_2_bits_instructionIndex;
  assign otherUnitDataQueueVec_2_enq_valid = vrfReadResults_2_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_2_deq_ready = dataDeqFire[2];
  wire                vrfReadDataPorts_3_valid_0 = otherTryReadVrf[3] | _storeUnit_vrfReadDataPorts_3_valid;
  wire [4:0]          vrfReadDataPorts_3_bits_vs_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_vs : _storeUnit_vrfReadDataPorts_3_bits_vs;
  wire [7:0]          vrfReadDataPorts_3_bits_offset_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_offset : _storeUnit_vrfReadDataPorts_3_bits_offset;
  wire [2:0]          vrfReadDataPorts_3_bits_instructionIndex_0 = otherTryReadVrf[3] ? _otherUnit_vrfReadDataPorts_bits_instructionIndex : _storeUnit_vrfReadDataPorts_3_bits_instructionIndex;
  assign otherUnitDataQueueVec_3_enq_valid = vrfReadResults_3_valid & ~otherUnitTargetQueue_empty;
  assign otherUnitDataQueueVec_3_deq_ready = dataDeqFire[3];
  wire [1:0]          otherUnit_vrfReadDataPorts_ready_lo = {vrfReadDataPorts_1_ready_0, vrfReadDataPorts_0_ready_0};
  wire [1:0]          otherUnit_vrfReadDataPorts_ready_hi = {vrfReadDataPorts_3_ready_0, vrfReadDataPorts_2_ready_0};
  wire                otherUnit_vrfReadDataPorts_ready = (|(otherTryReadVrf & {otherUnit_vrfReadDataPorts_ready_hi, otherUnit_vrfReadDataPorts_ready_lo})) & otherUnitTargetQueue_enq_ready;
  assign otherUnitTargetQueue_enq_valid = otherUnit_vrfReadDataPorts_ready & _otherUnit_vrfReadDataPorts_valid;
  wire [3:0]          otherUnitTargetQueue_deq_bits;
  wire [1:0]          otherUnit_vrfReadResults_valid_lo = {otherUnitDataQueueVec_1_deq_valid, otherUnitDataQueueVec_0_deq_valid};
  wire [1:0]          otherUnit_vrfReadResults_valid_hi = {otherUnitDataQueueVec_3_deq_valid, otherUnitDataQueueVec_2_deq_valid};
  assign otherUnitTargetQueue_deq_ready = otherUnitTargetQueue_deq_valid & (|(otherUnitTargetQueue_deq_bits & {otherUnit_vrfReadResults_valid_hi, otherUnit_vrfReadResults_valid_lo}));
  assign dataDeqFire = otherUnitTargetQueue_deq_ready ? otherUnitTargetQueue_deq_bits : 4'h0;
  wire [3:0]          otherTryToWrite = _otherUnit_vrfWritePort_valid ? _otherUnit_status_targetLane : 4'h0;
  wire [1:0]          otherUnit_vrfWritePort_ready_lo = {writeQueueVec_1_enq_ready, writeQueueVec_0_enq_ready};
  wire [1:0]          otherUnit_vrfWritePort_ready_hi = {writeQueueVec_3_enq_ready, writeQueueVec_2_enq_ready};
  assign writeQueueVec_0_enq_valid = otherTryToWrite[0] | _loadUnit_vrfWritePort_0_valid;
  assign writeQueueVec_0_enq_bits_data_vd = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_0_bits_vd;
  assign writeQueueVec_0_enq_bits_data_offset = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_0_bits_offset;
  assign writeQueueVec_0_enq_bits_data_mask = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_0_bits_mask;
  assign writeQueueVec_0_enq_bits_data_data = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_0_bits_data;
  assign writeQueueVec_0_enq_bits_data_last = otherTryToWrite[0] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_0_enq_bits_data_instructionIndex = otherTryToWrite[0] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_0_bits_instructionIndex;
  assign writeQueueVec_1_enq_valid = otherTryToWrite[1] | _loadUnit_vrfWritePort_1_valid;
  assign writeQueueVec_1_enq_bits_data_vd = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_1_bits_vd;
  assign writeQueueVec_1_enq_bits_data_offset = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_1_bits_offset;
  assign writeQueueVec_1_enq_bits_data_mask = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_1_bits_mask;
  assign writeQueueVec_1_enq_bits_data_data = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_1_bits_data;
  assign writeQueueVec_1_enq_bits_data_last = otherTryToWrite[1] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_1_enq_bits_data_instructionIndex = otherTryToWrite[1] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_1_bits_instructionIndex;
  assign writeQueueVec_2_enq_valid = otherTryToWrite[2] | _loadUnit_vrfWritePort_2_valid;
  assign writeQueueVec_2_enq_bits_data_vd = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_2_bits_vd;
  assign writeQueueVec_2_enq_bits_data_offset = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_2_bits_offset;
  assign writeQueueVec_2_enq_bits_data_mask = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_2_bits_mask;
  assign writeQueueVec_2_enq_bits_data_data = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_2_bits_data;
  assign writeQueueVec_2_enq_bits_data_last = otherTryToWrite[2] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_2_enq_bits_data_instructionIndex = otherTryToWrite[2] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_2_bits_instructionIndex;
  assign writeQueueVec_3_enq_valid = otherTryToWrite[3] | _loadUnit_vrfWritePort_3_valid;
  assign writeQueueVec_3_enq_bits_data_vd = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_vd : _loadUnit_vrfWritePort_3_bits_vd;
  assign writeQueueVec_3_enq_bits_data_offset = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_offset : _loadUnit_vrfWritePort_3_bits_offset;
  assign writeQueueVec_3_enq_bits_data_mask = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_mask : _loadUnit_vrfWritePort_3_bits_mask;
  assign writeQueueVec_3_enq_bits_data_data = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_data : _loadUnit_vrfWritePort_3_bits_data;
  assign writeQueueVec_3_enq_bits_data_last = otherTryToWrite[3] & _otherUnit_vrfWritePort_bits_last;
  assign writeQueueVec_3_enq_bits_data_instructionIndex = otherTryToWrite[3] ? _otherUnit_vrfWritePort_bits_instructionIndex : _loadUnit_vrfWritePort_3_bits_instructionIndex;
  wire [7:0]          _GEN_514 = {5'h0, _loadUnit_status_instructionIndex};
  wire [7:0]          _GEN_515 = {5'h0, _otherUnit_status_instructionIndex};
  wire [7:0]          dataInMSHR = (_loadUnit_status_idle ? 8'h0 : 8'h1 << _GEN_514) | (_otherUnit_status_idle | _otherUnit_status_isStore ? 8'h0 : 8'h1 << _GEN_515);
  reg  [6:0]          queueCount_0;
  reg  [6:0]          queueCount_1;
  reg  [6:0]          queueCount_2;
  reg  [6:0]          queueCount_3;
  reg  [6:0]          queueCount_4;
  reg  [6:0]          queueCount_5;
  reg  [6:0]          queueCount_6;
  reg  [6:0]          queueCount_7;
  wire [7:0]          enqOH = 8'h1 << writeQueueVec_0_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq = _probeWire_slots_0_writeValid_T ? enqOH : 8'h0;
  wire                writeIndexQueue_deq_valid;
  assign writeIndexQueue_deq_valid = ~_writeIndexQueue_fifo_empty;
  wire                writeIndexQueue_enq_ready = ~_writeIndexQueue_fifo_full;
  wire                writeIndexQueue_enq_valid;
  assign writeIndexQueue_enq_valid = writeQueueVec_0_deq_ready & writeQueueVec_0_deq_valid;
  wire [2:0]          writeIndexQueue_deq_bits;
  wire [7:0]          queueDeq = writeIndexQueue_deq_ready & writeIndexQueue_deq_valid ? 8'h1 << writeIndexQueue_deq_bits : 8'h0;
  wire [6:0]          counterUpdate = queueEnq[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_1 = queueEnq[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_2 = queueEnq[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_3 = queueEnq[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_4 = queueEnq[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_5 = queueEnq[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_6 = queueEnq[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_7 = queueEnq[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_0_lo_lo = {|queueCount_1, |queueCount_0};
  wire [1:0]          dataInWriteQueue_0_lo_hi = {|queueCount_3, |queueCount_2};
  wire [3:0]          dataInWriteQueue_0_lo = {dataInWriteQueue_0_lo_hi, dataInWriteQueue_0_lo_lo};
  wire [1:0]          dataInWriteQueue_0_hi_lo = {|queueCount_5, |queueCount_4};
  wire [1:0]          dataInWriteQueue_0_hi_hi = {|queueCount_7, |queueCount_6};
  wire [3:0]          dataInWriteQueue_0_hi = {dataInWriteQueue_0_hi_hi, dataInWriteQueue_0_hi_lo};
  reg  [6:0]          queueCount_0_1;
  reg  [6:0]          queueCount_1_1;
  reg  [6:0]          queueCount_2_1;
  reg  [6:0]          queueCount_3_1;
  reg  [6:0]          queueCount_4_1;
  reg  [6:0]          queueCount_5_1;
  reg  [6:0]          queueCount_6_1;
  reg  [6:0]          queueCount_7_1;
  wire [7:0]          enqOH_1 = 8'h1 << writeQueueVec_1_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq_1 = _probeWire_slots_1_writeValid_T ? enqOH_1 : 8'h0;
  wire                writeIndexQueue_1_deq_valid;
  assign writeIndexQueue_1_deq_valid = ~_writeIndexQueue_fifo_1_empty;
  wire                writeIndexQueue_1_enq_ready = ~_writeIndexQueue_fifo_1_full;
  wire                writeIndexQueue_1_enq_valid;
  assign writeIndexQueue_1_enq_valid = writeQueueVec_1_deq_ready & writeQueueVec_1_deq_valid;
  wire [2:0]          writeIndexQueue_1_deq_bits;
  wire [7:0]          queueDeq_1 = writeIndexQueue_1_deq_ready & writeIndexQueue_1_deq_valid ? 8'h1 << writeIndexQueue_1_deq_bits : 8'h0;
  wire [6:0]          counterUpdate_8 = queueEnq_1[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_9 = queueEnq_1[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_10 = queueEnq_1[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_11 = queueEnq_1[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_12 = queueEnq_1[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_13 = queueEnq_1[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_14 = queueEnq_1[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_15 = queueEnq_1[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_1_lo_lo = {|queueCount_1_1, |queueCount_0_1};
  wire [1:0]          dataInWriteQueue_1_lo_hi = {|queueCount_3_1, |queueCount_2_1};
  wire [3:0]          dataInWriteQueue_1_lo = {dataInWriteQueue_1_lo_hi, dataInWriteQueue_1_lo_lo};
  wire [1:0]          dataInWriteQueue_1_hi_lo = {|queueCount_5_1, |queueCount_4_1};
  wire [1:0]          dataInWriteQueue_1_hi_hi = {|queueCount_7_1, |queueCount_6_1};
  wire [3:0]          dataInWriteQueue_1_hi = {dataInWriteQueue_1_hi_hi, dataInWriteQueue_1_hi_lo};
  reg  [6:0]          queueCount_0_2;
  reg  [6:0]          queueCount_1_2;
  reg  [6:0]          queueCount_2_2;
  reg  [6:0]          queueCount_3_2;
  reg  [6:0]          queueCount_4_2;
  reg  [6:0]          queueCount_5_2;
  reg  [6:0]          queueCount_6_2;
  reg  [6:0]          queueCount_7_2;
  wire [7:0]          enqOH_2 = 8'h1 << writeQueueVec_2_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq_2 = _probeWire_slots_2_writeValid_T ? enqOH_2 : 8'h0;
  wire                writeIndexQueue_2_deq_valid;
  assign writeIndexQueue_2_deq_valid = ~_writeIndexQueue_fifo_2_empty;
  wire                writeIndexQueue_2_enq_ready = ~_writeIndexQueue_fifo_2_full;
  wire                writeIndexQueue_2_enq_valid;
  assign writeIndexQueue_2_enq_valid = writeQueueVec_2_deq_ready & writeQueueVec_2_deq_valid;
  wire [2:0]          writeIndexQueue_2_deq_bits;
  wire [7:0]          queueDeq_2 = writeIndexQueue_2_deq_ready & writeIndexQueue_2_deq_valid ? 8'h1 << writeIndexQueue_2_deq_bits : 8'h0;
  wire [6:0]          counterUpdate_16 = queueEnq_2[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_17 = queueEnq_2[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_18 = queueEnq_2[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_19 = queueEnq_2[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_20 = queueEnq_2[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_21 = queueEnq_2[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_22 = queueEnq_2[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_23 = queueEnq_2[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_2_lo_lo = {|queueCount_1_2, |queueCount_0_2};
  wire [1:0]          dataInWriteQueue_2_lo_hi = {|queueCount_3_2, |queueCount_2_2};
  wire [3:0]          dataInWriteQueue_2_lo = {dataInWriteQueue_2_lo_hi, dataInWriteQueue_2_lo_lo};
  wire [1:0]          dataInWriteQueue_2_hi_lo = {|queueCount_5_2, |queueCount_4_2};
  wire [1:0]          dataInWriteQueue_2_hi_hi = {|queueCount_7_2, |queueCount_6_2};
  wire [3:0]          dataInWriteQueue_2_hi = {dataInWriteQueue_2_hi_hi, dataInWriteQueue_2_hi_lo};
  reg  [6:0]          queueCount_0_3;
  reg  [6:0]          queueCount_1_3;
  reg  [6:0]          queueCount_2_3;
  reg  [6:0]          queueCount_3_3;
  reg  [6:0]          queueCount_4_3;
  reg  [6:0]          queueCount_5_3;
  reg  [6:0]          queueCount_6_3;
  reg  [6:0]          queueCount_7_3;
  wire [7:0]          enqOH_3 = 8'h1 << writeQueueVec_3_enq_bits_data_instructionIndex;
  wire [7:0]          queueEnq_3 = _probeWire_slots_3_writeValid_T ? enqOH_3 : 8'h0;
  wire                writeIndexQueue_3_deq_valid;
  assign writeIndexQueue_3_deq_valid = ~_writeIndexQueue_fifo_3_empty;
  wire                writeIndexQueue_3_enq_ready = ~_writeIndexQueue_fifo_3_full;
  wire                writeIndexQueue_3_enq_valid;
  assign writeIndexQueue_3_enq_valid = writeQueueVec_3_deq_ready & writeQueueVec_3_deq_valid;
  wire [2:0]          writeIndexQueue_3_deq_bits;
  wire [7:0]          queueDeq_3 = writeIndexQueue_3_deq_ready & writeIndexQueue_3_deq_valid ? 8'h1 << writeIndexQueue_3_deq_bits : 8'h0;
  wire [6:0]          counterUpdate_24 = queueEnq_3[0] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_25 = queueEnq_3[1] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_26 = queueEnq_3[2] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_27 = queueEnq_3[3] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_28 = queueEnq_3[4] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_29 = queueEnq_3[5] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_30 = queueEnq_3[6] ? 7'h1 : 7'h7F;
  wire [6:0]          counterUpdate_31 = queueEnq_3[7] ? 7'h1 : 7'h7F;
  wire [1:0]          dataInWriteQueue_3_lo_lo = {|queueCount_1_3, |queueCount_0_3};
  wire [1:0]          dataInWriteQueue_3_lo_hi = {|queueCount_3_3, |queueCount_2_3};
  wire [3:0]          dataInWriteQueue_3_lo = {dataInWriteQueue_3_lo_hi, dataInWriteQueue_3_lo_lo};
  wire [1:0]          dataInWriteQueue_3_hi_lo = {|queueCount_5_3, |queueCount_4_3};
  wire [1:0]          dataInWriteQueue_3_hi_hi = {|queueCount_7_3, |queueCount_6_3};
  wire [3:0]          dataInWriteQueue_3_hi = {dataInWriteQueue_3_hi_hi, dataInWriteQueue_3_hi_lo};
  wire                sourceQueue_deq_valid;
  assign sourceQueue_deq_valid = ~_sourceQueue_fifo_empty;
  wire                sourceQueue_enq_ready = ~_sourceQueue_fifo_full;
  wire                sourceQueue_enq_valid;
  wire                sourceQueue_deq_ready;
  wire                axi4Port_ar_valid_0 = _loadUnit_memRequest_valid & sourceQueue_enq_ready;
  wire                axi4Port_r_ready_0;
  assign sourceQueue_enq_valid = _loadUnit_memRequest_valid & axi4Port_ar_ready_0;
  assign sourceQueue_deq_ready = axi4Port_r_ready_0 & axi4Port_r_valid_0;
  assign dataQueue_deq_valid = ~_dataQueue_fifo_empty;
  wire                axi4Port_w_valid_0 = dataQueue_deq_valid;
  wire [127:0]        dataQueue_dataOut_data;
  wire [127:0]        axi4Port_w_bits_data_0 = dataQueue_deq_bits_data;
  wire [15:0]         dataQueue_dataOut_mask;
  wire [15:0]         axi4Port_w_bits_strb_0 = dataQueue_deq_bits_mask;
  wire [11:0]         dataQueue_dataOut_index;
  wire [31:0]         dataQueue_dataOut_address;
  wire [11:0]         dataQueue_enq_bits_index;
  wire [31:0]         dataQueue_enq_bits_address;
  wire [43:0]         dataQueue_dataIn_lo = {dataQueue_enq_bits_index, dataQueue_enq_bits_address};
  wire [127:0]        dataQueue_enq_bits_data;
  wire [15:0]         dataQueue_enq_bits_mask;
  wire [143:0]        dataQueue_dataIn_hi = {dataQueue_enq_bits_data, dataQueue_enq_bits_mask};
  wire [187:0]        dataQueue_dataIn = {dataQueue_dataIn_hi, dataQueue_dataIn_lo};
  assign dataQueue_dataOut_address = _dataQueue_fifo_data_out[31:0];
  assign dataQueue_dataOut_index = _dataQueue_fifo_data_out[43:32];
  assign dataQueue_dataOut_mask = _dataQueue_fifo_data_out[59:44];
  assign dataQueue_dataOut_data = _dataQueue_fifo_data_out[187:60];
  assign dataQueue_deq_bits_data = dataQueue_dataOut_data;
  assign dataQueue_deq_bits_mask = dataQueue_dataOut_mask;
  wire [11:0]         dataQueue_deq_bits_index = dataQueue_dataOut_index;
  wire [31:0]         dataQueue_deq_bits_address = dataQueue_dataOut_address;
  wire                dataQueue_enq_ready = ~_dataQueue_fifo_full;
  wire                dataQueue_enq_valid;
  wire                axi4Port_aw_valid_0 = _storeUnit_memRequest_valid & dataQueue_enq_ready;
  wire [1:0]          axi4Port_aw_bits_id_0 = _storeUnit_memRequest_bits_index[1:0];
  assign dataQueue_enq_valid = _storeUnit_memRequest_valid & axi4Port_aw_ready_0;
  wire                simpleSourceQueue_deq_valid;
  assign simpleSourceQueue_deq_valid = ~_simpleSourceQueue_fifo_empty;
  wire                simpleSourceQueue_enq_ready = ~_simpleSourceQueue_fifo_full;
  wire                simpleSourceQueue_enq_valid;
  wire                simpleSourceQueue_deq_ready;
  wire                simpleAccessPorts_ar_valid_0 = _otherUnit_memReadRequest_valid & simpleSourceQueue_enq_ready;
  wire                simpleAccessPorts_r_ready_0;
  assign simpleSourceQueue_enq_valid = _otherUnit_memReadRequest_valid & simpleAccessPorts_ar_ready_0;
  assign simpleSourceQueue_deq_ready = simpleAccessPorts_r_ready_0 & simpleAccessPorts_r_valid_0;
  assign simpleDataQueue_deq_valid = ~_simpleDataQueue_fifo_empty;
  wire                simpleAccessPorts_w_valid_0 = simpleDataQueue_deq_valid;
  wire [31:0]         simpleDataQueue_dataOut_data;
  wire [31:0]         simpleAccessPorts_w_bits_data_0 = simpleDataQueue_deq_bits_data;
  wire [3:0]          simpleDataQueue_dataOut_mask;
  wire [3:0]          simpleAccessPorts_w_bits_strb_0 = simpleDataQueue_deq_bits_mask;
  wire [7:0]          simpleDataQueue_dataOut_source;
  wire [31:0]         simpleDataQueue_dataOut_address;
  wire [1:0]          simpleDataQueue_dataOut_size;
  wire [31:0]         simpleDataQueue_enq_bits_address;
  wire [1:0]          simpleDataQueue_enq_bits_size;
  wire [33:0]         simpleDataQueue_dataIn_lo = {simpleDataQueue_enq_bits_address, simpleDataQueue_enq_bits_size};
  wire [31:0]         simpleDataQueue_enq_bits_data;
  wire [3:0]          simpleDataQueue_enq_bits_mask;
  wire [35:0]         simpleDataQueue_dataIn_hi_hi = {simpleDataQueue_enq_bits_data, simpleDataQueue_enq_bits_mask};
  wire [7:0]          simpleDataQueue_enq_bits_source;
  wire [43:0]         simpleDataQueue_dataIn_hi = {simpleDataQueue_dataIn_hi_hi, simpleDataQueue_enq_bits_source};
  wire [77:0]         simpleDataQueue_dataIn = {simpleDataQueue_dataIn_hi, simpleDataQueue_dataIn_lo};
  assign simpleDataQueue_dataOut_size = _simpleDataQueue_fifo_data_out[1:0];
  assign simpleDataQueue_dataOut_address = _simpleDataQueue_fifo_data_out[33:2];
  assign simpleDataQueue_dataOut_source = _simpleDataQueue_fifo_data_out[41:34];
  assign simpleDataQueue_dataOut_mask = _simpleDataQueue_fifo_data_out[45:42];
  assign simpleDataQueue_dataOut_data = _simpleDataQueue_fifo_data_out[77:46];
  assign simpleDataQueue_deq_bits_data = simpleDataQueue_dataOut_data;
  assign simpleDataQueue_deq_bits_mask = simpleDataQueue_dataOut_mask;
  wire [7:0]          simpleDataQueue_deq_bits_source = simpleDataQueue_dataOut_source;
  wire [31:0]         simpleDataQueue_deq_bits_address = simpleDataQueue_dataOut_address;
  wire [1:0]          simpleDataQueue_deq_bits_size = simpleDataQueue_dataOut_size;
  wire                simpleDataQueue_enq_ready = ~_simpleDataQueue_fifo_full;
  wire                simpleDataQueue_enq_valid;
  wire                simpleAccessPorts_aw_valid_0 = _otherUnit_memWriteRequest_valid & dataQueue_enq_ready;
  wire [2:0]          simpleAccessPorts_aw_bits_size_0 = {1'h0, _otherUnit_memWriteRequest_bits_size};
  wire [1:0]          simpleAccessPorts_aw_bits_id_0 = _otherUnit_memWriteRequest_bits_source[1:0];
  assign simpleDataQueue_enq_valid = _otherUnit_memWriteRequest_valid & simpleAccessPorts_aw_ready_0;
  wire [1:0]          tokenIO_offsetGroupRelease_lo = {_otherUnit_offsetRelease_1, _otherUnit_offsetRelease_0};
  wire [1:0]          tokenIO_offsetGroupRelease_hi = {_otherUnit_offsetRelease_3, _otherUnit_offsetRelease_2};
  wire                unitOrder =
    _loadUnit_status_instructionIndex == _storeUnit_status_instructionIndex | _loadUnit_status_instructionIndex[1:0] < _storeUnit_status_instructionIndex[1:0] ^ _loadUnit_status_instructionIndex[2] ^ _storeUnit_status_instructionIndex[2];
  wire                loadAddressConflict = _loadUnit_status_startAddress >= _storeUnit_status_startAddress & _loadUnit_status_startAddress <= _storeUnit_status_endAddress;
  wire                storeAddressConflict = _storeUnit_status_startAddress >= _loadUnit_status_startAddress & _storeUnit_status_startAddress <= _loadUnit_status_endAddress;
  wire                stallLoad = ~unitOrder & loadAddressConflict & ~_storeUnit_status_idle;
  wire                stallStore = unitOrder & storeAddressConflict & ~_loadUnit_status_idle;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      v0_32 <= 32'h0;
      v0_33 <= 32'h0;
      v0_34 <= 32'h0;
      v0_35 <= 32'h0;
      v0_36 <= 32'h0;
      v0_37 <= 32'h0;
      v0_38 <= 32'h0;
      v0_39 <= 32'h0;
      v0_40 <= 32'h0;
      v0_41 <= 32'h0;
      v0_42 <= 32'h0;
      v0_43 <= 32'h0;
      v0_44 <= 32'h0;
      v0_45 <= 32'h0;
      v0_46 <= 32'h0;
      v0_47 <= 32'h0;
      v0_48 <= 32'h0;
      v0_49 <= 32'h0;
      v0_50 <= 32'h0;
      v0_51 <= 32'h0;
      v0_52 <= 32'h0;
      v0_53 <= 32'h0;
      v0_54 <= 32'h0;
      v0_55 <= 32'h0;
      v0_56 <= 32'h0;
      v0_57 <= 32'h0;
      v0_58 <= 32'h0;
      v0_59 <= 32'h0;
      v0_60 <= 32'h0;
      v0_61 <= 32'h0;
      v0_62 <= 32'h0;
      v0_63 <= 32'h0;
      v0_64 <= 32'h0;
      v0_65 <= 32'h0;
      v0_66 <= 32'h0;
      v0_67 <= 32'h0;
      v0_68 <= 32'h0;
      v0_69 <= 32'h0;
      v0_70 <= 32'h0;
      v0_71 <= 32'h0;
      v0_72 <= 32'h0;
      v0_73 <= 32'h0;
      v0_74 <= 32'h0;
      v0_75 <= 32'h0;
      v0_76 <= 32'h0;
      v0_77 <= 32'h0;
      v0_78 <= 32'h0;
      v0_79 <= 32'h0;
      v0_80 <= 32'h0;
      v0_81 <= 32'h0;
      v0_82 <= 32'h0;
      v0_83 <= 32'h0;
      v0_84 <= 32'h0;
      v0_85 <= 32'h0;
      v0_86 <= 32'h0;
      v0_87 <= 32'h0;
      v0_88 <= 32'h0;
      v0_89 <= 32'h0;
      v0_90 <= 32'h0;
      v0_91 <= 32'h0;
      v0_92 <= 32'h0;
      v0_93 <= 32'h0;
      v0_94 <= 32'h0;
      v0_95 <= 32'h0;
      v0_96 <= 32'h0;
      v0_97 <= 32'h0;
      v0_98 <= 32'h0;
      v0_99 <= 32'h0;
      v0_100 <= 32'h0;
      v0_101 <= 32'h0;
      v0_102 <= 32'h0;
      v0_103 <= 32'h0;
      v0_104 <= 32'h0;
      v0_105 <= 32'h0;
      v0_106 <= 32'h0;
      v0_107 <= 32'h0;
      v0_108 <= 32'h0;
      v0_109 <= 32'h0;
      v0_110 <= 32'h0;
      v0_111 <= 32'h0;
      v0_112 <= 32'h0;
      v0_113 <= 32'h0;
      v0_114 <= 32'h0;
      v0_115 <= 32'h0;
      v0_116 <= 32'h0;
      v0_117 <= 32'h0;
      v0_118 <= 32'h0;
      v0_119 <= 32'h0;
      v0_120 <= 32'h0;
      v0_121 <= 32'h0;
      v0_122 <= 32'h0;
      v0_123 <= 32'h0;
      v0_124 <= 32'h0;
      v0_125 <= 32'h0;
      v0_126 <= 32'h0;
      v0_127 <= 32'h0;
      v0_128 <= 32'h0;
      v0_129 <= 32'h0;
      v0_130 <= 32'h0;
      v0_131 <= 32'h0;
      v0_132 <= 32'h0;
      v0_133 <= 32'h0;
      v0_134 <= 32'h0;
      v0_135 <= 32'h0;
      v0_136 <= 32'h0;
      v0_137 <= 32'h0;
      v0_138 <= 32'h0;
      v0_139 <= 32'h0;
      v0_140 <= 32'h0;
      v0_141 <= 32'h0;
      v0_142 <= 32'h0;
      v0_143 <= 32'h0;
      v0_144 <= 32'h0;
      v0_145 <= 32'h0;
      v0_146 <= 32'h0;
      v0_147 <= 32'h0;
      v0_148 <= 32'h0;
      v0_149 <= 32'h0;
      v0_150 <= 32'h0;
      v0_151 <= 32'h0;
      v0_152 <= 32'h0;
      v0_153 <= 32'h0;
      v0_154 <= 32'h0;
      v0_155 <= 32'h0;
      v0_156 <= 32'h0;
      v0_157 <= 32'h0;
      v0_158 <= 32'h0;
      v0_159 <= 32'h0;
      v0_160 <= 32'h0;
      v0_161 <= 32'h0;
      v0_162 <= 32'h0;
      v0_163 <= 32'h0;
      v0_164 <= 32'h0;
      v0_165 <= 32'h0;
      v0_166 <= 32'h0;
      v0_167 <= 32'h0;
      v0_168 <= 32'h0;
      v0_169 <= 32'h0;
      v0_170 <= 32'h0;
      v0_171 <= 32'h0;
      v0_172 <= 32'h0;
      v0_173 <= 32'h0;
      v0_174 <= 32'h0;
      v0_175 <= 32'h0;
      v0_176 <= 32'h0;
      v0_177 <= 32'h0;
      v0_178 <= 32'h0;
      v0_179 <= 32'h0;
      v0_180 <= 32'h0;
      v0_181 <= 32'h0;
      v0_182 <= 32'h0;
      v0_183 <= 32'h0;
      v0_184 <= 32'h0;
      v0_185 <= 32'h0;
      v0_186 <= 32'h0;
      v0_187 <= 32'h0;
      v0_188 <= 32'h0;
      v0_189 <= 32'h0;
      v0_190 <= 32'h0;
      v0_191 <= 32'h0;
      v0_192 <= 32'h0;
      v0_193 <= 32'h0;
      v0_194 <= 32'h0;
      v0_195 <= 32'h0;
      v0_196 <= 32'h0;
      v0_197 <= 32'h0;
      v0_198 <= 32'h0;
      v0_199 <= 32'h0;
      v0_200 <= 32'h0;
      v0_201 <= 32'h0;
      v0_202 <= 32'h0;
      v0_203 <= 32'h0;
      v0_204 <= 32'h0;
      v0_205 <= 32'h0;
      v0_206 <= 32'h0;
      v0_207 <= 32'h0;
      v0_208 <= 32'h0;
      v0_209 <= 32'h0;
      v0_210 <= 32'h0;
      v0_211 <= 32'h0;
      v0_212 <= 32'h0;
      v0_213 <= 32'h0;
      v0_214 <= 32'h0;
      v0_215 <= 32'h0;
      v0_216 <= 32'h0;
      v0_217 <= 32'h0;
      v0_218 <= 32'h0;
      v0_219 <= 32'h0;
      v0_220 <= 32'h0;
      v0_221 <= 32'h0;
      v0_222 <= 32'h0;
      v0_223 <= 32'h0;
      v0_224 <= 32'h0;
      v0_225 <= 32'h0;
      v0_226 <= 32'h0;
      v0_227 <= 32'h0;
      v0_228 <= 32'h0;
      v0_229 <= 32'h0;
      v0_230 <= 32'h0;
      v0_231 <= 32'h0;
      v0_232 <= 32'h0;
      v0_233 <= 32'h0;
      v0_234 <= 32'h0;
      v0_235 <= 32'h0;
      v0_236 <= 32'h0;
      v0_237 <= 32'h0;
      v0_238 <= 32'h0;
      v0_239 <= 32'h0;
      v0_240 <= 32'h0;
      v0_241 <= 32'h0;
      v0_242 <= 32'h0;
      v0_243 <= 32'h0;
      v0_244 <= 32'h0;
      v0_245 <= 32'h0;
      v0_246 <= 32'h0;
      v0_247 <= 32'h0;
      v0_248 <= 32'h0;
      v0_249 <= 32'h0;
      v0_250 <= 32'h0;
      v0_251 <= 32'h0;
      v0_252 <= 32'h0;
      v0_253 <= 32'h0;
      v0_254 <= 32'h0;
      v0_255 <= 32'h0;
      v0_256 <= 32'h0;
      v0_257 <= 32'h0;
      v0_258 <= 32'h0;
      v0_259 <= 32'h0;
      v0_260 <= 32'h0;
      v0_261 <= 32'h0;
      v0_262 <= 32'h0;
      v0_263 <= 32'h0;
      v0_264 <= 32'h0;
      v0_265 <= 32'h0;
      v0_266 <= 32'h0;
      v0_267 <= 32'h0;
      v0_268 <= 32'h0;
      v0_269 <= 32'h0;
      v0_270 <= 32'h0;
      v0_271 <= 32'h0;
      v0_272 <= 32'h0;
      v0_273 <= 32'h0;
      v0_274 <= 32'h0;
      v0_275 <= 32'h0;
      v0_276 <= 32'h0;
      v0_277 <= 32'h0;
      v0_278 <= 32'h0;
      v0_279 <= 32'h0;
      v0_280 <= 32'h0;
      v0_281 <= 32'h0;
      v0_282 <= 32'h0;
      v0_283 <= 32'h0;
      v0_284 <= 32'h0;
      v0_285 <= 32'h0;
      v0_286 <= 32'h0;
      v0_287 <= 32'h0;
      v0_288 <= 32'h0;
      v0_289 <= 32'h0;
      v0_290 <= 32'h0;
      v0_291 <= 32'h0;
      v0_292 <= 32'h0;
      v0_293 <= 32'h0;
      v0_294 <= 32'h0;
      v0_295 <= 32'h0;
      v0_296 <= 32'h0;
      v0_297 <= 32'h0;
      v0_298 <= 32'h0;
      v0_299 <= 32'h0;
      v0_300 <= 32'h0;
      v0_301 <= 32'h0;
      v0_302 <= 32'h0;
      v0_303 <= 32'h0;
      v0_304 <= 32'h0;
      v0_305 <= 32'h0;
      v0_306 <= 32'h0;
      v0_307 <= 32'h0;
      v0_308 <= 32'h0;
      v0_309 <= 32'h0;
      v0_310 <= 32'h0;
      v0_311 <= 32'h0;
      v0_312 <= 32'h0;
      v0_313 <= 32'h0;
      v0_314 <= 32'h0;
      v0_315 <= 32'h0;
      v0_316 <= 32'h0;
      v0_317 <= 32'h0;
      v0_318 <= 32'h0;
      v0_319 <= 32'h0;
      v0_320 <= 32'h0;
      v0_321 <= 32'h0;
      v0_322 <= 32'h0;
      v0_323 <= 32'h0;
      v0_324 <= 32'h0;
      v0_325 <= 32'h0;
      v0_326 <= 32'h0;
      v0_327 <= 32'h0;
      v0_328 <= 32'h0;
      v0_329 <= 32'h0;
      v0_330 <= 32'h0;
      v0_331 <= 32'h0;
      v0_332 <= 32'h0;
      v0_333 <= 32'h0;
      v0_334 <= 32'h0;
      v0_335 <= 32'h0;
      v0_336 <= 32'h0;
      v0_337 <= 32'h0;
      v0_338 <= 32'h0;
      v0_339 <= 32'h0;
      v0_340 <= 32'h0;
      v0_341 <= 32'h0;
      v0_342 <= 32'h0;
      v0_343 <= 32'h0;
      v0_344 <= 32'h0;
      v0_345 <= 32'h0;
      v0_346 <= 32'h0;
      v0_347 <= 32'h0;
      v0_348 <= 32'h0;
      v0_349 <= 32'h0;
      v0_350 <= 32'h0;
      v0_351 <= 32'h0;
      v0_352 <= 32'h0;
      v0_353 <= 32'h0;
      v0_354 <= 32'h0;
      v0_355 <= 32'h0;
      v0_356 <= 32'h0;
      v0_357 <= 32'h0;
      v0_358 <= 32'h0;
      v0_359 <= 32'h0;
      v0_360 <= 32'h0;
      v0_361 <= 32'h0;
      v0_362 <= 32'h0;
      v0_363 <= 32'h0;
      v0_364 <= 32'h0;
      v0_365 <= 32'h0;
      v0_366 <= 32'h0;
      v0_367 <= 32'h0;
      v0_368 <= 32'h0;
      v0_369 <= 32'h0;
      v0_370 <= 32'h0;
      v0_371 <= 32'h0;
      v0_372 <= 32'h0;
      v0_373 <= 32'h0;
      v0_374 <= 32'h0;
      v0_375 <= 32'h0;
      v0_376 <= 32'h0;
      v0_377 <= 32'h0;
      v0_378 <= 32'h0;
      v0_379 <= 32'h0;
      v0_380 <= 32'h0;
      v0_381 <= 32'h0;
      v0_382 <= 32'h0;
      v0_383 <= 32'h0;
      v0_384 <= 32'h0;
      v0_385 <= 32'h0;
      v0_386 <= 32'h0;
      v0_387 <= 32'h0;
      v0_388 <= 32'h0;
      v0_389 <= 32'h0;
      v0_390 <= 32'h0;
      v0_391 <= 32'h0;
      v0_392 <= 32'h0;
      v0_393 <= 32'h0;
      v0_394 <= 32'h0;
      v0_395 <= 32'h0;
      v0_396 <= 32'h0;
      v0_397 <= 32'h0;
      v0_398 <= 32'h0;
      v0_399 <= 32'h0;
      v0_400 <= 32'h0;
      v0_401 <= 32'h0;
      v0_402 <= 32'h0;
      v0_403 <= 32'h0;
      v0_404 <= 32'h0;
      v0_405 <= 32'h0;
      v0_406 <= 32'h0;
      v0_407 <= 32'h0;
      v0_408 <= 32'h0;
      v0_409 <= 32'h0;
      v0_410 <= 32'h0;
      v0_411 <= 32'h0;
      v0_412 <= 32'h0;
      v0_413 <= 32'h0;
      v0_414 <= 32'h0;
      v0_415 <= 32'h0;
      v0_416 <= 32'h0;
      v0_417 <= 32'h0;
      v0_418 <= 32'h0;
      v0_419 <= 32'h0;
      v0_420 <= 32'h0;
      v0_421 <= 32'h0;
      v0_422 <= 32'h0;
      v0_423 <= 32'h0;
      v0_424 <= 32'h0;
      v0_425 <= 32'h0;
      v0_426 <= 32'h0;
      v0_427 <= 32'h0;
      v0_428 <= 32'h0;
      v0_429 <= 32'h0;
      v0_430 <= 32'h0;
      v0_431 <= 32'h0;
      v0_432 <= 32'h0;
      v0_433 <= 32'h0;
      v0_434 <= 32'h0;
      v0_435 <= 32'h0;
      v0_436 <= 32'h0;
      v0_437 <= 32'h0;
      v0_438 <= 32'h0;
      v0_439 <= 32'h0;
      v0_440 <= 32'h0;
      v0_441 <= 32'h0;
      v0_442 <= 32'h0;
      v0_443 <= 32'h0;
      v0_444 <= 32'h0;
      v0_445 <= 32'h0;
      v0_446 <= 32'h0;
      v0_447 <= 32'h0;
      v0_448 <= 32'h0;
      v0_449 <= 32'h0;
      v0_450 <= 32'h0;
      v0_451 <= 32'h0;
      v0_452 <= 32'h0;
      v0_453 <= 32'h0;
      v0_454 <= 32'h0;
      v0_455 <= 32'h0;
      v0_456 <= 32'h0;
      v0_457 <= 32'h0;
      v0_458 <= 32'h0;
      v0_459 <= 32'h0;
      v0_460 <= 32'h0;
      v0_461 <= 32'h0;
      v0_462 <= 32'h0;
      v0_463 <= 32'h0;
      v0_464 <= 32'h0;
      v0_465 <= 32'h0;
      v0_466 <= 32'h0;
      v0_467 <= 32'h0;
      v0_468 <= 32'h0;
      v0_469 <= 32'h0;
      v0_470 <= 32'h0;
      v0_471 <= 32'h0;
      v0_472 <= 32'h0;
      v0_473 <= 32'h0;
      v0_474 <= 32'h0;
      v0_475 <= 32'h0;
      v0_476 <= 32'h0;
      v0_477 <= 32'h0;
      v0_478 <= 32'h0;
      v0_479 <= 32'h0;
      v0_480 <= 32'h0;
      v0_481 <= 32'h0;
      v0_482 <= 32'h0;
      v0_483 <= 32'h0;
      v0_484 <= 32'h0;
      v0_485 <= 32'h0;
      v0_486 <= 32'h0;
      v0_487 <= 32'h0;
      v0_488 <= 32'h0;
      v0_489 <= 32'h0;
      v0_490 <= 32'h0;
      v0_491 <= 32'h0;
      v0_492 <= 32'h0;
      v0_493 <= 32'h0;
      v0_494 <= 32'h0;
      v0_495 <= 32'h0;
      v0_496 <= 32'h0;
      v0_497 <= 32'h0;
      v0_498 <= 32'h0;
      v0_499 <= 32'h0;
      v0_500 <= 32'h0;
      v0_501 <= 32'h0;
      v0_502 <= 32'h0;
      v0_503 <= 32'h0;
      v0_504 <= 32'h0;
      v0_505 <= 32'h0;
      v0_506 <= 32'h0;
      v0_507 <= 32'h0;
      v0_508 <= 32'h0;
      v0_509 <= 32'h0;
      v0_510 <= 32'h0;
      v0_511 <= 32'h0;
      v0_512 <= 32'h0;
      v0_513 <= 32'h0;
      v0_514 <= 32'h0;
      v0_515 <= 32'h0;
      v0_516 <= 32'h0;
      v0_517 <= 32'h0;
      v0_518 <= 32'h0;
      v0_519 <= 32'h0;
      v0_520 <= 32'h0;
      v0_521 <= 32'h0;
      v0_522 <= 32'h0;
      v0_523 <= 32'h0;
      v0_524 <= 32'h0;
      v0_525 <= 32'h0;
      v0_526 <= 32'h0;
      v0_527 <= 32'h0;
      v0_528 <= 32'h0;
      v0_529 <= 32'h0;
      v0_530 <= 32'h0;
      v0_531 <= 32'h0;
      v0_532 <= 32'h0;
      v0_533 <= 32'h0;
      v0_534 <= 32'h0;
      v0_535 <= 32'h0;
      v0_536 <= 32'h0;
      v0_537 <= 32'h0;
      v0_538 <= 32'h0;
      v0_539 <= 32'h0;
      v0_540 <= 32'h0;
      v0_541 <= 32'h0;
      v0_542 <= 32'h0;
      v0_543 <= 32'h0;
      v0_544 <= 32'h0;
      v0_545 <= 32'h0;
      v0_546 <= 32'h0;
      v0_547 <= 32'h0;
      v0_548 <= 32'h0;
      v0_549 <= 32'h0;
      v0_550 <= 32'h0;
      v0_551 <= 32'h0;
      v0_552 <= 32'h0;
      v0_553 <= 32'h0;
      v0_554 <= 32'h0;
      v0_555 <= 32'h0;
      v0_556 <= 32'h0;
      v0_557 <= 32'h0;
      v0_558 <= 32'h0;
      v0_559 <= 32'h0;
      v0_560 <= 32'h0;
      v0_561 <= 32'h0;
      v0_562 <= 32'h0;
      v0_563 <= 32'h0;
      v0_564 <= 32'h0;
      v0_565 <= 32'h0;
      v0_566 <= 32'h0;
      v0_567 <= 32'h0;
      v0_568 <= 32'h0;
      v0_569 <= 32'h0;
      v0_570 <= 32'h0;
      v0_571 <= 32'h0;
      v0_572 <= 32'h0;
      v0_573 <= 32'h0;
      v0_574 <= 32'h0;
      v0_575 <= 32'h0;
      v0_576 <= 32'h0;
      v0_577 <= 32'h0;
      v0_578 <= 32'h0;
      v0_579 <= 32'h0;
      v0_580 <= 32'h0;
      v0_581 <= 32'h0;
      v0_582 <= 32'h0;
      v0_583 <= 32'h0;
      v0_584 <= 32'h0;
      v0_585 <= 32'h0;
      v0_586 <= 32'h0;
      v0_587 <= 32'h0;
      v0_588 <= 32'h0;
      v0_589 <= 32'h0;
      v0_590 <= 32'h0;
      v0_591 <= 32'h0;
      v0_592 <= 32'h0;
      v0_593 <= 32'h0;
      v0_594 <= 32'h0;
      v0_595 <= 32'h0;
      v0_596 <= 32'h0;
      v0_597 <= 32'h0;
      v0_598 <= 32'h0;
      v0_599 <= 32'h0;
      v0_600 <= 32'h0;
      v0_601 <= 32'h0;
      v0_602 <= 32'h0;
      v0_603 <= 32'h0;
      v0_604 <= 32'h0;
      v0_605 <= 32'h0;
      v0_606 <= 32'h0;
      v0_607 <= 32'h0;
      v0_608 <= 32'h0;
      v0_609 <= 32'h0;
      v0_610 <= 32'h0;
      v0_611 <= 32'h0;
      v0_612 <= 32'h0;
      v0_613 <= 32'h0;
      v0_614 <= 32'h0;
      v0_615 <= 32'h0;
      v0_616 <= 32'h0;
      v0_617 <= 32'h0;
      v0_618 <= 32'h0;
      v0_619 <= 32'h0;
      v0_620 <= 32'h0;
      v0_621 <= 32'h0;
      v0_622 <= 32'h0;
      v0_623 <= 32'h0;
      v0_624 <= 32'h0;
      v0_625 <= 32'h0;
      v0_626 <= 32'h0;
      v0_627 <= 32'h0;
      v0_628 <= 32'h0;
      v0_629 <= 32'h0;
      v0_630 <= 32'h0;
      v0_631 <= 32'h0;
      v0_632 <= 32'h0;
      v0_633 <= 32'h0;
      v0_634 <= 32'h0;
      v0_635 <= 32'h0;
      v0_636 <= 32'h0;
      v0_637 <= 32'h0;
      v0_638 <= 32'h0;
      v0_639 <= 32'h0;
      v0_640 <= 32'h0;
      v0_641 <= 32'h0;
      v0_642 <= 32'h0;
      v0_643 <= 32'h0;
      v0_644 <= 32'h0;
      v0_645 <= 32'h0;
      v0_646 <= 32'h0;
      v0_647 <= 32'h0;
      v0_648 <= 32'h0;
      v0_649 <= 32'h0;
      v0_650 <= 32'h0;
      v0_651 <= 32'h0;
      v0_652 <= 32'h0;
      v0_653 <= 32'h0;
      v0_654 <= 32'h0;
      v0_655 <= 32'h0;
      v0_656 <= 32'h0;
      v0_657 <= 32'h0;
      v0_658 <= 32'h0;
      v0_659 <= 32'h0;
      v0_660 <= 32'h0;
      v0_661 <= 32'h0;
      v0_662 <= 32'h0;
      v0_663 <= 32'h0;
      v0_664 <= 32'h0;
      v0_665 <= 32'h0;
      v0_666 <= 32'h0;
      v0_667 <= 32'h0;
      v0_668 <= 32'h0;
      v0_669 <= 32'h0;
      v0_670 <= 32'h0;
      v0_671 <= 32'h0;
      v0_672 <= 32'h0;
      v0_673 <= 32'h0;
      v0_674 <= 32'h0;
      v0_675 <= 32'h0;
      v0_676 <= 32'h0;
      v0_677 <= 32'h0;
      v0_678 <= 32'h0;
      v0_679 <= 32'h0;
      v0_680 <= 32'h0;
      v0_681 <= 32'h0;
      v0_682 <= 32'h0;
      v0_683 <= 32'h0;
      v0_684 <= 32'h0;
      v0_685 <= 32'h0;
      v0_686 <= 32'h0;
      v0_687 <= 32'h0;
      v0_688 <= 32'h0;
      v0_689 <= 32'h0;
      v0_690 <= 32'h0;
      v0_691 <= 32'h0;
      v0_692 <= 32'h0;
      v0_693 <= 32'h0;
      v0_694 <= 32'h0;
      v0_695 <= 32'h0;
      v0_696 <= 32'h0;
      v0_697 <= 32'h0;
      v0_698 <= 32'h0;
      v0_699 <= 32'h0;
      v0_700 <= 32'h0;
      v0_701 <= 32'h0;
      v0_702 <= 32'h0;
      v0_703 <= 32'h0;
      v0_704 <= 32'h0;
      v0_705 <= 32'h0;
      v0_706 <= 32'h0;
      v0_707 <= 32'h0;
      v0_708 <= 32'h0;
      v0_709 <= 32'h0;
      v0_710 <= 32'h0;
      v0_711 <= 32'h0;
      v0_712 <= 32'h0;
      v0_713 <= 32'h0;
      v0_714 <= 32'h0;
      v0_715 <= 32'h0;
      v0_716 <= 32'h0;
      v0_717 <= 32'h0;
      v0_718 <= 32'h0;
      v0_719 <= 32'h0;
      v0_720 <= 32'h0;
      v0_721 <= 32'h0;
      v0_722 <= 32'h0;
      v0_723 <= 32'h0;
      v0_724 <= 32'h0;
      v0_725 <= 32'h0;
      v0_726 <= 32'h0;
      v0_727 <= 32'h0;
      v0_728 <= 32'h0;
      v0_729 <= 32'h0;
      v0_730 <= 32'h0;
      v0_731 <= 32'h0;
      v0_732 <= 32'h0;
      v0_733 <= 32'h0;
      v0_734 <= 32'h0;
      v0_735 <= 32'h0;
      v0_736 <= 32'h0;
      v0_737 <= 32'h0;
      v0_738 <= 32'h0;
      v0_739 <= 32'h0;
      v0_740 <= 32'h0;
      v0_741 <= 32'h0;
      v0_742 <= 32'h0;
      v0_743 <= 32'h0;
      v0_744 <= 32'h0;
      v0_745 <= 32'h0;
      v0_746 <= 32'h0;
      v0_747 <= 32'h0;
      v0_748 <= 32'h0;
      v0_749 <= 32'h0;
      v0_750 <= 32'h0;
      v0_751 <= 32'h0;
      v0_752 <= 32'h0;
      v0_753 <= 32'h0;
      v0_754 <= 32'h0;
      v0_755 <= 32'h0;
      v0_756 <= 32'h0;
      v0_757 <= 32'h0;
      v0_758 <= 32'h0;
      v0_759 <= 32'h0;
      v0_760 <= 32'h0;
      v0_761 <= 32'h0;
      v0_762 <= 32'h0;
      v0_763 <= 32'h0;
      v0_764 <= 32'h0;
      v0_765 <= 32'h0;
      v0_766 <= 32'h0;
      v0_767 <= 32'h0;
      v0_768 <= 32'h0;
      v0_769 <= 32'h0;
      v0_770 <= 32'h0;
      v0_771 <= 32'h0;
      v0_772 <= 32'h0;
      v0_773 <= 32'h0;
      v0_774 <= 32'h0;
      v0_775 <= 32'h0;
      v0_776 <= 32'h0;
      v0_777 <= 32'h0;
      v0_778 <= 32'h0;
      v0_779 <= 32'h0;
      v0_780 <= 32'h0;
      v0_781 <= 32'h0;
      v0_782 <= 32'h0;
      v0_783 <= 32'h0;
      v0_784 <= 32'h0;
      v0_785 <= 32'h0;
      v0_786 <= 32'h0;
      v0_787 <= 32'h0;
      v0_788 <= 32'h0;
      v0_789 <= 32'h0;
      v0_790 <= 32'h0;
      v0_791 <= 32'h0;
      v0_792 <= 32'h0;
      v0_793 <= 32'h0;
      v0_794 <= 32'h0;
      v0_795 <= 32'h0;
      v0_796 <= 32'h0;
      v0_797 <= 32'h0;
      v0_798 <= 32'h0;
      v0_799 <= 32'h0;
      v0_800 <= 32'h0;
      v0_801 <= 32'h0;
      v0_802 <= 32'h0;
      v0_803 <= 32'h0;
      v0_804 <= 32'h0;
      v0_805 <= 32'h0;
      v0_806 <= 32'h0;
      v0_807 <= 32'h0;
      v0_808 <= 32'h0;
      v0_809 <= 32'h0;
      v0_810 <= 32'h0;
      v0_811 <= 32'h0;
      v0_812 <= 32'h0;
      v0_813 <= 32'h0;
      v0_814 <= 32'h0;
      v0_815 <= 32'h0;
      v0_816 <= 32'h0;
      v0_817 <= 32'h0;
      v0_818 <= 32'h0;
      v0_819 <= 32'h0;
      v0_820 <= 32'h0;
      v0_821 <= 32'h0;
      v0_822 <= 32'h0;
      v0_823 <= 32'h0;
      v0_824 <= 32'h0;
      v0_825 <= 32'h0;
      v0_826 <= 32'h0;
      v0_827 <= 32'h0;
      v0_828 <= 32'h0;
      v0_829 <= 32'h0;
      v0_830 <= 32'h0;
      v0_831 <= 32'h0;
      v0_832 <= 32'h0;
      v0_833 <= 32'h0;
      v0_834 <= 32'h0;
      v0_835 <= 32'h0;
      v0_836 <= 32'h0;
      v0_837 <= 32'h0;
      v0_838 <= 32'h0;
      v0_839 <= 32'h0;
      v0_840 <= 32'h0;
      v0_841 <= 32'h0;
      v0_842 <= 32'h0;
      v0_843 <= 32'h0;
      v0_844 <= 32'h0;
      v0_845 <= 32'h0;
      v0_846 <= 32'h0;
      v0_847 <= 32'h0;
      v0_848 <= 32'h0;
      v0_849 <= 32'h0;
      v0_850 <= 32'h0;
      v0_851 <= 32'h0;
      v0_852 <= 32'h0;
      v0_853 <= 32'h0;
      v0_854 <= 32'h0;
      v0_855 <= 32'h0;
      v0_856 <= 32'h0;
      v0_857 <= 32'h0;
      v0_858 <= 32'h0;
      v0_859 <= 32'h0;
      v0_860 <= 32'h0;
      v0_861 <= 32'h0;
      v0_862 <= 32'h0;
      v0_863 <= 32'h0;
      v0_864 <= 32'h0;
      v0_865 <= 32'h0;
      v0_866 <= 32'h0;
      v0_867 <= 32'h0;
      v0_868 <= 32'h0;
      v0_869 <= 32'h0;
      v0_870 <= 32'h0;
      v0_871 <= 32'h0;
      v0_872 <= 32'h0;
      v0_873 <= 32'h0;
      v0_874 <= 32'h0;
      v0_875 <= 32'h0;
      v0_876 <= 32'h0;
      v0_877 <= 32'h0;
      v0_878 <= 32'h0;
      v0_879 <= 32'h0;
      v0_880 <= 32'h0;
      v0_881 <= 32'h0;
      v0_882 <= 32'h0;
      v0_883 <= 32'h0;
      v0_884 <= 32'h0;
      v0_885 <= 32'h0;
      v0_886 <= 32'h0;
      v0_887 <= 32'h0;
      v0_888 <= 32'h0;
      v0_889 <= 32'h0;
      v0_890 <= 32'h0;
      v0_891 <= 32'h0;
      v0_892 <= 32'h0;
      v0_893 <= 32'h0;
      v0_894 <= 32'h0;
      v0_895 <= 32'h0;
      v0_896 <= 32'h0;
      v0_897 <= 32'h0;
      v0_898 <= 32'h0;
      v0_899 <= 32'h0;
      v0_900 <= 32'h0;
      v0_901 <= 32'h0;
      v0_902 <= 32'h0;
      v0_903 <= 32'h0;
      v0_904 <= 32'h0;
      v0_905 <= 32'h0;
      v0_906 <= 32'h0;
      v0_907 <= 32'h0;
      v0_908 <= 32'h0;
      v0_909 <= 32'h0;
      v0_910 <= 32'h0;
      v0_911 <= 32'h0;
      v0_912 <= 32'h0;
      v0_913 <= 32'h0;
      v0_914 <= 32'h0;
      v0_915 <= 32'h0;
      v0_916 <= 32'h0;
      v0_917 <= 32'h0;
      v0_918 <= 32'h0;
      v0_919 <= 32'h0;
      v0_920 <= 32'h0;
      v0_921 <= 32'h0;
      v0_922 <= 32'h0;
      v0_923 <= 32'h0;
      v0_924 <= 32'h0;
      v0_925 <= 32'h0;
      v0_926 <= 32'h0;
      v0_927 <= 32'h0;
      v0_928 <= 32'h0;
      v0_929 <= 32'h0;
      v0_930 <= 32'h0;
      v0_931 <= 32'h0;
      v0_932 <= 32'h0;
      v0_933 <= 32'h0;
      v0_934 <= 32'h0;
      v0_935 <= 32'h0;
      v0_936 <= 32'h0;
      v0_937 <= 32'h0;
      v0_938 <= 32'h0;
      v0_939 <= 32'h0;
      v0_940 <= 32'h0;
      v0_941 <= 32'h0;
      v0_942 <= 32'h0;
      v0_943 <= 32'h0;
      v0_944 <= 32'h0;
      v0_945 <= 32'h0;
      v0_946 <= 32'h0;
      v0_947 <= 32'h0;
      v0_948 <= 32'h0;
      v0_949 <= 32'h0;
      v0_950 <= 32'h0;
      v0_951 <= 32'h0;
      v0_952 <= 32'h0;
      v0_953 <= 32'h0;
      v0_954 <= 32'h0;
      v0_955 <= 32'h0;
      v0_956 <= 32'h0;
      v0_957 <= 32'h0;
      v0_958 <= 32'h0;
      v0_959 <= 32'h0;
      v0_960 <= 32'h0;
      v0_961 <= 32'h0;
      v0_962 <= 32'h0;
      v0_963 <= 32'h0;
      v0_964 <= 32'h0;
      v0_965 <= 32'h0;
      v0_966 <= 32'h0;
      v0_967 <= 32'h0;
      v0_968 <= 32'h0;
      v0_969 <= 32'h0;
      v0_970 <= 32'h0;
      v0_971 <= 32'h0;
      v0_972 <= 32'h0;
      v0_973 <= 32'h0;
      v0_974 <= 32'h0;
      v0_975 <= 32'h0;
      v0_976 <= 32'h0;
      v0_977 <= 32'h0;
      v0_978 <= 32'h0;
      v0_979 <= 32'h0;
      v0_980 <= 32'h0;
      v0_981 <= 32'h0;
      v0_982 <= 32'h0;
      v0_983 <= 32'h0;
      v0_984 <= 32'h0;
      v0_985 <= 32'h0;
      v0_986 <= 32'h0;
      v0_987 <= 32'h0;
      v0_988 <= 32'h0;
      v0_989 <= 32'h0;
      v0_990 <= 32'h0;
      v0_991 <= 32'h0;
      v0_992 <= 32'h0;
      v0_993 <= 32'h0;
      v0_994 <= 32'h0;
      v0_995 <= 32'h0;
      v0_996 <= 32'h0;
      v0_997 <= 32'h0;
      v0_998 <= 32'h0;
      v0_999 <= 32'h0;
      v0_1000 <= 32'h0;
      v0_1001 <= 32'h0;
      v0_1002 <= 32'h0;
      v0_1003 <= 32'h0;
      v0_1004 <= 32'h0;
      v0_1005 <= 32'h0;
      v0_1006 <= 32'h0;
      v0_1007 <= 32'h0;
      v0_1008 <= 32'h0;
      v0_1009 <= 32'h0;
      v0_1010 <= 32'h0;
      v0_1011 <= 32'h0;
      v0_1012 <= 32'h0;
      v0_1013 <= 32'h0;
      v0_1014 <= 32'h0;
      v0_1015 <= 32'h0;
      v0_1016 <= 32'h0;
      v0_1017 <= 32'h0;
      v0_1018 <= 32'h0;
      v0_1019 <= 32'h0;
      v0_1020 <= 32'h0;
      v0_1021 <= 32'h0;
      v0_1022 <= 32'h0;
      v0_1023 <= 32'h0;
      queueCount_0 <= 7'h0;
      queueCount_1 <= 7'h0;
      queueCount_2 <= 7'h0;
      queueCount_3 <= 7'h0;
      queueCount_4 <= 7'h0;
      queueCount_5 <= 7'h0;
      queueCount_6 <= 7'h0;
      queueCount_7 <= 7'h0;
      queueCount_0_1 <= 7'h0;
      queueCount_1_1 <= 7'h0;
      queueCount_2_1 <= 7'h0;
      queueCount_3_1 <= 7'h0;
      queueCount_4_1 <= 7'h0;
      queueCount_5_1 <= 7'h0;
      queueCount_6_1 <= 7'h0;
      queueCount_7_1 <= 7'h0;
      queueCount_0_2 <= 7'h0;
      queueCount_1_2 <= 7'h0;
      queueCount_2_2 <= 7'h0;
      queueCount_3_2 <= 7'h0;
      queueCount_4_2 <= 7'h0;
      queueCount_5_2 <= 7'h0;
      queueCount_6_2 <= 7'h0;
      queueCount_7_2 <= 7'h0;
      queueCount_0_3 <= 7'h0;
      queueCount_1_3 <= 7'h0;
      queueCount_2_3 <= 7'h0;
      queueCount_3_3 <= 7'h0;
      queueCount_4_3 <= 7'h0;
      queueCount_5_3 <= 7'h0;
      queueCount_6_3 <= 7'h0;
      queueCount_7_3 <= 7'h0;
    end
    else begin
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h0)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h0)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h0)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h0)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h1)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h1)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h1)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h1)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h2)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h2)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h2)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h2)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h3)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h3)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h3)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h3)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h4)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h4)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h4)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h4)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h5)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h5)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h5)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h5)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h6)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h6)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h6)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h6)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h7)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h7)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h7)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h7)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h8)
        v0_32 <= v0_32 & ~maskExt_32 | maskExt_32 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h8)
        v0_33 <= v0_33 & ~maskExt_33 | maskExt_33 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h8)
        v0_34 <= v0_34 & ~maskExt_34 | maskExt_34 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h8)
        v0_35 <= v0_35 & ~maskExt_35 | maskExt_35 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h9)
        v0_36 <= v0_36 & ~maskExt_36 | maskExt_36 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h9)
        v0_37 <= v0_37 & ~maskExt_37 | maskExt_37 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h9)
        v0_38 <= v0_38 & ~maskExt_38 | maskExt_38 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h9)
        v0_39 <= v0_39 & ~maskExt_39 | maskExt_39 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA)
        v0_40 <= v0_40 & ~maskExt_40 | maskExt_40 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA)
        v0_41 <= v0_41 & ~maskExt_41 | maskExt_41 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA)
        v0_42 <= v0_42 & ~maskExt_42 | maskExt_42 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA)
        v0_43 <= v0_43 & ~maskExt_43 | maskExt_43 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB)
        v0_44 <= v0_44 & ~maskExt_44 | maskExt_44 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB)
        v0_45 <= v0_45 & ~maskExt_45 | maskExt_45 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB)
        v0_46 <= v0_46 & ~maskExt_46 | maskExt_46 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB)
        v0_47 <= v0_47 & ~maskExt_47 | maskExt_47 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC)
        v0_48 <= v0_48 & ~maskExt_48 | maskExt_48 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC)
        v0_49 <= v0_49 & ~maskExt_49 | maskExt_49 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC)
        v0_50 <= v0_50 & ~maskExt_50 | maskExt_50 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC)
        v0_51 <= v0_51 & ~maskExt_51 | maskExt_51 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD)
        v0_52 <= v0_52 & ~maskExt_52 | maskExt_52 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD)
        v0_53 <= v0_53 & ~maskExt_53 | maskExt_53 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD)
        v0_54 <= v0_54 & ~maskExt_54 | maskExt_54 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD)
        v0_55 <= v0_55 & ~maskExt_55 | maskExt_55 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE)
        v0_56 <= v0_56 & ~maskExt_56 | maskExt_56 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE)
        v0_57 <= v0_57 & ~maskExt_57 | maskExt_57 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE)
        v0_58 <= v0_58 & ~maskExt_58 | maskExt_58 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE)
        v0_59 <= v0_59 & ~maskExt_59 | maskExt_59 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF)
        v0_60 <= v0_60 & ~maskExt_60 | maskExt_60 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF)
        v0_61 <= v0_61 & ~maskExt_61 | maskExt_61 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF)
        v0_62 <= v0_62 & ~maskExt_62 | maskExt_62 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF)
        v0_63 <= v0_63 & ~maskExt_63 | maskExt_63 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h10)
        v0_64 <= v0_64 & ~maskExt_64 | maskExt_64 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h10)
        v0_65 <= v0_65 & ~maskExt_65 | maskExt_65 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h10)
        v0_66 <= v0_66 & ~maskExt_66 | maskExt_66 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h10)
        v0_67 <= v0_67 & ~maskExt_67 | maskExt_67 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h11)
        v0_68 <= v0_68 & ~maskExt_68 | maskExt_68 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h11)
        v0_69 <= v0_69 & ~maskExt_69 | maskExt_69 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h11)
        v0_70 <= v0_70 & ~maskExt_70 | maskExt_70 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h11)
        v0_71 <= v0_71 & ~maskExt_71 | maskExt_71 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h12)
        v0_72 <= v0_72 & ~maskExt_72 | maskExt_72 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h12)
        v0_73 <= v0_73 & ~maskExt_73 | maskExt_73 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h12)
        v0_74 <= v0_74 & ~maskExt_74 | maskExt_74 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h12)
        v0_75 <= v0_75 & ~maskExt_75 | maskExt_75 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h13)
        v0_76 <= v0_76 & ~maskExt_76 | maskExt_76 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h13)
        v0_77 <= v0_77 & ~maskExt_77 | maskExt_77 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h13)
        v0_78 <= v0_78 & ~maskExt_78 | maskExt_78 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h13)
        v0_79 <= v0_79 & ~maskExt_79 | maskExt_79 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h14)
        v0_80 <= v0_80 & ~maskExt_80 | maskExt_80 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h14)
        v0_81 <= v0_81 & ~maskExt_81 | maskExt_81 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h14)
        v0_82 <= v0_82 & ~maskExt_82 | maskExt_82 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h14)
        v0_83 <= v0_83 & ~maskExt_83 | maskExt_83 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h15)
        v0_84 <= v0_84 & ~maskExt_84 | maskExt_84 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h15)
        v0_85 <= v0_85 & ~maskExt_85 | maskExt_85 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h15)
        v0_86 <= v0_86 & ~maskExt_86 | maskExt_86 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h15)
        v0_87 <= v0_87 & ~maskExt_87 | maskExt_87 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h16)
        v0_88 <= v0_88 & ~maskExt_88 | maskExt_88 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h16)
        v0_89 <= v0_89 & ~maskExt_89 | maskExt_89 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h16)
        v0_90 <= v0_90 & ~maskExt_90 | maskExt_90 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h16)
        v0_91 <= v0_91 & ~maskExt_91 | maskExt_91 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h17)
        v0_92 <= v0_92 & ~maskExt_92 | maskExt_92 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h17)
        v0_93 <= v0_93 & ~maskExt_93 | maskExt_93 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h17)
        v0_94 <= v0_94 & ~maskExt_94 | maskExt_94 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h17)
        v0_95 <= v0_95 & ~maskExt_95 | maskExt_95 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h18)
        v0_96 <= v0_96 & ~maskExt_96 | maskExt_96 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h18)
        v0_97 <= v0_97 & ~maskExt_97 | maskExt_97 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h18)
        v0_98 <= v0_98 & ~maskExt_98 | maskExt_98 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h18)
        v0_99 <= v0_99 & ~maskExt_99 | maskExt_99 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h19)
        v0_100 <= v0_100 & ~maskExt_100 | maskExt_100 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h19)
        v0_101 <= v0_101 & ~maskExt_101 | maskExt_101 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h19)
        v0_102 <= v0_102 & ~maskExt_102 | maskExt_102 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h19)
        v0_103 <= v0_103 & ~maskExt_103 | maskExt_103 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h1A)
        v0_104 <= v0_104 & ~maskExt_104 | maskExt_104 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h1A)
        v0_105 <= v0_105 & ~maskExt_105 | maskExt_105 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h1A)
        v0_106 <= v0_106 & ~maskExt_106 | maskExt_106 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h1A)
        v0_107 <= v0_107 & ~maskExt_107 | maskExt_107 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h1B)
        v0_108 <= v0_108 & ~maskExt_108 | maskExt_108 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h1B)
        v0_109 <= v0_109 & ~maskExt_109 | maskExt_109 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h1B)
        v0_110 <= v0_110 & ~maskExt_110 | maskExt_110 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h1B)
        v0_111 <= v0_111 & ~maskExt_111 | maskExt_111 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h1C)
        v0_112 <= v0_112 & ~maskExt_112 | maskExt_112 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h1C)
        v0_113 <= v0_113 & ~maskExt_113 | maskExt_113 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h1C)
        v0_114 <= v0_114 & ~maskExt_114 | maskExt_114 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h1C)
        v0_115 <= v0_115 & ~maskExt_115 | maskExt_115 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h1D)
        v0_116 <= v0_116 & ~maskExt_116 | maskExt_116 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h1D)
        v0_117 <= v0_117 & ~maskExt_117 | maskExt_117 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h1D)
        v0_118 <= v0_118 & ~maskExt_118 | maskExt_118 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h1D)
        v0_119 <= v0_119 & ~maskExt_119 | maskExt_119 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h1E)
        v0_120 <= v0_120 & ~maskExt_120 | maskExt_120 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h1E)
        v0_121 <= v0_121 & ~maskExt_121 | maskExt_121 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h1E)
        v0_122 <= v0_122 & ~maskExt_122 | maskExt_122 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h1E)
        v0_123 <= v0_123 & ~maskExt_123 | maskExt_123 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h1F)
        v0_124 <= v0_124 & ~maskExt_124 | maskExt_124 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h1F)
        v0_125 <= v0_125 & ~maskExt_125 | maskExt_125 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h1F)
        v0_126 <= v0_126 & ~maskExt_126 | maskExt_126 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h1F)
        v0_127 <= v0_127 & ~maskExt_127 | maskExt_127 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h20)
        v0_128 <= v0_128 & ~maskExt_128 | maskExt_128 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h20)
        v0_129 <= v0_129 & ~maskExt_129 | maskExt_129 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h20)
        v0_130 <= v0_130 & ~maskExt_130 | maskExt_130 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h20)
        v0_131 <= v0_131 & ~maskExt_131 | maskExt_131 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h21)
        v0_132 <= v0_132 & ~maskExt_132 | maskExt_132 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h21)
        v0_133 <= v0_133 & ~maskExt_133 | maskExt_133 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h21)
        v0_134 <= v0_134 & ~maskExt_134 | maskExt_134 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h21)
        v0_135 <= v0_135 & ~maskExt_135 | maskExt_135 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h22)
        v0_136 <= v0_136 & ~maskExt_136 | maskExt_136 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h22)
        v0_137 <= v0_137 & ~maskExt_137 | maskExt_137 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h22)
        v0_138 <= v0_138 & ~maskExt_138 | maskExt_138 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h22)
        v0_139 <= v0_139 & ~maskExt_139 | maskExt_139 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h23)
        v0_140 <= v0_140 & ~maskExt_140 | maskExt_140 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h23)
        v0_141 <= v0_141 & ~maskExt_141 | maskExt_141 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h23)
        v0_142 <= v0_142 & ~maskExt_142 | maskExt_142 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h23)
        v0_143 <= v0_143 & ~maskExt_143 | maskExt_143 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h24)
        v0_144 <= v0_144 & ~maskExt_144 | maskExt_144 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h24)
        v0_145 <= v0_145 & ~maskExt_145 | maskExt_145 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h24)
        v0_146 <= v0_146 & ~maskExt_146 | maskExt_146 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h24)
        v0_147 <= v0_147 & ~maskExt_147 | maskExt_147 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h25)
        v0_148 <= v0_148 & ~maskExt_148 | maskExt_148 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h25)
        v0_149 <= v0_149 & ~maskExt_149 | maskExt_149 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h25)
        v0_150 <= v0_150 & ~maskExt_150 | maskExt_150 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h25)
        v0_151 <= v0_151 & ~maskExt_151 | maskExt_151 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h26)
        v0_152 <= v0_152 & ~maskExt_152 | maskExt_152 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h26)
        v0_153 <= v0_153 & ~maskExt_153 | maskExt_153 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h26)
        v0_154 <= v0_154 & ~maskExt_154 | maskExt_154 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h26)
        v0_155 <= v0_155 & ~maskExt_155 | maskExt_155 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h27)
        v0_156 <= v0_156 & ~maskExt_156 | maskExt_156 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h27)
        v0_157 <= v0_157 & ~maskExt_157 | maskExt_157 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h27)
        v0_158 <= v0_158 & ~maskExt_158 | maskExt_158 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h27)
        v0_159 <= v0_159 & ~maskExt_159 | maskExt_159 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h28)
        v0_160 <= v0_160 & ~maskExt_160 | maskExt_160 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h28)
        v0_161 <= v0_161 & ~maskExt_161 | maskExt_161 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h28)
        v0_162 <= v0_162 & ~maskExt_162 | maskExt_162 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h28)
        v0_163 <= v0_163 & ~maskExt_163 | maskExt_163 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h29)
        v0_164 <= v0_164 & ~maskExt_164 | maskExt_164 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h29)
        v0_165 <= v0_165 & ~maskExt_165 | maskExt_165 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h29)
        v0_166 <= v0_166 & ~maskExt_166 | maskExt_166 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h29)
        v0_167 <= v0_167 & ~maskExt_167 | maskExt_167 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h2A)
        v0_168 <= v0_168 & ~maskExt_168 | maskExt_168 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h2A)
        v0_169 <= v0_169 & ~maskExt_169 | maskExt_169 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h2A)
        v0_170 <= v0_170 & ~maskExt_170 | maskExt_170 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h2A)
        v0_171 <= v0_171 & ~maskExt_171 | maskExt_171 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h2B)
        v0_172 <= v0_172 & ~maskExt_172 | maskExt_172 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h2B)
        v0_173 <= v0_173 & ~maskExt_173 | maskExt_173 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h2B)
        v0_174 <= v0_174 & ~maskExt_174 | maskExt_174 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h2B)
        v0_175 <= v0_175 & ~maskExt_175 | maskExt_175 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h2C)
        v0_176 <= v0_176 & ~maskExt_176 | maskExt_176 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h2C)
        v0_177 <= v0_177 & ~maskExt_177 | maskExt_177 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h2C)
        v0_178 <= v0_178 & ~maskExt_178 | maskExt_178 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h2C)
        v0_179 <= v0_179 & ~maskExt_179 | maskExt_179 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h2D)
        v0_180 <= v0_180 & ~maskExt_180 | maskExt_180 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h2D)
        v0_181 <= v0_181 & ~maskExt_181 | maskExt_181 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h2D)
        v0_182 <= v0_182 & ~maskExt_182 | maskExt_182 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h2D)
        v0_183 <= v0_183 & ~maskExt_183 | maskExt_183 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h2E)
        v0_184 <= v0_184 & ~maskExt_184 | maskExt_184 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h2E)
        v0_185 <= v0_185 & ~maskExt_185 | maskExt_185 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h2E)
        v0_186 <= v0_186 & ~maskExt_186 | maskExt_186 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h2E)
        v0_187 <= v0_187 & ~maskExt_187 | maskExt_187 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h2F)
        v0_188 <= v0_188 & ~maskExt_188 | maskExt_188 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h2F)
        v0_189 <= v0_189 & ~maskExt_189 | maskExt_189 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h2F)
        v0_190 <= v0_190 & ~maskExt_190 | maskExt_190 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h2F)
        v0_191 <= v0_191 & ~maskExt_191 | maskExt_191 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h30)
        v0_192 <= v0_192 & ~maskExt_192 | maskExt_192 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h30)
        v0_193 <= v0_193 & ~maskExt_193 | maskExt_193 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h30)
        v0_194 <= v0_194 & ~maskExt_194 | maskExt_194 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h30)
        v0_195 <= v0_195 & ~maskExt_195 | maskExt_195 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h31)
        v0_196 <= v0_196 & ~maskExt_196 | maskExt_196 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h31)
        v0_197 <= v0_197 & ~maskExt_197 | maskExt_197 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h31)
        v0_198 <= v0_198 & ~maskExt_198 | maskExt_198 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h31)
        v0_199 <= v0_199 & ~maskExt_199 | maskExt_199 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h32)
        v0_200 <= v0_200 & ~maskExt_200 | maskExt_200 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h32)
        v0_201 <= v0_201 & ~maskExt_201 | maskExt_201 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h32)
        v0_202 <= v0_202 & ~maskExt_202 | maskExt_202 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h32)
        v0_203 <= v0_203 & ~maskExt_203 | maskExt_203 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h33)
        v0_204 <= v0_204 & ~maskExt_204 | maskExt_204 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h33)
        v0_205 <= v0_205 & ~maskExt_205 | maskExt_205 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h33)
        v0_206 <= v0_206 & ~maskExt_206 | maskExt_206 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h33)
        v0_207 <= v0_207 & ~maskExt_207 | maskExt_207 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h34)
        v0_208 <= v0_208 & ~maskExt_208 | maskExt_208 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h34)
        v0_209 <= v0_209 & ~maskExt_209 | maskExt_209 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h34)
        v0_210 <= v0_210 & ~maskExt_210 | maskExt_210 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h34)
        v0_211 <= v0_211 & ~maskExt_211 | maskExt_211 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h35)
        v0_212 <= v0_212 & ~maskExt_212 | maskExt_212 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h35)
        v0_213 <= v0_213 & ~maskExt_213 | maskExt_213 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h35)
        v0_214 <= v0_214 & ~maskExt_214 | maskExt_214 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h35)
        v0_215 <= v0_215 & ~maskExt_215 | maskExt_215 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h36)
        v0_216 <= v0_216 & ~maskExt_216 | maskExt_216 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h36)
        v0_217 <= v0_217 & ~maskExt_217 | maskExt_217 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h36)
        v0_218 <= v0_218 & ~maskExt_218 | maskExt_218 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h36)
        v0_219 <= v0_219 & ~maskExt_219 | maskExt_219 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h37)
        v0_220 <= v0_220 & ~maskExt_220 | maskExt_220 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h37)
        v0_221 <= v0_221 & ~maskExt_221 | maskExt_221 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h37)
        v0_222 <= v0_222 & ~maskExt_222 | maskExt_222 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h37)
        v0_223 <= v0_223 & ~maskExt_223 | maskExt_223 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h38)
        v0_224 <= v0_224 & ~maskExt_224 | maskExt_224 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h38)
        v0_225 <= v0_225 & ~maskExt_225 | maskExt_225 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h38)
        v0_226 <= v0_226 & ~maskExt_226 | maskExt_226 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h38)
        v0_227 <= v0_227 & ~maskExt_227 | maskExt_227 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h39)
        v0_228 <= v0_228 & ~maskExt_228 | maskExt_228 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h39)
        v0_229 <= v0_229 & ~maskExt_229 | maskExt_229 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h39)
        v0_230 <= v0_230 & ~maskExt_230 | maskExt_230 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h39)
        v0_231 <= v0_231 & ~maskExt_231 | maskExt_231 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h3A)
        v0_232 <= v0_232 & ~maskExt_232 | maskExt_232 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h3A)
        v0_233 <= v0_233 & ~maskExt_233 | maskExt_233 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h3A)
        v0_234 <= v0_234 & ~maskExt_234 | maskExt_234 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h3A)
        v0_235 <= v0_235 & ~maskExt_235 | maskExt_235 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h3B)
        v0_236 <= v0_236 & ~maskExt_236 | maskExt_236 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h3B)
        v0_237 <= v0_237 & ~maskExt_237 | maskExt_237 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h3B)
        v0_238 <= v0_238 & ~maskExt_238 | maskExt_238 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h3B)
        v0_239 <= v0_239 & ~maskExt_239 | maskExt_239 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h3C)
        v0_240 <= v0_240 & ~maskExt_240 | maskExt_240 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h3C)
        v0_241 <= v0_241 & ~maskExt_241 | maskExt_241 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h3C)
        v0_242 <= v0_242 & ~maskExt_242 | maskExt_242 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h3C)
        v0_243 <= v0_243 & ~maskExt_243 | maskExt_243 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h3D)
        v0_244 <= v0_244 & ~maskExt_244 | maskExt_244 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h3D)
        v0_245 <= v0_245 & ~maskExt_245 | maskExt_245 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h3D)
        v0_246 <= v0_246 & ~maskExt_246 | maskExt_246 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h3D)
        v0_247 <= v0_247 & ~maskExt_247 | maskExt_247 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h3E)
        v0_248 <= v0_248 & ~maskExt_248 | maskExt_248 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h3E)
        v0_249 <= v0_249 & ~maskExt_249 | maskExt_249 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h3E)
        v0_250 <= v0_250 & ~maskExt_250 | maskExt_250 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h3E)
        v0_251 <= v0_251 & ~maskExt_251 | maskExt_251 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h3F)
        v0_252 <= v0_252 & ~maskExt_252 | maskExt_252 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h3F)
        v0_253 <= v0_253 & ~maskExt_253 | maskExt_253 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h3F)
        v0_254 <= v0_254 & ~maskExt_254 | maskExt_254 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h3F)
        v0_255 <= v0_255 & ~maskExt_255 | maskExt_255 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h40)
        v0_256 <= v0_256 & ~maskExt_256 | maskExt_256 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h40)
        v0_257 <= v0_257 & ~maskExt_257 | maskExt_257 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h40)
        v0_258 <= v0_258 & ~maskExt_258 | maskExt_258 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h40)
        v0_259 <= v0_259 & ~maskExt_259 | maskExt_259 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h41)
        v0_260 <= v0_260 & ~maskExt_260 | maskExt_260 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h41)
        v0_261 <= v0_261 & ~maskExt_261 | maskExt_261 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h41)
        v0_262 <= v0_262 & ~maskExt_262 | maskExt_262 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h41)
        v0_263 <= v0_263 & ~maskExt_263 | maskExt_263 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h42)
        v0_264 <= v0_264 & ~maskExt_264 | maskExt_264 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h42)
        v0_265 <= v0_265 & ~maskExt_265 | maskExt_265 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h42)
        v0_266 <= v0_266 & ~maskExt_266 | maskExt_266 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h42)
        v0_267 <= v0_267 & ~maskExt_267 | maskExt_267 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h43)
        v0_268 <= v0_268 & ~maskExt_268 | maskExt_268 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h43)
        v0_269 <= v0_269 & ~maskExt_269 | maskExt_269 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h43)
        v0_270 <= v0_270 & ~maskExt_270 | maskExt_270 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h43)
        v0_271 <= v0_271 & ~maskExt_271 | maskExt_271 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h44)
        v0_272 <= v0_272 & ~maskExt_272 | maskExt_272 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h44)
        v0_273 <= v0_273 & ~maskExt_273 | maskExt_273 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h44)
        v0_274 <= v0_274 & ~maskExt_274 | maskExt_274 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h44)
        v0_275 <= v0_275 & ~maskExt_275 | maskExt_275 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h45)
        v0_276 <= v0_276 & ~maskExt_276 | maskExt_276 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h45)
        v0_277 <= v0_277 & ~maskExt_277 | maskExt_277 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h45)
        v0_278 <= v0_278 & ~maskExt_278 | maskExt_278 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h45)
        v0_279 <= v0_279 & ~maskExt_279 | maskExt_279 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h46)
        v0_280 <= v0_280 & ~maskExt_280 | maskExt_280 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h46)
        v0_281 <= v0_281 & ~maskExt_281 | maskExt_281 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h46)
        v0_282 <= v0_282 & ~maskExt_282 | maskExt_282 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h46)
        v0_283 <= v0_283 & ~maskExt_283 | maskExt_283 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h47)
        v0_284 <= v0_284 & ~maskExt_284 | maskExt_284 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h47)
        v0_285 <= v0_285 & ~maskExt_285 | maskExt_285 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h47)
        v0_286 <= v0_286 & ~maskExt_286 | maskExt_286 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h47)
        v0_287 <= v0_287 & ~maskExt_287 | maskExt_287 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h48)
        v0_288 <= v0_288 & ~maskExt_288 | maskExt_288 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h48)
        v0_289 <= v0_289 & ~maskExt_289 | maskExt_289 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h48)
        v0_290 <= v0_290 & ~maskExt_290 | maskExt_290 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h48)
        v0_291 <= v0_291 & ~maskExt_291 | maskExt_291 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h49)
        v0_292 <= v0_292 & ~maskExt_292 | maskExt_292 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h49)
        v0_293 <= v0_293 & ~maskExt_293 | maskExt_293 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h49)
        v0_294 <= v0_294 & ~maskExt_294 | maskExt_294 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h49)
        v0_295 <= v0_295 & ~maskExt_295 | maskExt_295 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h4A)
        v0_296 <= v0_296 & ~maskExt_296 | maskExt_296 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h4A)
        v0_297 <= v0_297 & ~maskExt_297 | maskExt_297 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h4A)
        v0_298 <= v0_298 & ~maskExt_298 | maskExt_298 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h4A)
        v0_299 <= v0_299 & ~maskExt_299 | maskExt_299 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h4B)
        v0_300 <= v0_300 & ~maskExt_300 | maskExt_300 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h4B)
        v0_301 <= v0_301 & ~maskExt_301 | maskExt_301 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h4B)
        v0_302 <= v0_302 & ~maskExt_302 | maskExt_302 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h4B)
        v0_303 <= v0_303 & ~maskExt_303 | maskExt_303 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h4C)
        v0_304 <= v0_304 & ~maskExt_304 | maskExt_304 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h4C)
        v0_305 <= v0_305 & ~maskExt_305 | maskExt_305 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h4C)
        v0_306 <= v0_306 & ~maskExt_306 | maskExt_306 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h4C)
        v0_307 <= v0_307 & ~maskExt_307 | maskExt_307 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h4D)
        v0_308 <= v0_308 & ~maskExt_308 | maskExt_308 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h4D)
        v0_309 <= v0_309 & ~maskExt_309 | maskExt_309 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h4D)
        v0_310 <= v0_310 & ~maskExt_310 | maskExt_310 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h4D)
        v0_311 <= v0_311 & ~maskExt_311 | maskExt_311 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h4E)
        v0_312 <= v0_312 & ~maskExt_312 | maskExt_312 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h4E)
        v0_313 <= v0_313 & ~maskExt_313 | maskExt_313 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h4E)
        v0_314 <= v0_314 & ~maskExt_314 | maskExt_314 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h4E)
        v0_315 <= v0_315 & ~maskExt_315 | maskExt_315 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h4F)
        v0_316 <= v0_316 & ~maskExt_316 | maskExt_316 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h4F)
        v0_317 <= v0_317 & ~maskExt_317 | maskExt_317 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h4F)
        v0_318 <= v0_318 & ~maskExt_318 | maskExt_318 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h4F)
        v0_319 <= v0_319 & ~maskExt_319 | maskExt_319 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h50)
        v0_320 <= v0_320 & ~maskExt_320 | maskExt_320 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h50)
        v0_321 <= v0_321 & ~maskExt_321 | maskExt_321 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h50)
        v0_322 <= v0_322 & ~maskExt_322 | maskExt_322 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h50)
        v0_323 <= v0_323 & ~maskExt_323 | maskExt_323 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h51)
        v0_324 <= v0_324 & ~maskExt_324 | maskExt_324 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h51)
        v0_325 <= v0_325 & ~maskExt_325 | maskExt_325 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h51)
        v0_326 <= v0_326 & ~maskExt_326 | maskExt_326 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h51)
        v0_327 <= v0_327 & ~maskExt_327 | maskExt_327 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h52)
        v0_328 <= v0_328 & ~maskExt_328 | maskExt_328 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h52)
        v0_329 <= v0_329 & ~maskExt_329 | maskExt_329 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h52)
        v0_330 <= v0_330 & ~maskExt_330 | maskExt_330 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h52)
        v0_331 <= v0_331 & ~maskExt_331 | maskExt_331 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h53)
        v0_332 <= v0_332 & ~maskExt_332 | maskExt_332 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h53)
        v0_333 <= v0_333 & ~maskExt_333 | maskExt_333 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h53)
        v0_334 <= v0_334 & ~maskExt_334 | maskExt_334 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h53)
        v0_335 <= v0_335 & ~maskExt_335 | maskExt_335 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h54)
        v0_336 <= v0_336 & ~maskExt_336 | maskExt_336 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h54)
        v0_337 <= v0_337 & ~maskExt_337 | maskExt_337 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h54)
        v0_338 <= v0_338 & ~maskExt_338 | maskExt_338 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h54)
        v0_339 <= v0_339 & ~maskExt_339 | maskExt_339 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h55)
        v0_340 <= v0_340 & ~maskExt_340 | maskExt_340 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h55)
        v0_341 <= v0_341 & ~maskExt_341 | maskExt_341 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h55)
        v0_342 <= v0_342 & ~maskExt_342 | maskExt_342 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h55)
        v0_343 <= v0_343 & ~maskExt_343 | maskExt_343 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h56)
        v0_344 <= v0_344 & ~maskExt_344 | maskExt_344 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h56)
        v0_345 <= v0_345 & ~maskExt_345 | maskExt_345 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h56)
        v0_346 <= v0_346 & ~maskExt_346 | maskExt_346 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h56)
        v0_347 <= v0_347 & ~maskExt_347 | maskExt_347 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h57)
        v0_348 <= v0_348 & ~maskExt_348 | maskExt_348 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h57)
        v0_349 <= v0_349 & ~maskExt_349 | maskExt_349 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h57)
        v0_350 <= v0_350 & ~maskExt_350 | maskExt_350 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h57)
        v0_351 <= v0_351 & ~maskExt_351 | maskExt_351 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h58)
        v0_352 <= v0_352 & ~maskExt_352 | maskExt_352 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h58)
        v0_353 <= v0_353 & ~maskExt_353 | maskExt_353 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h58)
        v0_354 <= v0_354 & ~maskExt_354 | maskExt_354 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h58)
        v0_355 <= v0_355 & ~maskExt_355 | maskExt_355 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h59)
        v0_356 <= v0_356 & ~maskExt_356 | maskExt_356 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h59)
        v0_357 <= v0_357 & ~maskExt_357 | maskExt_357 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h59)
        v0_358 <= v0_358 & ~maskExt_358 | maskExt_358 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h59)
        v0_359 <= v0_359 & ~maskExt_359 | maskExt_359 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h5A)
        v0_360 <= v0_360 & ~maskExt_360 | maskExt_360 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h5A)
        v0_361 <= v0_361 & ~maskExt_361 | maskExt_361 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h5A)
        v0_362 <= v0_362 & ~maskExt_362 | maskExt_362 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h5A)
        v0_363 <= v0_363 & ~maskExt_363 | maskExt_363 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h5B)
        v0_364 <= v0_364 & ~maskExt_364 | maskExt_364 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h5B)
        v0_365 <= v0_365 & ~maskExt_365 | maskExt_365 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h5B)
        v0_366 <= v0_366 & ~maskExt_366 | maskExt_366 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h5B)
        v0_367 <= v0_367 & ~maskExt_367 | maskExt_367 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h5C)
        v0_368 <= v0_368 & ~maskExt_368 | maskExt_368 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h5C)
        v0_369 <= v0_369 & ~maskExt_369 | maskExt_369 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h5C)
        v0_370 <= v0_370 & ~maskExt_370 | maskExt_370 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h5C)
        v0_371 <= v0_371 & ~maskExt_371 | maskExt_371 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h5D)
        v0_372 <= v0_372 & ~maskExt_372 | maskExt_372 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h5D)
        v0_373 <= v0_373 & ~maskExt_373 | maskExt_373 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h5D)
        v0_374 <= v0_374 & ~maskExt_374 | maskExt_374 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h5D)
        v0_375 <= v0_375 & ~maskExt_375 | maskExt_375 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h5E)
        v0_376 <= v0_376 & ~maskExt_376 | maskExt_376 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h5E)
        v0_377 <= v0_377 & ~maskExt_377 | maskExt_377 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h5E)
        v0_378 <= v0_378 & ~maskExt_378 | maskExt_378 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h5E)
        v0_379 <= v0_379 & ~maskExt_379 | maskExt_379 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h5F)
        v0_380 <= v0_380 & ~maskExt_380 | maskExt_380 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h5F)
        v0_381 <= v0_381 & ~maskExt_381 | maskExt_381 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h5F)
        v0_382 <= v0_382 & ~maskExt_382 | maskExt_382 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h5F)
        v0_383 <= v0_383 & ~maskExt_383 | maskExt_383 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h60)
        v0_384 <= v0_384 & ~maskExt_384 | maskExt_384 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h60)
        v0_385 <= v0_385 & ~maskExt_385 | maskExt_385 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h60)
        v0_386 <= v0_386 & ~maskExt_386 | maskExt_386 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h60)
        v0_387 <= v0_387 & ~maskExt_387 | maskExt_387 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h61)
        v0_388 <= v0_388 & ~maskExt_388 | maskExt_388 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h61)
        v0_389 <= v0_389 & ~maskExt_389 | maskExt_389 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h61)
        v0_390 <= v0_390 & ~maskExt_390 | maskExt_390 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h61)
        v0_391 <= v0_391 & ~maskExt_391 | maskExt_391 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h62)
        v0_392 <= v0_392 & ~maskExt_392 | maskExt_392 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h62)
        v0_393 <= v0_393 & ~maskExt_393 | maskExt_393 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h62)
        v0_394 <= v0_394 & ~maskExt_394 | maskExt_394 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h62)
        v0_395 <= v0_395 & ~maskExt_395 | maskExt_395 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h63)
        v0_396 <= v0_396 & ~maskExt_396 | maskExt_396 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h63)
        v0_397 <= v0_397 & ~maskExt_397 | maskExt_397 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h63)
        v0_398 <= v0_398 & ~maskExt_398 | maskExt_398 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h63)
        v0_399 <= v0_399 & ~maskExt_399 | maskExt_399 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h64)
        v0_400 <= v0_400 & ~maskExt_400 | maskExt_400 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h64)
        v0_401 <= v0_401 & ~maskExt_401 | maskExt_401 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h64)
        v0_402 <= v0_402 & ~maskExt_402 | maskExt_402 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h64)
        v0_403 <= v0_403 & ~maskExt_403 | maskExt_403 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h65)
        v0_404 <= v0_404 & ~maskExt_404 | maskExt_404 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h65)
        v0_405 <= v0_405 & ~maskExt_405 | maskExt_405 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h65)
        v0_406 <= v0_406 & ~maskExt_406 | maskExt_406 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h65)
        v0_407 <= v0_407 & ~maskExt_407 | maskExt_407 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h66)
        v0_408 <= v0_408 & ~maskExt_408 | maskExt_408 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h66)
        v0_409 <= v0_409 & ~maskExt_409 | maskExt_409 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h66)
        v0_410 <= v0_410 & ~maskExt_410 | maskExt_410 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h66)
        v0_411 <= v0_411 & ~maskExt_411 | maskExt_411 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h67)
        v0_412 <= v0_412 & ~maskExt_412 | maskExt_412 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h67)
        v0_413 <= v0_413 & ~maskExt_413 | maskExt_413 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h67)
        v0_414 <= v0_414 & ~maskExt_414 | maskExt_414 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h67)
        v0_415 <= v0_415 & ~maskExt_415 | maskExt_415 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h68)
        v0_416 <= v0_416 & ~maskExt_416 | maskExt_416 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h68)
        v0_417 <= v0_417 & ~maskExt_417 | maskExt_417 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h68)
        v0_418 <= v0_418 & ~maskExt_418 | maskExt_418 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h68)
        v0_419 <= v0_419 & ~maskExt_419 | maskExt_419 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h69)
        v0_420 <= v0_420 & ~maskExt_420 | maskExt_420 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h69)
        v0_421 <= v0_421 & ~maskExt_421 | maskExt_421 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h69)
        v0_422 <= v0_422 & ~maskExt_422 | maskExt_422 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h69)
        v0_423 <= v0_423 & ~maskExt_423 | maskExt_423 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h6A)
        v0_424 <= v0_424 & ~maskExt_424 | maskExt_424 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h6A)
        v0_425 <= v0_425 & ~maskExt_425 | maskExt_425 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h6A)
        v0_426 <= v0_426 & ~maskExt_426 | maskExt_426 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h6A)
        v0_427 <= v0_427 & ~maskExt_427 | maskExt_427 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h6B)
        v0_428 <= v0_428 & ~maskExt_428 | maskExt_428 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h6B)
        v0_429 <= v0_429 & ~maskExt_429 | maskExt_429 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h6B)
        v0_430 <= v0_430 & ~maskExt_430 | maskExt_430 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h6B)
        v0_431 <= v0_431 & ~maskExt_431 | maskExt_431 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h6C)
        v0_432 <= v0_432 & ~maskExt_432 | maskExt_432 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h6C)
        v0_433 <= v0_433 & ~maskExt_433 | maskExt_433 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h6C)
        v0_434 <= v0_434 & ~maskExt_434 | maskExt_434 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h6C)
        v0_435 <= v0_435 & ~maskExt_435 | maskExt_435 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h6D)
        v0_436 <= v0_436 & ~maskExt_436 | maskExt_436 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h6D)
        v0_437 <= v0_437 & ~maskExt_437 | maskExt_437 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h6D)
        v0_438 <= v0_438 & ~maskExt_438 | maskExt_438 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h6D)
        v0_439 <= v0_439 & ~maskExt_439 | maskExt_439 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h6E)
        v0_440 <= v0_440 & ~maskExt_440 | maskExt_440 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h6E)
        v0_441 <= v0_441 & ~maskExt_441 | maskExt_441 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h6E)
        v0_442 <= v0_442 & ~maskExt_442 | maskExt_442 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h6E)
        v0_443 <= v0_443 & ~maskExt_443 | maskExt_443 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h6F)
        v0_444 <= v0_444 & ~maskExt_444 | maskExt_444 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h6F)
        v0_445 <= v0_445 & ~maskExt_445 | maskExt_445 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h6F)
        v0_446 <= v0_446 & ~maskExt_446 | maskExt_446 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h6F)
        v0_447 <= v0_447 & ~maskExt_447 | maskExt_447 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h70)
        v0_448 <= v0_448 & ~maskExt_448 | maskExt_448 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h70)
        v0_449 <= v0_449 & ~maskExt_449 | maskExt_449 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h70)
        v0_450 <= v0_450 & ~maskExt_450 | maskExt_450 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h70)
        v0_451 <= v0_451 & ~maskExt_451 | maskExt_451 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h71)
        v0_452 <= v0_452 & ~maskExt_452 | maskExt_452 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h71)
        v0_453 <= v0_453 & ~maskExt_453 | maskExt_453 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h71)
        v0_454 <= v0_454 & ~maskExt_454 | maskExt_454 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h71)
        v0_455 <= v0_455 & ~maskExt_455 | maskExt_455 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h72)
        v0_456 <= v0_456 & ~maskExt_456 | maskExt_456 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h72)
        v0_457 <= v0_457 & ~maskExt_457 | maskExt_457 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h72)
        v0_458 <= v0_458 & ~maskExt_458 | maskExt_458 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h72)
        v0_459 <= v0_459 & ~maskExt_459 | maskExt_459 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h73)
        v0_460 <= v0_460 & ~maskExt_460 | maskExt_460 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h73)
        v0_461 <= v0_461 & ~maskExt_461 | maskExt_461 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h73)
        v0_462 <= v0_462 & ~maskExt_462 | maskExt_462 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h73)
        v0_463 <= v0_463 & ~maskExt_463 | maskExt_463 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h74)
        v0_464 <= v0_464 & ~maskExt_464 | maskExt_464 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h74)
        v0_465 <= v0_465 & ~maskExt_465 | maskExt_465 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h74)
        v0_466 <= v0_466 & ~maskExt_466 | maskExt_466 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h74)
        v0_467 <= v0_467 & ~maskExt_467 | maskExt_467 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h75)
        v0_468 <= v0_468 & ~maskExt_468 | maskExt_468 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h75)
        v0_469 <= v0_469 & ~maskExt_469 | maskExt_469 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h75)
        v0_470 <= v0_470 & ~maskExt_470 | maskExt_470 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h75)
        v0_471 <= v0_471 & ~maskExt_471 | maskExt_471 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h76)
        v0_472 <= v0_472 & ~maskExt_472 | maskExt_472 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h76)
        v0_473 <= v0_473 & ~maskExt_473 | maskExt_473 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h76)
        v0_474 <= v0_474 & ~maskExt_474 | maskExt_474 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h76)
        v0_475 <= v0_475 & ~maskExt_475 | maskExt_475 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h77)
        v0_476 <= v0_476 & ~maskExt_476 | maskExt_476 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h77)
        v0_477 <= v0_477 & ~maskExt_477 | maskExt_477 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h77)
        v0_478 <= v0_478 & ~maskExt_478 | maskExt_478 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h77)
        v0_479 <= v0_479 & ~maskExt_479 | maskExt_479 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h78)
        v0_480 <= v0_480 & ~maskExt_480 | maskExt_480 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h78)
        v0_481 <= v0_481 & ~maskExt_481 | maskExt_481 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h78)
        v0_482 <= v0_482 & ~maskExt_482 | maskExt_482 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h78)
        v0_483 <= v0_483 & ~maskExt_483 | maskExt_483 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h79)
        v0_484 <= v0_484 & ~maskExt_484 | maskExt_484 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h79)
        v0_485 <= v0_485 & ~maskExt_485 | maskExt_485 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h79)
        v0_486 <= v0_486 & ~maskExt_486 | maskExt_486 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h79)
        v0_487 <= v0_487 & ~maskExt_487 | maskExt_487 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h7A)
        v0_488 <= v0_488 & ~maskExt_488 | maskExt_488 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h7A)
        v0_489 <= v0_489 & ~maskExt_489 | maskExt_489 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h7A)
        v0_490 <= v0_490 & ~maskExt_490 | maskExt_490 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h7A)
        v0_491 <= v0_491 & ~maskExt_491 | maskExt_491 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h7B)
        v0_492 <= v0_492 & ~maskExt_492 | maskExt_492 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h7B)
        v0_493 <= v0_493 & ~maskExt_493 | maskExt_493 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h7B)
        v0_494 <= v0_494 & ~maskExt_494 | maskExt_494 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h7B)
        v0_495 <= v0_495 & ~maskExt_495 | maskExt_495 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h7C)
        v0_496 <= v0_496 & ~maskExt_496 | maskExt_496 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h7C)
        v0_497 <= v0_497 & ~maskExt_497 | maskExt_497 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h7C)
        v0_498 <= v0_498 & ~maskExt_498 | maskExt_498 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h7C)
        v0_499 <= v0_499 & ~maskExt_499 | maskExt_499 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h7D)
        v0_500 <= v0_500 & ~maskExt_500 | maskExt_500 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h7D)
        v0_501 <= v0_501 & ~maskExt_501 | maskExt_501 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h7D)
        v0_502 <= v0_502 & ~maskExt_502 | maskExt_502 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h7D)
        v0_503 <= v0_503 & ~maskExt_503 | maskExt_503 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h7E)
        v0_504 <= v0_504 & ~maskExt_504 | maskExt_504 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h7E)
        v0_505 <= v0_505 & ~maskExt_505 | maskExt_505 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h7E)
        v0_506 <= v0_506 & ~maskExt_506 | maskExt_506 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h7E)
        v0_507 <= v0_507 & ~maskExt_507 | maskExt_507 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h7F)
        v0_508 <= v0_508 & ~maskExt_508 | maskExt_508 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h7F)
        v0_509 <= v0_509 & ~maskExt_509 | maskExt_509 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h7F)
        v0_510 <= v0_510 & ~maskExt_510 | maskExt_510 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h7F)
        v0_511 <= v0_511 & ~maskExt_511 | maskExt_511 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h80)
        v0_512 <= v0_512 & ~maskExt_512 | maskExt_512 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h80)
        v0_513 <= v0_513 & ~maskExt_513 | maskExt_513 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h80)
        v0_514 <= v0_514 & ~maskExt_514 | maskExt_514 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h80)
        v0_515 <= v0_515 & ~maskExt_515 | maskExt_515 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h81)
        v0_516 <= v0_516 & ~maskExt_516 | maskExt_516 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h81)
        v0_517 <= v0_517 & ~maskExt_517 | maskExt_517 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h81)
        v0_518 <= v0_518 & ~maskExt_518 | maskExt_518 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h81)
        v0_519 <= v0_519 & ~maskExt_519 | maskExt_519 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h82)
        v0_520 <= v0_520 & ~maskExt_520 | maskExt_520 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h82)
        v0_521 <= v0_521 & ~maskExt_521 | maskExt_521 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h82)
        v0_522 <= v0_522 & ~maskExt_522 | maskExt_522 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h82)
        v0_523 <= v0_523 & ~maskExt_523 | maskExt_523 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h83)
        v0_524 <= v0_524 & ~maskExt_524 | maskExt_524 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h83)
        v0_525 <= v0_525 & ~maskExt_525 | maskExt_525 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h83)
        v0_526 <= v0_526 & ~maskExt_526 | maskExt_526 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h83)
        v0_527 <= v0_527 & ~maskExt_527 | maskExt_527 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h84)
        v0_528 <= v0_528 & ~maskExt_528 | maskExt_528 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h84)
        v0_529 <= v0_529 & ~maskExt_529 | maskExt_529 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h84)
        v0_530 <= v0_530 & ~maskExt_530 | maskExt_530 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h84)
        v0_531 <= v0_531 & ~maskExt_531 | maskExt_531 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h85)
        v0_532 <= v0_532 & ~maskExt_532 | maskExt_532 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h85)
        v0_533 <= v0_533 & ~maskExt_533 | maskExt_533 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h85)
        v0_534 <= v0_534 & ~maskExt_534 | maskExt_534 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h85)
        v0_535 <= v0_535 & ~maskExt_535 | maskExt_535 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h86)
        v0_536 <= v0_536 & ~maskExt_536 | maskExt_536 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h86)
        v0_537 <= v0_537 & ~maskExt_537 | maskExt_537 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h86)
        v0_538 <= v0_538 & ~maskExt_538 | maskExt_538 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h86)
        v0_539 <= v0_539 & ~maskExt_539 | maskExt_539 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h87)
        v0_540 <= v0_540 & ~maskExt_540 | maskExt_540 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h87)
        v0_541 <= v0_541 & ~maskExt_541 | maskExt_541 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h87)
        v0_542 <= v0_542 & ~maskExt_542 | maskExt_542 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h87)
        v0_543 <= v0_543 & ~maskExt_543 | maskExt_543 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h88)
        v0_544 <= v0_544 & ~maskExt_544 | maskExt_544 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h88)
        v0_545 <= v0_545 & ~maskExt_545 | maskExt_545 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h88)
        v0_546 <= v0_546 & ~maskExt_546 | maskExt_546 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h88)
        v0_547 <= v0_547 & ~maskExt_547 | maskExt_547 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h89)
        v0_548 <= v0_548 & ~maskExt_548 | maskExt_548 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h89)
        v0_549 <= v0_549 & ~maskExt_549 | maskExt_549 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h89)
        v0_550 <= v0_550 & ~maskExt_550 | maskExt_550 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h89)
        v0_551 <= v0_551 & ~maskExt_551 | maskExt_551 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h8A)
        v0_552 <= v0_552 & ~maskExt_552 | maskExt_552 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h8A)
        v0_553 <= v0_553 & ~maskExt_553 | maskExt_553 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h8A)
        v0_554 <= v0_554 & ~maskExt_554 | maskExt_554 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h8A)
        v0_555 <= v0_555 & ~maskExt_555 | maskExt_555 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h8B)
        v0_556 <= v0_556 & ~maskExt_556 | maskExt_556 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h8B)
        v0_557 <= v0_557 & ~maskExt_557 | maskExt_557 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h8B)
        v0_558 <= v0_558 & ~maskExt_558 | maskExt_558 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h8B)
        v0_559 <= v0_559 & ~maskExt_559 | maskExt_559 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h8C)
        v0_560 <= v0_560 & ~maskExt_560 | maskExt_560 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h8C)
        v0_561 <= v0_561 & ~maskExt_561 | maskExt_561 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h8C)
        v0_562 <= v0_562 & ~maskExt_562 | maskExt_562 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h8C)
        v0_563 <= v0_563 & ~maskExt_563 | maskExt_563 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h8D)
        v0_564 <= v0_564 & ~maskExt_564 | maskExt_564 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h8D)
        v0_565 <= v0_565 & ~maskExt_565 | maskExt_565 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h8D)
        v0_566 <= v0_566 & ~maskExt_566 | maskExt_566 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h8D)
        v0_567 <= v0_567 & ~maskExt_567 | maskExt_567 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h8E)
        v0_568 <= v0_568 & ~maskExt_568 | maskExt_568 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h8E)
        v0_569 <= v0_569 & ~maskExt_569 | maskExt_569 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h8E)
        v0_570 <= v0_570 & ~maskExt_570 | maskExt_570 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h8E)
        v0_571 <= v0_571 & ~maskExt_571 | maskExt_571 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h8F)
        v0_572 <= v0_572 & ~maskExt_572 | maskExt_572 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h8F)
        v0_573 <= v0_573 & ~maskExt_573 | maskExt_573 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h8F)
        v0_574 <= v0_574 & ~maskExt_574 | maskExt_574 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h8F)
        v0_575 <= v0_575 & ~maskExt_575 | maskExt_575 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h90)
        v0_576 <= v0_576 & ~maskExt_576 | maskExt_576 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h90)
        v0_577 <= v0_577 & ~maskExt_577 | maskExt_577 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h90)
        v0_578 <= v0_578 & ~maskExt_578 | maskExt_578 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h90)
        v0_579 <= v0_579 & ~maskExt_579 | maskExt_579 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h91)
        v0_580 <= v0_580 & ~maskExt_580 | maskExt_580 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h91)
        v0_581 <= v0_581 & ~maskExt_581 | maskExt_581 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h91)
        v0_582 <= v0_582 & ~maskExt_582 | maskExt_582 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h91)
        v0_583 <= v0_583 & ~maskExt_583 | maskExt_583 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h92)
        v0_584 <= v0_584 & ~maskExt_584 | maskExt_584 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h92)
        v0_585 <= v0_585 & ~maskExt_585 | maskExt_585 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h92)
        v0_586 <= v0_586 & ~maskExt_586 | maskExt_586 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h92)
        v0_587 <= v0_587 & ~maskExt_587 | maskExt_587 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h93)
        v0_588 <= v0_588 & ~maskExt_588 | maskExt_588 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h93)
        v0_589 <= v0_589 & ~maskExt_589 | maskExt_589 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h93)
        v0_590 <= v0_590 & ~maskExt_590 | maskExt_590 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h93)
        v0_591 <= v0_591 & ~maskExt_591 | maskExt_591 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h94)
        v0_592 <= v0_592 & ~maskExt_592 | maskExt_592 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h94)
        v0_593 <= v0_593 & ~maskExt_593 | maskExt_593 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h94)
        v0_594 <= v0_594 & ~maskExt_594 | maskExt_594 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h94)
        v0_595 <= v0_595 & ~maskExt_595 | maskExt_595 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h95)
        v0_596 <= v0_596 & ~maskExt_596 | maskExt_596 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h95)
        v0_597 <= v0_597 & ~maskExt_597 | maskExt_597 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h95)
        v0_598 <= v0_598 & ~maskExt_598 | maskExt_598 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h95)
        v0_599 <= v0_599 & ~maskExt_599 | maskExt_599 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h96)
        v0_600 <= v0_600 & ~maskExt_600 | maskExt_600 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h96)
        v0_601 <= v0_601 & ~maskExt_601 | maskExt_601 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h96)
        v0_602 <= v0_602 & ~maskExt_602 | maskExt_602 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h96)
        v0_603 <= v0_603 & ~maskExt_603 | maskExt_603 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h97)
        v0_604 <= v0_604 & ~maskExt_604 | maskExt_604 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h97)
        v0_605 <= v0_605 & ~maskExt_605 | maskExt_605 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h97)
        v0_606 <= v0_606 & ~maskExt_606 | maskExt_606 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h97)
        v0_607 <= v0_607 & ~maskExt_607 | maskExt_607 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h98)
        v0_608 <= v0_608 & ~maskExt_608 | maskExt_608 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h98)
        v0_609 <= v0_609 & ~maskExt_609 | maskExt_609 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h98)
        v0_610 <= v0_610 & ~maskExt_610 | maskExt_610 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h98)
        v0_611 <= v0_611 & ~maskExt_611 | maskExt_611 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h99)
        v0_612 <= v0_612 & ~maskExt_612 | maskExt_612 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h99)
        v0_613 <= v0_613 & ~maskExt_613 | maskExt_613 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h99)
        v0_614 <= v0_614 & ~maskExt_614 | maskExt_614 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h99)
        v0_615 <= v0_615 & ~maskExt_615 | maskExt_615 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h9A)
        v0_616 <= v0_616 & ~maskExt_616 | maskExt_616 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h9A)
        v0_617 <= v0_617 & ~maskExt_617 | maskExt_617 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h9A)
        v0_618 <= v0_618 & ~maskExt_618 | maskExt_618 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h9A)
        v0_619 <= v0_619 & ~maskExt_619 | maskExt_619 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h9B)
        v0_620 <= v0_620 & ~maskExt_620 | maskExt_620 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h9B)
        v0_621 <= v0_621 & ~maskExt_621 | maskExt_621 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h9B)
        v0_622 <= v0_622 & ~maskExt_622 | maskExt_622 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h9B)
        v0_623 <= v0_623 & ~maskExt_623 | maskExt_623 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h9C)
        v0_624 <= v0_624 & ~maskExt_624 | maskExt_624 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h9C)
        v0_625 <= v0_625 & ~maskExt_625 | maskExt_625 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h9C)
        v0_626 <= v0_626 & ~maskExt_626 | maskExt_626 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h9C)
        v0_627 <= v0_627 & ~maskExt_627 | maskExt_627 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h9D)
        v0_628 <= v0_628 & ~maskExt_628 | maskExt_628 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h9D)
        v0_629 <= v0_629 & ~maskExt_629 | maskExt_629 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h9D)
        v0_630 <= v0_630 & ~maskExt_630 | maskExt_630 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h9D)
        v0_631 <= v0_631 & ~maskExt_631 | maskExt_631 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h9E)
        v0_632 <= v0_632 & ~maskExt_632 | maskExt_632 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h9E)
        v0_633 <= v0_633 & ~maskExt_633 | maskExt_633 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h9E)
        v0_634 <= v0_634 & ~maskExt_634 | maskExt_634 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h9E)
        v0_635 <= v0_635 & ~maskExt_635 | maskExt_635 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'h9F)
        v0_636 <= v0_636 & ~maskExt_636 | maskExt_636 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'h9F)
        v0_637 <= v0_637 & ~maskExt_637 | maskExt_637 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'h9F)
        v0_638 <= v0_638 & ~maskExt_638 | maskExt_638 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'h9F)
        v0_639 <= v0_639 & ~maskExt_639 | maskExt_639 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA0)
        v0_640 <= v0_640 & ~maskExt_640 | maskExt_640 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA0)
        v0_641 <= v0_641 & ~maskExt_641 | maskExt_641 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA0)
        v0_642 <= v0_642 & ~maskExt_642 | maskExt_642 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA0)
        v0_643 <= v0_643 & ~maskExt_643 | maskExt_643 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA1)
        v0_644 <= v0_644 & ~maskExt_644 | maskExt_644 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA1)
        v0_645 <= v0_645 & ~maskExt_645 | maskExt_645 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA1)
        v0_646 <= v0_646 & ~maskExt_646 | maskExt_646 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA1)
        v0_647 <= v0_647 & ~maskExt_647 | maskExt_647 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA2)
        v0_648 <= v0_648 & ~maskExt_648 | maskExt_648 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA2)
        v0_649 <= v0_649 & ~maskExt_649 | maskExt_649 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA2)
        v0_650 <= v0_650 & ~maskExt_650 | maskExt_650 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA2)
        v0_651 <= v0_651 & ~maskExt_651 | maskExt_651 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA3)
        v0_652 <= v0_652 & ~maskExt_652 | maskExt_652 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA3)
        v0_653 <= v0_653 & ~maskExt_653 | maskExt_653 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA3)
        v0_654 <= v0_654 & ~maskExt_654 | maskExt_654 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA3)
        v0_655 <= v0_655 & ~maskExt_655 | maskExt_655 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA4)
        v0_656 <= v0_656 & ~maskExt_656 | maskExt_656 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA4)
        v0_657 <= v0_657 & ~maskExt_657 | maskExt_657 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA4)
        v0_658 <= v0_658 & ~maskExt_658 | maskExt_658 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA4)
        v0_659 <= v0_659 & ~maskExt_659 | maskExt_659 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA5)
        v0_660 <= v0_660 & ~maskExt_660 | maskExt_660 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA5)
        v0_661 <= v0_661 & ~maskExt_661 | maskExt_661 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA5)
        v0_662 <= v0_662 & ~maskExt_662 | maskExt_662 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA5)
        v0_663 <= v0_663 & ~maskExt_663 | maskExt_663 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA6)
        v0_664 <= v0_664 & ~maskExt_664 | maskExt_664 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA6)
        v0_665 <= v0_665 & ~maskExt_665 | maskExt_665 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA6)
        v0_666 <= v0_666 & ~maskExt_666 | maskExt_666 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA6)
        v0_667 <= v0_667 & ~maskExt_667 | maskExt_667 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA7)
        v0_668 <= v0_668 & ~maskExt_668 | maskExt_668 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA7)
        v0_669 <= v0_669 & ~maskExt_669 | maskExt_669 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA7)
        v0_670 <= v0_670 & ~maskExt_670 | maskExt_670 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA7)
        v0_671 <= v0_671 & ~maskExt_671 | maskExt_671 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA8)
        v0_672 <= v0_672 & ~maskExt_672 | maskExt_672 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA8)
        v0_673 <= v0_673 & ~maskExt_673 | maskExt_673 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA8)
        v0_674 <= v0_674 & ~maskExt_674 | maskExt_674 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA8)
        v0_675 <= v0_675 & ~maskExt_675 | maskExt_675 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hA9)
        v0_676 <= v0_676 & ~maskExt_676 | maskExt_676 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hA9)
        v0_677 <= v0_677 & ~maskExt_677 | maskExt_677 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hA9)
        v0_678 <= v0_678 & ~maskExt_678 | maskExt_678 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hA9)
        v0_679 <= v0_679 & ~maskExt_679 | maskExt_679 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hAA)
        v0_680 <= v0_680 & ~maskExt_680 | maskExt_680 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hAA)
        v0_681 <= v0_681 & ~maskExt_681 | maskExt_681 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hAA)
        v0_682 <= v0_682 & ~maskExt_682 | maskExt_682 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hAA)
        v0_683 <= v0_683 & ~maskExt_683 | maskExt_683 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hAB)
        v0_684 <= v0_684 & ~maskExt_684 | maskExt_684 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hAB)
        v0_685 <= v0_685 & ~maskExt_685 | maskExt_685 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hAB)
        v0_686 <= v0_686 & ~maskExt_686 | maskExt_686 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hAB)
        v0_687 <= v0_687 & ~maskExt_687 | maskExt_687 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hAC)
        v0_688 <= v0_688 & ~maskExt_688 | maskExt_688 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hAC)
        v0_689 <= v0_689 & ~maskExt_689 | maskExt_689 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hAC)
        v0_690 <= v0_690 & ~maskExt_690 | maskExt_690 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hAC)
        v0_691 <= v0_691 & ~maskExt_691 | maskExt_691 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hAD)
        v0_692 <= v0_692 & ~maskExt_692 | maskExt_692 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hAD)
        v0_693 <= v0_693 & ~maskExt_693 | maskExt_693 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hAD)
        v0_694 <= v0_694 & ~maskExt_694 | maskExt_694 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hAD)
        v0_695 <= v0_695 & ~maskExt_695 | maskExt_695 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hAE)
        v0_696 <= v0_696 & ~maskExt_696 | maskExt_696 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hAE)
        v0_697 <= v0_697 & ~maskExt_697 | maskExt_697 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hAE)
        v0_698 <= v0_698 & ~maskExt_698 | maskExt_698 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hAE)
        v0_699 <= v0_699 & ~maskExt_699 | maskExt_699 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hAF)
        v0_700 <= v0_700 & ~maskExt_700 | maskExt_700 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hAF)
        v0_701 <= v0_701 & ~maskExt_701 | maskExt_701 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hAF)
        v0_702 <= v0_702 & ~maskExt_702 | maskExt_702 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hAF)
        v0_703 <= v0_703 & ~maskExt_703 | maskExt_703 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB0)
        v0_704 <= v0_704 & ~maskExt_704 | maskExt_704 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB0)
        v0_705 <= v0_705 & ~maskExt_705 | maskExt_705 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB0)
        v0_706 <= v0_706 & ~maskExt_706 | maskExt_706 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB0)
        v0_707 <= v0_707 & ~maskExt_707 | maskExt_707 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB1)
        v0_708 <= v0_708 & ~maskExt_708 | maskExt_708 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB1)
        v0_709 <= v0_709 & ~maskExt_709 | maskExt_709 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB1)
        v0_710 <= v0_710 & ~maskExt_710 | maskExt_710 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB1)
        v0_711 <= v0_711 & ~maskExt_711 | maskExt_711 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB2)
        v0_712 <= v0_712 & ~maskExt_712 | maskExt_712 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB2)
        v0_713 <= v0_713 & ~maskExt_713 | maskExt_713 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB2)
        v0_714 <= v0_714 & ~maskExt_714 | maskExt_714 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB2)
        v0_715 <= v0_715 & ~maskExt_715 | maskExt_715 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB3)
        v0_716 <= v0_716 & ~maskExt_716 | maskExt_716 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB3)
        v0_717 <= v0_717 & ~maskExt_717 | maskExt_717 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB3)
        v0_718 <= v0_718 & ~maskExt_718 | maskExt_718 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB3)
        v0_719 <= v0_719 & ~maskExt_719 | maskExt_719 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB4)
        v0_720 <= v0_720 & ~maskExt_720 | maskExt_720 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB4)
        v0_721 <= v0_721 & ~maskExt_721 | maskExt_721 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB4)
        v0_722 <= v0_722 & ~maskExt_722 | maskExt_722 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB4)
        v0_723 <= v0_723 & ~maskExt_723 | maskExt_723 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB5)
        v0_724 <= v0_724 & ~maskExt_724 | maskExt_724 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB5)
        v0_725 <= v0_725 & ~maskExt_725 | maskExt_725 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB5)
        v0_726 <= v0_726 & ~maskExt_726 | maskExt_726 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB5)
        v0_727 <= v0_727 & ~maskExt_727 | maskExt_727 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB6)
        v0_728 <= v0_728 & ~maskExt_728 | maskExt_728 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB6)
        v0_729 <= v0_729 & ~maskExt_729 | maskExt_729 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB6)
        v0_730 <= v0_730 & ~maskExt_730 | maskExt_730 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB6)
        v0_731 <= v0_731 & ~maskExt_731 | maskExt_731 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB7)
        v0_732 <= v0_732 & ~maskExt_732 | maskExt_732 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB7)
        v0_733 <= v0_733 & ~maskExt_733 | maskExt_733 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB7)
        v0_734 <= v0_734 & ~maskExt_734 | maskExt_734 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB7)
        v0_735 <= v0_735 & ~maskExt_735 | maskExt_735 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB8)
        v0_736 <= v0_736 & ~maskExt_736 | maskExt_736 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB8)
        v0_737 <= v0_737 & ~maskExt_737 | maskExt_737 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB8)
        v0_738 <= v0_738 & ~maskExt_738 | maskExt_738 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB8)
        v0_739 <= v0_739 & ~maskExt_739 | maskExt_739 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hB9)
        v0_740 <= v0_740 & ~maskExt_740 | maskExt_740 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hB9)
        v0_741 <= v0_741 & ~maskExt_741 | maskExt_741 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hB9)
        v0_742 <= v0_742 & ~maskExt_742 | maskExt_742 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hB9)
        v0_743 <= v0_743 & ~maskExt_743 | maskExt_743 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hBA)
        v0_744 <= v0_744 & ~maskExt_744 | maskExt_744 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hBA)
        v0_745 <= v0_745 & ~maskExt_745 | maskExt_745 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hBA)
        v0_746 <= v0_746 & ~maskExt_746 | maskExt_746 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hBA)
        v0_747 <= v0_747 & ~maskExt_747 | maskExt_747 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hBB)
        v0_748 <= v0_748 & ~maskExt_748 | maskExt_748 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hBB)
        v0_749 <= v0_749 & ~maskExt_749 | maskExt_749 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hBB)
        v0_750 <= v0_750 & ~maskExt_750 | maskExt_750 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hBB)
        v0_751 <= v0_751 & ~maskExt_751 | maskExt_751 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hBC)
        v0_752 <= v0_752 & ~maskExt_752 | maskExt_752 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hBC)
        v0_753 <= v0_753 & ~maskExt_753 | maskExt_753 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hBC)
        v0_754 <= v0_754 & ~maskExt_754 | maskExt_754 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hBC)
        v0_755 <= v0_755 & ~maskExt_755 | maskExt_755 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hBD)
        v0_756 <= v0_756 & ~maskExt_756 | maskExt_756 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hBD)
        v0_757 <= v0_757 & ~maskExt_757 | maskExt_757 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hBD)
        v0_758 <= v0_758 & ~maskExt_758 | maskExt_758 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hBD)
        v0_759 <= v0_759 & ~maskExt_759 | maskExt_759 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hBE)
        v0_760 <= v0_760 & ~maskExt_760 | maskExt_760 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hBE)
        v0_761 <= v0_761 & ~maskExt_761 | maskExt_761 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hBE)
        v0_762 <= v0_762 & ~maskExt_762 | maskExt_762 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hBE)
        v0_763 <= v0_763 & ~maskExt_763 | maskExt_763 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hBF)
        v0_764 <= v0_764 & ~maskExt_764 | maskExt_764 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hBF)
        v0_765 <= v0_765 & ~maskExt_765 | maskExt_765 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hBF)
        v0_766 <= v0_766 & ~maskExt_766 | maskExt_766 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hBF)
        v0_767 <= v0_767 & ~maskExt_767 | maskExt_767 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC0)
        v0_768 <= v0_768 & ~maskExt_768 | maskExt_768 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC0)
        v0_769 <= v0_769 & ~maskExt_769 | maskExt_769 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC0)
        v0_770 <= v0_770 & ~maskExt_770 | maskExt_770 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC0)
        v0_771 <= v0_771 & ~maskExt_771 | maskExt_771 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC1)
        v0_772 <= v0_772 & ~maskExt_772 | maskExt_772 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC1)
        v0_773 <= v0_773 & ~maskExt_773 | maskExt_773 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC1)
        v0_774 <= v0_774 & ~maskExt_774 | maskExt_774 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC1)
        v0_775 <= v0_775 & ~maskExt_775 | maskExt_775 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC2)
        v0_776 <= v0_776 & ~maskExt_776 | maskExt_776 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC2)
        v0_777 <= v0_777 & ~maskExt_777 | maskExt_777 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC2)
        v0_778 <= v0_778 & ~maskExt_778 | maskExt_778 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC2)
        v0_779 <= v0_779 & ~maskExt_779 | maskExt_779 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC3)
        v0_780 <= v0_780 & ~maskExt_780 | maskExt_780 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC3)
        v0_781 <= v0_781 & ~maskExt_781 | maskExt_781 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC3)
        v0_782 <= v0_782 & ~maskExt_782 | maskExt_782 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC3)
        v0_783 <= v0_783 & ~maskExt_783 | maskExt_783 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC4)
        v0_784 <= v0_784 & ~maskExt_784 | maskExt_784 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC4)
        v0_785 <= v0_785 & ~maskExt_785 | maskExt_785 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC4)
        v0_786 <= v0_786 & ~maskExt_786 | maskExt_786 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC4)
        v0_787 <= v0_787 & ~maskExt_787 | maskExt_787 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC5)
        v0_788 <= v0_788 & ~maskExt_788 | maskExt_788 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC5)
        v0_789 <= v0_789 & ~maskExt_789 | maskExt_789 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC5)
        v0_790 <= v0_790 & ~maskExt_790 | maskExt_790 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC5)
        v0_791 <= v0_791 & ~maskExt_791 | maskExt_791 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC6)
        v0_792 <= v0_792 & ~maskExt_792 | maskExt_792 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC6)
        v0_793 <= v0_793 & ~maskExt_793 | maskExt_793 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC6)
        v0_794 <= v0_794 & ~maskExt_794 | maskExt_794 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC6)
        v0_795 <= v0_795 & ~maskExt_795 | maskExt_795 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC7)
        v0_796 <= v0_796 & ~maskExt_796 | maskExt_796 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC7)
        v0_797 <= v0_797 & ~maskExt_797 | maskExt_797 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC7)
        v0_798 <= v0_798 & ~maskExt_798 | maskExt_798 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC7)
        v0_799 <= v0_799 & ~maskExt_799 | maskExt_799 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC8)
        v0_800 <= v0_800 & ~maskExt_800 | maskExt_800 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC8)
        v0_801 <= v0_801 & ~maskExt_801 | maskExt_801 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC8)
        v0_802 <= v0_802 & ~maskExt_802 | maskExt_802 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC8)
        v0_803 <= v0_803 & ~maskExt_803 | maskExt_803 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hC9)
        v0_804 <= v0_804 & ~maskExt_804 | maskExt_804 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hC9)
        v0_805 <= v0_805 & ~maskExt_805 | maskExt_805 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hC9)
        v0_806 <= v0_806 & ~maskExt_806 | maskExt_806 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hC9)
        v0_807 <= v0_807 & ~maskExt_807 | maskExt_807 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hCA)
        v0_808 <= v0_808 & ~maskExt_808 | maskExt_808 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hCA)
        v0_809 <= v0_809 & ~maskExt_809 | maskExt_809 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hCA)
        v0_810 <= v0_810 & ~maskExt_810 | maskExt_810 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hCA)
        v0_811 <= v0_811 & ~maskExt_811 | maskExt_811 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hCB)
        v0_812 <= v0_812 & ~maskExt_812 | maskExt_812 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hCB)
        v0_813 <= v0_813 & ~maskExt_813 | maskExt_813 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hCB)
        v0_814 <= v0_814 & ~maskExt_814 | maskExt_814 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hCB)
        v0_815 <= v0_815 & ~maskExt_815 | maskExt_815 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hCC)
        v0_816 <= v0_816 & ~maskExt_816 | maskExt_816 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hCC)
        v0_817 <= v0_817 & ~maskExt_817 | maskExt_817 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hCC)
        v0_818 <= v0_818 & ~maskExt_818 | maskExt_818 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hCC)
        v0_819 <= v0_819 & ~maskExt_819 | maskExt_819 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hCD)
        v0_820 <= v0_820 & ~maskExt_820 | maskExt_820 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hCD)
        v0_821 <= v0_821 & ~maskExt_821 | maskExt_821 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hCD)
        v0_822 <= v0_822 & ~maskExt_822 | maskExt_822 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hCD)
        v0_823 <= v0_823 & ~maskExt_823 | maskExt_823 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hCE)
        v0_824 <= v0_824 & ~maskExt_824 | maskExt_824 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hCE)
        v0_825 <= v0_825 & ~maskExt_825 | maskExt_825 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hCE)
        v0_826 <= v0_826 & ~maskExt_826 | maskExt_826 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hCE)
        v0_827 <= v0_827 & ~maskExt_827 | maskExt_827 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hCF)
        v0_828 <= v0_828 & ~maskExt_828 | maskExt_828 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hCF)
        v0_829 <= v0_829 & ~maskExt_829 | maskExt_829 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hCF)
        v0_830 <= v0_830 & ~maskExt_830 | maskExt_830 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hCF)
        v0_831 <= v0_831 & ~maskExt_831 | maskExt_831 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD0)
        v0_832 <= v0_832 & ~maskExt_832 | maskExt_832 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD0)
        v0_833 <= v0_833 & ~maskExt_833 | maskExt_833 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD0)
        v0_834 <= v0_834 & ~maskExt_834 | maskExt_834 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD0)
        v0_835 <= v0_835 & ~maskExt_835 | maskExt_835 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD1)
        v0_836 <= v0_836 & ~maskExt_836 | maskExt_836 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD1)
        v0_837 <= v0_837 & ~maskExt_837 | maskExt_837 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD1)
        v0_838 <= v0_838 & ~maskExt_838 | maskExt_838 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD1)
        v0_839 <= v0_839 & ~maskExt_839 | maskExt_839 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD2)
        v0_840 <= v0_840 & ~maskExt_840 | maskExt_840 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD2)
        v0_841 <= v0_841 & ~maskExt_841 | maskExt_841 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD2)
        v0_842 <= v0_842 & ~maskExt_842 | maskExt_842 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD2)
        v0_843 <= v0_843 & ~maskExt_843 | maskExt_843 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD3)
        v0_844 <= v0_844 & ~maskExt_844 | maskExt_844 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD3)
        v0_845 <= v0_845 & ~maskExt_845 | maskExt_845 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD3)
        v0_846 <= v0_846 & ~maskExt_846 | maskExt_846 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD3)
        v0_847 <= v0_847 & ~maskExt_847 | maskExt_847 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD4)
        v0_848 <= v0_848 & ~maskExt_848 | maskExt_848 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD4)
        v0_849 <= v0_849 & ~maskExt_849 | maskExt_849 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD4)
        v0_850 <= v0_850 & ~maskExt_850 | maskExt_850 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD4)
        v0_851 <= v0_851 & ~maskExt_851 | maskExt_851 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD5)
        v0_852 <= v0_852 & ~maskExt_852 | maskExt_852 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD5)
        v0_853 <= v0_853 & ~maskExt_853 | maskExt_853 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD5)
        v0_854 <= v0_854 & ~maskExt_854 | maskExt_854 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD5)
        v0_855 <= v0_855 & ~maskExt_855 | maskExt_855 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD6)
        v0_856 <= v0_856 & ~maskExt_856 | maskExt_856 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD6)
        v0_857 <= v0_857 & ~maskExt_857 | maskExt_857 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD6)
        v0_858 <= v0_858 & ~maskExt_858 | maskExt_858 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD6)
        v0_859 <= v0_859 & ~maskExt_859 | maskExt_859 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD7)
        v0_860 <= v0_860 & ~maskExt_860 | maskExt_860 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD7)
        v0_861 <= v0_861 & ~maskExt_861 | maskExt_861 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD7)
        v0_862 <= v0_862 & ~maskExt_862 | maskExt_862 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD7)
        v0_863 <= v0_863 & ~maskExt_863 | maskExt_863 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD8)
        v0_864 <= v0_864 & ~maskExt_864 | maskExt_864 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD8)
        v0_865 <= v0_865 & ~maskExt_865 | maskExt_865 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD8)
        v0_866 <= v0_866 & ~maskExt_866 | maskExt_866 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD8)
        v0_867 <= v0_867 & ~maskExt_867 | maskExt_867 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hD9)
        v0_868 <= v0_868 & ~maskExt_868 | maskExt_868 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hD9)
        v0_869 <= v0_869 & ~maskExt_869 | maskExt_869 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hD9)
        v0_870 <= v0_870 & ~maskExt_870 | maskExt_870 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hD9)
        v0_871 <= v0_871 & ~maskExt_871 | maskExt_871 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hDA)
        v0_872 <= v0_872 & ~maskExt_872 | maskExt_872 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hDA)
        v0_873 <= v0_873 & ~maskExt_873 | maskExt_873 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hDA)
        v0_874 <= v0_874 & ~maskExt_874 | maskExt_874 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hDA)
        v0_875 <= v0_875 & ~maskExt_875 | maskExt_875 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hDB)
        v0_876 <= v0_876 & ~maskExt_876 | maskExt_876 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hDB)
        v0_877 <= v0_877 & ~maskExt_877 | maskExt_877 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hDB)
        v0_878 <= v0_878 & ~maskExt_878 | maskExt_878 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hDB)
        v0_879 <= v0_879 & ~maskExt_879 | maskExt_879 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hDC)
        v0_880 <= v0_880 & ~maskExt_880 | maskExt_880 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hDC)
        v0_881 <= v0_881 & ~maskExt_881 | maskExt_881 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hDC)
        v0_882 <= v0_882 & ~maskExt_882 | maskExt_882 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hDC)
        v0_883 <= v0_883 & ~maskExt_883 | maskExt_883 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hDD)
        v0_884 <= v0_884 & ~maskExt_884 | maskExt_884 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hDD)
        v0_885 <= v0_885 & ~maskExt_885 | maskExt_885 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hDD)
        v0_886 <= v0_886 & ~maskExt_886 | maskExt_886 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hDD)
        v0_887 <= v0_887 & ~maskExt_887 | maskExt_887 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hDE)
        v0_888 <= v0_888 & ~maskExt_888 | maskExt_888 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hDE)
        v0_889 <= v0_889 & ~maskExt_889 | maskExt_889 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hDE)
        v0_890 <= v0_890 & ~maskExt_890 | maskExt_890 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hDE)
        v0_891 <= v0_891 & ~maskExt_891 | maskExt_891 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hDF)
        v0_892 <= v0_892 & ~maskExt_892 | maskExt_892 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hDF)
        v0_893 <= v0_893 & ~maskExt_893 | maskExt_893 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hDF)
        v0_894 <= v0_894 & ~maskExt_894 | maskExt_894 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hDF)
        v0_895 <= v0_895 & ~maskExt_895 | maskExt_895 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE0)
        v0_896 <= v0_896 & ~maskExt_896 | maskExt_896 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE0)
        v0_897 <= v0_897 & ~maskExt_897 | maskExt_897 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE0)
        v0_898 <= v0_898 & ~maskExt_898 | maskExt_898 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE0)
        v0_899 <= v0_899 & ~maskExt_899 | maskExt_899 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE1)
        v0_900 <= v0_900 & ~maskExt_900 | maskExt_900 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE1)
        v0_901 <= v0_901 & ~maskExt_901 | maskExt_901 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE1)
        v0_902 <= v0_902 & ~maskExt_902 | maskExt_902 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE1)
        v0_903 <= v0_903 & ~maskExt_903 | maskExt_903 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE2)
        v0_904 <= v0_904 & ~maskExt_904 | maskExt_904 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE2)
        v0_905 <= v0_905 & ~maskExt_905 | maskExt_905 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE2)
        v0_906 <= v0_906 & ~maskExt_906 | maskExt_906 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE2)
        v0_907 <= v0_907 & ~maskExt_907 | maskExt_907 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE3)
        v0_908 <= v0_908 & ~maskExt_908 | maskExt_908 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE3)
        v0_909 <= v0_909 & ~maskExt_909 | maskExt_909 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE3)
        v0_910 <= v0_910 & ~maskExt_910 | maskExt_910 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE3)
        v0_911 <= v0_911 & ~maskExt_911 | maskExt_911 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE4)
        v0_912 <= v0_912 & ~maskExt_912 | maskExt_912 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE4)
        v0_913 <= v0_913 & ~maskExt_913 | maskExt_913 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE4)
        v0_914 <= v0_914 & ~maskExt_914 | maskExt_914 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE4)
        v0_915 <= v0_915 & ~maskExt_915 | maskExt_915 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE5)
        v0_916 <= v0_916 & ~maskExt_916 | maskExt_916 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE5)
        v0_917 <= v0_917 & ~maskExt_917 | maskExt_917 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE5)
        v0_918 <= v0_918 & ~maskExt_918 | maskExt_918 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE5)
        v0_919 <= v0_919 & ~maskExt_919 | maskExt_919 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE6)
        v0_920 <= v0_920 & ~maskExt_920 | maskExt_920 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE6)
        v0_921 <= v0_921 & ~maskExt_921 | maskExt_921 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE6)
        v0_922 <= v0_922 & ~maskExt_922 | maskExt_922 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE6)
        v0_923 <= v0_923 & ~maskExt_923 | maskExt_923 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE7)
        v0_924 <= v0_924 & ~maskExt_924 | maskExt_924 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE7)
        v0_925 <= v0_925 & ~maskExt_925 | maskExt_925 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE7)
        v0_926 <= v0_926 & ~maskExt_926 | maskExt_926 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE7)
        v0_927 <= v0_927 & ~maskExt_927 | maskExt_927 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE8)
        v0_928 <= v0_928 & ~maskExt_928 | maskExt_928 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE8)
        v0_929 <= v0_929 & ~maskExt_929 | maskExt_929 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE8)
        v0_930 <= v0_930 & ~maskExt_930 | maskExt_930 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE8)
        v0_931 <= v0_931 & ~maskExt_931 | maskExt_931 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hE9)
        v0_932 <= v0_932 & ~maskExt_932 | maskExt_932 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hE9)
        v0_933 <= v0_933 & ~maskExt_933 | maskExt_933 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hE9)
        v0_934 <= v0_934 & ~maskExt_934 | maskExt_934 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hE9)
        v0_935 <= v0_935 & ~maskExt_935 | maskExt_935 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hEA)
        v0_936 <= v0_936 & ~maskExt_936 | maskExt_936 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hEA)
        v0_937 <= v0_937 & ~maskExt_937 | maskExt_937 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hEA)
        v0_938 <= v0_938 & ~maskExt_938 | maskExt_938 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hEA)
        v0_939 <= v0_939 & ~maskExt_939 | maskExt_939 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hEB)
        v0_940 <= v0_940 & ~maskExt_940 | maskExt_940 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hEB)
        v0_941 <= v0_941 & ~maskExt_941 | maskExt_941 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hEB)
        v0_942 <= v0_942 & ~maskExt_942 | maskExt_942 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hEB)
        v0_943 <= v0_943 & ~maskExt_943 | maskExt_943 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hEC)
        v0_944 <= v0_944 & ~maskExt_944 | maskExt_944 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hEC)
        v0_945 <= v0_945 & ~maskExt_945 | maskExt_945 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hEC)
        v0_946 <= v0_946 & ~maskExt_946 | maskExt_946 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hEC)
        v0_947 <= v0_947 & ~maskExt_947 | maskExt_947 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hED)
        v0_948 <= v0_948 & ~maskExt_948 | maskExt_948 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hED)
        v0_949 <= v0_949 & ~maskExt_949 | maskExt_949 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hED)
        v0_950 <= v0_950 & ~maskExt_950 | maskExt_950 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hED)
        v0_951 <= v0_951 & ~maskExt_951 | maskExt_951 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hEE)
        v0_952 <= v0_952 & ~maskExt_952 | maskExt_952 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hEE)
        v0_953 <= v0_953 & ~maskExt_953 | maskExt_953 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hEE)
        v0_954 <= v0_954 & ~maskExt_954 | maskExt_954 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hEE)
        v0_955 <= v0_955 & ~maskExt_955 | maskExt_955 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hEF)
        v0_956 <= v0_956 & ~maskExt_956 | maskExt_956 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hEF)
        v0_957 <= v0_957 & ~maskExt_957 | maskExt_957 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hEF)
        v0_958 <= v0_958 & ~maskExt_958 | maskExt_958 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hEF)
        v0_959 <= v0_959 & ~maskExt_959 | maskExt_959 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF0)
        v0_960 <= v0_960 & ~maskExt_960 | maskExt_960 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF0)
        v0_961 <= v0_961 & ~maskExt_961 | maskExt_961 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF0)
        v0_962 <= v0_962 & ~maskExt_962 | maskExt_962 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF0)
        v0_963 <= v0_963 & ~maskExt_963 | maskExt_963 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF1)
        v0_964 <= v0_964 & ~maskExt_964 | maskExt_964 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF1)
        v0_965 <= v0_965 & ~maskExt_965 | maskExt_965 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF1)
        v0_966 <= v0_966 & ~maskExt_966 | maskExt_966 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF1)
        v0_967 <= v0_967 & ~maskExt_967 | maskExt_967 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF2)
        v0_968 <= v0_968 & ~maskExt_968 | maskExt_968 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF2)
        v0_969 <= v0_969 & ~maskExt_969 | maskExt_969 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF2)
        v0_970 <= v0_970 & ~maskExt_970 | maskExt_970 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF2)
        v0_971 <= v0_971 & ~maskExt_971 | maskExt_971 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF3)
        v0_972 <= v0_972 & ~maskExt_972 | maskExt_972 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF3)
        v0_973 <= v0_973 & ~maskExt_973 | maskExt_973 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF3)
        v0_974 <= v0_974 & ~maskExt_974 | maskExt_974 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF3)
        v0_975 <= v0_975 & ~maskExt_975 | maskExt_975 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF4)
        v0_976 <= v0_976 & ~maskExt_976 | maskExt_976 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF4)
        v0_977 <= v0_977 & ~maskExt_977 | maskExt_977 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF4)
        v0_978 <= v0_978 & ~maskExt_978 | maskExt_978 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF4)
        v0_979 <= v0_979 & ~maskExt_979 | maskExt_979 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF5)
        v0_980 <= v0_980 & ~maskExt_980 | maskExt_980 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF5)
        v0_981 <= v0_981 & ~maskExt_981 | maskExt_981 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF5)
        v0_982 <= v0_982 & ~maskExt_982 | maskExt_982 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF5)
        v0_983 <= v0_983 & ~maskExt_983 | maskExt_983 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF6)
        v0_984 <= v0_984 & ~maskExt_984 | maskExt_984 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF6)
        v0_985 <= v0_985 & ~maskExt_985 | maskExt_985 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF6)
        v0_986 <= v0_986 & ~maskExt_986 | maskExt_986 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF6)
        v0_987 <= v0_987 & ~maskExt_987 | maskExt_987 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF7)
        v0_988 <= v0_988 & ~maskExt_988 | maskExt_988 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF7)
        v0_989 <= v0_989 & ~maskExt_989 | maskExt_989 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF7)
        v0_990 <= v0_990 & ~maskExt_990 | maskExt_990 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF7)
        v0_991 <= v0_991 & ~maskExt_991 | maskExt_991 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF8)
        v0_992 <= v0_992 & ~maskExt_992 | maskExt_992 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF8)
        v0_993 <= v0_993 & ~maskExt_993 | maskExt_993 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF8)
        v0_994 <= v0_994 & ~maskExt_994 | maskExt_994 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF8)
        v0_995 <= v0_995 & ~maskExt_995 | maskExt_995 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hF9)
        v0_996 <= v0_996 & ~maskExt_996 | maskExt_996 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hF9)
        v0_997 <= v0_997 & ~maskExt_997 | maskExt_997 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hF9)
        v0_998 <= v0_998 & ~maskExt_998 | maskExt_998 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hF9)
        v0_999 <= v0_999 & ~maskExt_999 | maskExt_999 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hFA)
        v0_1000 <= v0_1000 & ~maskExt_1000 | maskExt_1000 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hFA)
        v0_1001 <= v0_1001 & ~maskExt_1001 | maskExt_1001 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hFA)
        v0_1002 <= v0_1002 & ~maskExt_1002 | maskExt_1002 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hFA)
        v0_1003 <= v0_1003 & ~maskExt_1003 | maskExt_1003 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hFB)
        v0_1004 <= v0_1004 & ~maskExt_1004 | maskExt_1004 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hFB)
        v0_1005 <= v0_1005 & ~maskExt_1005 | maskExt_1005 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hFB)
        v0_1006 <= v0_1006 & ~maskExt_1006 | maskExt_1006 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hFB)
        v0_1007 <= v0_1007 & ~maskExt_1007 | maskExt_1007 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hFC)
        v0_1008 <= v0_1008 & ~maskExt_1008 | maskExt_1008 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hFC)
        v0_1009 <= v0_1009 & ~maskExt_1009 | maskExt_1009 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hFC)
        v0_1010 <= v0_1010 & ~maskExt_1010 | maskExt_1010 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hFC)
        v0_1011 <= v0_1011 & ~maskExt_1011 | maskExt_1011 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hFD)
        v0_1012 <= v0_1012 & ~maskExt_1012 | maskExt_1012 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hFD)
        v0_1013 <= v0_1013 & ~maskExt_1013 | maskExt_1013 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hFD)
        v0_1014 <= v0_1014 & ~maskExt_1014 | maskExt_1014 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hFD)
        v0_1015 <= v0_1015 & ~maskExt_1015 | maskExt_1015 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 8'hFE)
        v0_1016 <= v0_1016 & ~maskExt_1016 | maskExt_1016 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 8'hFE)
        v0_1017 <= v0_1017 & ~maskExt_1017 | maskExt_1017 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 8'hFE)
        v0_1018 <= v0_1018 & ~maskExt_1018 | maskExt_1018 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 8'hFE)
        v0_1019 <= v0_1019 & ~maskExt_1019 | maskExt_1019 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & (&v0UpdateVec_0_bits_offset))
        v0_1020 <= v0_1020 & ~maskExt_1020 | maskExt_1020 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & (&v0UpdateVec_1_bits_offset))
        v0_1021 <= v0_1021 & ~maskExt_1021 | maskExt_1021 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & (&v0UpdateVec_2_bits_offset))
        v0_1022 <= v0_1022 & ~maskExt_1022 | maskExt_1022 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & (&v0UpdateVec_3_bits_offset))
        v0_1023 <= v0_1023 & ~maskExt_1023 | maskExt_1023 & v0UpdateVec_3_bits_data;
      if (queueEnq[0] ^ queueDeq[0])
        queueCount_0 <= queueCount_0 + counterUpdate;
      if (queueEnq[1] ^ queueDeq[1])
        queueCount_1 <= queueCount_1 + counterUpdate_1;
      if (queueEnq[2] ^ queueDeq[2])
        queueCount_2 <= queueCount_2 + counterUpdate_2;
      if (queueEnq[3] ^ queueDeq[3])
        queueCount_3 <= queueCount_3 + counterUpdate_3;
      if (queueEnq[4] ^ queueDeq[4])
        queueCount_4 <= queueCount_4 + counterUpdate_4;
      if (queueEnq[5] ^ queueDeq[5])
        queueCount_5 <= queueCount_5 + counterUpdate_5;
      if (queueEnq[6] ^ queueDeq[6])
        queueCount_6 <= queueCount_6 + counterUpdate_6;
      if (queueEnq[7] ^ queueDeq[7])
        queueCount_7 <= queueCount_7 + counterUpdate_7;
      if (queueEnq_1[0] ^ queueDeq_1[0])
        queueCount_0_1 <= queueCount_0_1 + counterUpdate_8;
      if (queueEnq_1[1] ^ queueDeq_1[1])
        queueCount_1_1 <= queueCount_1_1 + counterUpdate_9;
      if (queueEnq_1[2] ^ queueDeq_1[2])
        queueCount_2_1 <= queueCount_2_1 + counterUpdate_10;
      if (queueEnq_1[3] ^ queueDeq_1[3])
        queueCount_3_1 <= queueCount_3_1 + counterUpdate_11;
      if (queueEnq_1[4] ^ queueDeq_1[4])
        queueCount_4_1 <= queueCount_4_1 + counterUpdate_12;
      if (queueEnq_1[5] ^ queueDeq_1[5])
        queueCount_5_1 <= queueCount_5_1 + counterUpdate_13;
      if (queueEnq_1[6] ^ queueDeq_1[6])
        queueCount_6_1 <= queueCount_6_1 + counterUpdate_14;
      if (queueEnq_1[7] ^ queueDeq_1[7])
        queueCount_7_1 <= queueCount_7_1 + counterUpdate_15;
      if (queueEnq_2[0] ^ queueDeq_2[0])
        queueCount_0_2 <= queueCount_0_2 + counterUpdate_16;
      if (queueEnq_2[1] ^ queueDeq_2[1])
        queueCount_1_2 <= queueCount_1_2 + counterUpdate_17;
      if (queueEnq_2[2] ^ queueDeq_2[2])
        queueCount_2_2 <= queueCount_2_2 + counterUpdate_18;
      if (queueEnq_2[3] ^ queueDeq_2[3])
        queueCount_3_2 <= queueCount_3_2 + counterUpdate_19;
      if (queueEnq_2[4] ^ queueDeq_2[4])
        queueCount_4_2 <= queueCount_4_2 + counterUpdate_20;
      if (queueEnq_2[5] ^ queueDeq_2[5])
        queueCount_5_2 <= queueCount_5_2 + counterUpdate_21;
      if (queueEnq_2[6] ^ queueDeq_2[6])
        queueCount_6_2 <= queueCount_6_2 + counterUpdate_22;
      if (queueEnq_2[7] ^ queueDeq_2[7])
        queueCount_7_2 <= queueCount_7_2 + counterUpdate_23;
      if (queueEnq_3[0] ^ queueDeq_3[0])
        queueCount_0_3 <= queueCount_0_3 + counterUpdate_24;
      if (queueEnq_3[1] ^ queueDeq_3[1])
        queueCount_1_3 <= queueCount_1_3 + counterUpdate_25;
      if (queueEnq_3[2] ^ queueDeq_3[2])
        queueCount_2_3 <= queueCount_2_3 + counterUpdate_26;
      if (queueEnq_3[3] ^ queueDeq_3[3])
        queueCount_3_3 <= queueCount_3_3 + counterUpdate_27;
      if (queueEnq_3[4] ^ queueDeq_3[4])
        queueCount_4_3 <= queueCount_4_3 + counterUpdate_28;
      if (queueEnq_3[5] ^ queueDeq_3[5])
        queueCount_5_3 <= queueCount_5_3 + counterUpdate_29;
      if (queueEnq_3[6] ^ queueDeq_3[6])
        queueCount_6_3 <= queueCount_6_3 + counterUpdate_30;
      if (queueEnq_3[7] ^ queueDeq_3[7])
        queueCount_7_3 <= queueCount_7_3 + counterUpdate_31;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:1030];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [10:0] i = 11'h0; i < 11'h407; i += 11'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[11'h0];
        v0_1 = _RANDOM[11'h1];
        v0_2 = _RANDOM[11'h2];
        v0_3 = _RANDOM[11'h3];
        v0_4 = _RANDOM[11'h4];
        v0_5 = _RANDOM[11'h5];
        v0_6 = _RANDOM[11'h6];
        v0_7 = _RANDOM[11'h7];
        v0_8 = _RANDOM[11'h8];
        v0_9 = _RANDOM[11'h9];
        v0_10 = _RANDOM[11'hA];
        v0_11 = _RANDOM[11'hB];
        v0_12 = _RANDOM[11'hC];
        v0_13 = _RANDOM[11'hD];
        v0_14 = _RANDOM[11'hE];
        v0_15 = _RANDOM[11'hF];
        v0_16 = _RANDOM[11'h10];
        v0_17 = _RANDOM[11'h11];
        v0_18 = _RANDOM[11'h12];
        v0_19 = _RANDOM[11'h13];
        v0_20 = _RANDOM[11'h14];
        v0_21 = _RANDOM[11'h15];
        v0_22 = _RANDOM[11'h16];
        v0_23 = _RANDOM[11'h17];
        v0_24 = _RANDOM[11'h18];
        v0_25 = _RANDOM[11'h19];
        v0_26 = _RANDOM[11'h1A];
        v0_27 = _RANDOM[11'h1B];
        v0_28 = _RANDOM[11'h1C];
        v0_29 = _RANDOM[11'h1D];
        v0_30 = _RANDOM[11'h1E];
        v0_31 = _RANDOM[11'h1F];
        v0_32 = _RANDOM[11'h20];
        v0_33 = _RANDOM[11'h21];
        v0_34 = _RANDOM[11'h22];
        v0_35 = _RANDOM[11'h23];
        v0_36 = _RANDOM[11'h24];
        v0_37 = _RANDOM[11'h25];
        v0_38 = _RANDOM[11'h26];
        v0_39 = _RANDOM[11'h27];
        v0_40 = _RANDOM[11'h28];
        v0_41 = _RANDOM[11'h29];
        v0_42 = _RANDOM[11'h2A];
        v0_43 = _RANDOM[11'h2B];
        v0_44 = _RANDOM[11'h2C];
        v0_45 = _RANDOM[11'h2D];
        v0_46 = _RANDOM[11'h2E];
        v0_47 = _RANDOM[11'h2F];
        v0_48 = _RANDOM[11'h30];
        v0_49 = _RANDOM[11'h31];
        v0_50 = _RANDOM[11'h32];
        v0_51 = _RANDOM[11'h33];
        v0_52 = _RANDOM[11'h34];
        v0_53 = _RANDOM[11'h35];
        v0_54 = _RANDOM[11'h36];
        v0_55 = _RANDOM[11'h37];
        v0_56 = _RANDOM[11'h38];
        v0_57 = _RANDOM[11'h39];
        v0_58 = _RANDOM[11'h3A];
        v0_59 = _RANDOM[11'h3B];
        v0_60 = _RANDOM[11'h3C];
        v0_61 = _RANDOM[11'h3D];
        v0_62 = _RANDOM[11'h3E];
        v0_63 = _RANDOM[11'h3F];
        v0_64 = _RANDOM[11'h40];
        v0_65 = _RANDOM[11'h41];
        v0_66 = _RANDOM[11'h42];
        v0_67 = _RANDOM[11'h43];
        v0_68 = _RANDOM[11'h44];
        v0_69 = _RANDOM[11'h45];
        v0_70 = _RANDOM[11'h46];
        v0_71 = _RANDOM[11'h47];
        v0_72 = _RANDOM[11'h48];
        v0_73 = _RANDOM[11'h49];
        v0_74 = _RANDOM[11'h4A];
        v0_75 = _RANDOM[11'h4B];
        v0_76 = _RANDOM[11'h4C];
        v0_77 = _RANDOM[11'h4D];
        v0_78 = _RANDOM[11'h4E];
        v0_79 = _RANDOM[11'h4F];
        v0_80 = _RANDOM[11'h50];
        v0_81 = _RANDOM[11'h51];
        v0_82 = _RANDOM[11'h52];
        v0_83 = _RANDOM[11'h53];
        v0_84 = _RANDOM[11'h54];
        v0_85 = _RANDOM[11'h55];
        v0_86 = _RANDOM[11'h56];
        v0_87 = _RANDOM[11'h57];
        v0_88 = _RANDOM[11'h58];
        v0_89 = _RANDOM[11'h59];
        v0_90 = _RANDOM[11'h5A];
        v0_91 = _RANDOM[11'h5B];
        v0_92 = _RANDOM[11'h5C];
        v0_93 = _RANDOM[11'h5D];
        v0_94 = _RANDOM[11'h5E];
        v0_95 = _RANDOM[11'h5F];
        v0_96 = _RANDOM[11'h60];
        v0_97 = _RANDOM[11'h61];
        v0_98 = _RANDOM[11'h62];
        v0_99 = _RANDOM[11'h63];
        v0_100 = _RANDOM[11'h64];
        v0_101 = _RANDOM[11'h65];
        v0_102 = _RANDOM[11'h66];
        v0_103 = _RANDOM[11'h67];
        v0_104 = _RANDOM[11'h68];
        v0_105 = _RANDOM[11'h69];
        v0_106 = _RANDOM[11'h6A];
        v0_107 = _RANDOM[11'h6B];
        v0_108 = _RANDOM[11'h6C];
        v0_109 = _RANDOM[11'h6D];
        v0_110 = _RANDOM[11'h6E];
        v0_111 = _RANDOM[11'h6F];
        v0_112 = _RANDOM[11'h70];
        v0_113 = _RANDOM[11'h71];
        v0_114 = _RANDOM[11'h72];
        v0_115 = _RANDOM[11'h73];
        v0_116 = _RANDOM[11'h74];
        v0_117 = _RANDOM[11'h75];
        v0_118 = _RANDOM[11'h76];
        v0_119 = _RANDOM[11'h77];
        v0_120 = _RANDOM[11'h78];
        v0_121 = _RANDOM[11'h79];
        v0_122 = _RANDOM[11'h7A];
        v0_123 = _RANDOM[11'h7B];
        v0_124 = _RANDOM[11'h7C];
        v0_125 = _RANDOM[11'h7D];
        v0_126 = _RANDOM[11'h7E];
        v0_127 = _RANDOM[11'h7F];
        v0_128 = _RANDOM[11'h80];
        v0_129 = _RANDOM[11'h81];
        v0_130 = _RANDOM[11'h82];
        v0_131 = _RANDOM[11'h83];
        v0_132 = _RANDOM[11'h84];
        v0_133 = _RANDOM[11'h85];
        v0_134 = _RANDOM[11'h86];
        v0_135 = _RANDOM[11'h87];
        v0_136 = _RANDOM[11'h88];
        v0_137 = _RANDOM[11'h89];
        v0_138 = _RANDOM[11'h8A];
        v0_139 = _RANDOM[11'h8B];
        v0_140 = _RANDOM[11'h8C];
        v0_141 = _RANDOM[11'h8D];
        v0_142 = _RANDOM[11'h8E];
        v0_143 = _RANDOM[11'h8F];
        v0_144 = _RANDOM[11'h90];
        v0_145 = _RANDOM[11'h91];
        v0_146 = _RANDOM[11'h92];
        v0_147 = _RANDOM[11'h93];
        v0_148 = _RANDOM[11'h94];
        v0_149 = _RANDOM[11'h95];
        v0_150 = _RANDOM[11'h96];
        v0_151 = _RANDOM[11'h97];
        v0_152 = _RANDOM[11'h98];
        v0_153 = _RANDOM[11'h99];
        v0_154 = _RANDOM[11'h9A];
        v0_155 = _RANDOM[11'h9B];
        v0_156 = _RANDOM[11'h9C];
        v0_157 = _RANDOM[11'h9D];
        v0_158 = _RANDOM[11'h9E];
        v0_159 = _RANDOM[11'h9F];
        v0_160 = _RANDOM[11'hA0];
        v0_161 = _RANDOM[11'hA1];
        v0_162 = _RANDOM[11'hA2];
        v0_163 = _RANDOM[11'hA3];
        v0_164 = _RANDOM[11'hA4];
        v0_165 = _RANDOM[11'hA5];
        v0_166 = _RANDOM[11'hA6];
        v0_167 = _RANDOM[11'hA7];
        v0_168 = _RANDOM[11'hA8];
        v0_169 = _RANDOM[11'hA9];
        v0_170 = _RANDOM[11'hAA];
        v0_171 = _RANDOM[11'hAB];
        v0_172 = _RANDOM[11'hAC];
        v0_173 = _RANDOM[11'hAD];
        v0_174 = _RANDOM[11'hAE];
        v0_175 = _RANDOM[11'hAF];
        v0_176 = _RANDOM[11'hB0];
        v0_177 = _RANDOM[11'hB1];
        v0_178 = _RANDOM[11'hB2];
        v0_179 = _RANDOM[11'hB3];
        v0_180 = _RANDOM[11'hB4];
        v0_181 = _RANDOM[11'hB5];
        v0_182 = _RANDOM[11'hB6];
        v0_183 = _RANDOM[11'hB7];
        v0_184 = _RANDOM[11'hB8];
        v0_185 = _RANDOM[11'hB9];
        v0_186 = _RANDOM[11'hBA];
        v0_187 = _RANDOM[11'hBB];
        v0_188 = _RANDOM[11'hBC];
        v0_189 = _RANDOM[11'hBD];
        v0_190 = _RANDOM[11'hBE];
        v0_191 = _RANDOM[11'hBF];
        v0_192 = _RANDOM[11'hC0];
        v0_193 = _RANDOM[11'hC1];
        v0_194 = _RANDOM[11'hC2];
        v0_195 = _RANDOM[11'hC3];
        v0_196 = _RANDOM[11'hC4];
        v0_197 = _RANDOM[11'hC5];
        v0_198 = _RANDOM[11'hC6];
        v0_199 = _RANDOM[11'hC7];
        v0_200 = _RANDOM[11'hC8];
        v0_201 = _RANDOM[11'hC9];
        v0_202 = _RANDOM[11'hCA];
        v0_203 = _RANDOM[11'hCB];
        v0_204 = _RANDOM[11'hCC];
        v0_205 = _RANDOM[11'hCD];
        v0_206 = _RANDOM[11'hCE];
        v0_207 = _RANDOM[11'hCF];
        v0_208 = _RANDOM[11'hD0];
        v0_209 = _RANDOM[11'hD1];
        v0_210 = _RANDOM[11'hD2];
        v0_211 = _RANDOM[11'hD3];
        v0_212 = _RANDOM[11'hD4];
        v0_213 = _RANDOM[11'hD5];
        v0_214 = _RANDOM[11'hD6];
        v0_215 = _RANDOM[11'hD7];
        v0_216 = _RANDOM[11'hD8];
        v0_217 = _RANDOM[11'hD9];
        v0_218 = _RANDOM[11'hDA];
        v0_219 = _RANDOM[11'hDB];
        v0_220 = _RANDOM[11'hDC];
        v0_221 = _RANDOM[11'hDD];
        v0_222 = _RANDOM[11'hDE];
        v0_223 = _RANDOM[11'hDF];
        v0_224 = _RANDOM[11'hE0];
        v0_225 = _RANDOM[11'hE1];
        v0_226 = _RANDOM[11'hE2];
        v0_227 = _RANDOM[11'hE3];
        v0_228 = _RANDOM[11'hE4];
        v0_229 = _RANDOM[11'hE5];
        v0_230 = _RANDOM[11'hE6];
        v0_231 = _RANDOM[11'hE7];
        v0_232 = _RANDOM[11'hE8];
        v0_233 = _RANDOM[11'hE9];
        v0_234 = _RANDOM[11'hEA];
        v0_235 = _RANDOM[11'hEB];
        v0_236 = _RANDOM[11'hEC];
        v0_237 = _RANDOM[11'hED];
        v0_238 = _RANDOM[11'hEE];
        v0_239 = _RANDOM[11'hEF];
        v0_240 = _RANDOM[11'hF0];
        v0_241 = _RANDOM[11'hF1];
        v0_242 = _RANDOM[11'hF2];
        v0_243 = _RANDOM[11'hF3];
        v0_244 = _RANDOM[11'hF4];
        v0_245 = _RANDOM[11'hF5];
        v0_246 = _RANDOM[11'hF6];
        v0_247 = _RANDOM[11'hF7];
        v0_248 = _RANDOM[11'hF8];
        v0_249 = _RANDOM[11'hF9];
        v0_250 = _RANDOM[11'hFA];
        v0_251 = _RANDOM[11'hFB];
        v0_252 = _RANDOM[11'hFC];
        v0_253 = _RANDOM[11'hFD];
        v0_254 = _RANDOM[11'hFE];
        v0_255 = _RANDOM[11'hFF];
        v0_256 = _RANDOM[11'h100];
        v0_257 = _RANDOM[11'h101];
        v0_258 = _RANDOM[11'h102];
        v0_259 = _RANDOM[11'h103];
        v0_260 = _RANDOM[11'h104];
        v0_261 = _RANDOM[11'h105];
        v0_262 = _RANDOM[11'h106];
        v0_263 = _RANDOM[11'h107];
        v0_264 = _RANDOM[11'h108];
        v0_265 = _RANDOM[11'h109];
        v0_266 = _RANDOM[11'h10A];
        v0_267 = _RANDOM[11'h10B];
        v0_268 = _RANDOM[11'h10C];
        v0_269 = _RANDOM[11'h10D];
        v0_270 = _RANDOM[11'h10E];
        v0_271 = _RANDOM[11'h10F];
        v0_272 = _RANDOM[11'h110];
        v0_273 = _RANDOM[11'h111];
        v0_274 = _RANDOM[11'h112];
        v0_275 = _RANDOM[11'h113];
        v0_276 = _RANDOM[11'h114];
        v0_277 = _RANDOM[11'h115];
        v0_278 = _RANDOM[11'h116];
        v0_279 = _RANDOM[11'h117];
        v0_280 = _RANDOM[11'h118];
        v0_281 = _RANDOM[11'h119];
        v0_282 = _RANDOM[11'h11A];
        v0_283 = _RANDOM[11'h11B];
        v0_284 = _RANDOM[11'h11C];
        v0_285 = _RANDOM[11'h11D];
        v0_286 = _RANDOM[11'h11E];
        v0_287 = _RANDOM[11'h11F];
        v0_288 = _RANDOM[11'h120];
        v0_289 = _RANDOM[11'h121];
        v0_290 = _RANDOM[11'h122];
        v0_291 = _RANDOM[11'h123];
        v0_292 = _RANDOM[11'h124];
        v0_293 = _RANDOM[11'h125];
        v0_294 = _RANDOM[11'h126];
        v0_295 = _RANDOM[11'h127];
        v0_296 = _RANDOM[11'h128];
        v0_297 = _RANDOM[11'h129];
        v0_298 = _RANDOM[11'h12A];
        v0_299 = _RANDOM[11'h12B];
        v0_300 = _RANDOM[11'h12C];
        v0_301 = _RANDOM[11'h12D];
        v0_302 = _RANDOM[11'h12E];
        v0_303 = _RANDOM[11'h12F];
        v0_304 = _RANDOM[11'h130];
        v0_305 = _RANDOM[11'h131];
        v0_306 = _RANDOM[11'h132];
        v0_307 = _RANDOM[11'h133];
        v0_308 = _RANDOM[11'h134];
        v0_309 = _RANDOM[11'h135];
        v0_310 = _RANDOM[11'h136];
        v0_311 = _RANDOM[11'h137];
        v0_312 = _RANDOM[11'h138];
        v0_313 = _RANDOM[11'h139];
        v0_314 = _RANDOM[11'h13A];
        v0_315 = _RANDOM[11'h13B];
        v0_316 = _RANDOM[11'h13C];
        v0_317 = _RANDOM[11'h13D];
        v0_318 = _RANDOM[11'h13E];
        v0_319 = _RANDOM[11'h13F];
        v0_320 = _RANDOM[11'h140];
        v0_321 = _RANDOM[11'h141];
        v0_322 = _RANDOM[11'h142];
        v0_323 = _RANDOM[11'h143];
        v0_324 = _RANDOM[11'h144];
        v0_325 = _RANDOM[11'h145];
        v0_326 = _RANDOM[11'h146];
        v0_327 = _RANDOM[11'h147];
        v0_328 = _RANDOM[11'h148];
        v0_329 = _RANDOM[11'h149];
        v0_330 = _RANDOM[11'h14A];
        v0_331 = _RANDOM[11'h14B];
        v0_332 = _RANDOM[11'h14C];
        v0_333 = _RANDOM[11'h14D];
        v0_334 = _RANDOM[11'h14E];
        v0_335 = _RANDOM[11'h14F];
        v0_336 = _RANDOM[11'h150];
        v0_337 = _RANDOM[11'h151];
        v0_338 = _RANDOM[11'h152];
        v0_339 = _RANDOM[11'h153];
        v0_340 = _RANDOM[11'h154];
        v0_341 = _RANDOM[11'h155];
        v0_342 = _RANDOM[11'h156];
        v0_343 = _RANDOM[11'h157];
        v0_344 = _RANDOM[11'h158];
        v0_345 = _RANDOM[11'h159];
        v0_346 = _RANDOM[11'h15A];
        v0_347 = _RANDOM[11'h15B];
        v0_348 = _RANDOM[11'h15C];
        v0_349 = _RANDOM[11'h15D];
        v0_350 = _RANDOM[11'h15E];
        v0_351 = _RANDOM[11'h15F];
        v0_352 = _RANDOM[11'h160];
        v0_353 = _RANDOM[11'h161];
        v0_354 = _RANDOM[11'h162];
        v0_355 = _RANDOM[11'h163];
        v0_356 = _RANDOM[11'h164];
        v0_357 = _RANDOM[11'h165];
        v0_358 = _RANDOM[11'h166];
        v0_359 = _RANDOM[11'h167];
        v0_360 = _RANDOM[11'h168];
        v0_361 = _RANDOM[11'h169];
        v0_362 = _RANDOM[11'h16A];
        v0_363 = _RANDOM[11'h16B];
        v0_364 = _RANDOM[11'h16C];
        v0_365 = _RANDOM[11'h16D];
        v0_366 = _RANDOM[11'h16E];
        v0_367 = _RANDOM[11'h16F];
        v0_368 = _RANDOM[11'h170];
        v0_369 = _RANDOM[11'h171];
        v0_370 = _RANDOM[11'h172];
        v0_371 = _RANDOM[11'h173];
        v0_372 = _RANDOM[11'h174];
        v0_373 = _RANDOM[11'h175];
        v0_374 = _RANDOM[11'h176];
        v0_375 = _RANDOM[11'h177];
        v0_376 = _RANDOM[11'h178];
        v0_377 = _RANDOM[11'h179];
        v0_378 = _RANDOM[11'h17A];
        v0_379 = _RANDOM[11'h17B];
        v0_380 = _RANDOM[11'h17C];
        v0_381 = _RANDOM[11'h17D];
        v0_382 = _RANDOM[11'h17E];
        v0_383 = _RANDOM[11'h17F];
        v0_384 = _RANDOM[11'h180];
        v0_385 = _RANDOM[11'h181];
        v0_386 = _RANDOM[11'h182];
        v0_387 = _RANDOM[11'h183];
        v0_388 = _RANDOM[11'h184];
        v0_389 = _RANDOM[11'h185];
        v0_390 = _RANDOM[11'h186];
        v0_391 = _RANDOM[11'h187];
        v0_392 = _RANDOM[11'h188];
        v0_393 = _RANDOM[11'h189];
        v0_394 = _RANDOM[11'h18A];
        v0_395 = _RANDOM[11'h18B];
        v0_396 = _RANDOM[11'h18C];
        v0_397 = _RANDOM[11'h18D];
        v0_398 = _RANDOM[11'h18E];
        v0_399 = _RANDOM[11'h18F];
        v0_400 = _RANDOM[11'h190];
        v0_401 = _RANDOM[11'h191];
        v0_402 = _RANDOM[11'h192];
        v0_403 = _RANDOM[11'h193];
        v0_404 = _RANDOM[11'h194];
        v0_405 = _RANDOM[11'h195];
        v0_406 = _RANDOM[11'h196];
        v0_407 = _RANDOM[11'h197];
        v0_408 = _RANDOM[11'h198];
        v0_409 = _RANDOM[11'h199];
        v0_410 = _RANDOM[11'h19A];
        v0_411 = _RANDOM[11'h19B];
        v0_412 = _RANDOM[11'h19C];
        v0_413 = _RANDOM[11'h19D];
        v0_414 = _RANDOM[11'h19E];
        v0_415 = _RANDOM[11'h19F];
        v0_416 = _RANDOM[11'h1A0];
        v0_417 = _RANDOM[11'h1A1];
        v0_418 = _RANDOM[11'h1A2];
        v0_419 = _RANDOM[11'h1A3];
        v0_420 = _RANDOM[11'h1A4];
        v0_421 = _RANDOM[11'h1A5];
        v0_422 = _RANDOM[11'h1A6];
        v0_423 = _RANDOM[11'h1A7];
        v0_424 = _RANDOM[11'h1A8];
        v0_425 = _RANDOM[11'h1A9];
        v0_426 = _RANDOM[11'h1AA];
        v0_427 = _RANDOM[11'h1AB];
        v0_428 = _RANDOM[11'h1AC];
        v0_429 = _RANDOM[11'h1AD];
        v0_430 = _RANDOM[11'h1AE];
        v0_431 = _RANDOM[11'h1AF];
        v0_432 = _RANDOM[11'h1B0];
        v0_433 = _RANDOM[11'h1B1];
        v0_434 = _RANDOM[11'h1B2];
        v0_435 = _RANDOM[11'h1B3];
        v0_436 = _RANDOM[11'h1B4];
        v0_437 = _RANDOM[11'h1B5];
        v0_438 = _RANDOM[11'h1B6];
        v0_439 = _RANDOM[11'h1B7];
        v0_440 = _RANDOM[11'h1B8];
        v0_441 = _RANDOM[11'h1B9];
        v0_442 = _RANDOM[11'h1BA];
        v0_443 = _RANDOM[11'h1BB];
        v0_444 = _RANDOM[11'h1BC];
        v0_445 = _RANDOM[11'h1BD];
        v0_446 = _RANDOM[11'h1BE];
        v0_447 = _RANDOM[11'h1BF];
        v0_448 = _RANDOM[11'h1C0];
        v0_449 = _RANDOM[11'h1C1];
        v0_450 = _RANDOM[11'h1C2];
        v0_451 = _RANDOM[11'h1C3];
        v0_452 = _RANDOM[11'h1C4];
        v0_453 = _RANDOM[11'h1C5];
        v0_454 = _RANDOM[11'h1C6];
        v0_455 = _RANDOM[11'h1C7];
        v0_456 = _RANDOM[11'h1C8];
        v0_457 = _RANDOM[11'h1C9];
        v0_458 = _RANDOM[11'h1CA];
        v0_459 = _RANDOM[11'h1CB];
        v0_460 = _RANDOM[11'h1CC];
        v0_461 = _RANDOM[11'h1CD];
        v0_462 = _RANDOM[11'h1CE];
        v0_463 = _RANDOM[11'h1CF];
        v0_464 = _RANDOM[11'h1D0];
        v0_465 = _RANDOM[11'h1D1];
        v0_466 = _RANDOM[11'h1D2];
        v0_467 = _RANDOM[11'h1D3];
        v0_468 = _RANDOM[11'h1D4];
        v0_469 = _RANDOM[11'h1D5];
        v0_470 = _RANDOM[11'h1D6];
        v0_471 = _RANDOM[11'h1D7];
        v0_472 = _RANDOM[11'h1D8];
        v0_473 = _RANDOM[11'h1D9];
        v0_474 = _RANDOM[11'h1DA];
        v0_475 = _RANDOM[11'h1DB];
        v0_476 = _RANDOM[11'h1DC];
        v0_477 = _RANDOM[11'h1DD];
        v0_478 = _RANDOM[11'h1DE];
        v0_479 = _RANDOM[11'h1DF];
        v0_480 = _RANDOM[11'h1E0];
        v0_481 = _RANDOM[11'h1E1];
        v0_482 = _RANDOM[11'h1E2];
        v0_483 = _RANDOM[11'h1E3];
        v0_484 = _RANDOM[11'h1E4];
        v0_485 = _RANDOM[11'h1E5];
        v0_486 = _RANDOM[11'h1E6];
        v0_487 = _RANDOM[11'h1E7];
        v0_488 = _RANDOM[11'h1E8];
        v0_489 = _RANDOM[11'h1E9];
        v0_490 = _RANDOM[11'h1EA];
        v0_491 = _RANDOM[11'h1EB];
        v0_492 = _RANDOM[11'h1EC];
        v0_493 = _RANDOM[11'h1ED];
        v0_494 = _RANDOM[11'h1EE];
        v0_495 = _RANDOM[11'h1EF];
        v0_496 = _RANDOM[11'h1F0];
        v0_497 = _RANDOM[11'h1F1];
        v0_498 = _RANDOM[11'h1F2];
        v0_499 = _RANDOM[11'h1F3];
        v0_500 = _RANDOM[11'h1F4];
        v0_501 = _RANDOM[11'h1F5];
        v0_502 = _RANDOM[11'h1F6];
        v0_503 = _RANDOM[11'h1F7];
        v0_504 = _RANDOM[11'h1F8];
        v0_505 = _RANDOM[11'h1F9];
        v0_506 = _RANDOM[11'h1FA];
        v0_507 = _RANDOM[11'h1FB];
        v0_508 = _RANDOM[11'h1FC];
        v0_509 = _RANDOM[11'h1FD];
        v0_510 = _RANDOM[11'h1FE];
        v0_511 = _RANDOM[11'h1FF];
        v0_512 = _RANDOM[11'h200];
        v0_513 = _RANDOM[11'h201];
        v0_514 = _RANDOM[11'h202];
        v0_515 = _RANDOM[11'h203];
        v0_516 = _RANDOM[11'h204];
        v0_517 = _RANDOM[11'h205];
        v0_518 = _RANDOM[11'h206];
        v0_519 = _RANDOM[11'h207];
        v0_520 = _RANDOM[11'h208];
        v0_521 = _RANDOM[11'h209];
        v0_522 = _RANDOM[11'h20A];
        v0_523 = _RANDOM[11'h20B];
        v0_524 = _RANDOM[11'h20C];
        v0_525 = _RANDOM[11'h20D];
        v0_526 = _RANDOM[11'h20E];
        v0_527 = _RANDOM[11'h20F];
        v0_528 = _RANDOM[11'h210];
        v0_529 = _RANDOM[11'h211];
        v0_530 = _RANDOM[11'h212];
        v0_531 = _RANDOM[11'h213];
        v0_532 = _RANDOM[11'h214];
        v0_533 = _RANDOM[11'h215];
        v0_534 = _RANDOM[11'h216];
        v0_535 = _RANDOM[11'h217];
        v0_536 = _RANDOM[11'h218];
        v0_537 = _RANDOM[11'h219];
        v0_538 = _RANDOM[11'h21A];
        v0_539 = _RANDOM[11'h21B];
        v0_540 = _RANDOM[11'h21C];
        v0_541 = _RANDOM[11'h21D];
        v0_542 = _RANDOM[11'h21E];
        v0_543 = _RANDOM[11'h21F];
        v0_544 = _RANDOM[11'h220];
        v0_545 = _RANDOM[11'h221];
        v0_546 = _RANDOM[11'h222];
        v0_547 = _RANDOM[11'h223];
        v0_548 = _RANDOM[11'h224];
        v0_549 = _RANDOM[11'h225];
        v0_550 = _RANDOM[11'h226];
        v0_551 = _RANDOM[11'h227];
        v0_552 = _RANDOM[11'h228];
        v0_553 = _RANDOM[11'h229];
        v0_554 = _RANDOM[11'h22A];
        v0_555 = _RANDOM[11'h22B];
        v0_556 = _RANDOM[11'h22C];
        v0_557 = _RANDOM[11'h22D];
        v0_558 = _RANDOM[11'h22E];
        v0_559 = _RANDOM[11'h22F];
        v0_560 = _RANDOM[11'h230];
        v0_561 = _RANDOM[11'h231];
        v0_562 = _RANDOM[11'h232];
        v0_563 = _RANDOM[11'h233];
        v0_564 = _RANDOM[11'h234];
        v0_565 = _RANDOM[11'h235];
        v0_566 = _RANDOM[11'h236];
        v0_567 = _RANDOM[11'h237];
        v0_568 = _RANDOM[11'h238];
        v0_569 = _RANDOM[11'h239];
        v0_570 = _RANDOM[11'h23A];
        v0_571 = _RANDOM[11'h23B];
        v0_572 = _RANDOM[11'h23C];
        v0_573 = _RANDOM[11'h23D];
        v0_574 = _RANDOM[11'h23E];
        v0_575 = _RANDOM[11'h23F];
        v0_576 = _RANDOM[11'h240];
        v0_577 = _RANDOM[11'h241];
        v0_578 = _RANDOM[11'h242];
        v0_579 = _RANDOM[11'h243];
        v0_580 = _RANDOM[11'h244];
        v0_581 = _RANDOM[11'h245];
        v0_582 = _RANDOM[11'h246];
        v0_583 = _RANDOM[11'h247];
        v0_584 = _RANDOM[11'h248];
        v0_585 = _RANDOM[11'h249];
        v0_586 = _RANDOM[11'h24A];
        v0_587 = _RANDOM[11'h24B];
        v0_588 = _RANDOM[11'h24C];
        v0_589 = _RANDOM[11'h24D];
        v0_590 = _RANDOM[11'h24E];
        v0_591 = _RANDOM[11'h24F];
        v0_592 = _RANDOM[11'h250];
        v0_593 = _RANDOM[11'h251];
        v0_594 = _RANDOM[11'h252];
        v0_595 = _RANDOM[11'h253];
        v0_596 = _RANDOM[11'h254];
        v0_597 = _RANDOM[11'h255];
        v0_598 = _RANDOM[11'h256];
        v0_599 = _RANDOM[11'h257];
        v0_600 = _RANDOM[11'h258];
        v0_601 = _RANDOM[11'h259];
        v0_602 = _RANDOM[11'h25A];
        v0_603 = _RANDOM[11'h25B];
        v0_604 = _RANDOM[11'h25C];
        v0_605 = _RANDOM[11'h25D];
        v0_606 = _RANDOM[11'h25E];
        v0_607 = _RANDOM[11'h25F];
        v0_608 = _RANDOM[11'h260];
        v0_609 = _RANDOM[11'h261];
        v0_610 = _RANDOM[11'h262];
        v0_611 = _RANDOM[11'h263];
        v0_612 = _RANDOM[11'h264];
        v0_613 = _RANDOM[11'h265];
        v0_614 = _RANDOM[11'h266];
        v0_615 = _RANDOM[11'h267];
        v0_616 = _RANDOM[11'h268];
        v0_617 = _RANDOM[11'h269];
        v0_618 = _RANDOM[11'h26A];
        v0_619 = _RANDOM[11'h26B];
        v0_620 = _RANDOM[11'h26C];
        v0_621 = _RANDOM[11'h26D];
        v0_622 = _RANDOM[11'h26E];
        v0_623 = _RANDOM[11'h26F];
        v0_624 = _RANDOM[11'h270];
        v0_625 = _RANDOM[11'h271];
        v0_626 = _RANDOM[11'h272];
        v0_627 = _RANDOM[11'h273];
        v0_628 = _RANDOM[11'h274];
        v0_629 = _RANDOM[11'h275];
        v0_630 = _RANDOM[11'h276];
        v0_631 = _RANDOM[11'h277];
        v0_632 = _RANDOM[11'h278];
        v0_633 = _RANDOM[11'h279];
        v0_634 = _RANDOM[11'h27A];
        v0_635 = _RANDOM[11'h27B];
        v0_636 = _RANDOM[11'h27C];
        v0_637 = _RANDOM[11'h27D];
        v0_638 = _RANDOM[11'h27E];
        v0_639 = _RANDOM[11'h27F];
        v0_640 = _RANDOM[11'h280];
        v0_641 = _RANDOM[11'h281];
        v0_642 = _RANDOM[11'h282];
        v0_643 = _RANDOM[11'h283];
        v0_644 = _RANDOM[11'h284];
        v0_645 = _RANDOM[11'h285];
        v0_646 = _RANDOM[11'h286];
        v0_647 = _RANDOM[11'h287];
        v0_648 = _RANDOM[11'h288];
        v0_649 = _RANDOM[11'h289];
        v0_650 = _RANDOM[11'h28A];
        v0_651 = _RANDOM[11'h28B];
        v0_652 = _RANDOM[11'h28C];
        v0_653 = _RANDOM[11'h28D];
        v0_654 = _RANDOM[11'h28E];
        v0_655 = _RANDOM[11'h28F];
        v0_656 = _RANDOM[11'h290];
        v0_657 = _RANDOM[11'h291];
        v0_658 = _RANDOM[11'h292];
        v0_659 = _RANDOM[11'h293];
        v0_660 = _RANDOM[11'h294];
        v0_661 = _RANDOM[11'h295];
        v0_662 = _RANDOM[11'h296];
        v0_663 = _RANDOM[11'h297];
        v0_664 = _RANDOM[11'h298];
        v0_665 = _RANDOM[11'h299];
        v0_666 = _RANDOM[11'h29A];
        v0_667 = _RANDOM[11'h29B];
        v0_668 = _RANDOM[11'h29C];
        v0_669 = _RANDOM[11'h29D];
        v0_670 = _RANDOM[11'h29E];
        v0_671 = _RANDOM[11'h29F];
        v0_672 = _RANDOM[11'h2A0];
        v0_673 = _RANDOM[11'h2A1];
        v0_674 = _RANDOM[11'h2A2];
        v0_675 = _RANDOM[11'h2A3];
        v0_676 = _RANDOM[11'h2A4];
        v0_677 = _RANDOM[11'h2A5];
        v0_678 = _RANDOM[11'h2A6];
        v0_679 = _RANDOM[11'h2A7];
        v0_680 = _RANDOM[11'h2A8];
        v0_681 = _RANDOM[11'h2A9];
        v0_682 = _RANDOM[11'h2AA];
        v0_683 = _RANDOM[11'h2AB];
        v0_684 = _RANDOM[11'h2AC];
        v0_685 = _RANDOM[11'h2AD];
        v0_686 = _RANDOM[11'h2AE];
        v0_687 = _RANDOM[11'h2AF];
        v0_688 = _RANDOM[11'h2B0];
        v0_689 = _RANDOM[11'h2B1];
        v0_690 = _RANDOM[11'h2B2];
        v0_691 = _RANDOM[11'h2B3];
        v0_692 = _RANDOM[11'h2B4];
        v0_693 = _RANDOM[11'h2B5];
        v0_694 = _RANDOM[11'h2B6];
        v0_695 = _RANDOM[11'h2B7];
        v0_696 = _RANDOM[11'h2B8];
        v0_697 = _RANDOM[11'h2B9];
        v0_698 = _RANDOM[11'h2BA];
        v0_699 = _RANDOM[11'h2BB];
        v0_700 = _RANDOM[11'h2BC];
        v0_701 = _RANDOM[11'h2BD];
        v0_702 = _RANDOM[11'h2BE];
        v0_703 = _RANDOM[11'h2BF];
        v0_704 = _RANDOM[11'h2C0];
        v0_705 = _RANDOM[11'h2C1];
        v0_706 = _RANDOM[11'h2C2];
        v0_707 = _RANDOM[11'h2C3];
        v0_708 = _RANDOM[11'h2C4];
        v0_709 = _RANDOM[11'h2C5];
        v0_710 = _RANDOM[11'h2C6];
        v0_711 = _RANDOM[11'h2C7];
        v0_712 = _RANDOM[11'h2C8];
        v0_713 = _RANDOM[11'h2C9];
        v0_714 = _RANDOM[11'h2CA];
        v0_715 = _RANDOM[11'h2CB];
        v0_716 = _RANDOM[11'h2CC];
        v0_717 = _RANDOM[11'h2CD];
        v0_718 = _RANDOM[11'h2CE];
        v0_719 = _RANDOM[11'h2CF];
        v0_720 = _RANDOM[11'h2D0];
        v0_721 = _RANDOM[11'h2D1];
        v0_722 = _RANDOM[11'h2D2];
        v0_723 = _RANDOM[11'h2D3];
        v0_724 = _RANDOM[11'h2D4];
        v0_725 = _RANDOM[11'h2D5];
        v0_726 = _RANDOM[11'h2D6];
        v0_727 = _RANDOM[11'h2D7];
        v0_728 = _RANDOM[11'h2D8];
        v0_729 = _RANDOM[11'h2D9];
        v0_730 = _RANDOM[11'h2DA];
        v0_731 = _RANDOM[11'h2DB];
        v0_732 = _RANDOM[11'h2DC];
        v0_733 = _RANDOM[11'h2DD];
        v0_734 = _RANDOM[11'h2DE];
        v0_735 = _RANDOM[11'h2DF];
        v0_736 = _RANDOM[11'h2E0];
        v0_737 = _RANDOM[11'h2E1];
        v0_738 = _RANDOM[11'h2E2];
        v0_739 = _RANDOM[11'h2E3];
        v0_740 = _RANDOM[11'h2E4];
        v0_741 = _RANDOM[11'h2E5];
        v0_742 = _RANDOM[11'h2E6];
        v0_743 = _RANDOM[11'h2E7];
        v0_744 = _RANDOM[11'h2E8];
        v0_745 = _RANDOM[11'h2E9];
        v0_746 = _RANDOM[11'h2EA];
        v0_747 = _RANDOM[11'h2EB];
        v0_748 = _RANDOM[11'h2EC];
        v0_749 = _RANDOM[11'h2ED];
        v0_750 = _RANDOM[11'h2EE];
        v0_751 = _RANDOM[11'h2EF];
        v0_752 = _RANDOM[11'h2F0];
        v0_753 = _RANDOM[11'h2F1];
        v0_754 = _RANDOM[11'h2F2];
        v0_755 = _RANDOM[11'h2F3];
        v0_756 = _RANDOM[11'h2F4];
        v0_757 = _RANDOM[11'h2F5];
        v0_758 = _RANDOM[11'h2F6];
        v0_759 = _RANDOM[11'h2F7];
        v0_760 = _RANDOM[11'h2F8];
        v0_761 = _RANDOM[11'h2F9];
        v0_762 = _RANDOM[11'h2FA];
        v0_763 = _RANDOM[11'h2FB];
        v0_764 = _RANDOM[11'h2FC];
        v0_765 = _RANDOM[11'h2FD];
        v0_766 = _RANDOM[11'h2FE];
        v0_767 = _RANDOM[11'h2FF];
        v0_768 = _RANDOM[11'h300];
        v0_769 = _RANDOM[11'h301];
        v0_770 = _RANDOM[11'h302];
        v0_771 = _RANDOM[11'h303];
        v0_772 = _RANDOM[11'h304];
        v0_773 = _RANDOM[11'h305];
        v0_774 = _RANDOM[11'h306];
        v0_775 = _RANDOM[11'h307];
        v0_776 = _RANDOM[11'h308];
        v0_777 = _RANDOM[11'h309];
        v0_778 = _RANDOM[11'h30A];
        v0_779 = _RANDOM[11'h30B];
        v0_780 = _RANDOM[11'h30C];
        v0_781 = _RANDOM[11'h30D];
        v0_782 = _RANDOM[11'h30E];
        v0_783 = _RANDOM[11'h30F];
        v0_784 = _RANDOM[11'h310];
        v0_785 = _RANDOM[11'h311];
        v0_786 = _RANDOM[11'h312];
        v0_787 = _RANDOM[11'h313];
        v0_788 = _RANDOM[11'h314];
        v0_789 = _RANDOM[11'h315];
        v0_790 = _RANDOM[11'h316];
        v0_791 = _RANDOM[11'h317];
        v0_792 = _RANDOM[11'h318];
        v0_793 = _RANDOM[11'h319];
        v0_794 = _RANDOM[11'h31A];
        v0_795 = _RANDOM[11'h31B];
        v0_796 = _RANDOM[11'h31C];
        v0_797 = _RANDOM[11'h31D];
        v0_798 = _RANDOM[11'h31E];
        v0_799 = _RANDOM[11'h31F];
        v0_800 = _RANDOM[11'h320];
        v0_801 = _RANDOM[11'h321];
        v0_802 = _RANDOM[11'h322];
        v0_803 = _RANDOM[11'h323];
        v0_804 = _RANDOM[11'h324];
        v0_805 = _RANDOM[11'h325];
        v0_806 = _RANDOM[11'h326];
        v0_807 = _RANDOM[11'h327];
        v0_808 = _RANDOM[11'h328];
        v0_809 = _RANDOM[11'h329];
        v0_810 = _RANDOM[11'h32A];
        v0_811 = _RANDOM[11'h32B];
        v0_812 = _RANDOM[11'h32C];
        v0_813 = _RANDOM[11'h32D];
        v0_814 = _RANDOM[11'h32E];
        v0_815 = _RANDOM[11'h32F];
        v0_816 = _RANDOM[11'h330];
        v0_817 = _RANDOM[11'h331];
        v0_818 = _RANDOM[11'h332];
        v0_819 = _RANDOM[11'h333];
        v0_820 = _RANDOM[11'h334];
        v0_821 = _RANDOM[11'h335];
        v0_822 = _RANDOM[11'h336];
        v0_823 = _RANDOM[11'h337];
        v0_824 = _RANDOM[11'h338];
        v0_825 = _RANDOM[11'h339];
        v0_826 = _RANDOM[11'h33A];
        v0_827 = _RANDOM[11'h33B];
        v0_828 = _RANDOM[11'h33C];
        v0_829 = _RANDOM[11'h33D];
        v0_830 = _RANDOM[11'h33E];
        v0_831 = _RANDOM[11'h33F];
        v0_832 = _RANDOM[11'h340];
        v0_833 = _RANDOM[11'h341];
        v0_834 = _RANDOM[11'h342];
        v0_835 = _RANDOM[11'h343];
        v0_836 = _RANDOM[11'h344];
        v0_837 = _RANDOM[11'h345];
        v0_838 = _RANDOM[11'h346];
        v0_839 = _RANDOM[11'h347];
        v0_840 = _RANDOM[11'h348];
        v0_841 = _RANDOM[11'h349];
        v0_842 = _RANDOM[11'h34A];
        v0_843 = _RANDOM[11'h34B];
        v0_844 = _RANDOM[11'h34C];
        v0_845 = _RANDOM[11'h34D];
        v0_846 = _RANDOM[11'h34E];
        v0_847 = _RANDOM[11'h34F];
        v0_848 = _RANDOM[11'h350];
        v0_849 = _RANDOM[11'h351];
        v0_850 = _RANDOM[11'h352];
        v0_851 = _RANDOM[11'h353];
        v0_852 = _RANDOM[11'h354];
        v0_853 = _RANDOM[11'h355];
        v0_854 = _RANDOM[11'h356];
        v0_855 = _RANDOM[11'h357];
        v0_856 = _RANDOM[11'h358];
        v0_857 = _RANDOM[11'h359];
        v0_858 = _RANDOM[11'h35A];
        v0_859 = _RANDOM[11'h35B];
        v0_860 = _RANDOM[11'h35C];
        v0_861 = _RANDOM[11'h35D];
        v0_862 = _RANDOM[11'h35E];
        v0_863 = _RANDOM[11'h35F];
        v0_864 = _RANDOM[11'h360];
        v0_865 = _RANDOM[11'h361];
        v0_866 = _RANDOM[11'h362];
        v0_867 = _RANDOM[11'h363];
        v0_868 = _RANDOM[11'h364];
        v0_869 = _RANDOM[11'h365];
        v0_870 = _RANDOM[11'h366];
        v0_871 = _RANDOM[11'h367];
        v0_872 = _RANDOM[11'h368];
        v0_873 = _RANDOM[11'h369];
        v0_874 = _RANDOM[11'h36A];
        v0_875 = _RANDOM[11'h36B];
        v0_876 = _RANDOM[11'h36C];
        v0_877 = _RANDOM[11'h36D];
        v0_878 = _RANDOM[11'h36E];
        v0_879 = _RANDOM[11'h36F];
        v0_880 = _RANDOM[11'h370];
        v0_881 = _RANDOM[11'h371];
        v0_882 = _RANDOM[11'h372];
        v0_883 = _RANDOM[11'h373];
        v0_884 = _RANDOM[11'h374];
        v0_885 = _RANDOM[11'h375];
        v0_886 = _RANDOM[11'h376];
        v0_887 = _RANDOM[11'h377];
        v0_888 = _RANDOM[11'h378];
        v0_889 = _RANDOM[11'h379];
        v0_890 = _RANDOM[11'h37A];
        v0_891 = _RANDOM[11'h37B];
        v0_892 = _RANDOM[11'h37C];
        v0_893 = _RANDOM[11'h37D];
        v0_894 = _RANDOM[11'h37E];
        v0_895 = _RANDOM[11'h37F];
        v0_896 = _RANDOM[11'h380];
        v0_897 = _RANDOM[11'h381];
        v0_898 = _RANDOM[11'h382];
        v0_899 = _RANDOM[11'h383];
        v0_900 = _RANDOM[11'h384];
        v0_901 = _RANDOM[11'h385];
        v0_902 = _RANDOM[11'h386];
        v0_903 = _RANDOM[11'h387];
        v0_904 = _RANDOM[11'h388];
        v0_905 = _RANDOM[11'h389];
        v0_906 = _RANDOM[11'h38A];
        v0_907 = _RANDOM[11'h38B];
        v0_908 = _RANDOM[11'h38C];
        v0_909 = _RANDOM[11'h38D];
        v0_910 = _RANDOM[11'h38E];
        v0_911 = _RANDOM[11'h38F];
        v0_912 = _RANDOM[11'h390];
        v0_913 = _RANDOM[11'h391];
        v0_914 = _RANDOM[11'h392];
        v0_915 = _RANDOM[11'h393];
        v0_916 = _RANDOM[11'h394];
        v0_917 = _RANDOM[11'h395];
        v0_918 = _RANDOM[11'h396];
        v0_919 = _RANDOM[11'h397];
        v0_920 = _RANDOM[11'h398];
        v0_921 = _RANDOM[11'h399];
        v0_922 = _RANDOM[11'h39A];
        v0_923 = _RANDOM[11'h39B];
        v0_924 = _RANDOM[11'h39C];
        v0_925 = _RANDOM[11'h39D];
        v0_926 = _RANDOM[11'h39E];
        v0_927 = _RANDOM[11'h39F];
        v0_928 = _RANDOM[11'h3A0];
        v0_929 = _RANDOM[11'h3A1];
        v0_930 = _RANDOM[11'h3A2];
        v0_931 = _RANDOM[11'h3A3];
        v0_932 = _RANDOM[11'h3A4];
        v0_933 = _RANDOM[11'h3A5];
        v0_934 = _RANDOM[11'h3A6];
        v0_935 = _RANDOM[11'h3A7];
        v0_936 = _RANDOM[11'h3A8];
        v0_937 = _RANDOM[11'h3A9];
        v0_938 = _RANDOM[11'h3AA];
        v0_939 = _RANDOM[11'h3AB];
        v0_940 = _RANDOM[11'h3AC];
        v0_941 = _RANDOM[11'h3AD];
        v0_942 = _RANDOM[11'h3AE];
        v0_943 = _RANDOM[11'h3AF];
        v0_944 = _RANDOM[11'h3B0];
        v0_945 = _RANDOM[11'h3B1];
        v0_946 = _RANDOM[11'h3B2];
        v0_947 = _RANDOM[11'h3B3];
        v0_948 = _RANDOM[11'h3B4];
        v0_949 = _RANDOM[11'h3B5];
        v0_950 = _RANDOM[11'h3B6];
        v0_951 = _RANDOM[11'h3B7];
        v0_952 = _RANDOM[11'h3B8];
        v0_953 = _RANDOM[11'h3B9];
        v0_954 = _RANDOM[11'h3BA];
        v0_955 = _RANDOM[11'h3BB];
        v0_956 = _RANDOM[11'h3BC];
        v0_957 = _RANDOM[11'h3BD];
        v0_958 = _RANDOM[11'h3BE];
        v0_959 = _RANDOM[11'h3BF];
        v0_960 = _RANDOM[11'h3C0];
        v0_961 = _RANDOM[11'h3C1];
        v0_962 = _RANDOM[11'h3C2];
        v0_963 = _RANDOM[11'h3C3];
        v0_964 = _RANDOM[11'h3C4];
        v0_965 = _RANDOM[11'h3C5];
        v0_966 = _RANDOM[11'h3C6];
        v0_967 = _RANDOM[11'h3C7];
        v0_968 = _RANDOM[11'h3C8];
        v0_969 = _RANDOM[11'h3C9];
        v0_970 = _RANDOM[11'h3CA];
        v0_971 = _RANDOM[11'h3CB];
        v0_972 = _RANDOM[11'h3CC];
        v0_973 = _RANDOM[11'h3CD];
        v0_974 = _RANDOM[11'h3CE];
        v0_975 = _RANDOM[11'h3CF];
        v0_976 = _RANDOM[11'h3D0];
        v0_977 = _RANDOM[11'h3D1];
        v0_978 = _RANDOM[11'h3D2];
        v0_979 = _RANDOM[11'h3D3];
        v0_980 = _RANDOM[11'h3D4];
        v0_981 = _RANDOM[11'h3D5];
        v0_982 = _RANDOM[11'h3D6];
        v0_983 = _RANDOM[11'h3D7];
        v0_984 = _RANDOM[11'h3D8];
        v0_985 = _RANDOM[11'h3D9];
        v0_986 = _RANDOM[11'h3DA];
        v0_987 = _RANDOM[11'h3DB];
        v0_988 = _RANDOM[11'h3DC];
        v0_989 = _RANDOM[11'h3DD];
        v0_990 = _RANDOM[11'h3DE];
        v0_991 = _RANDOM[11'h3DF];
        v0_992 = _RANDOM[11'h3E0];
        v0_993 = _RANDOM[11'h3E1];
        v0_994 = _RANDOM[11'h3E2];
        v0_995 = _RANDOM[11'h3E3];
        v0_996 = _RANDOM[11'h3E4];
        v0_997 = _RANDOM[11'h3E5];
        v0_998 = _RANDOM[11'h3E6];
        v0_999 = _RANDOM[11'h3E7];
        v0_1000 = _RANDOM[11'h3E8];
        v0_1001 = _RANDOM[11'h3E9];
        v0_1002 = _RANDOM[11'h3EA];
        v0_1003 = _RANDOM[11'h3EB];
        v0_1004 = _RANDOM[11'h3EC];
        v0_1005 = _RANDOM[11'h3ED];
        v0_1006 = _RANDOM[11'h3EE];
        v0_1007 = _RANDOM[11'h3EF];
        v0_1008 = _RANDOM[11'h3F0];
        v0_1009 = _RANDOM[11'h3F1];
        v0_1010 = _RANDOM[11'h3F2];
        v0_1011 = _RANDOM[11'h3F3];
        v0_1012 = _RANDOM[11'h3F4];
        v0_1013 = _RANDOM[11'h3F5];
        v0_1014 = _RANDOM[11'h3F6];
        v0_1015 = _RANDOM[11'h3F7];
        v0_1016 = _RANDOM[11'h3F8];
        v0_1017 = _RANDOM[11'h3F9];
        v0_1018 = _RANDOM[11'h3FA];
        v0_1019 = _RANDOM[11'h3FB];
        v0_1020 = _RANDOM[11'h3FC];
        v0_1021 = _RANDOM[11'h3FD];
        v0_1022 = _RANDOM[11'h3FE];
        v0_1023 = _RANDOM[11'h3FF];
        queueCount_0 = _RANDOM[11'h400][6:0];
        queueCount_1 = _RANDOM[11'h400][13:7];
        queueCount_2 = _RANDOM[11'h400][20:14];
        queueCount_3 = _RANDOM[11'h400][27:21];
        queueCount_4 = {_RANDOM[11'h400][31:28], _RANDOM[11'h401][2:0]};
        queueCount_5 = _RANDOM[11'h401][9:3];
        queueCount_6 = _RANDOM[11'h401][16:10];
        queueCount_7 = _RANDOM[11'h401][23:17];
        queueCount_0_1 = _RANDOM[11'h401][30:24];
        queueCount_1_1 = {_RANDOM[11'h401][31], _RANDOM[11'h402][5:0]};
        queueCount_2_1 = _RANDOM[11'h402][12:6];
        queueCount_3_1 = _RANDOM[11'h402][19:13];
        queueCount_4_1 = _RANDOM[11'h402][26:20];
        queueCount_5_1 = {_RANDOM[11'h402][31:27], _RANDOM[11'h403][1:0]};
        queueCount_6_1 = _RANDOM[11'h403][8:2];
        queueCount_7_1 = _RANDOM[11'h403][15:9];
        queueCount_0_2 = _RANDOM[11'h403][22:16];
        queueCount_1_2 = _RANDOM[11'h403][29:23];
        queueCount_2_2 = {_RANDOM[11'h403][31:30], _RANDOM[11'h404][4:0]};
        queueCount_3_2 = _RANDOM[11'h404][11:5];
        queueCount_4_2 = _RANDOM[11'h404][18:12];
        queueCount_5_2 = _RANDOM[11'h404][25:19];
        queueCount_6_2 = {_RANDOM[11'h404][31:26], _RANDOM[11'h405][0]};
        queueCount_7_2 = _RANDOM[11'h405][7:1];
        queueCount_0_3 = _RANDOM[11'h405][14:8];
        queueCount_1_3 = _RANDOM[11'h405][21:15];
        queueCount_2_3 = _RANDOM[11'h405][28:22];
        queueCount_3_3 = {_RANDOM[11'h405][31:29], _RANDOM[11'h406][3:0]};
        queueCount_4_3 = _RANDOM[11'h406][10:4];
        queueCount_5_3 = _RANDOM[11'h406][17:11];
        queueCount_6_3 = _RANDOM[11'h406][24:18];
        queueCount_7_3 = _RANDOM[11'h406][31:25];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire [11:0]         sourceQueue_deq_bits;
  wire [31:0]         axi4Port_aw_bits_addr_0;
  assign axi4Port_aw_bits_addr_0 = _storeUnit_memRequest_bits_address;
  assign dataQueue_enq_bits_index = _storeUnit_memRequest_bits_index;
  assign dataQueue_enq_bits_address = _storeUnit_memRequest_bits_address;
  wire [6:0]          simpleSourceQueue_deq_bits;
  wire [31:0]         simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_addr_0 = _otherUnit_memWriteRequest_bits_address;
  wire [3:0]          otherUnitTargetQueue_enq_bits;
  assign otherUnitTargetQueue_enq_bits = _otherUnit_status_targetLane;
  assign simpleDataQueue_enq_bits_source = _otherUnit_memWriteRequest_bits_source;
  assign simpleDataQueue_enq_bits_address = _otherUnit_memWriteRequest_bits_address;
  assign simpleDataQueue_enq_bits_size = _otherUnit_memWriteRequest_bits_size;
  wire                writeQueueVec_0_empty;
  assign writeQueueVec_0_empty = _writeQueueVec_fifo_empty;
  wire                writeQueueVec_0_full;
  assign writeQueueVec_0_full = _writeQueueVec_fifo_full;
  wire                writeQueueVec_1_empty;
  assign writeQueueVec_1_empty = _writeQueueVec_fifo_1_empty;
  wire                writeQueueVec_1_full;
  assign writeQueueVec_1_full = _writeQueueVec_fifo_1_full;
  wire                writeQueueVec_2_empty;
  assign writeQueueVec_2_empty = _writeQueueVec_fifo_2_empty;
  wire                writeQueueVec_2_full;
  assign writeQueueVec_2_full = _writeQueueVec_fifo_2_full;
  wire                writeQueueVec_3_empty;
  assign writeQueueVec_3_empty = _writeQueueVec_fifo_3_empty;
  wire                writeQueueVec_3_full;
  assign writeQueueVec_3_full = _writeQueueVec_fifo_3_full;
  assign otherUnitTargetQueue_empty = _otherUnitTargetQueue_fifo_empty;
  wire                otherUnitTargetQueue_full;
  assign otherUnitTargetQueue_full = _otherUnitTargetQueue_fifo_full;
  wire                otherUnitDataQueueVec_0_empty;
  assign otherUnitDataQueueVec_0_empty = _otherUnitDataQueueVec_fifo_empty;
  wire                otherUnitDataQueueVec_0_full;
  assign otherUnitDataQueueVec_0_full = _otherUnitDataQueueVec_fifo_full;
  wire                otherUnitDataQueueVec_1_empty;
  assign otherUnitDataQueueVec_1_empty = _otherUnitDataQueueVec_fifo_1_empty;
  wire                otherUnitDataQueueVec_1_full;
  assign otherUnitDataQueueVec_1_full = _otherUnitDataQueueVec_fifo_1_full;
  wire                otherUnitDataQueueVec_2_empty;
  assign otherUnitDataQueueVec_2_empty = _otherUnitDataQueueVec_fifo_2_empty;
  wire                otherUnitDataQueueVec_2_full;
  assign otherUnitDataQueueVec_2_full = _otherUnitDataQueueVec_fifo_2_full;
  wire                otherUnitDataQueueVec_3_empty;
  assign otherUnitDataQueueVec_3_empty = _otherUnitDataQueueVec_fifo_3_empty;
  wire                otherUnitDataQueueVec_3_full;
  assign otherUnitDataQueueVec_3_full = _otherUnitDataQueueVec_fifo_3_full;
  wire                writeIndexQueue_empty;
  assign writeIndexQueue_empty = _writeIndexQueue_fifo_empty;
  wire                writeIndexQueue_full;
  assign writeIndexQueue_full = _writeIndexQueue_fifo_full;
  wire                writeIndexQueue_1_empty;
  assign writeIndexQueue_1_empty = _writeIndexQueue_fifo_1_empty;
  wire                writeIndexQueue_1_full;
  assign writeIndexQueue_1_full = _writeIndexQueue_fifo_1_full;
  wire                writeIndexQueue_2_empty;
  assign writeIndexQueue_2_empty = _writeIndexQueue_fifo_2_empty;
  wire                writeIndexQueue_2_full;
  assign writeIndexQueue_2_full = _writeIndexQueue_fifo_2_full;
  wire                writeIndexQueue_3_empty;
  assign writeIndexQueue_3_empty = _writeIndexQueue_fifo_3_empty;
  wire                writeIndexQueue_3_full;
  assign writeIndexQueue_3_full = _writeIndexQueue_fifo_3_full;
  wire                sourceQueue_empty;
  assign sourceQueue_empty = _sourceQueue_fifo_empty;
  wire                sourceQueue_full;
  assign sourceQueue_full = _sourceQueue_fifo_full;
  wire                dataQueue_empty;
  assign dataQueue_empty = _dataQueue_fifo_empty;
  wire                dataQueue_full;
  assign dataQueue_full = _dataQueue_fifo_full;
  wire                simpleSourceQueue_empty;
  assign simpleSourceQueue_empty = _simpleSourceQueue_fifo_empty;
  wire                simpleSourceQueue_full;
  assign simpleSourceQueue_full = _simpleSourceQueue_fifo_full;
  wire                simpleDataQueue_empty;
  assign simpleDataQueue_empty = _simpleDataQueue_fifo_empty;
  wire                simpleDataQueue_full;
  assign simpleDataQueue_full = _simpleDataQueue_fifo_full;
  LoadUnit loadUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_0),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_511[maskSelect]),
    .maskSelect_valid                                       (_loadUnit_maskSelect_valid),
    .maskSelect_bits                                        (_loadUnit_maskSelect_bits),
    .addressConflict                                        (stallLoad),
    .memRequest_ready                                       (sourceQueue_enq_ready & axi4Port_ar_ready_0),
    .memRequest_valid                                       (_loadUnit_memRequest_valid),
    .memRequest_bits_src                                    (sourceQueue_enq_bits),
    .memRequest_bits_address                                (axi4Port_ar_bits_addr_0),
    .memResponse_ready                                      (axi4Port_r_ready_0),
    .memResponse_valid                                      (axi4Port_r_valid_0),
    .memResponse_bits_data                                  (axi4Port_r_bits_data_0),
    .memResponse_bits_index                                 (sourceQueue_deq_bits),
    .status_idle                                            (_loadUnit_status_idle),
    .status_last                                            (_loadUnit_status_last),
    .status_instructionIndex                                (_loadUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_loadUnit_status_startAddress),
    .status_endAddress                                      (_loadUnit_status_endAddress),
    .vrfWritePort_0_ready                                   (writeQueueVec_0_enq_ready & ~(otherTryToWrite[0])),
    .vrfWritePort_0_valid                                   (_loadUnit_vrfWritePort_0_valid),
    .vrfWritePort_0_bits_vd                                 (_loadUnit_vrfWritePort_0_bits_vd),
    .vrfWritePort_0_bits_offset                             (_loadUnit_vrfWritePort_0_bits_offset),
    .vrfWritePort_0_bits_mask                               (_loadUnit_vrfWritePort_0_bits_mask),
    .vrfWritePort_0_bits_data                               (_loadUnit_vrfWritePort_0_bits_data),
    .vrfWritePort_0_bits_instructionIndex                   (_loadUnit_vrfWritePort_0_bits_instructionIndex),
    .vrfWritePort_1_ready                                   (writeQueueVec_1_enq_ready & ~(otherTryToWrite[1])),
    .vrfWritePort_1_valid                                   (_loadUnit_vrfWritePort_1_valid),
    .vrfWritePort_1_bits_vd                                 (_loadUnit_vrfWritePort_1_bits_vd),
    .vrfWritePort_1_bits_offset                             (_loadUnit_vrfWritePort_1_bits_offset),
    .vrfWritePort_1_bits_mask                               (_loadUnit_vrfWritePort_1_bits_mask),
    .vrfWritePort_1_bits_data                               (_loadUnit_vrfWritePort_1_bits_data),
    .vrfWritePort_1_bits_instructionIndex                   (_loadUnit_vrfWritePort_1_bits_instructionIndex),
    .vrfWritePort_2_ready                                   (writeQueueVec_2_enq_ready & ~(otherTryToWrite[2])),
    .vrfWritePort_2_valid                                   (_loadUnit_vrfWritePort_2_valid),
    .vrfWritePort_2_bits_vd                                 (_loadUnit_vrfWritePort_2_bits_vd),
    .vrfWritePort_2_bits_offset                             (_loadUnit_vrfWritePort_2_bits_offset),
    .vrfWritePort_2_bits_mask                               (_loadUnit_vrfWritePort_2_bits_mask),
    .vrfWritePort_2_bits_data                               (_loadUnit_vrfWritePort_2_bits_data),
    .vrfWritePort_2_bits_instructionIndex                   (_loadUnit_vrfWritePort_2_bits_instructionIndex),
    .vrfWritePort_3_ready                                   (writeQueueVec_3_enq_ready & ~(otherTryToWrite[3])),
    .vrfWritePort_3_valid                                   (_loadUnit_vrfWritePort_3_valid),
    .vrfWritePort_3_bits_vd                                 (_loadUnit_vrfWritePort_3_bits_vd),
    .vrfWritePort_3_bits_offset                             (_loadUnit_vrfWritePort_3_bits_offset),
    .vrfWritePort_3_bits_mask                               (_loadUnit_vrfWritePort_3_bits_mask),
    .vrfWritePort_3_bits_data                               (_loadUnit_vrfWritePort_3_bits_data),
    .vrfWritePort_3_bits_instructionIndex                   (_loadUnit_vrfWritePort_3_bits_instructionIndex)
  );
  StoreUnit storeUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_1),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .maskInput                                              (_GEN_512[maskSelect_1]),
    .maskSelect_valid                                       (_storeUnit_maskSelect_valid),
    .maskSelect_bits                                        (_storeUnit_maskSelect_bits),
    .memRequest_ready                                       (axi4Port_aw_ready_0 & dataQueue_enq_ready),
    .memRequest_valid                                       (_storeUnit_memRequest_valid),
    .memRequest_bits_data                                   (dataQueue_enq_bits_data),
    .memRequest_bits_mask                                   (dataQueue_enq_bits_mask),
    .memRequest_bits_index                                  (_storeUnit_memRequest_bits_index),
    .memRequest_bits_address                                (_storeUnit_memRequest_bits_address),
    .status_idle                                            (_storeUnit_status_idle),
    .status_last                                            (_storeUnit_status_last),
    .status_instructionIndex                                (_storeUnit_status_instructionIndex),
    .status_changeMaskGroup                                 (/* unused */),
    .status_startAddress                                    (_storeUnit_status_startAddress),
    .status_endAddress                                      (_storeUnit_status_endAddress),
    .vrfReadDataPorts_0_ready                               (vrfReadDataPorts_0_ready_0 & ~(otherTryReadVrf[0])),
    .vrfReadDataPorts_0_valid                               (_storeUnit_vrfReadDataPorts_0_valid),
    .vrfReadDataPorts_0_bits_vs                             (_storeUnit_vrfReadDataPorts_0_bits_vs),
    .vrfReadDataPorts_0_bits_offset                         (_storeUnit_vrfReadDataPorts_0_bits_offset),
    .vrfReadDataPorts_0_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_0_bits_instructionIndex),
    .vrfReadDataPorts_1_ready                               (vrfReadDataPorts_1_ready_0 & ~(otherTryReadVrf[1])),
    .vrfReadDataPorts_1_valid                               (_storeUnit_vrfReadDataPorts_1_valid),
    .vrfReadDataPorts_1_bits_vs                             (_storeUnit_vrfReadDataPorts_1_bits_vs),
    .vrfReadDataPorts_1_bits_offset                         (_storeUnit_vrfReadDataPorts_1_bits_offset),
    .vrfReadDataPorts_1_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_1_bits_instructionIndex),
    .vrfReadDataPorts_2_ready                               (vrfReadDataPorts_2_ready_0 & ~(otherTryReadVrf[2])),
    .vrfReadDataPorts_2_valid                               (_storeUnit_vrfReadDataPorts_2_valid),
    .vrfReadDataPorts_2_bits_vs                             (_storeUnit_vrfReadDataPorts_2_bits_vs),
    .vrfReadDataPorts_2_bits_offset                         (_storeUnit_vrfReadDataPorts_2_bits_offset),
    .vrfReadDataPorts_2_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_2_bits_instructionIndex),
    .vrfReadDataPorts_3_ready                               (vrfReadDataPorts_3_ready_0 & ~(otherTryReadVrf[3])),
    .vrfReadDataPorts_3_valid                               (_storeUnit_vrfReadDataPorts_3_valid),
    .vrfReadDataPorts_3_bits_vs                             (_storeUnit_vrfReadDataPorts_3_bits_vs),
    .vrfReadDataPorts_3_bits_offset                         (_storeUnit_vrfReadDataPorts_3_bits_offset),
    .vrfReadDataPorts_3_bits_instructionIndex               (_storeUnit_vrfReadDataPorts_3_bits_instructionIndex),
    .vrfReadResults_0_valid                                 (vrfReadResults_0_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_0_bits                                  (vrfReadResults_0_bits),
    .vrfReadResults_1_valid                                 (vrfReadResults_1_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_1_bits                                  (vrfReadResults_1_bits),
    .vrfReadResults_2_valid                                 (vrfReadResults_2_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_2_bits                                  (vrfReadResults_2_bits),
    .vrfReadResults_3_valid                                 (vrfReadResults_3_valid & otherUnitTargetQueue_empty),
    .vrfReadResults_3_bits                                  (vrfReadResults_3_bits),
    .storeResponse                                          (axi4Port_b_valid_0)
  );
  SimpleAccessUnit otherUnit (
    .clock                                                  (clock),
    .reset                                                  (reset),
    .lsuRequest_valid                                       (reqEnq_2),
    .lsuRequest_bits_instructionInformation_nf              (request_bits_instructionInformation_nf_0),
    .lsuRequest_bits_instructionInformation_mew             (request_bits_instructionInformation_mew_0),
    .lsuRequest_bits_instructionInformation_mop             (request_bits_instructionInformation_mop_0),
    .lsuRequest_bits_instructionInformation_lumop           (request_bits_instructionInformation_lumop_0),
    .lsuRequest_bits_instructionInformation_eew             (request_bits_instructionInformation_eew_0),
    .lsuRequest_bits_instructionInformation_vs3             (request_bits_instructionInformation_vs3_0),
    .lsuRequest_bits_instructionInformation_isStore         (request_bits_instructionInformation_isStore_0),
    .lsuRequest_bits_instructionInformation_maskedLoadStore (request_bits_instructionInformation_maskedLoadStore_0),
    .lsuRequest_bits_rs1Data                                (request_bits_rs1Data_0),
    .lsuRequest_bits_rs2Data                                (request_bits_rs2Data_0),
    .lsuRequest_bits_instructionIndex                       (request_bits_instructionIndex_0),
    .vrfReadDataPorts_ready                                 (otherUnit_vrfReadDataPorts_ready),
    .vrfReadDataPorts_valid                                 (_otherUnit_vrfReadDataPorts_valid),
    .vrfReadDataPorts_bits_vs                               (_otherUnit_vrfReadDataPorts_bits_vs),
    .vrfReadDataPorts_bits_offset                           (_otherUnit_vrfReadDataPorts_bits_offset),
    .vrfReadDataPorts_bits_instructionIndex                 (_otherUnit_vrfReadDataPorts_bits_instructionIndex),
    .vrfReadResults_valid                                   (otherUnitTargetQueue_deq_ready),
    .vrfReadResults_bits
      ((otherUnitTargetQueue_deq_bits[0] ? otherUnitDataQueueVec_0_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[1] ? otherUnitDataQueueVec_1_deq_bits : 32'h0)
       | (otherUnitTargetQueue_deq_bits[2] ? otherUnitDataQueueVec_2_deq_bits : 32'h0) | (otherUnitTargetQueue_deq_bits[3] ? otherUnitDataQueueVec_3_deq_bits : 32'h0)),
    .offsetReadResult_0_valid                               (offsetReadResult_0_valid),
    .offsetReadResult_0_bits                                (offsetReadResult_0_bits),
    .offsetReadResult_1_valid                               (offsetReadResult_1_valid),
    .offsetReadResult_1_bits                                (offsetReadResult_1_bits),
    .offsetReadResult_2_valid                               (offsetReadResult_2_valid),
    .offsetReadResult_2_bits                                (offsetReadResult_2_bits),
    .offsetReadResult_3_valid                               (offsetReadResult_3_valid),
    .offsetReadResult_3_bits                                (offsetReadResult_3_bits),
    .maskInput                                              (_GEN_513[maskSelect_2]),
    .maskSelect_valid                                       (_otherUnit_maskSelect_valid),
    .maskSelect_bits                                        (_otherUnit_maskSelect_bits),
    .memReadRequest_ready                                   (simpleSourceQueue_enq_ready & simpleAccessPorts_ar_ready_0),
    .memReadRequest_valid                                   (_otherUnit_memReadRequest_valid),
    .memReadRequest_bits_address                            (simpleAccessPorts_ar_bits_addr_0),
    .memReadRequest_bits_source                             (simpleSourceQueue_enq_bits),
    .memReadResponse_ready                                  (simpleAccessPorts_r_ready_0),
    .memReadResponse_valid                                  (simpleAccessPorts_r_valid_0),
    .memReadResponse_bits_data                              (simpleAccessPorts_r_bits_data_0),
    .memReadResponse_bits_source                            (simpleSourceQueue_deq_bits),
    .memWriteRequest_ready                                  (simpleAccessPorts_aw_ready_0 & simpleDataQueue_enq_ready),
    .memWriteRequest_valid                                  (_otherUnit_memWriteRequest_valid),
    .memWriteRequest_bits_data                              (simpleDataQueue_enq_bits_data),
    .memWriteRequest_bits_mask                              (simpleDataQueue_enq_bits_mask),
    .memWriteRequest_bits_source                            (_otherUnit_memWriteRequest_bits_source),
    .memWriteRequest_bits_address                           (_otherUnit_memWriteRequest_bits_address),
    .memWriteRequest_bits_size                              (_otherUnit_memWriteRequest_bits_size),
    .vrfWritePort_ready                                     (|(_otherUnit_status_targetLane & {otherUnit_vrfWritePort_ready_hi, otherUnit_vrfWritePort_ready_lo})),
    .vrfWritePort_valid                                     (_otherUnit_vrfWritePort_valid),
    .vrfWritePort_bits_vd                                   (_otherUnit_vrfWritePort_bits_vd),
    .vrfWritePort_bits_offset                               (_otherUnit_vrfWritePort_bits_offset),
    .vrfWritePort_bits_mask                                 (_otherUnit_vrfWritePort_bits_mask),
    .vrfWritePort_bits_data                                 (_otherUnit_vrfWritePort_bits_data),
    .vrfWritePort_bits_last                                 (_otherUnit_vrfWritePort_bits_last),
    .vrfWritePort_bits_instructionIndex                     (_otherUnit_vrfWritePort_bits_instructionIndex),
    .csrInterface_vl                                        (csrInterface_vl),
    .csrInterface_vStart                                    (csrInterface_vStart),
    .csrInterface_vlmul                                     (csrInterface_vlmul),
    .csrInterface_vSew                                      (csrInterface_vSew),
    .csrInterface_vxrm                                      (csrInterface_vxrm),
    .csrInterface_vta                                       (csrInterface_vta),
    .csrInterface_vma                                       (csrInterface_vma),
    .status_idle                                            (_otherUnit_status_idle),
    .status_last                                            (_otherUnit_status_last),
    .status_instructionIndex                                (_otherUnit_status_instructionIndex),
    .status_targetLane                                      (_otherUnit_status_targetLane),
    .status_isStore                                         (_otherUnit_status_isStore),
    .offsetRelease_0                                        (_otherUnit_offsetRelease_0),
    .offsetRelease_1                                        (_otherUnit_offsetRelease_1),
    .offsetRelease_2                                        (_otherUnit_offsetRelease_2),
    .offsetRelease_3                                        (_otherUnit_offsetRelease_3)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(57)
  ) writeQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_0_writeValid_T & ~(_writeQueueVec_fifo_empty & writeQueueVec_0_deq_ready))),
    .pop_req_n    (~(writeQueueVec_0_deq_ready & ~_writeQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn),
    .empty        (_writeQueueVec_fifo_empty),
    .almost_empty (writeQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_0_almostFull),
    .full         (_writeQueueVec_fifo_full),
    .error        (_writeQueueVec_fifo_error),
    .data_out     (_writeQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(57)
  ) writeQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_1_writeValid_T & ~(_writeQueueVec_fifo_1_empty & writeQueueVec_1_deq_ready))),
    .pop_req_n    (~(writeQueueVec_1_deq_ready & ~_writeQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_1),
    .empty        (_writeQueueVec_fifo_1_empty),
    .almost_empty (writeQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_1_almostFull),
    .full         (_writeQueueVec_fifo_1_full),
    .error        (_writeQueueVec_fifo_1_error),
    .data_out     (_writeQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(57)
  ) writeQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_2_writeValid_T & ~(_writeQueueVec_fifo_2_empty & writeQueueVec_2_deq_ready))),
    .pop_req_n    (~(writeQueueVec_2_deq_ready & ~_writeQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_2),
    .empty        (_writeQueueVec_fifo_2_empty),
    .almost_empty (writeQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_2_almostFull),
    .full         (_writeQueueVec_fifo_2_full),
    .error        (_writeQueueVec_fifo_2_error),
    .data_out     (_writeQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(96),
    .err_mode(2),
    .rst_mode(3),
    .width(57)
  ) writeQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(_probeWire_slots_3_writeValid_T & ~(_writeQueueVec_fifo_3_empty & writeQueueVec_3_deq_ready))),
    .pop_req_n    (~(writeQueueVec_3_deq_ready & ~_writeQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueueVec_dataIn_3),
    .empty        (_writeQueueVec_fifo_3_empty),
    .almost_empty (writeQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueueVec_3_almostFull),
    .full         (_writeQueueVec_fifo_3_full),
    .error        (_writeQueueVec_fifo_3_error),
    .data_out     (_writeQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(4)
  ) otherUnitTargetQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitTargetQueue_enq_ready & otherUnitTargetQueue_enq_valid)),
    .pop_req_n    (~(otherUnitTargetQueue_deq_ready & ~_otherUnitTargetQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitTargetQueue_enq_bits),
    .empty        (_otherUnitTargetQueue_fifo_empty),
    .almost_empty (otherUnitTargetQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitTargetQueue_almostFull),
    .full         (_otherUnitTargetQueue_fifo_full),
    .error        (_otherUnitTargetQueue_fifo_error),
    .data_out     (otherUnitTargetQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_0_enq_ready & otherUnitDataQueueVec_0_enq_valid & ~(_otherUnitDataQueueVec_fifo_empty & otherUnitDataQueueVec_0_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_0_deq_ready & ~_otherUnitDataQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_0_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_empty),
    .almost_empty (otherUnitDataQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_0_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_full),
    .error        (_otherUnitDataQueueVec_fifo_error),
    .data_out     (_otherUnitDataQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_1_enq_ready & otherUnitDataQueueVec_1_enq_valid & ~(_otherUnitDataQueueVec_fifo_1_empty & otherUnitDataQueueVec_1_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_1_deq_ready & ~_otherUnitDataQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_1_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_1_empty),
    .almost_empty (otherUnitDataQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_1_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_1_full),
    .error        (_otherUnitDataQueueVec_fifo_1_error),
    .data_out     (_otherUnitDataQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_2_enq_ready & otherUnitDataQueueVec_2_enq_valid & ~(_otherUnitDataQueueVec_fifo_2_empty & otherUnitDataQueueVec_2_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_2_deq_ready & ~_otherUnitDataQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_2_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_2_empty),
    .almost_empty (otherUnitDataQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_2_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_2_full),
    .error        (_otherUnitDataQueueVec_fifo_2_error),
    .data_out     (_otherUnitDataQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) otherUnitDataQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(otherUnitDataQueueVec_3_enq_ready & otherUnitDataQueueVec_3_enq_valid & ~(_otherUnitDataQueueVec_fifo_3_empty & otherUnitDataQueueVec_3_deq_ready))),
    .pop_req_n    (~(otherUnitDataQueueVec_3_deq_ready & ~_otherUnitDataQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (otherUnitDataQueueVec_3_enq_bits),
    .empty        (_otherUnitDataQueueVec_fifo_3_empty),
    .almost_empty (otherUnitDataQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (otherUnitDataQueueVec_3_almostFull),
    .full         (_otherUnitDataQueueVec_fifo_3_full),
    .error        (_otherUnitDataQueueVec_fifo_3_error),
    .data_out     (_otherUnitDataQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_enq_ready & writeIndexQueue_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_deq_ready & ~_writeIndexQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_enq_bits),
    .empty        (_writeIndexQueue_fifo_empty),
    .almost_empty (writeIndexQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_almostFull),
    .full         (_writeIndexQueue_fifo_full),
    .error        (_writeIndexQueue_fifo_error),
    .data_out     (writeIndexQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_1_enq_ready & writeIndexQueue_1_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_1_deq_ready & ~_writeIndexQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_1_enq_bits),
    .empty        (_writeIndexQueue_fifo_1_empty),
    .almost_empty (writeIndexQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_1_almostFull),
    .full         (_writeIndexQueue_fifo_1_full),
    .error        (_writeIndexQueue_fifo_1_error),
    .data_out     (writeIndexQueue_1_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_2_enq_ready & writeIndexQueue_2_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_2_deq_ready & ~_writeIndexQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_2_enq_bits),
    .empty        (_writeIndexQueue_fifo_2_empty),
    .almost_empty (writeIndexQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_2_almostFull),
    .full         (_writeIndexQueue_fifo_2_full),
    .error        (_writeIndexQueue_fifo_2_error),
    .data_out     (writeIndexQueue_2_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(3)
  ) writeIndexQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeIndexQueue_3_enq_ready & writeIndexQueue_3_enq_valid)),
    .pop_req_n    (~(writeIndexQueue_3_deq_ready & ~_writeIndexQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeIndexQueue_3_enq_bits),
    .empty        (_writeIndexQueue_fifo_3_empty),
    .almost_empty (writeIndexQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeIndexQueue_3_almostFull),
    .full         (_writeIndexQueue_fifo_3_full),
    .error        (_writeIndexQueue_fifo_3_error),
    .data_out     (writeIndexQueue_3_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) sourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(sourceQueue_enq_ready & sourceQueue_enq_valid)),
    .pop_req_n    (~(sourceQueue_deq_ready & ~_sourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (sourceQueue_enq_bits),
    .empty        (_sourceQueue_fifo_empty),
    .almost_empty (sourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (sourceQueue_almostFull),
    .full         (_sourceQueue_fifo_full),
    .error        (_sourceQueue_fifo_error),
    .data_out     (sourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(188)
  ) dataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(dataQueue_enq_ready & dataQueue_enq_valid)),
    .pop_req_n    (~(dataQueue_deq_ready & ~_dataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (dataQueue_dataIn),
    .empty        (_dataQueue_fifo_empty),
    .almost_empty (dataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (dataQueue_almostFull),
    .full         (_dataQueue_fifo_full),
    .error        (_dataQueue_fifo_error),
    .data_out     (_dataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(7)
  ) simpleSourceQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleSourceQueue_enq_ready & simpleSourceQueue_enq_valid)),
    .pop_req_n    (~(simpleSourceQueue_deq_ready & ~_simpleSourceQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleSourceQueue_enq_bits),
    .empty        (_simpleSourceQueue_fifo_empty),
    .almost_empty (simpleSourceQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleSourceQueue_almostFull),
    .full         (_simpleSourceQueue_fifo_full),
    .error        (_simpleSourceQueue_fifo_error),
    .data_out     (simpleSourceQueue_deq_bits)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(2),
    .err_mode(2),
    .rst_mode(3),
    .width(78)
  ) simpleDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(simpleDataQueue_enq_ready & simpleDataQueue_enq_valid)),
    .pop_req_n    (~(simpleDataQueue_deq_ready & ~_simpleDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (simpleDataQueue_dataIn),
    .empty        (_simpleDataQueue_fifo_empty),
    .almost_empty (simpleDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (simpleDataQueue_almostFull),
    .full         (_simpleDataQueue_fifo_full),
    .error        (_simpleDataQueue_fifo_error),
    .data_out     (_simpleDataQueue_fifo_data_out)
  );
  assign request_ready = request_ready_0;
  assign axi4Port_aw_valid = axi4Port_aw_valid_0;
  assign axi4Port_aw_bits_id = axi4Port_aw_bits_id_0;
  assign axi4Port_aw_bits_addr = axi4Port_aw_bits_addr_0;
  assign axi4Port_w_valid = axi4Port_w_valid_0;
  assign axi4Port_w_bits_data = axi4Port_w_bits_data_0;
  assign axi4Port_w_bits_strb = axi4Port_w_bits_strb_0;
  assign axi4Port_ar_valid = axi4Port_ar_valid_0;
  assign axi4Port_ar_bits_addr = axi4Port_ar_bits_addr_0;
  assign axi4Port_r_ready = axi4Port_r_ready_0;
  assign simpleAccessPorts_aw_valid = simpleAccessPorts_aw_valid_0;
  assign simpleAccessPorts_aw_bits_id = simpleAccessPorts_aw_bits_id_0;
  assign simpleAccessPorts_aw_bits_addr = simpleAccessPorts_aw_bits_addr_0;
  assign simpleAccessPorts_aw_bits_size = simpleAccessPorts_aw_bits_size_0;
  assign simpleAccessPorts_w_valid = simpleAccessPorts_w_valid_0;
  assign simpleAccessPorts_w_bits_data = simpleAccessPorts_w_bits_data_0;
  assign simpleAccessPorts_w_bits_strb = simpleAccessPorts_w_bits_strb_0;
  assign simpleAccessPorts_ar_valid = simpleAccessPorts_ar_valid_0;
  assign simpleAccessPorts_ar_bits_addr = simpleAccessPorts_ar_bits_addr_0;
  assign simpleAccessPorts_r_ready = simpleAccessPorts_r_ready_0;
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_offset = vrfReadDataPorts_0_bits_offset_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_offset = vrfReadDataPorts_1_bits_offset_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_offset = vrfReadDataPorts_2_bits_offset_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_offset = vrfReadDataPorts_3_bits_offset_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_offset = vrfWritePort_0_bits_offset_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_last = vrfWritePort_0_bits_last_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_offset = vrfWritePort_1_bits_offset_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_last = vrfWritePort_1_bits_last_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_offset = vrfWritePort_2_bits_offset_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_last = vrfWritePort_2_bits_last_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_offset = vrfWritePort_3_bits_offset_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_last = vrfWritePort_3_bits_last_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
  assign dataInWriteQueue_0 = {dataInWriteQueue_0_hi, dataInWriteQueue_0_lo} | dataInMSHR;
  assign dataInWriteQueue_1 = {dataInWriteQueue_1_hi, dataInWriteQueue_1_lo} | dataInMSHR;
  assign dataInWriteQueue_2 = {dataInWriteQueue_2_hi, dataInWriteQueue_2_lo} | dataInMSHR;
  assign dataInWriteQueue_3 = {dataInWriteQueue_3_hi, dataInWriteQueue_3_lo} | dataInMSHR;
  assign lastReport = (_loadUnit_status_last ? 8'h1 << _GEN_514 : 8'h0) | (_storeUnit_status_last ? 8'h1 << _storeUnit_status_instructionIndex : 8'h0) | (_otherUnit_status_last ? 8'h1 << _GEN_515 : 8'h0);
  assign tokenIO_offsetGroupRelease = {tokenIO_offsetGroupRelease_hi, tokenIO_offsetGroupRelease_lo};
endmodule

