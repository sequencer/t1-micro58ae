
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskUnit(
  input         clock,
                reset,
                instReq_valid,
  input  [2:0]  instReq_bits_instructionIndex,
  input         instReq_bits_decodeResult_orderReduce,
                instReq_bits_decodeResult_floatMul,
  input  [1:0]  instReq_bits_decodeResult_fpExecutionType,
  input         instReq_bits_decodeResult_float,
                instReq_bits_decodeResult_specialSlot,
  input  [4:0]  instReq_bits_decodeResult_topUop,
  input         instReq_bits_decodeResult_popCount,
                instReq_bits_decodeResult_ffo,
                instReq_bits_decodeResult_average,
                instReq_bits_decodeResult_reverse,
                instReq_bits_decodeResult_dontNeedExecuteInLane,
                instReq_bits_decodeResult_scheduler,
                instReq_bits_decodeResult_sReadVD,
                instReq_bits_decodeResult_vtype,
                instReq_bits_decodeResult_sWrite,
                instReq_bits_decodeResult_crossRead,
                instReq_bits_decodeResult_crossWrite,
                instReq_bits_decodeResult_maskUnit,
                instReq_bits_decodeResult_special,
                instReq_bits_decodeResult_saturate,
                instReq_bits_decodeResult_vwmacc,
                instReq_bits_decodeResult_readOnly,
                instReq_bits_decodeResult_maskSource,
                instReq_bits_decodeResult_maskDestination,
                instReq_bits_decodeResult_maskLogic,
  input  [3:0]  instReq_bits_decodeResult_uop,
  input         instReq_bits_decodeResult_iota,
                instReq_bits_decodeResult_mv,
                instReq_bits_decodeResult_extend,
                instReq_bits_decodeResult_unOrderWrite,
                instReq_bits_decodeResult_compress,
                instReq_bits_decodeResult_gather16,
                instReq_bits_decodeResult_gather,
                instReq_bits_decodeResult_slid,
                instReq_bits_decodeResult_targetRd,
                instReq_bits_decodeResult_widenReduce,
                instReq_bits_decodeResult_red,
                instReq_bits_decodeResult_nr,
                instReq_bits_decodeResult_itype,
                instReq_bits_decodeResult_unsigned1,
                instReq_bits_decodeResult_unsigned0,
                instReq_bits_decodeResult_other,
                instReq_bits_decodeResult_multiCycle,
                instReq_bits_decodeResult_divider,
                instReq_bits_decodeResult_multiplier,
                instReq_bits_decodeResult_shift,
                instReq_bits_decodeResult_adder,
                instReq_bits_decodeResult_logic,
  input  [31:0] instReq_bits_readFromScala,
  input  [1:0]  instReq_bits_sew,
  input  [2:0]  instReq_bits_vlmul,
  input         instReq_bits_maskType,
  input  [2:0]  instReq_bits_vxrm,
  input  [4:0]  instReq_bits_vs2,
                instReq_bits_vs1,
                instReq_bits_vd,
  input  [10:0] instReq_bits_vl,
  input         exeReq_0_valid,
  input  [31:0] exeReq_0_bits_source1,
                exeReq_0_bits_source2,
  input  [2:0]  exeReq_0_bits_index,
  input         exeReq_0_bits_ffo,
                exeReq_0_bits_fpReduceValid,
                exeReq_1_valid,
  input  [31:0] exeReq_1_bits_source1,
                exeReq_1_bits_source2,
  input  [2:0]  exeReq_1_bits_index,
  input         exeReq_1_bits_ffo,
                exeReq_1_bits_fpReduceValid,
                exeReq_2_valid,
  input  [31:0] exeReq_2_bits_source1,
                exeReq_2_bits_source2,
  input  [2:0]  exeReq_2_bits_index,
  input         exeReq_2_bits_ffo,
                exeReq_2_bits_fpReduceValid,
                exeReq_3_valid,
  input  [31:0] exeReq_3_bits_source1,
                exeReq_3_bits_source2,
  input  [2:0]  exeReq_3_bits_index,
  input         exeReq_3_bits_ffo,
                exeReq_3_bits_fpReduceValid,
                exeReq_4_valid,
  input  [31:0] exeReq_4_bits_source1,
                exeReq_4_bits_source2,
  input  [2:0]  exeReq_4_bits_index,
  input         exeReq_4_bits_ffo,
                exeReq_4_bits_fpReduceValid,
                exeReq_5_valid,
  input  [31:0] exeReq_5_bits_source1,
                exeReq_5_bits_source2,
  input  [2:0]  exeReq_5_bits_index,
  input         exeReq_5_bits_ffo,
                exeReq_5_bits_fpReduceValid,
                exeReq_6_valid,
  input  [31:0] exeReq_6_bits_source1,
                exeReq_6_bits_source2,
  input  [2:0]  exeReq_6_bits_index,
  input         exeReq_6_bits_ffo,
                exeReq_6_bits_fpReduceValid,
                exeReq_7_valid,
  input  [31:0] exeReq_7_bits_source1,
                exeReq_7_bits_source2,
  input  [2:0]  exeReq_7_bits_index,
  input         exeReq_7_bits_ffo,
                exeReq_7_bits_fpReduceValid,
                exeReq_8_valid,
  input  [31:0] exeReq_8_bits_source1,
                exeReq_8_bits_source2,
  input  [2:0]  exeReq_8_bits_index,
  input         exeReq_8_bits_ffo,
                exeReq_8_bits_fpReduceValid,
                exeReq_9_valid,
  input  [31:0] exeReq_9_bits_source1,
                exeReq_9_bits_source2,
  input  [2:0]  exeReq_9_bits_index,
  input         exeReq_9_bits_ffo,
                exeReq_9_bits_fpReduceValid,
                exeReq_10_valid,
  input  [31:0] exeReq_10_bits_source1,
                exeReq_10_bits_source2,
  input  [2:0]  exeReq_10_bits_index,
  input         exeReq_10_bits_ffo,
                exeReq_10_bits_fpReduceValid,
                exeReq_11_valid,
  input  [31:0] exeReq_11_bits_source1,
                exeReq_11_bits_source2,
  input  [2:0]  exeReq_11_bits_index,
  input         exeReq_11_bits_ffo,
                exeReq_11_bits_fpReduceValid,
                exeReq_12_valid,
  input  [31:0] exeReq_12_bits_source1,
                exeReq_12_bits_source2,
  input  [2:0]  exeReq_12_bits_index,
  input         exeReq_12_bits_ffo,
                exeReq_12_bits_fpReduceValid,
                exeReq_13_valid,
  input  [31:0] exeReq_13_bits_source1,
                exeReq_13_bits_source2,
  input  [2:0]  exeReq_13_bits_index,
  input         exeReq_13_bits_ffo,
                exeReq_13_bits_fpReduceValid,
                exeReq_14_valid,
  input  [31:0] exeReq_14_bits_source1,
                exeReq_14_bits_source2,
  input  [2:0]  exeReq_14_bits_index,
  input         exeReq_14_bits_ffo,
                exeReq_14_bits_fpReduceValid,
                exeReq_15_valid,
  input  [31:0] exeReq_15_bits_source1,
                exeReq_15_bits_source2,
  input  [2:0]  exeReq_15_bits_index,
  input         exeReq_15_bits_ffo,
                exeReq_15_bits_fpReduceValid,
                exeResp_0_ready,
  output        exeResp_0_valid,
  output [4:0]  exeResp_0_bits_vd,
  output        exeResp_0_bits_offset,
  output [3:0]  exeResp_0_bits_mask,
  output [31:0] exeResp_0_bits_data,
  output [2:0]  exeResp_0_bits_instructionIndex,
  input         exeResp_1_ready,
  output        exeResp_1_valid,
  output [4:0]  exeResp_1_bits_vd,
  output        exeResp_1_bits_offset,
  output [3:0]  exeResp_1_bits_mask,
  output [31:0] exeResp_1_bits_data,
  output [2:0]  exeResp_1_bits_instructionIndex,
  input         exeResp_2_ready,
  output        exeResp_2_valid,
  output [4:0]  exeResp_2_bits_vd,
  output        exeResp_2_bits_offset,
  output [3:0]  exeResp_2_bits_mask,
  output [31:0] exeResp_2_bits_data,
  output [2:0]  exeResp_2_bits_instructionIndex,
  input         exeResp_3_ready,
  output        exeResp_3_valid,
  output [4:0]  exeResp_3_bits_vd,
  output        exeResp_3_bits_offset,
  output [3:0]  exeResp_3_bits_mask,
  output [31:0] exeResp_3_bits_data,
  output [2:0]  exeResp_3_bits_instructionIndex,
  input         exeResp_4_ready,
  output        exeResp_4_valid,
  output [4:0]  exeResp_4_bits_vd,
  output        exeResp_4_bits_offset,
  output [3:0]  exeResp_4_bits_mask,
  output [31:0] exeResp_4_bits_data,
  output [2:0]  exeResp_4_bits_instructionIndex,
  input         exeResp_5_ready,
  output        exeResp_5_valid,
  output [4:0]  exeResp_5_bits_vd,
  output        exeResp_5_bits_offset,
  output [3:0]  exeResp_5_bits_mask,
  output [31:0] exeResp_5_bits_data,
  output [2:0]  exeResp_5_bits_instructionIndex,
  input         exeResp_6_ready,
  output        exeResp_6_valid,
  output [4:0]  exeResp_6_bits_vd,
  output        exeResp_6_bits_offset,
  output [3:0]  exeResp_6_bits_mask,
  output [31:0] exeResp_6_bits_data,
  output [2:0]  exeResp_6_bits_instructionIndex,
  input         exeResp_7_ready,
  output        exeResp_7_valid,
  output [4:0]  exeResp_7_bits_vd,
  output        exeResp_7_bits_offset,
  output [3:0]  exeResp_7_bits_mask,
  output [31:0] exeResp_7_bits_data,
  output [2:0]  exeResp_7_bits_instructionIndex,
  input         exeResp_8_ready,
  output        exeResp_8_valid,
  output [4:0]  exeResp_8_bits_vd,
  output        exeResp_8_bits_offset,
  output [3:0]  exeResp_8_bits_mask,
  output [31:0] exeResp_8_bits_data,
  output [2:0]  exeResp_8_bits_instructionIndex,
  input         exeResp_9_ready,
  output        exeResp_9_valid,
  output [4:0]  exeResp_9_bits_vd,
  output        exeResp_9_bits_offset,
  output [3:0]  exeResp_9_bits_mask,
  output [31:0] exeResp_9_bits_data,
  output [2:0]  exeResp_9_bits_instructionIndex,
  input         exeResp_10_ready,
  output        exeResp_10_valid,
  output [4:0]  exeResp_10_bits_vd,
  output        exeResp_10_bits_offset,
  output [3:0]  exeResp_10_bits_mask,
  output [31:0] exeResp_10_bits_data,
  output [2:0]  exeResp_10_bits_instructionIndex,
  input         exeResp_11_ready,
  output        exeResp_11_valid,
  output [4:0]  exeResp_11_bits_vd,
  output        exeResp_11_bits_offset,
  output [3:0]  exeResp_11_bits_mask,
  output [31:0] exeResp_11_bits_data,
  output [2:0]  exeResp_11_bits_instructionIndex,
  input         exeResp_12_ready,
  output        exeResp_12_valid,
  output [4:0]  exeResp_12_bits_vd,
  output        exeResp_12_bits_offset,
  output [3:0]  exeResp_12_bits_mask,
  output [31:0] exeResp_12_bits_data,
  output [2:0]  exeResp_12_bits_instructionIndex,
  input         exeResp_13_ready,
  output        exeResp_13_valid,
  output [4:0]  exeResp_13_bits_vd,
  output        exeResp_13_bits_offset,
  output [3:0]  exeResp_13_bits_mask,
  output [31:0] exeResp_13_bits_data,
  output [2:0]  exeResp_13_bits_instructionIndex,
  input         exeResp_14_ready,
  output        exeResp_14_valid,
  output [4:0]  exeResp_14_bits_vd,
  output        exeResp_14_bits_offset,
  output [3:0]  exeResp_14_bits_mask,
  output [31:0] exeResp_14_bits_data,
  output [2:0]  exeResp_14_bits_instructionIndex,
  input         exeResp_15_ready,
  output        exeResp_15_valid,
  output [4:0]  exeResp_15_bits_vd,
  output        exeResp_15_bits_offset,
  output [3:0]  exeResp_15_bits_mask,
  output [31:0] exeResp_15_bits_data,
  output [2:0]  exeResp_15_bits_instructionIndex,
  input         writeRelease_0,
                writeRelease_1,
                writeRelease_2,
                writeRelease_3,
                writeRelease_4,
                writeRelease_5,
                writeRelease_6,
                writeRelease_7,
                writeRelease_8,
                writeRelease_9,
                writeRelease_10,
                writeRelease_11,
                writeRelease_12,
                writeRelease_13,
                writeRelease_14,
                writeRelease_15,
  output        tokenIO_0_maskRequestRelease,
                tokenIO_1_maskRequestRelease,
                tokenIO_2_maskRequestRelease,
                tokenIO_3_maskRequestRelease,
                tokenIO_4_maskRequestRelease,
                tokenIO_5_maskRequestRelease,
                tokenIO_6_maskRequestRelease,
                tokenIO_7_maskRequestRelease,
                tokenIO_8_maskRequestRelease,
                tokenIO_9_maskRequestRelease,
                tokenIO_10_maskRequestRelease,
                tokenIO_11_maskRequestRelease,
                tokenIO_12_maskRequestRelease,
                tokenIO_13_maskRequestRelease,
                tokenIO_14_maskRequestRelease,
                tokenIO_15_maskRequestRelease,
  input         readChannel_0_ready,
  output        readChannel_0_valid,
  output [4:0]  readChannel_0_bits_vs,
  output        readChannel_0_bits_offset,
  output [2:0]  readChannel_0_bits_instructionIndex,
  input         readChannel_1_ready,
  output        readChannel_1_valid,
  output [4:0]  readChannel_1_bits_vs,
  output        readChannel_1_bits_offset,
  output [2:0]  readChannel_1_bits_instructionIndex,
  input         readChannel_2_ready,
  output        readChannel_2_valid,
  output [4:0]  readChannel_2_bits_vs,
  output        readChannel_2_bits_offset,
  output [2:0]  readChannel_2_bits_instructionIndex,
  input         readChannel_3_ready,
  output        readChannel_3_valid,
  output [4:0]  readChannel_3_bits_vs,
  output        readChannel_3_bits_offset,
  output [2:0]  readChannel_3_bits_instructionIndex,
  input         readChannel_4_ready,
  output        readChannel_4_valid,
  output [4:0]  readChannel_4_bits_vs,
  output        readChannel_4_bits_offset,
  output [2:0]  readChannel_4_bits_instructionIndex,
  input         readChannel_5_ready,
  output        readChannel_5_valid,
  output [4:0]  readChannel_5_bits_vs,
  output        readChannel_5_bits_offset,
  output [2:0]  readChannel_5_bits_instructionIndex,
  input         readChannel_6_ready,
  output        readChannel_6_valid,
  output [4:0]  readChannel_6_bits_vs,
  output        readChannel_6_bits_offset,
  output [2:0]  readChannel_6_bits_instructionIndex,
  input         readChannel_7_ready,
  output        readChannel_7_valid,
  output [4:0]  readChannel_7_bits_vs,
  output        readChannel_7_bits_offset,
  output [2:0]  readChannel_7_bits_instructionIndex,
  input         readChannel_8_ready,
  output        readChannel_8_valid,
  output [4:0]  readChannel_8_bits_vs,
  output        readChannel_8_bits_offset,
  output [2:0]  readChannel_8_bits_instructionIndex,
  input         readChannel_9_ready,
  output        readChannel_9_valid,
  output [4:0]  readChannel_9_bits_vs,
  output        readChannel_9_bits_offset,
  output [2:0]  readChannel_9_bits_instructionIndex,
  input         readChannel_10_ready,
  output        readChannel_10_valid,
  output [4:0]  readChannel_10_bits_vs,
  output        readChannel_10_bits_offset,
  output [2:0]  readChannel_10_bits_instructionIndex,
  input         readChannel_11_ready,
  output        readChannel_11_valid,
  output [4:0]  readChannel_11_bits_vs,
  output        readChannel_11_bits_offset,
  output [2:0]  readChannel_11_bits_instructionIndex,
  input         readChannel_12_ready,
  output        readChannel_12_valid,
  output [4:0]  readChannel_12_bits_vs,
  output        readChannel_12_bits_offset,
  output [2:0]  readChannel_12_bits_instructionIndex,
  input         readChannel_13_ready,
  output        readChannel_13_valid,
  output [4:0]  readChannel_13_bits_vs,
  output        readChannel_13_bits_offset,
  output [2:0]  readChannel_13_bits_instructionIndex,
  input         readChannel_14_ready,
  output        readChannel_14_valid,
  output [4:0]  readChannel_14_bits_vs,
  output        readChannel_14_bits_offset,
  output [2:0]  readChannel_14_bits_instructionIndex,
  input         readChannel_15_ready,
  output        readChannel_15_valid,
  output [4:0]  readChannel_15_bits_vs,
  output        readChannel_15_bits_offset,
  output [2:0]  readChannel_15_bits_instructionIndex,
  input         readResult_0_valid,
  input  [31:0] readResult_0_bits,
  input         readResult_1_valid,
  input  [31:0] readResult_1_bits,
  input         readResult_2_valid,
  input  [31:0] readResult_2_bits,
  input         readResult_3_valid,
  input  [31:0] readResult_3_bits,
  input         readResult_4_valid,
  input  [31:0] readResult_4_bits,
  input         readResult_5_valid,
  input  [31:0] readResult_5_bits,
  input         readResult_6_valid,
  input  [31:0] readResult_6_bits,
  input         readResult_7_valid,
  input  [31:0] readResult_7_bits,
  input         readResult_8_valid,
  input  [31:0] readResult_8_bits,
  input         readResult_9_valid,
  input  [31:0] readResult_9_bits,
  input         readResult_10_valid,
  input  [31:0] readResult_10_bits,
  input         readResult_11_valid,
  input  [31:0] readResult_11_bits,
  input         readResult_12_valid,
  input  [31:0] readResult_12_bits,
  input         readResult_13_valid,
  input  [31:0] readResult_13_bits,
  input         readResult_14_valid,
  input  [31:0] readResult_14_bits,
  input         readResult_15_valid,
  input  [31:0] readResult_15_bits,
  output [7:0]  lastReport,
  output [31:0] laneMaskInput_0,
                laneMaskInput_1,
                laneMaskInput_2,
                laneMaskInput_3,
                laneMaskInput_4,
                laneMaskInput_5,
                laneMaskInput_6,
                laneMaskInput_7,
                laneMaskInput_8,
                laneMaskInput_9,
                laneMaskInput_10,
                laneMaskInput_11,
                laneMaskInput_12,
                laneMaskInput_13,
                laneMaskInput_14,
                laneMaskInput_15,
  input  [4:0]  laneMaskSelect_0,
                laneMaskSelect_1,
                laneMaskSelect_2,
                laneMaskSelect_3,
                laneMaskSelect_4,
                laneMaskSelect_5,
                laneMaskSelect_6,
                laneMaskSelect_7,
                laneMaskSelect_8,
                laneMaskSelect_9,
                laneMaskSelect_10,
                laneMaskSelect_11,
                laneMaskSelect_12,
                laneMaskSelect_13,
                laneMaskSelect_14,
                laneMaskSelect_15,
  input  [1:0]  laneMaskSewSelect_0,
                laneMaskSewSelect_1,
                laneMaskSewSelect_2,
                laneMaskSewSelect_3,
                laneMaskSewSelect_4,
                laneMaskSewSelect_5,
                laneMaskSewSelect_6,
                laneMaskSewSelect_7,
                laneMaskSewSelect_8,
                laneMaskSewSelect_9,
                laneMaskSewSelect_10,
                laneMaskSewSelect_11,
                laneMaskSewSelect_12,
                laneMaskSewSelect_13,
                laneMaskSewSelect_14,
                laneMaskSewSelect_15,
  input         v0UpdateVec_0_valid,
  input  [31:0] v0UpdateVec_0_bits_data,
  input         v0UpdateVec_0_bits_offset,
  input  [3:0]  v0UpdateVec_0_bits_mask,
  input         v0UpdateVec_1_valid,
  input  [31:0] v0UpdateVec_1_bits_data,
  input         v0UpdateVec_1_bits_offset,
  input  [3:0]  v0UpdateVec_1_bits_mask,
  input         v0UpdateVec_2_valid,
  input  [31:0] v0UpdateVec_2_bits_data,
  input         v0UpdateVec_2_bits_offset,
  input  [3:0]  v0UpdateVec_2_bits_mask,
  input         v0UpdateVec_3_valid,
  input  [31:0] v0UpdateVec_3_bits_data,
  input         v0UpdateVec_3_bits_offset,
  input  [3:0]  v0UpdateVec_3_bits_mask,
  input         v0UpdateVec_4_valid,
  input  [31:0] v0UpdateVec_4_bits_data,
  input         v0UpdateVec_4_bits_offset,
  input  [3:0]  v0UpdateVec_4_bits_mask,
  input         v0UpdateVec_5_valid,
  input  [31:0] v0UpdateVec_5_bits_data,
  input         v0UpdateVec_5_bits_offset,
  input  [3:0]  v0UpdateVec_5_bits_mask,
  input         v0UpdateVec_6_valid,
  input  [31:0] v0UpdateVec_6_bits_data,
  input         v0UpdateVec_6_bits_offset,
  input  [3:0]  v0UpdateVec_6_bits_mask,
  input         v0UpdateVec_7_valid,
  input  [31:0] v0UpdateVec_7_bits_data,
  input         v0UpdateVec_7_bits_offset,
  input  [3:0]  v0UpdateVec_7_bits_mask,
  input         v0UpdateVec_8_valid,
  input  [31:0] v0UpdateVec_8_bits_data,
  input         v0UpdateVec_8_bits_offset,
  input  [3:0]  v0UpdateVec_8_bits_mask,
  input         v0UpdateVec_9_valid,
  input  [31:0] v0UpdateVec_9_bits_data,
  input         v0UpdateVec_9_bits_offset,
  input  [3:0]  v0UpdateVec_9_bits_mask,
  input         v0UpdateVec_10_valid,
  input  [31:0] v0UpdateVec_10_bits_data,
  input         v0UpdateVec_10_bits_offset,
  input  [3:0]  v0UpdateVec_10_bits_mask,
  input         v0UpdateVec_11_valid,
  input  [31:0] v0UpdateVec_11_bits_data,
  input         v0UpdateVec_11_bits_offset,
  input  [3:0]  v0UpdateVec_11_bits_mask,
  input         v0UpdateVec_12_valid,
  input  [31:0] v0UpdateVec_12_bits_data,
  input         v0UpdateVec_12_bits_offset,
  input  [3:0]  v0UpdateVec_12_bits_mask,
  input         v0UpdateVec_13_valid,
  input  [31:0] v0UpdateVec_13_bits_data,
  input         v0UpdateVec_13_bits_offset,
  input  [3:0]  v0UpdateVec_13_bits_mask,
  input         v0UpdateVec_14_valid,
  input  [31:0] v0UpdateVec_14_bits_data,
  input         v0UpdateVec_14_bits_offset,
  input  [3:0]  v0UpdateVec_14_bits_mask,
  input         v0UpdateVec_15_valid,
  input  [31:0] v0UpdateVec_15_bits_data,
  input         v0UpdateVec_15_bits_offset,
  input  [3:0]  v0UpdateVec_15_bits_mask,
  output [31:0] writeRDData,
  input         gatherData_ready,
  output        gatherData_valid,
  output [31:0] gatherData_bits,
  input         gatherRead
);

  wire              readCrossBar_input_15_valid;
  wire              readCrossBar_input_14_valid;
  wire              readCrossBar_input_13_valid;
  wire              readCrossBar_input_12_valid;
  wire              readCrossBar_input_11_valid;
  wire              readCrossBar_input_10_valid;
  wire              readCrossBar_input_9_valid;
  wire              readCrossBar_input_8_valid;
  wire              readCrossBar_input_7_valid;
  wire              readCrossBar_input_6_valid;
  wire              readCrossBar_input_5_valid;
  wire              readCrossBar_input_4_valid;
  wire              readCrossBar_input_3_valid;
  wire              readCrossBar_input_2_valid;
  wire              readCrossBar_input_1_valid;
  wire              readCrossBar_input_0_valid;
  wire              _writeQueue_fifo_15_empty;
  wire              _writeQueue_fifo_15_full;
  wire              _writeQueue_fifo_15_error;
  wire [49:0]       _writeQueue_fifo_15_data_out;
  wire              _writeQueue_fifo_14_empty;
  wire              _writeQueue_fifo_14_full;
  wire              _writeQueue_fifo_14_error;
  wire [49:0]       _writeQueue_fifo_14_data_out;
  wire              _writeQueue_fifo_13_empty;
  wire              _writeQueue_fifo_13_full;
  wire              _writeQueue_fifo_13_error;
  wire [49:0]       _writeQueue_fifo_13_data_out;
  wire              _writeQueue_fifo_12_empty;
  wire              _writeQueue_fifo_12_full;
  wire              _writeQueue_fifo_12_error;
  wire [49:0]       _writeQueue_fifo_12_data_out;
  wire              _writeQueue_fifo_11_empty;
  wire              _writeQueue_fifo_11_full;
  wire              _writeQueue_fifo_11_error;
  wire [49:0]       _writeQueue_fifo_11_data_out;
  wire              _writeQueue_fifo_10_empty;
  wire              _writeQueue_fifo_10_full;
  wire              _writeQueue_fifo_10_error;
  wire [49:0]       _writeQueue_fifo_10_data_out;
  wire              _writeQueue_fifo_9_empty;
  wire              _writeQueue_fifo_9_full;
  wire              _writeQueue_fifo_9_error;
  wire [49:0]       _writeQueue_fifo_9_data_out;
  wire              _writeQueue_fifo_8_empty;
  wire              _writeQueue_fifo_8_full;
  wire              _writeQueue_fifo_8_error;
  wire [49:0]       _writeQueue_fifo_8_data_out;
  wire              _writeQueue_fifo_7_empty;
  wire              _writeQueue_fifo_7_full;
  wire              _writeQueue_fifo_7_error;
  wire [49:0]       _writeQueue_fifo_7_data_out;
  wire              _writeQueue_fifo_6_empty;
  wire              _writeQueue_fifo_6_full;
  wire              _writeQueue_fifo_6_error;
  wire [49:0]       _writeQueue_fifo_6_data_out;
  wire              _writeQueue_fifo_5_empty;
  wire              _writeQueue_fifo_5_full;
  wire              _writeQueue_fifo_5_error;
  wire [49:0]       _writeQueue_fifo_5_data_out;
  wire              _writeQueue_fifo_4_empty;
  wire              _writeQueue_fifo_4_full;
  wire              _writeQueue_fifo_4_error;
  wire [49:0]       _writeQueue_fifo_4_data_out;
  wire              _writeQueue_fifo_3_empty;
  wire              _writeQueue_fifo_3_full;
  wire              _writeQueue_fifo_3_error;
  wire [49:0]       _writeQueue_fifo_3_data_out;
  wire              _writeQueue_fifo_2_empty;
  wire              _writeQueue_fifo_2_full;
  wire              _writeQueue_fifo_2_error;
  wire [49:0]       _writeQueue_fifo_2_data_out;
  wire              _writeQueue_fifo_1_empty;
  wire              _writeQueue_fifo_1_full;
  wire              _writeQueue_fifo_1_error;
  wire [49:0]       _writeQueue_fifo_1_data_out;
  wire              _writeQueue_fifo_empty;
  wire              _writeQueue_fifo_full;
  wire              _writeQueue_fifo_error;
  wire [49:0]       _writeQueue_fifo_data_out;
  wire [511:0]      _extendUnit_out;
  wire              _reduceUnit_in_ready;
  wire              _reduceUnit_out_valid;
  wire [31:0]       _reduceUnit_out_bits_data;
  wire [3:0]        _reduceUnit_out_bits_mask;
  wire              _compressUnit_out_compressValid;
  wire [31:0]       _compressUnit_writeData;
  wire              _compressUnit_stageValid;
  wire              _readData_readDataQueue_fifo_15_empty;
  wire              _readData_readDataQueue_fifo_15_full;
  wire              _readData_readDataQueue_fifo_15_error;
  wire [31:0]       _readData_readDataQueue_fifo_15_data_out;
  wire              _readData_readDataQueue_fifo_14_empty;
  wire              _readData_readDataQueue_fifo_14_full;
  wire              _readData_readDataQueue_fifo_14_error;
  wire [31:0]       _readData_readDataQueue_fifo_14_data_out;
  wire              _readData_readDataQueue_fifo_13_empty;
  wire              _readData_readDataQueue_fifo_13_full;
  wire              _readData_readDataQueue_fifo_13_error;
  wire [31:0]       _readData_readDataQueue_fifo_13_data_out;
  wire              _readData_readDataQueue_fifo_12_empty;
  wire              _readData_readDataQueue_fifo_12_full;
  wire              _readData_readDataQueue_fifo_12_error;
  wire [31:0]       _readData_readDataQueue_fifo_12_data_out;
  wire              _readData_readDataQueue_fifo_11_empty;
  wire              _readData_readDataQueue_fifo_11_full;
  wire              _readData_readDataQueue_fifo_11_error;
  wire [31:0]       _readData_readDataQueue_fifo_11_data_out;
  wire              _readData_readDataQueue_fifo_10_empty;
  wire              _readData_readDataQueue_fifo_10_full;
  wire              _readData_readDataQueue_fifo_10_error;
  wire [31:0]       _readData_readDataQueue_fifo_10_data_out;
  wire              _readData_readDataQueue_fifo_9_empty;
  wire              _readData_readDataQueue_fifo_9_full;
  wire              _readData_readDataQueue_fifo_9_error;
  wire [31:0]       _readData_readDataQueue_fifo_9_data_out;
  wire              _readData_readDataQueue_fifo_8_empty;
  wire              _readData_readDataQueue_fifo_8_full;
  wire              _readData_readDataQueue_fifo_8_error;
  wire [31:0]       _readData_readDataQueue_fifo_8_data_out;
  wire              _readData_readDataQueue_fifo_7_empty;
  wire              _readData_readDataQueue_fifo_7_full;
  wire              _readData_readDataQueue_fifo_7_error;
  wire [31:0]       _readData_readDataQueue_fifo_7_data_out;
  wire              _readData_readDataQueue_fifo_6_empty;
  wire              _readData_readDataQueue_fifo_6_full;
  wire              _readData_readDataQueue_fifo_6_error;
  wire [31:0]       _readData_readDataQueue_fifo_6_data_out;
  wire              _readData_readDataQueue_fifo_5_empty;
  wire              _readData_readDataQueue_fifo_5_full;
  wire              _readData_readDataQueue_fifo_5_error;
  wire [31:0]       _readData_readDataQueue_fifo_5_data_out;
  wire              _readData_readDataQueue_fifo_4_empty;
  wire              _readData_readDataQueue_fifo_4_full;
  wire              _readData_readDataQueue_fifo_4_error;
  wire [31:0]       _readData_readDataQueue_fifo_4_data_out;
  wire              _readData_readDataQueue_fifo_3_empty;
  wire              _readData_readDataQueue_fifo_3_full;
  wire              _readData_readDataQueue_fifo_3_error;
  wire [31:0]       _readData_readDataQueue_fifo_3_data_out;
  wire              _readData_readDataQueue_fifo_2_empty;
  wire              _readData_readDataQueue_fifo_2_full;
  wire              _readData_readDataQueue_fifo_2_error;
  wire [31:0]       _readData_readDataQueue_fifo_2_data_out;
  wire              _readData_readDataQueue_fifo_1_empty;
  wire              _readData_readDataQueue_fifo_1_full;
  wire              _readData_readDataQueue_fifo_1_error;
  wire [31:0]       _readData_readDataQueue_fifo_1_data_out;
  wire              _readData_readDataQueue_fifo_empty;
  wire              _readData_readDataQueue_fifo_full;
  wire              _readData_readDataQueue_fifo_error;
  wire [31:0]       _readData_readDataQueue_fifo_data_out;
  wire              _readMessageQueue_fifo_15_empty;
  wire              _readMessageQueue_fifo_15_full;
  wire              _readMessageQueue_fifo_15_error;
  wire [17:0]       _readMessageQueue_fifo_15_data_out;
  wire              _readMessageQueue_fifo_14_empty;
  wire              _readMessageQueue_fifo_14_full;
  wire              _readMessageQueue_fifo_14_error;
  wire [17:0]       _readMessageQueue_fifo_14_data_out;
  wire              _readMessageQueue_fifo_13_empty;
  wire              _readMessageQueue_fifo_13_full;
  wire              _readMessageQueue_fifo_13_error;
  wire [17:0]       _readMessageQueue_fifo_13_data_out;
  wire              _readMessageQueue_fifo_12_empty;
  wire              _readMessageQueue_fifo_12_full;
  wire              _readMessageQueue_fifo_12_error;
  wire [17:0]       _readMessageQueue_fifo_12_data_out;
  wire              _readMessageQueue_fifo_11_empty;
  wire              _readMessageQueue_fifo_11_full;
  wire              _readMessageQueue_fifo_11_error;
  wire [17:0]       _readMessageQueue_fifo_11_data_out;
  wire              _readMessageQueue_fifo_10_empty;
  wire              _readMessageQueue_fifo_10_full;
  wire              _readMessageQueue_fifo_10_error;
  wire [17:0]       _readMessageQueue_fifo_10_data_out;
  wire              _readMessageQueue_fifo_9_empty;
  wire              _readMessageQueue_fifo_9_full;
  wire              _readMessageQueue_fifo_9_error;
  wire [17:0]       _readMessageQueue_fifo_9_data_out;
  wire              _readMessageQueue_fifo_8_empty;
  wire              _readMessageQueue_fifo_8_full;
  wire              _readMessageQueue_fifo_8_error;
  wire [17:0]       _readMessageQueue_fifo_8_data_out;
  wire              _readMessageQueue_fifo_7_empty;
  wire              _readMessageQueue_fifo_7_full;
  wire              _readMessageQueue_fifo_7_error;
  wire [17:0]       _readMessageQueue_fifo_7_data_out;
  wire              _readMessageQueue_fifo_6_empty;
  wire              _readMessageQueue_fifo_6_full;
  wire              _readMessageQueue_fifo_6_error;
  wire [17:0]       _readMessageQueue_fifo_6_data_out;
  wire              _readMessageQueue_fifo_5_empty;
  wire              _readMessageQueue_fifo_5_full;
  wire              _readMessageQueue_fifo_5_error;
  wire [17:0]       _readMessageQueue_fifo_5_data_out;
  wire              _readMessageQueue_fifo_4_empty;
  wire              _readMessageQueue_fifo_4_full;
  wire              _readMessageQueue_fifo_4_error;
  wire [17:0]       _readMessageQueue_fifo_4_data_out;
  wire              _readMessageQueue_fifo_3_empty;
  wire              _readMessageQueue_fifo_3_full;
  wire              _readMessageQueue_fifo_3_error;
  wire [17:0]       _readMessageQueue_fifo_3_data_out;
  wire              _readMessageQueue_fifo_2_empty;
  wire              _readMessageQueue_fifo_2_full;
  wire              _readMessageQueue_fifo_2_error;
  wire [17:0]       _readMessageQueue_fifo_2_data_out;
  wire              _readMessageQueue_fifo_1_empty;
  wire              _readMessageQueue_fifo_1_full;
  wire              _readMessageQueue_fifo_1_error;
  wire [17:0]       _readMessageQueue_fifo_1_data_out;
  wire              _readMessageQueue_fifo_empty;
  wire              _readMessageQueue_fifo_full;
  wire              _readMessageQueue_fifo_error;
  wire [17:0]       _readMessageQueue_fifo_data_out;
  wire              _reorderQueueVec_fifo_15_empty;
  wire              _reorderQueueVec_fifo_15_full;
  wire              _reorderQueueVec_fifo_15_error;
  wire [47:0]       _reorderQueueVec_fifo_15_data_out;
  wire              _reorderQueueVec_fifo_14_empty;
  wire              _reorderQueueVec_fifo_14_full;
  wire              _reorderQueueVec_fifo_14_error;
  wire [47:0]       _reorderQueueVec_fifo_14_data_out;
  wire              _reorderQueueVec_fifo_13_empty;
  wire              _reorderQueueVec_fifo_13_full;
  wire              _reorderQueueVec_fifo_13_error;
  wire [47:0]       _reorderQueueVec_fifo_13_data_out;
  wire              _reorderQueueVec_fifo_12_empty;
  wire              _reorderQueueVec_fifo_12_full;
  wire              _reorderQueueVec_fifo_12_error;
  wire [47:0]       _reorderQueueVec_fifo_12_data_out;
  wire              _reorderQueueVec_fifo_11_empty;
  wire              _reorderQueueVec_fifo_11_full;
  wire              _reorderQueueVec_fifo_11_error;
  wire [47:0]       _reorderQueueVec_fifo_11_data_out;
  wire              _reorderQueueVec_fifo_10_empty;
  wire              _reorderQueueVec_fifo_10_full;
  wire              _reorderQueueVec_fifo_10_error;
  wire [47:0]       _reorderQueueVec_fifo_10_data_out;
  wire              _reorderQueueVec_fifo_9_empty;
  wire              _reorderQueueVec_fifo_9_full;
  wire              _reorderQueueVec_fifo_9_error;
  wire [47:0]       _reorderQueueVec_fifo_9_data_out;
  wire              _reorderQueueVec_fifo_8_empty;
  wire              _reorderQueueVec_fifo_8_full;
  wire              _reorderQueueVec_fifo_8_error;
  wire [47:0]       _reorderQueueVec_fifo_8_data_out;
  wire              _reorderQueueVec_fifo_7_empty;
  wire              _reorderQueueVec_fifo_7_full;
  wire              _reorderQueueVec_fifo_7_error;
  wire [47:0]       _reorderQueueVec_fifo_7_data_out;
  wire              _reorderQueueVec_fifo_6_empty;
  wire              _reorderQueueVec_fifo_6_full;
  wire              _reorderQueueVec_fifo_6_error;
  wire [47:0]       _reorderQueueVec_fifo_6_data_out;
  wire              _reorderQueueVec_fifo_5_empty;
  wire              _reorderQueueVec_fifo_5_full;
  wire              _reorderQueueVec_fifo_5_error;
  wire [47:0]       _reorderQueueVec_fifo_5_data_out;
  wire              _reorderQueueVec_fifo_4_empty;
  wire              _reorderQueueVec_fifo_4_full;
  wire              _reorderQueueVec_fifo_4_error;
  wire [47:0]       _reorderQueueVec_fifo_4_data_out;
  wire              _reorderQueueVec_fifo_3_empty;
  wire              _reorderQueueVec_fifo_3_full;
  wire              _reorderQueueVec_fifo_3_error;
  wire [47:0]       _reorderQueueVec_fifo_3_data_out;
  wire              _reorderQueueVec_fifo_2_empty;
  wire              _reorderQueueVec_fifo_2_full;
  wire              _reorderQueueVec_fifo_2_error;
  wire [47:0]       _reorderQueueVec_fifo_2_data_out;
  wire              _reorderQueueVec_fifo_1_empty;
  wire              _reorderQueueVec_fifo_1_full;
  wire              _reorderQueueVec_fifo_1_error;
  wire [47:0]       _reorderQueueVec_fifo_1_data_out;
  wire              _reorderQueueVec_fifo_empty;
  wire              _reorderQueueVec_fifo_full;
  wire              _reorderQueueVec_fifo_error;
  wire [47:0]       _reorderQueueVec_fifo_data_out;
  wire              _compressUnitResultQueue_fifo_empty;
  wire              _compressUnitResultQueue_fifo_full;
  wire              _compressUnitResultQueue_fifo_error;
  wire [597:0]      _compressUnitResultQueue_fifo_data_out;
  wire              _readWaitQueue_fifo_empty;
  wire              _readWaitQueue_fifo_full;
  wire              _readWaitQueue_fifo_error;
  wire [55:0]       _readWaitQueue_fifo_data_out;
  wire              _readCrossBar_input_0_ready;
  wire              _readCrossBar_input_1_ready;
  wire              _readCrossBar_input_2_ready;
  wire              _readCrossBar_input_3_ready;
  wire              _readCrossBar_input_4_ready;
  wire              _readCrossBar_input_5_ready;
  wire              _readCrossBar_input_6_ready;
  wire              _readCrossBar_input_7_ready;
  wire              _readCrossBar_input_8_ready;
  wire              _readCrossBar_input_9_ready;
  wire              _readCrossBar_input_10_ready;
  wire              _readCrossBar_input_11_ready;
  wire              _readCrossBar_input_12_ready;
  wire              _readCrossBar_input_13_ready;
  wire              _readCrossBar_input_14_ready;
  wire              _readCrossBar_input_15_ready;
  wire              _readCrossBar_output_0_valid;
  wire [4:0]        _readCrossBar_output_0_bits_vs;
  wire              _readCrossBar_output_0_bits_offset;
  wire [3:0]        _readCrossBar_output_0_bits_writeIndex;
  wire              _readCrossBar_output_1_valid;
  wire [4:0]        _readCrossBar_output_1_bits_vs;
  wire              _readCrossBar_output_1_bits_offset;
  wire [3:0]        _readCrossBar_output_1_bits_writeIndex;
  wire              _readCrossBar_output_2_valid;
  wire [4:0]        _readCrossBar_output_2_bits_vs;
  wire              _readCrossBar_output_2_bits_offset;
  wire [3:0]        _readCrossBar_output_2_bits_writeIndex;
  wire              _readCrossBar_output_3_valid;
  wire [4:0]        _readCrossBar_output_3_bits_vs;
  wire              _readCrossBar_output_3_bits_offset;
  wire [3:0]        _readCrossBar_output_3_bits_writeIndex;
  wire              _readCrossBar_output_4_valid;
  wire [4:0]        _readCrossBar_output_4_bits_vs;
  wire              _readCrossBar_output_4_bits_offset;
  wire [3:0]        _readCrossBar_output_4_bits_writeIndex;
  wire              _readCrossBar_output_5_valid;
  wire [4:0]        _readCrossBar_output_5_bits_vs;
  wire              _readCrossBar_output_5_bits_offset;
  wire [3:0]        _readCrossBar_output_5_bits_writeIndex;
  wire              _readCrossBar_output_6_valid;
  wire [4:0]        _readCrossBar_output_6_bits_vs;
  wire              _readCrossBar_output_6_bits_offset;
  wire [3:0]        _readCrossBar_output_6_bits_writeIndex;
  wire              _readCrossBar_output_7_valid;
  wire [4:0]        _readCrossBar_output_7_bits_vs;
  wire              _readCrossBar_output_7_bits_offset;
  wire [3:0]        _readCrossBar_output_7_bits_writeIndex;
  wire              _readCrossBar_output_8_valid;
  wire [4:0]        _readCrossBar_output_8_bits_vs;
  wire              _readCrossBar_output_8_bits_offset;
  wire [3:0]        _readCrossBar_output_8_bits_writeIndex;
  wire              _readCrossBar_output_9_valid;
  wire [4:0]        _readCrossBar_output_9_bits_vs;
  wire              _readCrossBar_output_9_bits_offset;
  wire [3:0]        _readCrossBar_output_9_bits_writeIndex;
  wire              _readCrossBar_output_10_valid;
  wire [4:0]        _readCrossBar_output_10_bits_vs;
  wire              _readCrossBar_output_10_bits_offset;
  wire [3:0]        _readCrossBar_output_10_bits_writeIndex;
  wire              _readCrossBar_output_11_valid;
  wire [4:0]        _readCrossBar_output_11_bits_vs;
  wire              _readCrossBar_output_11_bits_offset;
  wire [3:0]        _readCrossBar_output_11_bits_writeIndex;
  wire              _readCrossBar_output_12_valid;
  wire [4:0]        _readCrossBar_output_12_bits_vs;
  wire              _readCrossBar_output_12_bits_offset;
  wire [3:0]        _readCrossBar_output_12_bits_writeIndex;
  wire              _readCrossBar_output_13_valid;
  wire [4:0]        _readCrossBar_output_13_bits_vs;
  wire              _readCrossBar_output_13_bits_offset;
  wire [3:0]        _readCrossBar_output_13_bits_writeIndex;
  wire              _readCrossBar_output_14_valid;
  wire [4:0]        _readCrossBar_output_14_bits_vs;
  wire              _readCrossBar_output_14_bits_offset;
  wire [3:0]        _readCrossBar_output_14_bits_writeIndex;
  wire              _readCrossBar_output_15_valid;
  wire [4:0]        _readCrossBar_output_15_bits_vs;
  wire              _readCrossBar_output_15_bits_offset;
  wire [3:0]        _readCrossBar_output_15_bits_writeIndex;
  wire              _accessCountQueue_fifo_empty;
  wire              _accessCountQueue_fifo_full;
  wire              _accessCountQueue_fifo_error;
  wire [79:0]       _accessCountQueue_fifo_data_out;
  wire              _slideAddressGen_indexDeq_valid;
  wire [15:0]       _slideAddressGen_indexDeq_bits_needRead;
  wire [15:0]       _slideAddressGen_indexDeq_bits_elementValid;
  wire [15:0]       _slideAddressGen_indexDeq_bits_replaceVs1;
  wire [15:0]       _slideAddressGen_indexDeq_bits_readOffset;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_0;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_1;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_2;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_3;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_4;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_5;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_6;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_7;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_8;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_9;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_10;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_11;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_12;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_13;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_14;
  wire [3:0]        _slideAddressGen_indexDeq_bits_accessLane_15;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_0;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_1;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_2;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_3;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_4;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_5;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_6;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_7;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_8;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_9;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_10;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_11;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_12;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_13;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_14;
  wire [2:0]        _slideAddressGen_indexDeq_bits_vsGrowth_15;
  wire [6:0]        _slideAddressGen_indexDeq_bits_executeGroup;
  wire [31:0]       _slideAddressGen_indexDeq_bits_readDataOffset;
  wire              _slideAddressGen_indexDeq_bits_last;
  wire [6:0]        _slideAddressGen_slideGroupOut;
  wire              _exeRequestQueue_queue_fifo_15_empty;
  wire              _exeRequestQueue_queue_fifo_15_full;
  wire              _exeRequestQueue_queue_fifo_15_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_15_data_out;
  wire              _exeRequestQueue_queue_fifo_14_empty;
  wire              _exeRequestQueue_queue_fifo_14_full;
  wire              _exeRequestQueue_queue_fifo_14_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_14_data_out;
  wire              _exeRequestQueue_queue_fifo_13_empty;
  wire              _exeRequestQueue_queue_fifo_13_full;
  wire              _exeRequestQueue_queue_fifo_13_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_13_data_out;
  wire              _exeRequestQueue_queue_fifo_12_empty;
  wire              _exeRequestQueue_queue_fifo_12_full;
  wire              _exeRequestQueue_queue_fifo_12_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_12_data_out;
  wire              _exeRequestQueue_queue_fifo_11_empty;
  wire              _exeRequestQueue_queue_fifo_11_full;
  wire              _exeRequestQueue_queue_fifo_11_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_11_data_out;
  wire              _exeRequestQueue_queue_fifo_10_empty;
  wire              _exeRequestQueue_queue_fifo_10_full;
  wire              _exeRequestQueue_queue_fifo_10_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_10_data_out;
  wire              _exeRequestQueue_queue_fifo_9_empty;
  wire              _exeRequestQueue_queue_fifo_9_full;
  wire              _exeRequestQueue_queue_fifo_9_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_9_data_out;
  wire              _exeRequestQueue_queue_fifo_8_empty;
  wire              _exeRequestQueue_queue_fifo_8_full;
  wire              _exeRequestQueue_queue_fifo_8_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_8_data_out;
  wire              _exeRequestQueue_queue_fifo_7_empty;
  wire              _exeRequestQueue_queue_fifo_7_full;
  wire              _exeRequestQueue_queue_fifo_7_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_7_data_out;
  wire              _exeRequestQueue_queue_fifo_6_empty;
  wire              _exeRequestQueue_queue_fifo_6_full;
  wire              _exeRequestQueue_queue_fifo_6_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_6_data_out;
  wire              _exeRequestQueue_queue_fifo_5_empty;
  wire              _exeRequestQueue_queue_fifo_5_full;
  wire              _exeRequestQueue_queue_fifo_5_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_5_data_out;
  wire              _exeRequestQueue_queue_fifo_4_empty;
  wire              _exeRequestQueue_queue_fifo_4_full;
  wire              _exeRequestQueue_queue_fifo_4_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_4_data_out;
  wire              _exeRequestQueue_queue_fifo_3_empty;
  wire              _exeRequestQueue_queue_fifo_3_full;
  wire              _exeRequestQueue_queue_fifo_3_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_3_data_out;
  wire              _exeRequestQueue_queue_fifo_2_empty;
  wire              _exeRequestQueue_queue_fifo_2_full;
  wire              _exeRequestQueue_queue_fifo_2_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_2_data_out;
  wire              _exeRequestQueue_queue_fifo_1_empty;
  wire              _exeRequestQueue_queue_fifo_1_full;
  wire              _exeRequestQueue_queue_fifo_1_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_1_data_out;
  wire              _exeRequestQueue_queue_fifo_empty;
  wire              _exeRequestQueue_queue_fifo_full;
  wire              _exeRequestQueue_queue_fifo_error;
  wire [68:0]       _exeRequestQueue_queue_fifo_data_out;
  wire              _maskedWrite_in_0_ready;
  wire              _maskedWrite_in_1_ready;
  wire              _maskedWrite_in_2_ready;
  wire              _maskedWrite_in_3_ready;
  wire              _maskedWrite_in_4_ready;
  wire              _maskedWrite_in_5_ready;
  wire              _maskedWrite_in_6_ready;
  wire              _maskedWrite_in_7_ready;
  wire              _maskedWrite_in_8_ready;
  wire              _maskedWrite_in_9_ready;
  wire              _maskedWrite_in_10_ready;
  wire              _maskedWrite_in_11_ready;
  wire              _maskedWrite_in_12_ready;
  wire              _maskedWrite_in_13_ready;
  wire              _maskedWrite_in_14_ready;
  wire              _maskedWrite_in_15_ready;
  wire              _maskedWrite_out_0_valid;
  wire              _maskedWrite_out_0_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_0_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_0_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_0_bits_writeData_groupCounter;
  wire              _maskedWrite_out_1_valid;
  wire              _maskedWrite_out_1_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_1_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_1_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_1_bits_writeData_groupCounter;
  wire              _maskedWrite_out_2_valid;
  wire              _maskedWrite_out_2_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_2_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_2_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_2_bits_writeData_groupCounter;
  wire              _maskedWrite_out_3_valid;
  wire              _maskedWrite_out_3_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_3_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_3_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_3_bits_writeData_groupCounter;
  wire              _maskedWrite_out_4_valid;
  wire              _maskedWrite_out_4_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_4_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_4_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_4_bits_writeData_groupCounter;
  wire              _maskedWrite_out_5_valid;
  wire              _maskedWrite_out_5_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_5_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_5_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_5_bits_writeData_groupCounter;
  wire              _maskedWrite_out_6_valid;
  wire              _maskedWrite_out_6_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_6_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_6_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_6_bits_writeData_groupCounter;
  wire              _maskedWrite_out_7_valid;
  wire              _maskedWrite_out_7_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_7_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_7_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_7_bits_writeData_groupCounter;
  wire              _maskedWrite_out_8_valid;
  wire              _maskedWrite_out_8_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_8_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_8_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_8_bits_writeData_groupCounter;
  wire              _maskedWrite_out_9_valid;
  wire              _maskedWrite_out_9_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_9_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_9_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_9_bits_writeData_groupCounter;
  wire              _maskedWrite_out_10_valid;
  wire              _maskedWrite_out_10_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_10_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_10_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_10_bits_writeData_groupCounter;
  wire              _maskedWrite_out_11_valid;
  wire              _maskedWrite_out_11_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_11_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_11_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_11_bits_writeData_groupCounter;
  wire              _maskedWrite_out_12_valid;
  wire              _maskedWrite_out_12_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_12_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_12_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_12_bits_writeData_groupCounter;
  wire              _maskedWrite_out_13_valid;
  wire              _maskedWrite_out_13_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_13_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_13_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_13_bits_writeData_groupCounter;
  wire              _maskedWrite_out_14_valid;
  wire              _maskedWrite_out_14_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_14_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_14_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_14_bits_writeData_groupCounter;
  wire              _maskedWrite_out_15_valid;
  wire              _maskedWrite_out_15_bits_ffoByOther;
  wire [31:0]       _maskedWrite_out_15_bits_writeData_data;
  wire [3:0]        _maskedWrite_out_15_bits_writeData_mask;
  wire [4:0]        _maskedWrite_out_15_bits_writeData_groupCounter;
  wire              _maskedWrite_readChannel_0_valid;
  wire [4:0]        _maskedWrite_readChannel_0_bits_vs;
  wire              _maskedWrite_readChannel_0_bits_offset;
  wire              _maskedWrite_readChannel_1_valid;
  wire [4:0]        _maskedWrite_readChannel_1_bits_vs;
  wire              _maskedWrite_readChannel_1_bits_offset;
  wire              _maskedWrite_readChannel_2_valid;
  wire [4:0]        _maskedWrite_readChannel_2_bits_vs;
  wire              _maskedWrite_readChannel_2_bits_offset;
  wire              _maskedWrite_readChannel_3_valid;
  wire [4:0]        _maskedWrite_readChannel_3_bits_vs;
  wire              _maskedWrite_readChannel_3_bits_offset;
  wire              _maskedWrite_readChannel_4_valid;
  wire [4:0]        _maskedWrite_readChannel_4_bits_vs;
  wire              _maskedWrite_readChannel_4_bits_offset;
  wire              _maskedWrite_readChannel_5_valid;
  wire [4:0]        _maskedWrite_readChannel_5_bits_vs;
  wire              _maskedWrite_readChannel_5_bits_offset;
  wire              _maskedWrite_readChannel_6_valid;
  wire [4:0]        _maskedWrite_readChannel_6_bits_vs;
  wire              _maskedWrite_readChannel_6_bits_offset;
  wire              _maskedWrite_readChannel_7_valid;
  wire [4:0]        _maskedWrite_readChannel_7_bits_vs;
  wire              _maskedWrite_readChannel_7_bits_offset;
  wire              _maskedWrite_readChannel_8_valid;
  wire [4:0]        _maskedWrite_readChannel_8_bits_vs;
  wire              _maskedWrite_readChannel_8_bits_offset;
  wire              _maskedWrite_readChannel_9_valid;
  wire [4:0]        _maskedWrite_readChannel_9_bits_vs;
  wire              _maskedWrite_readChannel_9_bits_offset;
  wire              _maskedWrite_readChannel_10_valid;
  wire [4:0]        _maskedWrite_readChannel_10_bits_vs;
  wire              _maskedWrite_readChannel_10_bits_offset;
  wire              _maskedWrite_readChannel_11_valid;
  wire [4:0]        _maskedWrite_readChannel_11_bits_vs;
  wire              _maskedWrite_readChannel_11_bits_offset;
  wire              _maskedWrite_readChannel_12_valid;
  wire [4:0]        _maskedWrite_readChannel_12_bits_vs;
  wire              _maskedWrite_readChannel_12_bits_offset;
  wire              _maskedWrite_readChannel_13_valid;
  wire [4:0]        _maskedWrite_readChannel_13_bits_vs;
  wire              _maskedWrite_readChannel_13_bits_offset;
  wire              _maskedWrite_readChannel_14_valid;
  wire [4:0]        _maskedWrite_readChannel_14_bits_vs;
  wire              _maskedWrite_readChannel_14_bits_offset;
  wire              _maskedWrite_readChannel_15_valid;
  wire [4:0]        _maskedWrite_readChannel_15_bits_vs;
  wire              _maskedWrite_readChannel_15_bits_offset;
  wire              _maskedWrite_stageClear;
  wire              writeQueue_15_almostFull;
  wire              writeQueue_15_almostEmpty;
  wire              writeQueue_14_almostFull;
  wire              writeQueue_14_almostEmpty;
  wire              writeQueue_13_almostFull;
  wire              writeQueue_13_almostEmpty;
  wire              writeQueue_12_almostFull;
  wire              writeQueue_12_almostEmpty;
  wire              writeQueue_11_almostFull;
  wire              writeQueue_11_almostEmpty;
  wire              writeQueue_10_almostFull;
  wire              writeQueue_10_almostEmpty;
  wire              writeQueue_9_almostFull;
  wire              writeQueue_9_almostEmpty;
  wire              writeQueue_8_almostFull;
  wire              writeQueue_8_almostEmpty;
  wire              writeQueue_7_almostFull;
  wire              writeQueue_7_almostEmpty;
  wire              writeQueue_6_almostFull;
  wire              writeQueue_6_almostEmpty;
  wire              writeQueue_5_almostFull;
  wire              writeQueue_5_almostEmpty;
  wire              writeQueue_4_almostFull;
  wire              writeQueue_4_almostEmpty;
  wire              writeQueue_3_almostFull;
  wire              writeQueue_3_almostEmpty;
  wire              writeQueue_2_almostFull;
  wire              writeQueue_2_almostEmpty;
  wire              writeQueue_1_almostFull;
  wire              writeQueue_1_almostEmpty;
  wire              writeQueue_0_almostFull;
  wire              writeQueue_0_almostEmpty;
  wire              readData_readDataQueue_15_almostFull;
  wire              readData_readDataQueue_15_almostEmpty;
  wire              readData_readDataQueue_14_almostFull;
  wire              readData_readDataQueue_14_almostEmpty;
  wire              readData_readDataQueue_13_almostFull;
  wire              readData_readDataQueue_13_almostEmpty;
  wire              readData_readDataQueue_12_almostFull;
  wire              readData_readDataQueue_12_almostEmpty;
  wire              readData_readDataQueue_11_almostFull;
  wire              readData_readDataQueue_11_almostEmpty;
  wire              readData_readDataQueue_10_almostFull;
  wire              readData_readDataQueue_10_almostEmpty;
  wire              readData_readDataQueue_9_almostFull;
  wire              readData_readDataQueue_9_almostEmpty;
  wire              readData_readDataQueue_8_almostFull;
  wire              readData_readDataQueue_8_almostEmpty;
  wire              readData_readDataQueue_7_almostFull;
  wire              readData_readDataQueue_7_almostEmpty;
  wire              readData_readDataQueue_6_almostFull;
  wire              readData_readDataQueue_6_almostEmpty;
  wire              readData_readDataQueue_5_almostFull;
  wire              readData_readDataQueue_5_almostEmpty;
  wire              readData_readDataQueue_4_almostFull;
  wire              readData_readDataQueue_4_almostEmpty;
  wire              readData_readDataQueue_3_almostFull;
  wire              readData_readDataQueue_3_almostEmpty;
  wire              readData_readDataQueue_2_almostFull;
  wire              readData_readDataQueue_2_almostEmpty;
  wire              readData_readDataQueue_1_almostFull;
  wire              readData_readDataQueue_1_almostEmpty;
  wire              readData_readDataQueue_almostFull;
  wire              readData_readDataQueue_almostEmpty;
  wire              readMessageQueue_15_almostFull;
  wire              readMessageQueue_15_almostEmpty;
  wire              readMessageQueue_14_almostFull;
  wire              readMessageQueue_14_almostEmpty;
  wire              readMessageQueue_13_almostFull;
  wire              readMessageQueue_13_almostEmpty;
  wire              readMessageQueue_12_almostFull;
  wire              readMessageQueue_12_almostEmpty;
  wire              readMessageQueue_11_almostFull;
  wire              readMessageQueue_11_almostEmpty;
  wire              readMessageQueue_10_almostFull;
  wire              readMessageQueue_10_almostEmpty;
  wire              readMessageQueue_9_almostFull;
  wire              readMessageQueue_9_almostEmpty;
  wire              readMessageQueue_8_almostFull;
  wire              readMessageQueue_8_almostEmpty;
  wire              readMessageQueue_7_almostFull;
  wire              readMessageQueue_7_almostEmpty;
  wire              readMessageQueue_6_almostFull;
  wire              readMessageQueue_6_almostEmpty;
  wire              readMessageQueue_5_almostFull;
  wire              readMessageQueue_5_almostEmpty;
  wire              readMessageQueue_4_almostFull;
  wire              readMessageQueue_4_almostEmpty;
  wire              readMessageQueue_3_almostFull;
  wire              readMessageQueue_3_almostEmpty;
  wire              readMessageQueue_2_almostFull;
  wire              readMessageQueue_2_almostEmpty;
  wire              readMessageQueue_1_almostFull;
  wire              readMessageQueue_1_almostEmpty;
  wire              readMessageQueue_almostFull;
  wire              readMessageQueue_almostEmpty;
  wire              reorderQueueVec_15_almostFull;
  wire              reorderQueueVec_15_almostEmpty;
  wire              reorderQueueVec_14_almostFull;
  wire              reorderQueueVec_14_almostEmpty;
  wire              reorderQueueVec_13_almostFull;
  wire              reorderQueueVec_13_almostEmpty;
  wire              reorderQueueVec_12_almostFull;
  wire              reorderQueueVec_12_almostEmpty;
  wire              reorderQueueVec_11_almostFull;
  wire              reorderQueueVec_11_almostEmpty;
  wire              reorderQueueVec_10_almostFull;
  wire              reorderQueueVec_10_almostEmpty;
  wire              reorderQueueVec_9_almostFull;
  wire              reorderQueueVec_9_almostEmpty;
  wire              reorderQueueVec_8_almostFull;
  wire              reorderQueueVec_8_almostEmpty;
  wire              reorderQueueVec_7_almostFull;
  wire              reorderQueueVec_7_almostEmpty;
  wire              reorderQueueVec_6_almostFull;
  wire              reorderQueueVec_6_almostEmpty;
  wire              reorderQueueVec_5_almostFull;
  wire              reorderQueueVec_5_almostEmpty;
  wire              reorderQueueVec_4_almostFull;
  wire              reorderQueueVec_4_almostEmpty;
  wire              reorderQueueVec_3_almostFull;
  wire              reorderQueueVec_3_almostEmpty;
  wire              reorderQueueVec_2_almostFull;
  wire              reorderQueueVec_2_almostEmpty;
  wire              reorderQueueVec_1_almostFull;
  wire              reorderQueueVec_1_almostEmpty;
  wire              reorderQueueVec_0_almostFull;
  wire              reorderQueueVec_0_almostEmpty;
  wire              compressUnitResultQueue_almostFull;
  wire              compressUnitResultQueue_almostEmpty;
  wire              readWaitQueue_almostFull;
  wire              readWaitQueue_almostEmpty;
  wire              accessCountQueue_almostFull;
  wire              accessCountQueue_almostEmpty;
  wire              exeRequestQueue_15_almostFull;
  wire              exeRequestQueue_15_almostEmpty;
  wire              exeRequestQueue_14_almostFull;
  wire              exeRequestQueue_14_almostEmpty;
  wire              exeRequestQueue_13_almostFull;
  wire              exeRequestQueue_13_almostEmpty;
  wire              exeRequestQueue_12_almostFull;
  wire              exeRequestQueue_12_almostEmpty;
  wire              exeRequestQueue_11_almostFull;
  wire              exeRequestQueue_11_almostEmpty;
  wire              exeRequestQueue_10_almostFull;
  wire              exeRequestQueue_10_almostEmpty;
  wire              exeRequestQueue_9_almostFull;
  wire              exeRequestQueue_9_almostEmpty;
  wire              exeRequestQueue_8_almostFull;
  wire              exeRequestQueue_8_almostEmpty;
  wire              exeRequestQueue_7_almostFull;
  wire              exeRequestQueue_7_almostEmpty;
  wire              exeRequestQueue_6_almostFull;
  wire              exeRequestQueue_6_almostEmpty;
  wire              exeRequestQueue_5_almostFull;
  wire              exeRequestQueue_5_almostEmpty;
  wire              exeRequestQueue_4_almostFull;
  wire              exeRequestQueue_4_almostEmpty;
  wire              exeRequestQueue_3_almostFull;
  wire              exeRequestQueue_3_almostEmpty;
  wire              exeRequestQueue_2_almostFull;
  wire              exeRequestQueue_2_almostEmpty;
  wire              exeRequestQueue_1_almostFull;
  wire              exeRequestQueue_1_almostEmpty;
  wire              exeRequestQueue_0_almostFull;
  wire              exeRequestQueue_0_almostEmpty;
  wire [31:0]       reorderQueueVec_15_deq_bits_data;
  wire [31:0]       reorderQueueVec_14_deq_bits_data;
  wire [31:0]       reorderQueueVec_13_deq_bits_data;
  wire [31:0]       reorderQueueVec_12_deq_bits_data;
  wire [31:0]       reorderQueueVec_11_deq_bits_data;
  wire [31:0]       reorderQueueVec_10_deq_bits_data;
  wire [31:0]       reorderQueueVec_9_deq_bits_data;
  wire [31:0]       reorderQueueVec_8_deq_bits_data;
  wire [31:0]       reorderQueueVec_7_deq_bits_data;
  wire [31:0]       reorderQueueVec_6_deq_bits_data;
  wire [31:0]       reorderQueueVec_5_deq_bits_data;
  wire [31:0]       reorderQueueVec_4_deq_bits_data;
  wire [31:0]       reorderQueueVec_3_deq_bits_data;
  wire [31:0]       reorderQueueVec_2_deq_bits_data;
  wire [31:0]       reorderQueueVec_1_deq_bits_data;
  wire [31:0]       reorderQueueVec_0_deq_bits_data;
  wire [4:0]        accessCountEnq_15;
  wire [4:0]        accessCountEnq_14;
  wire [4:0]        accessCountEnq_13;
  wire [4:0]        accessCountEnq_12;
  wire [4:0]        accessCountEnq_11;
  wire [4:0]        accessCountEnq_10;
  wire [4:0]        accessCountEnq_9;
  wire [4:0]        accessCountEnq_8;
  wire [4:0]        accessCountEnq_7;
  wire [4:0]        accessCountEnq_6;
  wire [4:0]        accessCountEnq_5;
  wire [4:0]        accessCountEnq_4;
  wire [4:0]        accessCountEnq_3;
  wire [4:0]        accessCountEnq_2;
  wire [4:0]        accessCountEnq_1;
  wire [4:0]        accessCountEnq_0;
  wire              exeResp_0_ready_0 = exeResp_0_ready;
  wire              exeResp_1_ready_0 = exeResp_1_ready;
  wire              exeResp_2_ready_0 = exeResp_2_ready;
  wire              exeResp_3_ready_0 = exeResp_3_ready;
  wire              exeResp_4_ready_0 = exeResp_4_ready;
  wire              exeResp_5_ready_0 = exeResp_5_ready;
  wire              exeResp_6_ready_0 = exeResp_6_ready;
  wire              exeResp_7_ready_0 = exeResp_7_ready;
  wire              exeResp_8_ready_0 = exeResp_8_ready;
  wire              exeResp_9_ready_0 = exeResp_9_ready;
  wire              exeResp_10_ready_0 = exeResp_10_ready;
  wire              exeResp_11_ready_0 = exeResp_11_ready;
  wire              exeResp_12_ready_0 = exeResp_12_ready;
  wire              exeResp_13_ready_0 = exeResp_13_ready;
  wire              exeResp_14_ready_0 = exeResp_14_ready;
  wire              exeResp_15_ready_0 = exeResp_15_ready;
  wire              readChannel_0_ready_0 = readChannel_0_ready;
  wire              readChannel_1_ready_0 = readChannel_1_ready;
  wire              readChannel_2_ready_0 = readChannel_2_ready;
  wire              readChannel_3_ready_0 = readChannel_3_ready;
  wire              readChannel_4_ready_0 = readChannel_4_ready;
  wire              readChannel_5_ready_0 = readChannel_5_ready;
  wire              readChannel_6_ready_0 = readChannel_6_ready;
  wire              readChannel_7_ready_0 = readChannel_7_ready;
  wire              readChannel_8_ready_0 = readChannel_8_ready;
  wire              readChannel_9_ready_0 = readChannel_9_ready;
  wire              readChannel_10_ready_0 = readChannel_10_ready;
  wire              readChannel_11_ready_0 = readChannel_11_ready;
  wire              readChannel_12_ready_0 = readChannel_12_ready;
  wire              readChannel_13_ready_0 = readChannel_13_ready;
  wire              readChannel_14_ready_0 = readChannel_14_ready;
  wire              readChannel_15_ready_0 = readChannel_15_ready;
  wire              gatherData_ready_0 = gatherData_ready;
  wire              exeRequestQueue_0_enq_valid = exeReq_0_valid;
  wire [31:0]       exeRequestQueue_0_enq_bits_source1 = exeReq_0_bits_source1;
  wire [31:0]       exeRequestQueue_0_enq_bits_source2 = exeReq_0_bits_source2;
  wire [2:0]        exeRequestQueue_0_enq_bits_index = exeReq_0_bits_index;
  wire              exeRequestQueue_0_enq_bits_ffo = exeReq_0_bits_ffo;
  wire              exeRequestQueue_0_enq_bits_fpReduceValid = exeReq_0_bits_fpReduceValid;
  wire              exeRequestQueue_1_enq_valid = exeReq_1_valid;
  wire [31:0]       exeRequestQueue_1_enq_bits_source1 = exeReq_1_bits_source1;
  wire [31:0]       exeRequestQueue_1_enq_bits_source2 = exeReq_1_bits_source2;
  wire [2:0]        exeRequestQueue_1_enq_bits_index = exeReq_1_bits_index;
  wire              exeRequestQueue_1_enq_bits_ffo = exeReq_1_bits_ffo;
  wire              exeRequestQueue_1_enq_bits_fpReduceValid = exeReq_1_bits_fpReduceValid;
  wire              exeRequestQueue_2_enq_valid = exeReq_2_valid;
  wire [31:0]       exeRequestQueue_2_enq_bits_source1 = exeReq_2_bits_source1;
  wire [31:0]       exeRequestQueue_2_enq_bits_source2 = exeReq_2_bits_source2;
  wire [2:0]        exeRequestQueue_2_enq_bits_index = exeReq_2_bits_index;
  wire              exeRequestQueue_2_enq_bits_ffo = exeReq_2_bits_ffo;
  wire              exeRequestQueue_2_enq_bits_fpReduceValid = exeReq_2_bits_fpReduceValid;
  wire              exeRequestQueue_3_enq_valid = exeReq_3_valid;
  wire [31:0]       exeRequestQueue_3_enq_bits_source1 = exeReq_3_bits_source1;
  wire [31:0]       exeRequestQueue_3_enq_bits_source2 = exeReq_3_bits_source2;
  wire [2:0]        exeRequestQueue_3_enq_bits_index = exeReq_3_bits_index;
  wire              exeRequestQueue_3_enq_bits_ffo = exeReq_3_bits_ffo;
  wire              exeRequestQueue_3_enq_bits_fpReduceValid = exeReq_3_bits_fpReduceValid;
  wire              exeRequestQueue_4_enq_valid = exeReq_4_valid;
  wire [31:0]       exeRequestQueue_4_enq_bits_source1 = exeReq_4_bits_source1;
  wire [31:0]       exeRequestQueue_4_enq_bits_source2 = exeReq_4_bits_source2;
  wire [2:0]        exeRequestQueue_4_enq_bits_index = exeReq_4_bits_index;
  wire              exeRequestQueue_4_enq_bits_ffo = exeReq_4_bits_ffo;
  wire              exeRequestQueue_4_enq_bits_fpReduceValid = exeReq_4_bits_fpReduceValid;
  wire              exeRequestQueue_5_enq_valid = exeReq_5_valid;
  wire [31:0]       exeRequestQueue_5_enq_bits_source1 = exeReq_5_bits_source1;
  wire [31:0]       exeRequestQueue_5_enq_bits_source2 = exeReq_5_bits_source2;
  wire [2:0]        exeRequestQueue_5_enq_bits_index = exeReq_5_bits_index;
  wire              exeRequestQueue_5_enq_bits_ffo = exeReq_5_bits_ffo;
  wire              exeRequestQueue_5_enq_bits_fpReduceValid = exeReq_5_bits_fpReduceValid;
  wire              exeRequestQueue_6_enq_valid = exeReq_6_valid;
  wire [31:0]       exeRequestQueue_6_enq_bits_source1 = exeReq_6_bits_source1;
  wire [31:0]       exeRequestQueue_6_enq_bits_source2 = exeReq_6_bits_source2;
  wire [2:0]        exeRequestQueue_6_enq_bits_index = exeReq_6_bits_index;
  wire              exeRequestQueue_6_enq_bits_ffo = exeReq_6_bits_ffo;
  wire              exeRequestQueue_6_enq_bits_fpReduceValid = exeReq_6_bits_fpReduceValid;
  wire              exeRequestQueue_7_enq_valid = exeReq_7_valid;
  wire [31:0]       exeRequestQueue_7_enq_bits_source1 = exeReq_7_bits_source1;
  wire [31:0]       exeRequestQueue_7_enq_bits_source2 = exeReq_7_bits_source2;
  wire [2:0]        exeRequestQueue_7_enq_bits_index = exeReq_7_bits_index;
  wire              exeRequestQueue_7_enq_bits_ffo = exeReq_7_bits_ffo;
  wire              exeRequestQueue_7_enq_bits_fpReduceValid = exeReq_7_bits_fpReduceValid;
  wire              exeRequestQueue_8_enq_valid = exeReq_8_valid;
  wire [31:0]       exeRequestQueue_8_enq_bits_source1 = exeReq_8_bits_source1;
  wire [31:0]       exeRequestQueue_8_enq_bits_source2 = exeReq_8_bits_source2;
  wire [2:0]        exeRequestQueue_8_enq_bits_index = exeReq_8_bits_index;
  wire              exeRequestQueue_8_enq_bits_ffo = exeReq_8_bits_ffo;
  wire              exeRequestQueue_8_enq_bits_fpReduceValid = exeReq_8_bits_fpReduceValid;
  wire              exeRequestQueue_9_enq_valid = exeReq_9_valid;
  wire [31:0]       exeRequestQueue_9_enq_bits_source1 = exeReq_9_bits_source1;
  wire [31:0]       exeRequestQueue_9_enq_bits_source2 = exeReq_9_bits_source2;
  wire [2:0]        exeRequestQueue_9_enq_bits_index = exeReq_9_bits_index;
  wire              exeRequestQueue_9_enq_bits_ffo = exeReq_9_bits_ffo;
  wire              exeRequestQueue_9_enq_bits_fpReduceValid = exeReq_9_bits_fpReduceValid;
  wire              exeRequestQueue_10_enq_valid = exeReq_10_valid;
  wire [31:0]       exeRequestQueue_10_enq_bits_source1 = exeReq_10_bits_source1;
  wire [31:0]       exeRequestQueue_10_enq_bits_source2 = exeReq_10_bits_source2;
  wire [2:0]        exeRequestQueue_10_enq_bits_index = exeReq_10_bits_index;
  wire              exeRequestQueue_10_enq_bits_ffo = exeReq_10_bits_ffo;
  wire              exeRequestQueue_10_enq_bits_fpReduceValid = exeReq_10_bits_fpReduceValid;
  wire              exeRequestQueue_11_enq_valid = exeReq_11_valid;
  wire [31:0]       exeRequestQueue_11_enq_bits_source1 = exeReq_11_bits_source1;
  wire [31:0]       exeRequestQueue_11_enq_bits_source2 = exeReq_11_bits_source2;
  wire [2:0]        exeRequestQueue_11_enq_bits_index = exeReq_11_bits_index;
  wire              exeRequestQueue_11_enq_bits_ffo = exeReq_11_bits_ffo;
  wire              exeRequestQueue_11_enq_bits_fpReduceValid = exeReq_11_bits_fpReduceValid;
  wire              exeRequestQueue_12_enq_valid = exeReq_12_valid;
  wire [31:0]       exeRequestQueue_12_enq_bits_source1 = exeReq_12_bits_source1;
  wire [31:0]       exeRequestQueue_12_enq_bits_source2 = exeReq_12_bits_source2;
  wire [2:0]        exeRequestQueue_12_enq_bits_index = exeReq_12_bits_index;
  wire              exeRequestQueue_12_enq_bits_ffo = exeReq_12_bits_ffo;
  wire              exeRequestQueue_12_enq_bits_fpReduceValid = exeReq_12_bits_fpReduceValid;
  wire              exeRequestQueue_13_enq_valid = exeReq_13_valid;
  wire [31:0]       exeRequestQueue_13_enq_bits_source1 = exeReq_13_bits_source1;
  wire [31:0]       exeRequestQueue_13_enq_bits_source2 = exeReq_13_bits_source2;
  wire [2:0]        exeRequestQueue_13_enq_bits_index = exeReq_13_bits_index;
  wire              exeRequestQueue_13_enq_bits_ffo = exeReq_13_bits_ffo;
  wire              exeRequestQueue_13_enq_bits_fpReduceValid = exeReq_13_bits_fpReduceValid;
  wire              exeRequestQueue_14_enq_valid = exeReq_14_valid;
  wire [31:0]       exeRequestQueue_14_enq_bits_source1 = exeReq_14_bits_source1;
  wire [31:0]       exeRequestQueue_14_enq_bits_source2 = exeReq_14_bits_source2;
  wire [2:0]        exeRequestQueue_14_enq_bits_index = exeReq_14_bits_index;
  wire              exeRequestQueue_14_enq_bits_ffo = exeReq_14_bits_ffo;
  wire              exeRequestQueue_14_enq_bits_fpReduceValid = exeReq_14_bits_fpReduceValid;
  wire              exeRequestQueue_15_enq_valid = exeReq_15_valid;
  wire [31:0]       exeRequestQueue_15_enq_bits_source1 = exeReq_15_bits_source1;
  wire [31:0]       exeRequestQueue_15_enq_bits_source2 = exeReq_15_bits_source2;
  wire [2:0]        exeRequestQueue_15_enq_bits_index = exeReq_15_bits_index;
  wire              exeRequestQueue_15_enq_bits_ffo = exeReq_15_bits_ffo;
  wire              exeRequestQueue_15_enq_bits_fpReduceValid = exeReq_15_bits_fpReduceValid;
  wire              reorderQueueVec_0_enq_valid = readResult_0_valid;
  wire              reorderQueueVec_1_enq_valid = readResult_1_valid;
  wire              reorderQueueVec_2_enq_valid = readResult_2_valid;
  wire              reorderQueueVec_3_enq_valid = readResult_3_valid;
  wire              reorderQueueVec_4_enq_valid = readResult_4_valid;
  wire              reorderQueueVec_5_enq_valid = readResult_5_valid;
  wire              reorderQueueVec_6_enq_valid = readResult_6_valid;
  wire              reorderQueueVec_7_enq_valid = readResult_7_valid;
  wire              reorderQueueVec_8_enq_valid = readResult_8_valid;
  wire              reorderQueueVec_9_enq_valid = readResult_9_valid;
  wire              reorderQueueVec_10_enq_valid = readResult_10_valid;
  wire              reorderQueueVec_11_enq_valid = readResult_11_valid;
  wire              reorderQueueVec_12_enq_valid = readResult_12_valid;
  wire              reorderQueueVec_13_enq_valid = readResult_13_valid;
  wire              reorderQueueVec_14_enq_valid = readResult_14_valid;
  wire              reorderQueueVec_15_enq_valid = readResult_15_valid;
  wire              readMessageQueue_deq_ready = readResult_0_valid;
  wire              readMessageQueue_1_deq_ready = readResult_1_valid;
  wire              readMessageQueue_2_deq_ready = readResult_2_valid;
  wire              readMessageQueue_3_deq_ready = readResult_3_valid;
  wire              readMessageQueue_4_deq_ready = readResult_4_valid;
  wire              readMessageQueue_5_deq_ready = readResult_5_valid;
  wire              readMessageQueue_6_deq_ready = readResult_6_valid;
  wire              readMessageQueue_7_deq_ready = readResult_7_valid;
  wire              readMessageQueue_8_deq_ready = readResult_8_valid;
  wire              readMessageQueue_9_deq_ready = readResult_9_valid;
  wire              readMessageQueue_10_deq_ready = readResult_10_valid;
  wire              readMessageQueue_11_deq_ready = readResult_11_valid;
  wire              readMessageQueue_12_deq_ready = readResult_12_valid;
  wire              readMessageQueue_13_deq_ready = readResult_13_valid;
  wire              readMessageQueue_14_deq_ready = readResult_14_valid;
  wire              readMessageQueue_15_deq_ready = readResult_15_valid;
  wire [7:0]        checkVec_checkResult_lo_lo_lo_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_lo_lo_hi_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_lo_hi_lo_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_lo_hi_hi_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_hi_lo_lo_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_hi_lo_hi_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_hi_hi_lo_14 = 8'hFF;
  wire [7:0]        checkVec_checkResult_hi_hi_hi_14 = 8'hFF;
  wire [1:0]        checkVec_checkResultVec_0_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_1_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_2_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_3_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_4_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_5_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_6_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_7_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_8_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_9_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_10_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_11_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_12_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_13_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_14_1_2 = 2'h0;
  wire [1:0]        checkVec_checkResultVec_15_1_2 = 2'h0;
  wire [15:0]       checkVec_checkResult_lo_lo_14 = 16'hFFFF;
  wire [15:0]       checkVec_checkResult_lo_hi_14 = 16'hFFFF;
  wire [15:0]       checkVec_checkResult_hi_lo_14 = 16'hFFFF;
  wire [15:0]       checkVec_checkResult_hi_hi_14 = 16'hFFFF;
  wire [31:0]       checkVec_checkResult_lo_14 = 32'hFFFFFFFF;
  wire [31:0]       checkVec_checkResult_hi_14 = 32'hFFFFFFFF;
  wire [63:0]       checkVec_2_0 = 64'hFFFFFFFFFFFFFFFF;
  wire [7:0]        checkVec_checkResult_lo_lo_15 = 8'h0;
  wire [7:0]        checkVec_checkResult_lo_hi_15 = 8'h0;
  wire [7:0]        checkVec_checkResult_hi_lo_15 = 8'h0;
  wire [7:0]        checkVec_checkResult_hi_hi_15 = 8'h0;
  wire [3:0]        readVS1Req_requestIndex = 4'h0;
  wire [3:0]        checkVec_checkResult_lo_lo_lo_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_lo_lo_hi_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_lo_hi_lo_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_lo_hi_hi_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_hi_lo_lo_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_hi_lo_hi_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_hi_hi_lo_15 = 4'h0;
  wire [3:0]        checkVec_checkResult_hi_hi_hi_15 = 4'h0;
  wire [3:0]        selectExecuteReq_0_bits_requestIndex = 4'h0;
  wire [3:0]        selectExecuteReq_1_bits_requestIndex = 4'h1;
  wire [3:0]        selectExecuteReq_2_bits_requestIndex = 4'h2;
  wire [3:0]        selectExecuteReq_3_bits_requestIndex = 4'h3;
  wire [3:0]        selectExecuteReq_4_bits_requestIndex = 4'h4;
  wire [3:0]        selectExecuteReq_5_bits_requestIndex = 4'h5;
  wire [3:0]        selectExecuteReq_6_bits_requestIndex = 4'h6;
  wire [3:0]        selectExecuteReq_7_bits_requestIndex = 4'h7;
  wire [3:0]        selectExecuteReq_8_bits_requestIndex = 4'h8;
  wire [3:0]        selectExecuteReq_9_bits_requestIndex = 4'h9;
  wire [3:0]        selectExecuteReq_10_bits_requestIndex = 4'hA;
  wire [3:0]        selectExecuteReq_11_bits_requestIndex = 4'hB;
  wire [3:0]        selectExecuteReq_12_bits_requestIndex = 4'hC;
  wire [3:0]        selectExecuteReq_13_bits_requestIndex = 4'hD;
  wire [3:0]        selectExecuteReq_14_bits_requestIndex = 4'hE;
  wire [3:0]        selectExecuteReq_15_bits_requestIndex = 4'hF;
  wire [15:0]       checkVec_checkResult_lo_15 = 16'h0;
  wire [15:0]       checkVec_checkResult_hi_15 = 16'h0;
  wire              vs1Split_0_2 = 1'h1;
  wire              vs1Split_1_2 = 1'h1;
  wire [31:0]       checkVec_2_1 = 32'h0;
  wire [1:0]        readChannel_0_bits_readSource = 2'h2;
  wire [1:0]        readChannel_1_bits_readSource = 2'h2;
  wire [1:0]        readChannel_2_bits_readSource = 2'h2;
  wire [1:0]        readChannel_3_bits_readSource = 2'h2;
  wire [1:0]        readChannel_4_bits_readSource = 2'h2;
  wire [1:0]        readChannel_5_bits_readSource = 2'h2;
  wire [1:0]        readChannel_6_bits_readSource = 2'h2;
  wire [1:0]        readChannel_7_bits_readSource = 2'h2;
  wire [1:0]        readChannel_8_bits_readSource = 2'h2;
  wire [1:0]        readChannel_9_bits_readSource = 2'h2;
  wire [1:0]        readChannel_10_bits_readSource = 2'h2;
  wire [1:0]        readChannel_11_bits_readSource = 2'h2;
  wire [1:0]        readChannel_12_bits_readSource = 2'h2;
  wire [1:0]        readChannel_13_bits_readSource = 2'h2;
  wire [1:0]        readChannel_14_bits_readSource = 2'h2;
  wire [1:0]        readChannel_15_bits_readSource = 2'h2;
  wire              exeResp_0_bits_last = 1'h0;
  wire              exeResp_1_bits_last = 1'h0;
  wire              exeResp_2_bits_last = 1'h0;
  wire              exeResp_3_bits_last = 1'h0;
  wire              exeResp_4_bits_last = 1'h0;
  wire              exeResp_5_bits_last = 1'h0;
  wire              exeResp_6_bits_last = 1'h0;
  wire              exeResp_7_bits_last = 1'h0;
  wire              exeResp_8_bits_last = 1'h0;
  wire              exeResp_9_bits_last = 1'h0;
  wire              exeResp_10_bits_last = 1'h0;
  wire              exeResp_11_bits_last = 1'h0;
  wire              exeResp_12_bits_last = 1'h0;
  wire              exeResp_13_bits_last = 1'h0;
  wire              exeResp_14_bits_last = 1'h0;
  wire              exeResp_15_bits_last = 1'h0;
  wire              writeRequest_0_ffoByOther = 1'h0;
  wire              writeRequest_1_ffoByOther = 1'h0;
  wire              writeRequest_2_ffoByOther = 1'h0;
  wire              writeRequest_3_ffoByOther = 1'h0;
  wire              writeRequest_4_ffoByOther = 1'h0;
  wire              writeRequest_5_ffoByOther = 1'h0;
  wire              writeRequest_6_ffoByOther = 1'h0;
  wire              writeRequest_7_ffoByOther = 1'h0;
  wire              writeRequest_8_ffoByOther = 1'h0;
  wire              writeRequest_9_ffoByOther = 1'h0;
  wire              writeRequest_10_ffoByOther = 1'h0;
  wire              writeRequest_11_ffoByOther = 1'h0;
  wire              writeRequest_12_ffoByOther = 1'h0;
  wire              writeRequest_13_ffoByOther = 1'h0;
  wire              writeRequest_14_ffoByOther = 1'h0;
  wire              writeRequest_15_ffoByOther = 1'h0;
  wire              writeQueue_0_deq_ready = exeResp_0_ready_0;
  wire              writeQueue_0_deq_valid;
  wire [3:0]        writeQueue_0_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_0_deq_bits_writeData_data;
  wire              writeQueue_1_deq_ready = exeResp_1_ready_0;
  wire              writeQueue_1_deq_valid;
  wire [3:0]        writeQueue_1_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_1_deq_bits_writeData_data;
  wire              writeQueue_2_deq_ready = exeResp_2_ready_0;
  wire              writeQueue_2_deq_valid;
  wire [3:0]        writeQueue_2_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_2_deq_bits_writeData_data;
  wire              writeQueue_3_deq_ready = exeResp_3_ready_0;
  wire              writeQueue_3_deq_valid;
  wire [3:0]        writeQueue_3_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_3_deq_bits_writeData_data;
  wire              writeQueue_4_deq_ready = exeResp_4_ready_0;
  wire              writeQueue_4_deq_valid;
  wire [3:0]        writeQueue_4_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_4_deq_bits_writeData_data;
  wire              writeQueue_5_deq_ready = exeResp_5_ready_0;
  wire              writeQueue_5_deq_valid;
  wire [3:0]        writeQueue_5_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_5_deq_bits_writeData_data;
  wire              writeQueue_6_deq_ready = exeResp_6_ready_0;
  wire              writeQueue_6_deq_valid;
  wire [3:0]        writeQueue_6_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_6_deq_bits_writeData_data;
  wire              writeQueue_7_deq_ready = exeResp_7_ready_0;
  wire              writeQueue_7_deq_valid;
  wire [3:0]        writeQueue_7_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_7_deq_bits_writeData_data;
  wire              writeQueue_8_deq_ready = exeResp_8_ready_0;
  wire              writeQueue_8_deq_valid;
  wire [3:0]        writeQueue_8_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_8_deq_bits_writeData_data;
  wire              writeQueue_9_deq_ready = exeResp_9_ready_0;
  wire              writeQueue_9_deq_valid;
  wire [3:0]        writeQueue_9_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_9_deq_bits_writeData_data;
  wire              writeQueue_10_deq_ready = exeResp_10_ready_0;
  wire              writeQueue_10_deq_valid;
  wire [3:0]        writeQueue_10_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_10_deq_bits_writeData_data;
  wire              writeQueue_11_deq_ready = exeResp_11_ready_0;
  wire              writeQueue_11_deq_valid;
  wire [3:0]        writeQueue_11_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_11_deq_bits_writeData_data;
  wire              writeQueue_12_deq_ready = exeResp_12_ready_0;
  wire              writeQueue_12_deq_valid;
  wire [3:0]        writeQueue_12_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_12_deq_bits_writeData_data;
  wire              writeQueue_13_deq_ready = exeResp_13_ready_0;
  wire              writeQueue_13_deq_valid;
  wire [3:0]        writeQueue_13_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_13_deq_bits_writeData_data;
  wire              writeQueue_14_deq_ready = exeResp_14_ready_0;
  wire              writeQueue_14_deq_valid;
  wire [3:0]        writeQueue_14_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_14_deq_bits_writeData_data;
  wire              writeQueue_15_deq_ready = exeResp_15_ready_0;
  wire              writeQueue_15_deq_valid;
  wire [3:0]        writeQueue_15_deq_bits_writeData_mask;
  wire [31:0]       writeQueue_15_deq_bits_writeData_data;
  wire              gatherResponse;
  reg  [31:0]       v0_0;
  reg  [31:0]       v0_1;
  reg  [31:0]       v0_2;
  reg  [31:0]       v0_3;
  reg  [31:0]       v0_4;
  reg  [31:0]       v0_5;
  reg  [31:0]       v0_6;
  reg  [31:0]       v0_7;
  reg  [31:0]       v0_8;
  reg  [31:0]       v0_9;
  reg  [31:0]       v0_10;
  reg  [31:0]       v0_11;
  reg  [31:0]       v0_12;
  reg  [31:0]       v0_13;
  reg  [31:0]       v0_14;
  reg  [31:0]       v0_15;
  reg  [31:0]       v0_16;
  reg  [31:0]       v0_17;
  reg  [31:0]       v0_18;
  reg  [31:0]       v0_19;
  reg  [31:0]       v0_20;
  reg  [31:0]       v0_21;
  reg  [31:0]       v0_22;
  reg  [31:0]       v0_23;
  reg  [31:0]       v0_24;
  reg  [31:0]       v0_25;
  reg  [31:0]       v0_26;
  reg  [31:0]       v0_27;
  reg  [31:0]       v0_28;
  reg  [31:0]       v0_29;
  reg  [31:0]       v0_30;
  reg  [31:0]       v0_31;
  wire [15:0]       maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]       maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]       maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]       maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]       maskExt_lo_4 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_4 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]       maskExt_lo_5 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_5 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]       maskExt_lo_6 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_6 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]       maskExt_lo_7 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_7 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]       maskExt_lo_8 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_8 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]       maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]       maskExt_lo_9 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_9 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]       maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]       maskExt_lo_10 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_10 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]       maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]       maskExt_lo_11 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_11 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]       maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]       maskExt_lo_12 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_12 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]       maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]       maskExt_lo_13 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_13 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]       maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]       maskExt_lo_14 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_14 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]       maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]       maskExt_lo_15 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_15 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]       maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]       maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]       maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]       maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]       maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]       maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]       maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]       maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]       maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]       maskExt_lo_20 = {{8{v0UpdateVec_4_bits_mask[1]}}, {8{v0UpdateVec_4_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_20 = {{8{v0UpdateVec_4_bits_mask[3]}}, {8{v0UpdateVec_4_bits_mask[2]}}};
  wire [31:0]       maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]       maskExt_lo_21 = {{8{v0UpdateVec_5_bits_mask[1]}}, {8{v0UpdateVec_5_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_21 = {{8{v0UpdateVec_5_bits_mask[3]}}, {8{v0UpdateVec_5_bits_mask[2]}}};
  wire [31:0]       maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]       maskExt_lo_22 = {{8{v0UpdateVec_6_bits_mask[1]}}, {8{v0UpdateVec_6_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_22 = {{8{v0UpdateVec_6_bits_mask[3]}}, {8{v0UpdateVec_6_bits_mask[2]}}};
  wire [31:0]       maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]       maskExt_lo_23 = {{8{v0UpdateVec_7_bits_mask[1]}}, {8{v0UpdateVec_7_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_23 = {{8{v0UpdateVec_7_bits_mask[3]}}, {8{v0UpdateVec_7_bits_mask[2]}}};
  wire [31:0]       maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]       maskExt_lo_24 = {{8{v0UpdateVec_8_bits_mask[1]}}, {8{v0UpdateVec_8_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_24 = {{8{v0UpdateVec_8_bits_mask[3]}}, {8{v0UpdateVec_8_bits_mask[2]}}};
  wire [31:0]       maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]       maskExt_lo_25 = {{8{v0UpdateVec_9_bits_mask[1]}}, {8{v0UpdateVec_9_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_25 = {{8{v0UpdateVec_9_bits_mask[3]}}, {8{v0UpdateVec_9_bits_mask[2]}}};
  wire [31:0]       maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]       maskExt_lo_26 = {{8{v0UpdateVec_10_bits_mask[1]}}, {8{v0UpdateVec_10_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_26 = {{8{v0UpdateVec_10_bits_mask[3]}}, {8{v0UpdateVec_10_bits_mask[2]}}};
  wire [31:0]       maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]       maskExt_lo_27 = {{8{v0UpdateVec_11_bits_mask[1]}}, {8{v0UpdateVec_11_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_27 = {{8{v0UpdateVec_11_bits_mask[3]}}, {8{v0UpdateVec_11_bits_mask[2]}}};
  wire [31:0]       maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]       maskExt_lo_28 = {{8{v0UpdateVec_12_bits_mask[1]}}, {8{v0UpdateVec_12_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_28 = {{8{v0UpdateVec_12_bits_mask[3]}}, {8{v0UpdateVec_12_bits_mask[2]}}};
  wire [31:0]       maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]       maskExt_lo_29 = {{8{v0UpdateVec_13_bits_mask[1]}}, {8{v0UpdateVec_13_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_29 = {{8{v0UpdateVec_13_bits_mask[3]}}, {8{v0UpdateVec_13_bits_mask[2]}}};
  wire [31:0]       maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]       maskExt_lo_30 = {{8{v0UpdateVec_14_bits_mask[1]}}, {8{v0UpdateVec_14_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_30 = {{8{v0UpdateVec_14_bits_mask[3]}}, {8{v0UpdateVec_14_bits_mask[2]}}};
  wire [31:0]       maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]       maskExt_lo_31 = {{8{v0UpdateVec_15_bits_mask[1]}}, {8{v0UpdateVec_15_bits_mask[0]}}};
  wire [15:0]       maskExt_hi_31 = {{8{v0UpdateVec_15_bits_mask[3]}}, {8{v0UpdateVec_15_bits_mask[2]}}};
  wire [31:0]       maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [63:0]       _GEN = {v0_1, v0_0};
  wire [63:0]       regroupV0_lo_lo_lo_lo;
  assign regroupV0_lo_lo_lo_lo = _GEN;
  wire [63:0]       regroupV0_lo_lo_lo_lo_1;
  assign regroupV0_lo_lo_lo_lo_1 = _GEN;
  wire [63:0]       regroupV0_lo_lo_lo_lo_18;
  assign regroupV0_lo_lo_lo_lo_18 = _GEN;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo = _GEN;
  wire [63:0]       selectReadStageMask_lo_lo_lo_lo;
  assign selectReadStageMask_lo_lo_lo_lo = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_1 = _GEN;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_2 = _GEN;
  wire [63:0]       maskForDestination_lo_lo_lo_lo;
  assign maskForDestination_lo_lo_lo_lo = _GEN;
  wire [63:0]       _GEN_0 = {v0_3, v0_2};
  wire [63:0]       regroupV0_lo_lo_lo_hi;
  assign regroupV0_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       regroupV0_lo_lo_lo_hi_1;
  assign regroupV0_lo_lo_lo_hi_1 = _GEN_0;
  wire [63:0]       regroupV0_lo_lo_lo_hi_18;
  assign regroupV0_lo_lo_lo_hi_18 = _GEN_0;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       selectReadStageMask_lo_lo_lo_hi;
  assign selectReadStageMask_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_1 = _GEN_0;
  wire [63:0]       maskSplit_maskSelect_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_2 = _GEN_0;
  wire [63:0]       maskForDestination_lo_lo_lo_hi;
  assign maskForDestination_lo_lo_lo_hi = _GEN_0;
  wire [127:0]      regroupV0_lo_lo_lo = {regroupV0_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo};
  wire [63:0]       _GEN_1 = {v0_5, v0_4};
  wire [63:0]       regroupV0_lo_lo_hi_lo;
  assign regroupV0_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       regroupV0_lo_lo_hi_lo_1;
  assign regroupV0_lo_lo_hi_lo_1 = _GEN_1;
  wire [63:0]       regroupV0_lo_lo_hi_lo_18;
  assign regroupV0_lo_lo_hi_lo_18 = _GEN_1;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       selectReadStageMask_lo_lo_hi_lo;
  assign selectReadStageMask_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_1 = _GEN_1;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_2 = _GEN_1;
  wire [63:0]       maskForDestination_lo_lo_hi_lo;
  assign maskForDestination_lo_lo_hi_lo = _GEN_1;
  wire [63:0]       _GEN_2 = {v0_7, v0_6};
  wire [63:0]       regroupV0_lo_lo_hi_hi;
  assign regroupV0_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       regroupV0_lo_lo_hi_hi_1;
  assign regroupV0_lo_lo_hi_hi_1 = _GEN_2;
  wire [63:0]       regroupV0_lo_lo_hi_hi_18;
  assign regroupV0_lo_lo_hi_hi_18 = _GEN_2;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       selectReadStageMask_lo_lo_hi_hi;
  assign selectReadStageMask_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_1 = _GEN_2;
  wire [63:0]       maskSplit_maskSelect_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_2 = _GEN_2;
  wire [63:0]       maskForDestination_lo_lo_hi_hi;
  assign maskForDestination_lo_lo_hi_hi = _GEN_2;
  wire [127:0]      regroupV0_lo_lo_hi = {regroupV0_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo};
  wire [255:0]      regroupV0_lo_lo = {regroupV0_lo_lo_hi, regroupV0_lo_lo_lo};
  wire [63:0]       _GEN_3 = {v0_9, v0_8};
  wire [63:0]       regroupV0_lo_hi_lo_lo;
  assign regroupV0_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       regroupV0_lo_hi_lo_lo_1;
  assign regroupV0_lo_hi_lo_lo_1 = _GEN_3;
  wire [63:0]       regroupV0_lo_hi_lo_lo_18;
  assign regroupV0_lo_hi_lo_lo_18 = _GEN_3;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       selectReadStageMask_lo_hi_lo_lo;
  assign selectReadStageMask_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_1 = _GEN_3;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_2 = _GEN_3;
  wire [63:0]       maskForDestination_lo_hi_lo_lo;
  assign maskForDestination_lo_hi_lo_lo = _GEN_3;
  wire [63:0]       _GEN_4 = {v0_11, v0_10};
  wire [63:0]       regroupV0_lo_hi_lo_hi;
  assign regroupV0_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       regroupV0_lo_hi_lo_hi_1;
  assign regroupV0_lo_hi_lo_hi_1 = _GEN_4;
  wire [63:0]       regroupV0_lo_hi_lo_hi_18;
  assign regroupV0_lo_hi_lo_hi_18 = _GEN_4;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       selectReadStageMask_lo_hi_lo_hi;
  assign selectReadStageMask_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi = _GEN_4;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_1 = _GEN_4;
  wire [63:0]       maskSplit_maskSelect_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_2 = _GEN_4;
  wire [63:0]       maskForDestination_lo_hi_lo_hi;
  assign maskForDestination_lo_hi_lo_hi = _GEN_4;
  wire [127:0]      regroupV0_lo_hi_lo = {regroupV0_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo};
  wire [63:0]       _GEN_5 = {v0_13, v0_12};
  wire [63:0]       regroupV0_lo_hi_hi_lo;
  assign regroupV0_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       regroupV0_lo_hi_hi_lo_1;
  assign regroupV0_lo_hi_hi_lo_1 = _GEN_5;
  wire [63:0]       regroupV0_lo_hi_hi_lo_18;
  assign regroupV0_lo_hi_hi_lo_18 = _GEN_5;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       selectReadStageMask_lo_hi_hi_lo;
  assign selectReadStageMask_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_1 = _GEN_5;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_2 = _GEN_5;
  wire [63:0]       maskForDestination_lo_hi_hi_lo;
  assign maskForDestination_lo_hi_hi_lo = _GEN_5;
  wire [63:0]       _GEN_6 = {v0_15, v0_14};
  wire [63:0]       regroupV0_lo_hi_hi_hi;
  assign regroupV0_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       regroupV0_lo_hi_hi_hi_1;
  assign regroupV0_lo_hi_hi_hi_1 = _GEN_6;
  wire [63:0]       regroupV0_lo_hi_hi_hi_18;
  assign regroupV0_lo_hi_hi_hi_18 = _GEN_6;
  wire [63:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       selectReadStageMask_lo_hi_hi_hi;
  assign selectReadStageMask_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi = _GEN_6;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_1 = _GEN_6;
  wire [63:0]       maskSplit_maskSelect_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_2 = _GEN_6;
  wire [63:0]       maskForDestination_lo_hi_hi_hi;
  assign maskForDestination_lo_hi_hi_hi = _GEN_6;
  wire [127:0]      regroupV0_lo_hi_hi = {regroupV0_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo};
  wire [255:0]      regroupV0_lo_hi = {regroupV0_lo_hi_hi, regroupV0_lo_hi_lo};
  wire [511:0]      regroupV0_lo = {regroupV0_lo_hi, regroupV0_lo_lo};
  wire [63:0]       _GEN_7 = {v0_17, v0_16};
  wire [63:0]       regroupV0_hi_lo_lo_lo;
  assign regroupV0_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       regroupV0_hi_lo_lo_lo_1;
  assign regroupV0_hi_lo_lo_lo_1 = _GEN_7;
  wire [63:0]       regroupV0_hi_lo_lo_lo_18;
  assign regroupV0_hi_lo_lo_lo_18 = _GEN_7;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       selectReadStageMask_hi_lo_lo_lo;
  assign selectReadStageMask_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_1 = _GEN_7;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_2 = _GEN_7;
  wire [63:0]       maskForDestination_hi_lo_lo_lo;
  assign maskForDestination_hi_lo_lo_lo = _GEN_7;
  wire [63:0]       _GEN_8 = {v0_19, v0_18};
  wire [63:0]       regroupV0_hi_lo_lo_hi;
  assign regroupV0_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       regroupV0_hi_lo_lo_hi_1;
  assign regroupV0_hi_lo_lo_hi_1 = _GEN_8;
  wire [63:0]       regroupV0_hi_lo_lo_hi_18;
  assign regroupV0_hi_lo_lo_hi_18 = _GEN_8;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       selectReadStageMask_hi_lo_lo_hi;
  assign selectReadStageMask_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi = _GEN_8;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_1 = _GEN_8;
  wire [63:0]       maskSplit_maskSelect_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_2 = _GEN_8;
  wire [63:0]       maskForDestination_hi_lo_lo_hi;
  assign maskForDestination_hi_lo_lo_hi = _GEN_8;
  wire [127:0]      regroupV0_hi_lo_lo = {regroupV0_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo};
  wire [63:0]       _GEN_9 = {v0_21, v0_20};
  wire [63:0]       regroupV0_hi_lo_hi_lo;
  assign regroupV0_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       regroupV0_hi_lo_hi_lo_1;
  assign regroupV0_hi_lo_hi_lo_1 = _GEN_9;
  wire [63:0]       regroupV0_hi_lo_hi_lo_18;
  assign regroupV0_hi_lo_hi_lo_18 = _GEN_9;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       selectReadStageMask_hi_lo_hi_lo;
  assign selectReadStageMask_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_1 = _GEN_9;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_2 = _GEN_9;
  wire [63:0]       maskForDestination_hi_lo_hi_lo;
  assign maskForDestination_hi_lo_hi_lo = _GEN_9;
  wire [63:0]       _GEN_10 = {v0_23, v0_22};
  wire [63:0]       regroupV0_hi_lo_hi_hi;
  assign regroupV0_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       regroupV0_hi_lo_hi_hi_1;
  assign regroupV0_hi_lo_hi_hi_1 = _GEN_10;
  wire [63:0]       regroupV0_hi_lo_hi_hi_18;
  assign regroupV0_hi_lo_hi_hi_18 = _GEN_10;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       selectReadStageMask_hi_lo_hi_hi;
  assign selectReadStageMask_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi = _GEN_10;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_1 = _GEN_10;
  wire [63:0]       maskSplit_maskSelect_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_2 = _GEN_10;
  wire [63:0]       maskForDestination_hi_lo_hi_hi;
  assign maskForDestination_hi_lo_hi_hi = _GEN_10;
  wire [127:0]      regroupV0_hi_lo_hi = {regroupV0_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo};
  wire [255:0]      regroupV0_hi_lo = {regroupV0_hi_lo_hi, regroupV0_hi_lo_lo};
  wire [63:0]       _GEN_11 = {v0_25, v0_24};
  wire [63:0]       regroupV0_hi_hi_lo_lo;
  assign regroupV0_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       regroupV0_hi_hi_lo_lo_1;
  assign regroupV0_hi_hi_lo_lo_1 = _GEN_11;
  wire [63:0]       regroupV0_hi_hi_lo_lo_18;
  assign regroupV0_hi_hi_lo_lo_18 = _GEN_11;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       selectReadStageMask_hi_hi_lo_lo;
  assign selectReadStageMask_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_1 = _GEN_11;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_2 = _GEN_11;
  wire [63:0]       maskForDestination_hi_hi_lo_lo;
  assign maskForDestination_hi_hi_lo_lo = _GEN_11;
  wire [63:0]       _GEN_12 = {v0_27, v0_26};
  wire [63:0]       regroupV0_hi_hi_lo_hi;
  assign regroupV0_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       regroupV0_hi_hi_lo_hi_1;
  assign regroupV0_hi_hi_lo_hi_1 = _GEN_12;
  wire [63:0]       regroupV0_hi_hi_lo_hi_18;
  assign regroupV0_hi_hi_lo_hi_18 = _GEN_12;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       selectReadStageMask_hi_hi_lo_hi;
  assign selectReadStageMask_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi = _GEN_12;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_1 = _GEN_12;
  wire [63:0]       maskSplit_maskSelect_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_2 = _GEN_12;
  wire [63:0]       maskForDestination_hi_hi_lo_hi;
  assign maskForDestination_hi_hi_lo_hi = _GEN_12;
  wire [127:0]      regroupV0_hi_hi_lo = {regroupV0_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo};
  wire [63:0]       _GEN_13 = {v0_29, v0_28};
  wire [63:0]       regroupV0_hi_hi_hi_lo;
  assign regroupV0_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       regroupV0_hi_hi_hi_lo_1;
  assign regroupV0_hi_hi_hi_lo_1 = _GEN_13;
  wire [63:0]       regroupV0_hi_hi_hi_lo_18;
  assign regroupV0_hi_hi_hi_lo_18 = _GEN_13;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       selectReadStageMask_hi_hi_hi_lo;
  assign selectReadStageMask_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_1 = _GEN_13;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_2 = _GEN_13;
  wire [63:0]       maskForDestination_hi_hi_hi_lo;
  assign maskForDestination_hi_hi_hi_lo = _GEN_13;
  wire [63:0]       _GEN_14 = {v0_31, v0_30};
  wire [63:0]       regroupV0_hi_hi_hi_hi;
  assign regroupV0_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       regroupV0_hi_hi_hi_hi_1;
  assign regroupV0_hi_hi_hi_hi_1 = _GEN_14;
  wire [63:0]       regroupV0_hi_hi_hi_hi_18;
  assign regroupV0_hi_hi_hi_hi_18 = _GEN_14;
  wire [63:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       selectReadStageMask_hi_hi_hi_hi;
  assign selectReadStageMask_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi = _GEN_14;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_1 = _GEN_14;
  wire [63:0]       maskSplit_maskSelect_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_2 = _GEN_14;
  wire [63:0]       maskForDestination_hi_hi_hi_hi;
  assign maskForDestination_hi_hi_hi_hi = _GEN_14;
  wire [127:0]      regroupV0_hi_hi_hi = {regroupV0_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo};
  wire [255:0]      regroupV0_hi_hi = {regroupV0_hi_hi_hi, regroupV0_hi_hi_lo};
  wire [511:0]      regroupV0_hi = {regroupV0_hi_hi, regroupV0_hi_lo};
  wire [7:0]        regroupV0_lo_lo_lo_1 = {regroupV0_lo[67:64], regroupV0_lo[3:0]};
  wire [7:0]        regroupV0_lo_lo_hi_1 = {regroupV0_lo[195:192], regroupV0_lo[131:128]};
  wire [15:0]       regroupV0_lo_lo_1 = {regroupV0_lo_lo_hi_1, regroupV0_lo_lo_lo_1};
  wire [7:0]        regroupV0_lo_hi_lo_1 = {regroupV0_lo[323:320], regroupV0_lo[259:256]};
  wire [7:0]        regroupV0_lo_hi_hi_1 = {regroupV0_lo[451:448], regroupV0_lo[387:384]};
  wire [15:0]       regroupV0_lo_hi_1 = {regroupV0_lo_hi_hi_1, regroupV0_lo_hi_lo_1};
  wire [31:0]       regroupV0_lo_1 = {regroupV0_lo_hi_1, regroupV0_lo_lo_1};
  wire [7:0]        regroupV0_hi_lo_lo_1 = {regroupV0_hi[67:64], regroupV0_hi[3:0]};
  wire [7:0]        regroupV0_hi_lo_hi_1 = {regroupV0_hi[195:192], regroupV0_hi[131:128]};
  wire [15:0]       regroupV0_hi_lo_1 = {regroupV0_hi_lo_hi_1, regroupV0_hi_lo_lo_1};
  wire [7:0]        regroupV0_hi_hi_lo_1 = {regroupV0_hi[323:320], regroupV0_hi[259:256]};
  wire [7:0]        regroupV0_hi_hi_hi_1 = {regroupV0_hi[451:448], regroupV0_hi[387:384]};
  wire [15:0]       regroupV0_hi_hi_1 = {regroupV0_hi_hi_hi_1, regroupV0_hi_hi_lo_1};
  wire [31:0]       regroupV0_hi_1 = {regroupV0_hi_hi_1, regroupV0_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_lo_2 = {regroupV0_lo[71:68], regroupV0_lo[7:4]};
  wire [7:0]        regroupV0_lo_lo_hi_2 = {regroupV0_lo[199:196], regroupV0_lo[135:132]};
  wire [15:0]       regroupV0_lo_lo_2 = {regroupV0_lo_lo_hi_2, regroupV0_lo_lo_lo_2};
  wire [7:0]        regroupV0_lo_hi_lo_2 = {regroupV0_lo[327:324], regroupV0_lo[263:260]};
  wire [7:0]        regroupV0_lo_hi_hi_2 = {regroupV0_lo[455:452], regroupV0_lo[391:388]};
  wire [15:0]       regroupV0_lo_hi_2 = {regroupV0_lo_hi_hi_2, regroupV0_lo_hi_lo_2};
  wire [31:0]       regroupV0_lo_2 = {regroupV0_lo_hi_2, regroupV0_lo_lo_2};
  wire [7:0]        regroupV0_hi_lo_lo_2 = {regroupV0_hi[71:68], regroupV0_hi[7:4]};
  wire [7:0]        regroupV0_hi_lo_hi_2 = {regroupV0_hi[199:196], regroupV0_hi[135:132]};
  wire [15:0]       regroupV0_hi_lo_2 = {regroupV0_hi_lo_hi_2, regroupV0_hi_lo_lo_2};
  wire [7:0]        regroupV0_hi_hi_lo_2 = {regroupV0_hi[327:324], regroupV0_hi[263:260]};
  wire [7:0]        regroupV0_hi_hi_hi_2 = {regroupV0_hi[455:452], regroupV0_hi[391:388]};
  wire [15:0]       regroupV0_hi_hi_2 = {regroupV0_hi_hi_hi_2, regroupV0_hi_hi_lo_2};
  wire [31:0]       regroupV0_hi_2 = {regroupV0_hi_hi_2, regroupV0_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_lo_3 = {regroupV0_lo[75:72], regroupV0_lo[11:8]};
  wire [7:0]        regroupV0_lo_lo_hi_3 = {regroupV0_lo[203:200], regroupV0_lo[139:136]};
  wire [15:0]       regroupV0_lo_lo_3 = {regroupV0_lo_lo_hi_3, regroupV0_lo_lo_lo_3};
  wire [7:0]        regroupV0_lo_hi_lo_3 = {regroupV0_lo[331:328], regroupV0_lo[267:264]};
  wire [7:0]        regroupV0_lo_hi_hi_3 = {regroupV0_lo[459:456], regroupV0_lo[395:392]};
  wire [15:0]       regroupV0_lo_hi_3 = {regroupV0_lo_hi_hi_3, regroupV0_lo_hi_lo_3};
  wire [31:0]       regroupV0_lo_3 = {regroupV0_lo_hi_3, regroupV0_lo_lo_3};
  wire [7:0]        regroupV0_hi_lo_lo_3 = {regroupV0_hi[75:72], regroupV0_hi[11:8]};
  wire [7:0]        regroupV0_hi_lo_hi_3 = {regroupV0_hi[203:200], regroupV0_hi[139:136]};
  wire [15:0]       regroupV0_hi_lo_3 = {regroupV0_hi_lo_hi_3, regroupV0_hi_lo_lo_3};
  wire [7:0]        regroupV0_hi_hi_lo_3 = {regroupV0_hi[331:328], regroupV0_hi[267:264]};
  wire [7:0]        regroupV0_hi_hi_hi_3 = {regroupV0_hi[459:456], regroupV0_hi[395:392]};
  wire [15:0]       regroupV0_hi_hi_3 = {regroupV0_hi_hi_hi_3, regroupV0_hi_hi_lo_3};
  wire [31:0]       regroupV0_hi_3 = {regroupV0_hi_hi_3, regroupV0_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_lo_4 = {regroupV0_lo[79:76], regroupV0_lo[15:12]};
  wire [7:0]        regroupV0_lo_lo_hi_4 = {regroupV0_lo[207:204], regroupV0_lo[143:140]};
  wire [15:0]       regroupV0_lo_lo_4 = {regroupV0_lo_lo_hi_4, regroupV0_lo_lo_lo_4};
  wire [7:0]        regroupV0_lo_hi_lo_4 = {regroupV0_lo[335:332], regroupV0_lo[271:268]};
  wire [7:0]        regroupV0_lo_hi_hi_4 = {regroupV0_lo[463:460], regroupV0_lo[399:396]};
  wire [15:0]       regroupV0_lo_hi_4 = {regroupV0_lo_hi_hi_4, regroupV0_lo_hi_lo_4};
  wire [31:0]       regroupV0_lo_4 = {regroupV0_lo_hi_4, regroupV0_lo_lo_4};
  wire [7:0]        regroupV0_hi_lo_lo_4 = {regroupV0_hi[79:76], regroupV0_hi[15:12]};
  wire [7:0]        regroupV0_hi_lo_hi_4 = {regroupV0_hi[207:204], regroupV0_hi[143:140]};
  wire [15:0]       regroupV0_hi_lo_4 = {regroupV0_hi_lo_hi_4, regroupV0_hi_lo_lo_4};
  wire [7:0]        regroupV0_hi_hi_lo_4 = {regroupV0_hi[335:332], regroupV0_hi[271:268]};
  wire [7:0]        regroupV0_hi_hi_hi_4 = {regroupV0_hi[463:460], regroupV0_hi[399:396]};
  wire [15:0]       regroupV0_hi_hi_4 = {regroupV0_hi_hi_hi_4, regroupV0_hi_hi_lo_4};
  wire [31:0]       regroupV0_hi_4 = {regroupV0_hi_hi_4, regroupV0_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_lo_5 = {regroupV0_lo[83:80], regroupV0_lo[19:16]};
  wire [7:0]        regroupV0_lo_lo_hi_5 = {regroupV0_lo[211:208], regroupV0_lo[147:144]};
  wire [15:0]       regroupV0_lo_lo_5 = {regroupV0_lo_lo_hi_5, regroupV0_lo_lo_lo_5};
  wire [7:0]        regroupV0_lo_hi_lo_5 = {regroupV0_lo[339:336], regroupV0_lo[275:272]};
  wire [7:0]        regroupV0_lo_hi_hi_5 = {regroupV0_lo[467:464], regroupV0_lo[403:400]};
  wire [15:0]       regroupV0_lo_hi_5 = {regroupV0_lo_hi_hi_5, regroupV0_lo_hi_lo_5};
  wire [31:0]       regroupV0_lo_5 = {regroupV0_lo_hi_5, regroupV0_lo_lo_5};
  wire [7:0]        regroupV0_hi_lo_lo_5 = {regroupV0_hi[83:80], regroupV0_hi[19:16]};
  wire [7:0]        regroupV0_hi_lo_hi_5 = {regroupV0_hi[211:208], regroupV0_hi[147:144]};
  wire [15:0]       regroupV0_hi_lo_5 = {regroupV0_hi_lo_hi_5, regroupV0_hi_lo_lo_5};
  wire [7:0]        regroupV0_hi_hi_lo_5 = {regroupV0_hi[339:336], regroupV0_hi[275:272]};
  wire [7:0]        regroupV0_hi_hi_hi_5 = {regroupV0_hi[467:464], regroupV0_hi[403:400]};
  wire [15:0]       regroupV0_hi_hi_5 = {regroupV0_hi_hi_hi_5, regroupV0_hi_hi_lo_5};
  wire [31:0]       regroupV0_hi_5 = {regroupV0_hi_hi_5, regroupV0_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_lo_6 = {regroupV0_lo[87:84], regroupV0_lo[23:20]};
  wire [7:0]        regroupV0_lo_lo_hi_6 = {regroupV0_lo[215:212], regroupV0_lo[151:148]};
  wire [15:0]       regroupV0_lo_lo_6 = {regroupV0_lo_lo_hi_6, regroupV0_lo_lo_lo_6};
  wire [7:0]        regroupV0_lo_hi_lo_6 = {regroupV0_lo[343:340], regroupV0_lo[279:276]};
  wire [7:0]        regroupV0_lo_hi_hi_6 = {regroupV0_lo[471:468], regroupV0_lo[407:404]};
  wire [15:0]       regroupV0_lo_hi_6 = {regroupV0_lo_hi_hi_6, regroupV0_lo_hi_lo_6};
  wire [31:0]       regroupV0_lo_6 = {regroupV0_lo_hi_6, regroupV0_lo_lo_6};
  wire [7:0]        regroupV0_hi_lo_lo_6 = {regroupV0_hi[87:84], regroupV0_hi[23:20]};
  wire [7:0]        regroupV0_hi_lo_hi_6 = {regroupV0_hi[215:212], regroupV0_hi[151:148]};
  wire [15:0]       regroupV0_hi_lo_6 = {regroupV0_hi_lo_hi_6, regroupV0_hi_lo_lo_6};
  wire [7:0]        regroupV0_hi_hi_lo_6 = {regroupV0_hi[343:340], regroupV0_hi[279:276]};
  wire [7:0]        regroupV0_hi_hi_hi_6 = {regroupV0_hi[471:468], regroupV0_hi[407:404]};
  wire [15:0]       regroupV0_hi_hi_6 = {regroupV0_hi_hi_hi_6, regroupV0_hi_hi_lo_6};
  wire [31:0]       regroupV0_hi_6 = {regroupV0_hi_hi_6, regroupV0_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_lo_7 = {regroupV0_lo[91:88], regroupV0_lo[27:24]};
  wire [7:0]        regroupV0_lo_lo_hi_7 = {regroupV0_lo[219:216], regroupV0_lo[155:152]};
  wire [15:0]       regroupV0_lo_lo_7 = {regroupV0_lo_lo_hi_7, regroupV0_lo_lo_lo_7};
  wire [7:0]        regroupV0_lo_hi_lo_7 = {regroupV0_lo[347:344], regroupV0_lo[283:280]};
  wire [7:0]        regroupV0_lo_hi_hi_7 = {regroupV0_lo[475:472], regroupV0_lo[411:408]};
  wire [15:0]       regroupV0_lo_hi_7 = {regroupV0_lo_hi_hi_7, regroupV0_lo_hi_lo_7};
  wire [31:0]       regroupV0_lo_7 = {regroupV0_lo_hi_7, regroupV0_lo_lo_7};
  wire [7:0]        regroupV0_hi_lo_lo_7 = {regroupV0_hi[91:88], regroupV0_hi[27:24]};
  wire [7:0]        regroupV0_hi_lo_hi_7 = {regroupV0_hi[219:216], regroupV0_hi[155:152]};
  wire [15:0]       regroupV0_hi_lo_7 = {regroupV0_hi_lo_hi_7, regroupV0_hi_lo_lo_7};
  wire [7:0]        regroupV0_hi_hi_lo_7 = {regroupV0_hi[347:344], regroupV0_hi[283:280]};
  wire [7:0]        regroupV0_hi_hi_hi_7 = {regroupV0_hi[475:472], regroupV0_hi[411:408]};
  wire [15:0]       regroupV0_hi_hi_7 = {regroupV0_hi_hi_hi_7, regroupV0_hi_hi_lo_7};
  wire [31:0]       regroupV0_hi_7 = {regroupV0_hi_hi_7, regroupV0_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_lo_8 = {regroupV0_lo[95:92], regroupV0_lo[31:28]};
  wire [7:0]        regroupV0_lo_lo_hi_8 = {regroupV0_lo[223:220], regroupV0_lo[159:156]};
  wire [15:0]       regroupV0_lo_lo_8 = {regroupV0_lo_lo_hi_8, regroupV0_lo_lo_lo_8};
  wire [7:0]        regroupV0_lo_hi_lo_8 = {regroupV0_lo[351:348], regroupV0_lo[287:284]};
  wire [7:0]        regroupV0_lo_hi_hi_8 = {regroupV0_lo[479:476], regroupV0_lo[415:412]};
  wire [15:0]       regroupV0_lo_hi_8 = {regroupV0_lo_hi_hi_8, regroupV0_lo_hi_lo_8};
  wire [31:0]       regroupV0_lo_8 = {regroupV0_lo_hi_8, regroupV0_lo_lo_8};
  wire [7:0]        regroupV0_hi_lo_lo_8 = {regroupV0_hi[95:92], regroupV0_hi[31:28]};
  wire [7:0]        regroupV0_hi_lo_hi_8 = {regroupV0_hi[223:220], regroupV0_hi[159:156]};
  wire [15:0]       regroupV0_hi_lo_8 = {regroupV0_hi_lo_hi_8, regroupV0_hi_lo_lo_8};
  wire [7:0]        regroupV0_hi_hi_lo_8 = {regroupV0_hi[351:348], regroupV0_hi[287:284]};
  wire [7:0]        regroupV0_hi_hi_hi_8 = {regroupV0_hi[479:476], regroupV0_hi[415:412]};
  wire [15:0]       regroupV0_hi_hi_8 = {regroupV0_hi_hi_hi_8, regroupV0_hi_hi_lo_8};
  wire [31:0]       regroupV0_hi_8 = {regroupV0_hi_hi_8, regroupV0_hi_lo_8};
  wire [7:0]        regroupV0_lo_lo_lo_9 = {regroupV0_lo[99:96], regroupV0_lo[35:32]};
  wire [7:0]        regroupV0_lo_lo_hi_9 = {regroupV0_lo[227:224], regroupV0_lo[163:160]};
  wire [15:0]       regroupV0_lo_lo_9 = {regroupV0_lo_lo_hi_9, regroupV0_lo_lo_lo_9};
  wire [7:0]        regroupV0_lo_hi_lo_9 = {regroupV0_lo[355:352], regroupV0_lo[291:288]};
  wire [7:0]        regroupV0_lo_hi_hi_9 = {regroupV0_lo[483:480], regroupV0_lo[419:416]};
  wire [15:0]       regroupV0_lo_hi_9 = {regroupV0_lo_hi_hi_9, regroupV0_lo_hi_lo_9};
  wire [31:0]       regroupV0_lo_9 = {regroupV0_lo_hi_9, regroupV0_lo_lo_9};
  wire [7:0]        regroupV0_hi_lo_lo_9 = {regroupV0_hi[99:96], regroupV0_hi[35:32]};
  wire [7:0]        regroupV0_hi_lo_hi_9 = {regroupV0_hi[227:224], regroupV0_hi[163:160]};
  wire [15:0]       regroupV0_hi_lo_9 = {regroupV0_hi_lo_hi_9, regroupV0_hi_lo_lo_9};
  wire [7:0]        regroupV0_hi_hi_lo_9 = {regroupV0_hi[355:352], regroupV0_hi[291:288]};
  wire [7:0]        regroupV0_hi_hi_hi_9 = {regroupV0_hi[483:480], regroupV0_hi[419:416]};
  wire [15:0]       regroupV0_hi_hi_9 = {regroupV0_hi_hi_hi_9, regroupV0_hi_hi_lo_9};
  wire [31:0]       regroupV0_hi_9 = {regroupV0_hi_hi_9, regroupV0_hi_lo_9};
  wire [7:0]        regroupV0_lo_lo_lo_10 = {regroupV0_lo[103:100], regroupV0_lo[39:36]};
  wire [7:0]        regroupV0_lo_lo_hi_10 = {regroupV0_lo[231:228], regroupV0_lo[167:164]};
  wire [15:0]       regroupV0_lo_lo_10 = {regroupV0_lo_lo_hi_10, regroupV0_lo_lo_lo_10};
  wire [7:0]        regroupV0_lo_hi_lo_10 = {regroupV0_lo[359:356], regroupV0_lo[295:292]};
  wire [7:0]        regroupV0_lo_hi_hi_10 = {regroupV0_lo[487:484], regroupV0_lo[423:420]};
  wire [15:0]       regroupV0_lo_hi_10 = {regroupV0_lo_hi_hi_10, regroupV0_lo_hi_lo_10};
  wire [31:0]       regroupV0_lo_10 = {regroupV0_lo_hi_10, regroupV0_lo_lo_10};
  wire [7:0]        regroupV0_hi_lo_lo_10 = {regroupV0_hi[103:100], regroupV0_hi[39:36]};
  wire [7:0]        regroupV0_hi_lo_hi_10 = {regroupV0_hi[231:228], regroupV0_hi[167:164]};
  wire [15:0]       regroupV0_hi_lo_10 = {regroupV0_hi_lo_hi_10, regroupV0_hi_lo_lo_10};
  wire [7:0]        regroupV0_hi_hi_lo_10 = {regroupV0_hi[359:356], regroupV0_hi[295:292]};
  wire [7:0]        regroupV0_hi_hi_hi_10 = {regroupV0_hi[487:484], regroupV0_hi[423:420]};
  wire [15:0]       regroupV0_hi_hi_10 = {regroupV0_hi_hi_hi_10, regroupV0_hi_hi_lo_10};
  wire [31:0]       regroupV0_hi_10 = {regroupV0_hi_hi_10, regroupV0_hi_lo_10};
  wire [7:0]        regroupV0_lo_lo_lo_11 = {regroupV0_lo[107:104], regroupV0_lo[43:40]};
  wire [7:0]        regroupV0_lo_lo_hi_11 = {regroupV0_lo[235:232], regroupV0_lo[171:168]};
  wire [15:0]       regroupV0_lo_lo_11 = {regroupV0_lo_lo_hi_11, regroupV0_lo_lo_lo_11};
  wire [7:0]        regroupV0_lo_hi_lo_11 = {regroupV0_lo[363:360], regroupV0_lo[299:296]};
  wire [7:0]        regroupV0_lo_hi_hi_11 = {regroupV0_lo[491:488], regroupV0_lo[427:424]};
  wire [15:0]       regroupV0_lo_hi_11 = {regroupV0_lo_hi_hi_11, regroupV0_lo_hi_lo_11};
  wire [31:0]       regroupV0_lo_11 = {regroupV0_lo_hi_11, regroupV0_lo_lo_11};
  wire [7:0]        regroupV0_hi_lo_lo_11 = {regroupV0_hi[107:104], regroupV0_hi[43:40]};
  wire [7:0]        regroupV0_hi_lo_hi_11 = {regroupV0_hi[235:232], regroupV0_hi[171:168]};
  wire [15:0]       regroupV0_hi_lo_11 = {regroupV0_hi_lo_hi_11, regroupV0_hi_lo_lo_11};
  wire [7:0]        regroupV0_hi_hi_lo_11 = {regroupV0_hi[363:360], regroupV0_hi[299:296]};
  wire [7:0]        regroupV0_hi_hi_hi_11 = {regroupV0_hi[491:488], regroupV0_hi[427:424]};
  wire [15:0]       regroupV0_hi_hi_11 = {regroupV0_hi_hi_hi_11, regroupV0_hi_hi_lo_11};
  wire [31:0]       regroupV0_hi_11 = {regroupV0_hi_hi_11, regroupV0_hi_lo_11};
  wire [7:0]        regroupV0_lo_lo_lo_12 = {regroupV0_lo[111:108], regroupV0_lo[47:44]};
  wire [7:0]        regroupV0_lo_lo_hi_12 = {regroupV0_lo[239:236], regroupV0_lo[175:172]};
  wire [15:0]       regroupV0_lo_lo_12 = {regroupV0_lo_lo_hi_12, regroupV0_lo_lo_lo_12};
  wire [7:0]        regroupV0_lo_hi_lo_12 = {regroupV0_lo[367:364], regroupV0_lo[303:300]};
  wire [7:0]        regroupV0_lo_hi_hi_12 = {regroupV0_lo[495:492], regroupV0_lo[431:428]};
  wire [15:0]       regroupV0_lo_hi_12 = {regroupV0_lo_hi_hi_12, regroupV0_lo_hi_lo_12};
  wire [31:0]       regroupV0_lo_12 = {regroupV0_lo_hi_12, regroupV0_lo_lo_12};
  wire [7:0]        regroupV0_hi_lo_lo_12 = {regroupV0_hi[111:108], regroupV0_hi[47:44]};
  wire [7:0]        regroupV0_hi_lo_hi_12 = {regroupV0_hi[239:236], regroupV0_hi[175:172]};
  wire [15:0]       regroupV0_hi_lo_12 = {regroupV0_hi_lo_hi_12, regroupV0_hi_lo_lo_12};
  wire [7:0]        regroupV0_hi_hi_lo_12 = {regroupV0_hi[367:364], regroupV0_hi[303:300]};
  wire [7:0]        regroupV0_hi_hi_hi_12 = {regroupV0_hi[495:492], regroupV0_hi[431:428]};
  wire [15:0]       regroupV0_hi_hi_12 = {regroupV0_hi_hi_hi_12, regroupV0_hi_hi_lo_12};
  wire [31:0]       regroupV0_hi_12 = {regroupV0_hi_hi_12, regroupV0_hi_lo_12};
  wire [7:0]        regroupV0_lo_lo_lo_13 = {regroupV0_lo[115:112], regroupV0_lo[51:48]};
  wire [7:0]        regroupV0_lo_lo_hi_13 = {regroupV0_lo[243:240], regroupV0_lo[179:176]};
  wire [15:0]       regroupV0_lo_lo_13 = {regroupV0_lo_lo_hi_13, regroupV0_lo_lo_lo_13};
  wire [7:0]        regroupV0_lo_hi_lo_13 = {regroupV0_lo[371:368], regroupV0_lo[307:304]};
  wire [7:0]        regroupV0_lo_hi_hi_13 = {regroupV0_lo[499:496], regroupV0_lo[435:432]};
  wire [15:0]       regroupV0_lo_hi_13 = {regroupV0_lo_hi_hi_13, regroupV0_lo_hi_lo_13};
  wire [31:0]       regroupV0_lo_13 = {regroupV0_lo_hi_13, regroupV0_lo_lo_13};
  wire [7:0]        regroupV0_hi_lo_lo_13 = {regroupV0_hi[115:112], regroupV0_hi[51:48]};
  wire [7:0]        regroupV0_hi_lo_hi_13 = {regroupV0_hi[243:240], regroupV0_hi[179:176]};
  wire [15:0]       regroupV0_hi_lo_13 = {regroupV0_hi_lo_hi_13, regroupV0_hi_lo_lo_13};
  wire [7:0]        regroupV0_hi_hi_lo_13 = {regroupV0_hi[371:368], regroupV0_hi[307:304]};
  wire [7:0]        regroupV0_hi_hi_hi_13 = {regroupV0_hi[499:496], regroupV0_hi[435:432]};
  wire [15:0]       regroupV0_hi_hi_13 = {regroupV0_hi_hi_hi_13, regroupV0_hi_hi_lo_13};
  wire [31:0]       regroupV0_hi_13 = {regroupV0_hi_hi_13, regroupV0_hi_lo_13};
  wire [7:0]        regroupV0_lo_lo_lo_14 = {regroupV0_lo[119:116], regroupV0_lo[55:52]};
  wire [7:0]        regroupV0_lo_lo_hi_14 = {regroupV0_lo[247:244], regroupV0_lo[183:180]};
  wire [15:0]       regroupV0_lo_lo_14 = {regroupV0_lo_lo_hi_14, regroupV0_lo_lo_lo_14};
  wire [7:0]        regroupV0_lo_hi_lo_14 = {regroupV0_lo[375:372], regroupV0_lo[311:308]};
  wire [7:0]        regroupV0_lo_hi_hi_14 = {regroupV0_lo[503:500], regroupV0_lo[439:436]};
  wire [15:0]       regroupV0_lo_hi_14 = {regroupV0_lo_hi_hi_14, regroupV0_lo_hi_lo_14};
  wire [31:0]       regroupV0_lo_14 = {regroupV0_lo_hi_14, regroupV0_lo_lo_14};
  wire [7:0]        regroupV0_hi_lo_lo_14 = {regroupV0_hi[119:116], regroupV0_hi[55:52]};
  wire [7:0]        regroupV0_hi_lo_hi_14 = {regroupV0_hi[247:244], regroupV0_hi[183:180]};
  wire [15:0]       regroupV0_hi_lo_14 = {regroupV0_hi_lo_hi_14, regroupV0_hi_lo_lo_14};
  wire [7:0]        regroupV0_hi_hi_lo_14 = {regroupV0_hi[375:372], regroupV0_hi[311:308]};
  wire [7:0]        regroupV0_hi_hi_hi_14 = {regroupV0_hi[503:500], regroupV0_hi[439:436]};
  wire [15:0]       regroupV0_hi_hi_14 = {regroupV0_hi_hi_hi_14, regroupV0_hi_hi_lo_14};
  wire [31:0]       regroupV0_hi_14 = {regroupV0_hi_hi_14, regroupV0_hi_lo_14};
  wire [7:0]        regroupV0_lo_lo_lo_15 = {regroupV0_lo[123:120], regroupV0_lo[59:56]};
  wire [7:0]        regroupV0_lo_lo_hi_15 = {regroupV0_lo[251:248], regroupV0_lo[187:184]};
  wire [15:0]       regroupV0_lo_lo_15 = {regroupV0_lo_lo_hi_15, regroupV0_lo_lo_lo_15};
  wire [7:0]        regroupV0_lo_hi_lo_15 = {regroupV0_lo[379:376], regroupV0_lo[315:312]};
  wire [7:0]        regroupV0_lo_hi_hi_15 = {regroupV0_lo[507:504], regroupV0_lo[443:440]};
  wire [15:0]       regroupV0_lo_hi_15 = {regroupV0_lo_hi_hi_15, regroupV0_lo_hi_lo_15};
  wire [31:0]       regroupV0_lo_15 = {regroupV0_lo_hi_15, regroupV0_lo_lo_15};
  wire [7:0]        regroupV0_hi_lo_lo_15 = {regroupV0_hi[123:120], regroupV0_hi[59:56]};
  wire [7:0]        regroupV0_hi_lo_hi_15 = {regroupV0_hi[251:248], regroupV0_hi[187:184]};
  wire [15:0]       regroupV0_hi_lo_15 = {regroupV0_hi_lo_hi_15, regroupV0_hi_lo_lo_15};
  wire [7:0]        regroupV0_hi_hi_lo_15 = {regroupV0_hi[379:376], regroupV0_hi[315:312]};
  wire [7:0]        regroupV0_hi_hi_hi_15 = {regroupV0_hi[507:504], regroupV0_hi[443:440]};
  wire [15:0]       regroupV0_hi_hi_15 = {regroupV0_hi_hi_hi_15, regroupV0_hi_hi_lo_15};
  wire [31:0]       regroupV0_hi_15 = {regroupV0_hi_hi_15, regroupV0_hi_lo_15};
  wire [7:0]        regroupV0_lo_lo_lo_16 = {regroupV0_lo[127:124], regroupV0_lo[63:60]};
  wire [7:0]        regroupV0_lo_lo_hi_16 = {regroupV0_lo[255:252], regroupV0_lo[191:188]};
  wire [15:0]       regroupV0_lo_lo_16 = {regroupV0_lo_lo_hi_16, regroupV0_lo_lo_lo_16};
  wire [7:0]        regroupV0_lo_hi_lo_16 = {regroupV0_lo[383:380], regroupV0_lo[319:316]};
  wire [7:0]        regroupV0_lo_hi_hi_16 = {regroupV0_lo[511:508], regroupV0_lo[447:444]};
  wire [15:0]       regroupV0_lo_hi_16 = {regroupV0_lo_hi_hi_16, regroupV0_lo_hi_lo_16};
  wire [31:0]       regroupV0_lo_16 = {regroupV0_lo_hi_16, regroupV0_lo_lo_16};
  wire [7:0]        regroupV0_hi_lo_lo_16 = {regroupV0_hi[127:124], regroupV0_hi[63:60]};
  wire [7:0]        regroupV0_hi_lo_hi_16 = {regroupV0_hi[255:252], regroupV0_hi[191:188]};
  wire [15:0]       regroupV0_hi_lo_16 = {regroupV0_hi_lo_hi_16, regroupV0_hi_lo_lo_16};
  wire [7:0]        regroupV0_hi_hi_lo_16 = {regroupV0_hi[383:380], regroupV0_hi[319:316]};
  wire [7:0]        regroupV0_hi_hi_hi_16 = {regroupV0_hi[511:508], regroupV0_hi[447:444]};
  wire [15:0]       regroupV0_hi_hi_16 = {regroupV0_hi_hi_hi_16, regroupV0_hi_hi_lo_16};
  wire [31:0]       regroupV0_hi_16 = {regroupV0_hi_hi_16, regroupV0_hi_lo_16};
  wire [127:0]      regroupV0_lo_lo_lo_17 = {regroupV0_hi_2, regroupV0_lo_2, regroupV0_hi_1, regroupV0_lo_1};
  wire [127:0]      regroupV0_lo_lo_hi_17 = {regroupV0_hi_4, regroupV0_lo_4, regroupV0_hi_3, regroupV0_lo_3};
  wire [255:0]      regroupV0_lo_lo_17 = {regroupV0_lo_lo_hi_17, regroupV0_lo_lo_lo_17};
  wire [127:0]      regroupV0_lo_hi_lo_17 = {regroupV0_hi_6, regroupV0_lo_6, regroupV0_hi_5, regroupV0_lo_5};
  wire [127:0]      regroupV0_lo_hi_hi_17 = {regroupV0_hi_8, regroupV0_lo_8, regroupV0_hi_7, regroupV0_lo_7};
  wire [255:0]      regroupV0_lo_hi_17 = {regroupV0_lo_hi_hi_17, regroupV0_lo_hi_lo_17};
  wire [511:0]      regroupV0_lo_17 = {regroupV0_lo_hi_17, regroupV0_lo_lo_17};
  wire [127:0]      regroupV0_hi_lo_lo_17 = {regroupV0_hi_10, regroupV0_lo_10, regroupV0_hi_9, regroupV0_lo_9};
  wire [127:0]      regroupV0_hi_lo_hi_17 = {regroupV0_hi_12, regroupV0_lo_12, regroupV0_hi_11, regroupV0_lo_11};
  wire [255:0]      regroupV0_hi_lo_17 = {regroupV0_hi_lo_hi_17, regroupV0_hi_lo_lo_17};
  wire [127:0]      regroupV0_hi_hi_lo_17 = {regroupV0_hi_14, regroupV0_lo_14, regroupV0_hi_13, regroupV0_lo_13};
  wire [127:0]      regroupV0_hi_hi_hi_17 = {regroupV0_hi_16, regroupV0_lo_16, regroupV0_hi_15, regroupV0_lo_15};
  wire [255:0]      regroupV0_hi_hi_17 = {regroupV0_hi_hi_hi_17, regroupV0_hi_hi_lo_17};
  wire [511:0]      regroupV0_hi_17 = {regroupV0_hi_hi_17, regroupV0_hi_lo_17};
  wire [1023:0]     regroupV0_0 = {regroupV0_hi_17, regroupV0_lo_17};
  wire [127:0]      regroupV0_lo_lo_lo_18 = {regroupV0_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_1};
  wire [127:0]      regroupV0_lo_lo_hi_18 = {regroupV0_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_1};
  wire [255:0]      regroupV0_lo_lo_18 = {regroupV0_lo_lo_hi_18, regroupV0_lo_lo_lo_18};
  wire [127:0]      regroupV0_lo_hi_lo_18 = {regroupV0_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_1};
  wire [127:0]      regroupV0_lo_hi_hi_18 = {regroupV0_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_1};
  wire [255:0]      regroupV0_lo_hi_18 = {regroupV0_lo_hi_hi_18, regroupV0_lo_hi_lo_18};
  wire [511:0]      regroupV0_lo_18 = {regroupV0_lo_hi_18, regroupV0_lo_lo_18};
  wire [127:0]      regroupV0_hi_lo_lo_18 = {regroupV0_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_1};
  wire [127:0]      regroupV0_hi_lo_hi_18 = {regroupV0_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_1};
  wire [255:0]      regroupV0_hi_lo_18 = {regroupV0_hi_lo_hi_18, regroupV0_hi_lo_lo_18};
  wire [127:0]      regroupV0_hi_hi_lo_18 = {regroupV0_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_1};
  wire [127:0]      regroupV0_hi_hi_hi_18 = {regroupV0_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_1};
  wire [255:0]      regroupV0_hi_hi_18 = {regroupV0_hi_hi_hi_18, regroupV0_hi_hi_lo_18};
  wire [511:0]      regroupV0_hi_18 = {regroupV0_hi_hi_18, regroupV0_hi_lo_18};
  wire [3:0]        regroupV0_lo_lo_lo_lo_2 = {regroupV0_lo_18[33:32], regroupV0_lo_18[1:0]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_2 = {regroupV0_lo_18[97:96], regroupV0_lo_18[65:64]};
  wire [7:0]        regroupV0_lo_lo_lo_19 = {regroupV0_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_2};
  wire [3:0]        regroupV0_lo_lo_hi_lo_2 = {regroupV0_lo_18[161:160], regroupV0_lo_18[129:128]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_2 = {regroupV0_lo_18[225:224], regroupV0_lo_18[193:192]};
  wire [7:0]        regroupV0_lo_lo_hi_19 = {regroupV0_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_2};
  wire [15:0]       regroupV0_lo_lo_19 = {regroupV0_lo_lo_hi_19, regroupV0_lo_lo_lo_19};
  wire [3:0]        regroupV0_lo_hi_lo_lo_2 = {regroupV0_lo_18[289:288], regroupV0_lo_18[257:256]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_2 = {regroupV0_lo_18[353:352], regroupV0_lo_18[321:320]};
  wire [7:0]        regroupV0_lo_hi_lo_19 = {regroupV0_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_2};
  wire [3:0]        regroupV0_lo_hi_hi_lo_2 = {regroupV0_lo_18[417:416], regroupV0_lo_18[385:384]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_2 = {regroupV0_lo_18[481:480], regroupV0_lo_18[449:448]};
  wire [7:0]        regroupV0_lo_hi_hi_19 = {regroupV0_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_2};
  wire [15:0]       regroupV0_lo_hi_19 = {regroupV0_lo_hi_hi_19, regroupV0_lo_hi_lo_19};
  wire [31:0]       regroupV0_lo_19 = {regroupV0_lo_hi_19, regroupV0_lo_lo_19};
  wire [3:0]        regroupV0_hi_lo_lo_lo_2 = {regroupV0_hi_18[33:32], regroupV0_hi_18[1:0]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_2 = {regroupV0_hi_18[97:96], regroupV0_hi_18[65:64]};
  wire [7:0]        regroupV0_hi_lo_lo_19 = {regroupV0_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_2};
  wire [3:0]        regroupV0_hi_lo_hi_lo_2 = {regroupV0_hi_18[161:160], regroupV0_hi_18[129:128]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_2 = {regroupV0_hi_18[225:224], regroupV0_hi_18[193:192]};
  wire [7:0]        regroupV0_hi_lo_hi_19 = {regroupV0_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_2};
  wire [15:0]       regroupV0_hi_lo_19 = {regroupV0_hi_lo_hi_19, regroupV0_hi_lo_lo_19};
  wire [3:0]        regroupV0_hi_hi_lo_lo_2 = {regroupV0_hi_18[289:288], regroupV0_hi_18[257:256]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_2 = {regroupV0_hi_18[353:352], regroupV0_hi_18[321:320]};
  wire [7:0]        regroupV0_hi_hi_lo_19 = {regroupV0_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_2};
  wire [3:0]        regroupV0_hi_hi_hi_lo_2 = {regroupV0_hi_18[417:416], regroupV0_hi_18[385:384]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_2 = {regroupV0_hi_18[481:480], regroupV0_hi_18[449:448]};
  wire [7:0]        regroupV0_hi_hi_hi_19 = {regroupV0_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_2};
  wire [15:0]       regroupV0_hi_hi_19 = {regroupV0_hi_hi_hi_19, regroupV0_hi_hi_lo_19};
  wire [31:0]       regroupV0_hi_19 = {regroupV0_hi_hi_19, regroupV0_hi_lo_19};
  wire [3:0]        regroupV0_lo_lo_lo_lo_3 = {regroupV0_lo_18[35:34], regroupV0_lo_18[3:2]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_3 = {regroupV0_lo_18[99:98], regroupV0_lo_18[67:66]};
  wire [7:0]        regroupV0_lo_lo_lo_20 = {regroupV0_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_3};
  wire [3:0]        regroupV0_lo_lo_hi_lo_3 = {regroupV0_lo_18[163:162], regroupV0_lo_18[131:130]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_3 = {regroupV0_lo_18[227:226], regroupV0_lo_18[195:194]};
  wire [7:0]        regroupV0_lo_lo_hi_20 = {regroupV0_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_3};
  wire [15:0]       regroupV0_lo_lo_20 = {regroupV0_lo_lo_hi_20, regroupV0_lo_lo_lo_20};
  wire [3:0]        regroupV0_lo_hi_lo_lo_3 = {regroupV0_lo_18[291:290], regroupV0_lo_18[259:258]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_3 = {regroupV0_lo_18[355:354], regroupV0_lo_18[323:322]};
  wire [7:0]        regroupV0_lo_hi_lo_20 = {regroupV0_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_3};
  wire [3:0]        regroupV0_lo_hi_hi_lo_3 = {regroupV0_lo_18[419:418], regroupV0_lo_18[387:386]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_3 = {regroupV0_lo_18[483:482], regroupV0_lo_18[451:450]};
  wire [7:0]        regroupV0_lo_hi_hi_20 = {regroupV0_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_3};
  wire [15:0]       regroupV0_lo_hi_20 = {regroupV0_lo_hi_hi_20, regroupV0_lo_hi_lo_20};
  wire [31:0]       regroupV0_lo_20 = {regroupV0_lo_hi_20, regroupV0_lo_lo_20};
  wire [3:0]        regroupV0_hi_lo_lo_lo_3 = {regroupV0_hi_18[35:34], regroupV0_hi_18[3:2]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_3 = {regroupV0_hi_18[99:98], regroupV0_hi_18[67:66]};
  wire [7:0]        regroupV0_hi_lo_lo_20 = {regroupV0_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_3};
  wire [3:0]        regroupV0_hi_lo_hi_lo_3 = {regroupV0_hi_18[163:162], regroupV0_hi_18[131:130]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_3 = {regroupV0_hi_18[227:226], regroupV0_hi_18[195:194]};
  wire [7:0]        regroupV0_hi_lo_hi_20 = {regroupV0_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_3};
  wire [15:0]       regroupV0_hi_lo_20 = {regroupV0_hi_lo_hi_20, regroupV0_hi_lo_lo_20};
  wire [3:0]        regroupV0_hi_hi_lo_lo_3 = {regroupV0_hi_18[291:290], regroupV0_hi_18[259:258]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_3 = {regroupV0_hi_18[355:354], regroupV0_hi_18[323:322]};
  wire [7:0]        regroupV0_hi_hi_lo_20 = {regroupV0_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_3};
  wire [3:0]        regroupV0_hi_hi_hi_lo_3 = {regroupV0_hi_18[419:418], regroupV0_hi_18[387:386]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_3 = {regroupV0_hi_18[483:482], regroupV0_hi_18[451:450]};
  wire [7:0]        regroupV0_hi_hi_hi_20 = {regroupV0_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_3};
  wire [15:0]       regroupV0_hi_hi_20 = {regroupV0_hi_hi_hi_20, regroupV0_hi_hi_lo_20};
  wire [31:0]       regroupV0_hi_20 = {regroupV0_hi_hi_20, regroupV0_hi_lo_20};
  wire [3:0]        regroupV0_lo_lo_lo_lo_4 = {regroupV0_lo_18[37:36], regroupV0_lo_18[5:4]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_4 = {regroupV0_lo_18[101:100], regroupV0_lo_18[69:68]};
  wire [7:0]        regroupV0_lo_lo_lo_21 = {regroupV0_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_4};
  wire [3:0]        regroupV0_lo_lo_hi_lo_4 = {regroupV0_lo_18[165:164], regroupV0_lo_18[133:132]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_4 = {regroupV0_lo_18[229:228], regroupV0_lo_18[197:196]};
  wire [7:0]        regroupV0_lo_lo_hi_21 = {regroupV0_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_4};
  wire [15:0]       regroupV0_lo_lo_21 = {regroupV0_lo_lo_hi_21, regroupV0_lo_lo_lo_21};
  wire [3:0]        regroupV0_lo_hi_lo_lo_4 = {regroupV0_lo_18[293:292], regroupV0_lo_18[261:260]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_4 = {regroupV0_lo_18[357:356], regroupV0_lo_18[325:324]};
  wire [7:0]        regroupV0_lo_hi_lo_21 = {regroupV0_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_4};
  wire [3:0]        regroupV0_lo_hi_hi_lo_4 = {regroupV0_lo_18[421:420], regroupV0_lo_18[389:388]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_4 = {regroupV0_lo_18[485:484], regroupV0_lo_18[453:452]};
  wire [7:0]        regroupV0_lo_hi_hi_21 = {regroupV0_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_4};
  wire [15:0]       regroupV0_lo_hi_21 = {regroupV0_lo_hi_hi_21, regroupV0_lo_hi_lo_21};
  wire [31:0]       regroupV0_lo_21 = {regroupV0_lo_hi_21, regroupV0_lo_lo_21};
  wire [3:0]        regroupV0_hi_lo_lo_lo_4 = {regroupV0_hi_18[37:36], regroupV0_hi_18[5:4]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_4 = {regroupV0_hi_18[101:100], regroupV0_hi_18[69:68]};
  wire [7:0]        regroupV0_hi_lo_lo_21 = {regroupV0_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_4};
  wire [3:0]        regroupV0_hi_lo_hi_lo_4 = {regroupV0_hi_18[165:164], regroupV0_hi_18[133:132]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_4 = {regroupV0_hi_18[229:228], regroupV0_hi_18[197:196]};
  wire [7:0]        regroupV0_hi_lo_hi_21 = {regroupV0_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_4};
  wire [15:0]       regroupV0_hi_lo_21 = {regroupV0_hi_lo_hi_21, regroupV0_hi_lo_lo_21};
  wire [3:0]        regroupV0_hi_hi_lo_lo_4 = {regroupV0_hi_18[293:292], regroupV0_hi_18[261:260]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_4 = {regroupV0_hi_18[357:356], regroupV0_hi_18[325:324]};
  wire [7:0]        regroupV0_hi_hi_lo_21 = {regroupV0_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_4};
  wire [3:0]        regroupV0_hi_hi_hi_lo_4 = {regroupV0_hi_18[421:420], regroupV0_hi_18[389:388]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_4 = {regroupV0_hi_18[485:484], regroupV0_hi_18[453:452]};
  wire [7:0]        regroupV0_hi_hi_hi_21 = {regroupV0_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_4};
  wire [15:0]       regroupV0_hi_hi_21 = {regroupV0_hi_hi_hi_21, regroupV0_hi_hi_lo_21};
  wire [31:0]       regroupV0_hi_21 = {regroupV0_hi_hi_21, regroupV0_hi_lo_21};
  wire [3:0]        regroupV0_lo_lo_lo_lo_5 = {regroupV0_lo_18[39:38], regroupV0_lo_18[7:6]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_5 = {regroupV0_lo_18[103:102], regroupV0_lo_18[71:70]};
  wire [7:0]        regroupV0_lo_lo_lo_22 = {regroupV0_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_5};
  wire [3:0]        regroupV0_lo_lo_hi_lo_5 = {regroupV0_lo_18[167:166], regroupV0_lo_18[135:134]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_5 = {regroupV0_lo_18[231:230], regroupV0_lo_18[199:198]};
  wire [7:0]        regroupV0_lo_lo_hi_22 = {regroupV0_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_5};
  wire [15:0]       regroupV0_lo_lo_22 = {regroupV0_lo_lo_hi_22, regroupV0_lo_lo_lo_22};
  wire [3:0]        regroupV0_lo_hi_lo_lo_5 = {regroupV0_lo_18[295:294], regroupV0_lo_18[263:262]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_5 = {regroupV0_lo_18[359:358], regroupV0_lo_18[327:326]};
  wire [7:0]        regroupV0_lo_hi_lo_22 = {regroupV0_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_5};
  wire [3:0]        regroupV0_lo_hi_hi_lo_5 = {regroupV0_lo_18[423:422], regroupV0_lo_18[391:390]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_5 = {regroupV0_lo_18[487:486], regroupV0_lo_18[455:454]};
  wire [7:0]        regroupV0_lo_hi_hi_22 = {regroupV0_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_5};
  wire [15:0]       regroupV0_lo_hi_22 = {regroupV0_lo_hi_hi_22, regroupV0_lo_hi_lo_22};
  wire [31:0]       regroupV0_lo_22 = {regroupV0_lo_hi_22, regroupV0_lo_lo_22};
  wire [3:0]        regroupV0_hi_lo_lo_lo_5 = {regroupV0_hi_18[39:38], regroupV0_hi_18[7:6]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_5 = {regroupV0_hi_18[103:102], regroupV0_hi_18[71:70]};
  wire [7:0]        regroupV0_hi_lo_lo_22 = {regroupV0_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_5};
  wire [3:0]        regroupV0_hi_lo_hi_lo_5 = {regroupV0_hi_18[167:166], regroupV0_hi_18[135:134]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_5 = {regroupV0_hi_18[231:230], regroupV0_hi_18[199:198]};
  wire [7:0]        regroupV0_hi_lo_hi_22 = {regroupV0_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_5};
  wire [15:0]       regroupV0_hi_lo_22 = {regroupV0_hi_lo_hi_22, regroupV0_hi_lo_lo_22};
  wire [3:0]        regroupV0_hi_hi_lo_lo_5 = {regroupV0_hi_18[295:294], regroupV0_hi_18[263:262]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_5 = {regroupV0_hi_18[359:358], regroupV0_hi_18[327:326]};
  wire [7:0]        regroupV0_hi_hi_lo_22 = {regroupV0_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_5};
  wire [3:0]        regroupV0_hi_hi_hi_lo_5 = {regroupV0_hi_18[423:422], regroupV0_hi_18[391:390]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_5 = {regroupV0_hi_18[487:486], regroupV0_hi_18[455:454]};
  wire [7:0]        regroupV0_hi_hi_hi_22 = {regroupV0_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_5};
  wire [15:0]       regroupV0_hi_hi_22 = {regroupV0_hi_hi_hi_22, regroupV0_hi_hi_lo_22};
  wire [31:0]       regroupV0_hi_22 = {regroupV0_hi_hi_22, regroupV0_hi_lo_22};
  wire [3:0]        regroupV0_lo_lo_lo_lo_6 = {regroupV0_lo_18[41:40], regroupV0_lo_18[9:8]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_6 = {regroupV0_lo_18[105:104], regroupV0_lo_18[73:72]};
  wire [7:0]        regroupV0_lo_lo_lo_23 = {regroupV0_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_6};
  wire [3:0]        regroupV0_lo_lo_hi_lo_6 = {regroupV0_lo_18[169:168], regroupV0_lo_18[137:136]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_6 = {regroupV0_lo_18[233:232], regroupV0_lo_18[201:200]};
  wire [7:0]        regroupV0_lo_lo_hi_23 = {regroupV0_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_6};
  wire [15:0]       regroupV0_lo_lo_23 = {regroupV0_lo_lo_hi_23, regroupV0_lo_lo_lo_23};
  wire [3:0]        regroupV0_lo_hi_lo_lo_6 = {regroupV0_lo_18[297:296], regroupV0_lo_18[265:264]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_6 = {regroupV0_lo_18[361:360], regroupV0_lo_18[329:328]};
  wire [7:0]        regroupV0_lo_hi_lo_23 = {regroupV0_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_6};
  wire [3:0]        regroupV0_lo_hi_hi_lo_6 = {regroupV0_lo_18[425:424], regroupV0_lo_18[393:392]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_6 = {regroupV0_lo_18[489:488], regroupV0_lo_18[457:456]};
  wire [7:0]        regroupV0_lo_hi_hi_23 = {regroupV0_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_6};
  wire [15:0]       regroupV0_lo_hi_23 = {regroupV0_lo_hi_hi_23, regroupV0_lo_hi_lo_23};
  wire [31:0]       regroupV0_lo_23 = {regroupV0_lo_hi_23, regroupV0_lo_lo_23};
  wire [3:0]        regroupV0_hi_lo_lo_lo_6 = {regroupV0_hi_18[41:40], regroupV0_hi_18[9:8]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_6 = {regroupV0_hi_18[105:104], regroupV0_hi_18[73:72]};
  wire [7:0]        regroupV0_hi_lo_lo_23 = {regroupV0_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_6};
  wire [3:0]        regroupV0_hi_lo_hi_lo_6 = {regroupV0_hi_18[169:168], regroupV0_hi_18[137:136]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_6 = {regroupV0_hi_18[233:232], regroupV0_hi_18[201:200]};
  wire [7:0]        regroupV0_hi_lo_hi_23 = {regroupV0_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_6};
  wire [15:0]       regroupV0_hi_lo_23 = {regroupV0_hi_lo_hi_23, regroupV0_hi_lo_lo_23};
  wire [3:0]        regroupV0_hi_hi_lo_lo_6 = {regroupV0_hi_18[297:296], regroupV0_hi_18[265:264]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_6 = {regroupV0_hi_18[361:360], regroupV0_hi_18[329:328]};
  wire [7:0]        regroupV0_hi_hi_lo_23 = {regroupV0_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_6};
  wire [3:0]        regroupV0_hi_hi_hi_lo_6 = {regroupV0_hi_18[425:424], regroupV0_hi_18[393:392]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_6 = {regroupV0_hi_18[489:488], regroupV0_hi_18[457:456]};
  wire [7:0]        regroupV0_hi_hi_hi_23 = {regroupV0_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_6};
  wire [15:0]       regroupV0_hi_hi_23 = {regroupV0_hi_hi_hi_23, regroupV0_hi_hi_lo_23};
  wire [31:0]       regroupV0_hi_23 = {regroupV0_hi_hi_23, regroupV0_hi_lo_23};
  wire [3:0]        regroupV0_lo_lo_lo_lo_7 = {regroupV0_lo_18[43:42], regroupV0_lo_18[11:10]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_7 = {regroupV0_lo_18[107:106], regroupV0_lo_18[75:74]};
  wire [7:0]        regroupV0_lo_lo_lo_24 = {regroupV0_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_7};
  wire [3:0]        regroupV0_lo_lo_hi_lo_7 = {regroupV0_lo_18[171:170], regroupV0_lo_18[139:138]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_7 = {regroupV0_lo_18[235:234], regroupV0_lo_18[203:202]};
  wire [7:0]        regroupV0_lo_lo_hi_24 = {regroupV0_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_7};
  wire [15:0]       regroupV0_lo_lo_24 = {regroupV0_lo_lo_hi_24, regroupV0_lo_lo_lo_24};
  wire [3:0]        regroupV0_lo_hi_lo_lo_7 = {regroupV0_lo_18[299:298], regroupV0_lo_18[267:266]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_7 = {regroupV0_lo_18[363:362], regroupV0_lo_18[331:330]};
  wire [7:0]        regroupV0_lo_hi_lo_24 = {regroupV0_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_7};
  wire [3:0]        regroupV0_lo_hi_hi_lo_7 = {regroupV0_lo_18[427:426], regroupV0_lo_18[395:394]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_7 = {regroupV0_lo_18[491:490], regroupV0_lo_18[459:458]};
  wire [7:0]        regroupV0_lo_hi_hi_24 = {regroupV0_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_7};
  wire [15:0]       regroupV0_lo_hi_24 = {regroupV0_lo_hi_hi_24, regroupV0_lo_hi_lo_24};
  wire [31:0]       regroupV0_lo_24 = {regroupV0_lo_hi_24, regroupV0_lo_lo_24};
  wire [3:0]        regroupV0_hi_lo_lo_lo_7 = {regroupV0_hi_18[43:42], regroupV0_hi_18[11:10]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_7 = {regroupV0_hi_18[107:106], regroupV0_hi_18[75:74]};
  wire [7:0]        regroupV0_hi_lo_lo_24 = {regroupV0_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_7};
  wire [3:0]        regroupV0_hi_lo_hi_lo_7 = {regroupV0_hi_18[171:170], regroupV0_hi_18[139:138]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_7 = {regroupV0_hi_18[235:234], regroupV0_hi_18[203:202]};
  wire [7:0]        regroupV0_hi_lo_hi_24 = {regroupV0_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_7};
  wire [15:0]       regroupV0_hi_lo_24 = {regroupV0_hi_lo_hi_24, regroupV0_hi_lo_lo_24};
  wire [3:0]        regroupV0_hi_hi_lo_lo_7 = {regroupV0_hi_18[299:298], regroupV0_hi_18[267:266]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_7 = {regroupV0_hi_18[363:362], regroupV0_hi_18[331:330]};
  wire [7:0]        regroupV0_hi_hi_lo_24 = {regroupV0_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_7};
  wire [3:0]        regroupV0_hi_hi_hi_lo_7 = {regroupV0_hi_18[427:426], regroupV0_hi_18[395:394]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_7 = {regroupV0_hi_18[491:490], regroupV0_hi_18[459:458]};
  wire [7:0]        regroupV0_hi_hi_hi_24 = {regroupV0_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_7};
  wire [15:0]       regroupV0_hi_hi_24 = {regroupV0_hi_hi_hi_24, regroupV0_hi_hi_lo_24};
  wire [31:0]       regroupV0_hi_24 = {regroupV0_hi_hi_24, regroupV0_hi_lo_24};
  wire [3:0]        regroupV0_lo_lo_lo_lo_8 = {regroupV0_lo_18[45:44], regroupV0_lo_18[13:12]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_8 = {regroupV0_lo_18[109:108], regroupV0_lo_18[77:76]};
  wire [7:0]        regroupV0_lo_lo_lo_25 = {regroupV0_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_8};
  wire [3:0]        regroupV0_lo_lo_hi_lo_8 = {regroupV0_lo_18[173:172], regroupV0_lo_18[141:140]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_8 = {regroupV0_lo_18[237:236], regroupV0_lo_18[205:204]};
  wire [7:0]        regroupV0_lo_lo_hi_25 = {regroupV0_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_8};
  wire [15:0]       regroupV0_lo_lo_25 = {regroupV0_lo_lo_hi_25, regroupV0_lo_lo_lo_25};
  wire [3:0]        regroupV0_lo_hi_lo_lo_8 = {regroupV0_lo_18[301:300], regroupV0_lo_18[269:268]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_8 = {regroupV0_lo_18[365:364], regroupV0_lo_18[333:332]};
  wire [7:0]        regroupV0_lo_hi_lo_25 = {regroupV0_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_8};
  wire [3:0]        regroupV0_lo_hi_hi_lo_8 = {regroupV0_lo_18[429:428], regroupV0_lo_18[397:396]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_8 = {regroupV0_lo_18[493:492], regroupV0_lo_18[461:460]};
  wire [7:0]        regroupV0_lo_hi_hi_25 = {regroupV0_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_8};
  wire [15:0]       regroupV0_lo_hi_25 = {regroupV0_lo_hi_hi_25, regroupV0_lo_hi_lo_25};
  wire [31:0]       regroupV0_lo_25 = {regroupV0_lo_hi_25, regroupV0_lo_lo_25};
  wire [3:0]        regroupV0_hi_lo_lo_lo_8 = {regroupV0_hi_18[45:44], regroupV0_hi_18[13:12]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_8 = {regroupV0_hi_18[109:108], regroupV0_hi_18[77:76]};
  wire [7:0]        regroupV0_hi_lo_lo_25 = {regroupV0_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_8};
  wire [3:0]        regroupV0_hi_lo_hi_lo_8 = {regroupV0_hi_18[173:172], regroupV0_hi_18[141:140]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_8 = {regroupV0_hi_18[237:236], regroupV0_hi_18[205:204]};
  wire [7:0]        regroupV0_hi_lo_hi_25 = {regroupV0_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_8};
  wire [15:0]       regroupV0_hi_lo_25 = {regroupV0_hi_lo_hi_25, regroupV0_hi_lo_lo_25};
  wire [3:0]        regroupV0_hi_hi_lo_lo_8 = {regroupV0_hi_18[301:300], regroupV0_hi_18[269:268]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_8 = {regroupV0_hi_18[365:364], regroupV0_hi_18[333:332]};
  wire [7:0]        regroupV0_hi_hi_lo_25 = {regroupV0_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_8};
  wire [3:0]        regroupV0_hi_hi_hi_lo_8 = {regroupV0_hi_18[429:428], regroupV0_hi_18[397:396]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_8 = {regroupV0_hi_18[493:492], regroupV0_hi_18[461:460]};
  wire [7:0]        regroupV0_hi_hi_hi_25 = {regroupV0_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_8};
  wire [15:0]       regroupV0_hi_hi_25 = {regroupV0_hi_hi_hi_25, regroupV0_hi_hi_lo_25};
  wire [31:0]       regroupV0_hi_25 = {regroupV0_hi_hi_25, regroupV0_hi_lo_25};
  wire [3:0]        regroupV0_lo_lo_lo_lo_9 = {regroupV0_lo_18[47:46], regroupV0_lo_18[15:14]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_9 = {regroupV0_lo_18[111:110], regroupV0_lo_18[79:78]};
  wire [7:0]        regroupV0_lo_lo_lo_26 = {regroupV0_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_9};
  wire [3:0]        regroupV0_lo_lo_hi_lo_9 = {regroupV0_lo_18[175:174], regroupV0_lo_18[143:142]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_9 = {regroupV0_lo_18[239:238], regroupV0_lo_18[207:206]};
  wire [7:0]        regroupV0_lo_lo_hi_26 = {regroupV0_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_9};
  wire [15:0]       regroupV0_lo_lo_26 = {regroupV0_lo_lo_hi_26, regroupV0_lo_lo_lo_26};
  wire [3:0]        regroupV0_lo_hi_lo_lo_9 = {regroupV0_lo_18[303:302], regroupV0_lo_18[271:270]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_9 = {regroupV0_lo_18[367:366], regroupV0_lo_18[335:334]};
  wire [7:0]        regroupV0_lo_hi_lo_26 = {regroupV0_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_9};
  wire [3:0]        regroupV0_lo_hi_hi_lo_9 = {regroupV0_lo_18[431:430], regroupV0_lo_18[399:398]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_9 = {regroupV0_lo_18[495:494], regroupV0_lo_18[463:462]};
  wire [7:0]        regroupV0_lo_hi_hi_26 = {regroupV0_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_9};
  wire [15:0]       regroupV0_lo_hi_26 = {regroupV0_lo_hi_hi_26, regroupV0_lo_hi_lo_26};
  wire [31:0]       regroupV0_lo_26 = {regroupV0_lo_hi_26, regroupV0_lo_lo_26};
  wire [3:0]        regroupV0_hi_lo_lo_lo_9 = {regroupV0_hi_18[47:46], regroupV0_hi_18[15:14]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_9 = {regroupV0_hi_18[111:110], regroupV0_hi_18[79:78]};
  wire [7:0]        regroupV0_hi_lo_lo_26 = {regroupV0_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_9};
  wire [3:0]        regroupV0_hi_lo_hi_lo_9 = {regroupV0_hi_18[175:174], regroupV0_hi_18[143:142]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_9 = {regroupV0_hi_18[239:238], regroupV0_hi_18[207:206]};
  wire [7:0]        regroupV0_hi_lo_hi_26 = {regroupV0_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_9};
  wire [15:0]       regroupV0_hi_lo_26 = {regroupV0_hi_lo_hi_26, regroupV0_hi_lo_lo_26};
  wire [3:0]        regroupV0_hi_hi_lo_lo_9 = {regroupV0_hi_18[303:302], regroupV0_hi_18[271:270]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_9 = {regroupV0_hi_18[367:366], regroupV0_hi_18[335:334]};
  wire [7:0]        regroupV0_hi_hi_lo_26 = {regroupV0_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_9};
  wire [3:0]        regroupV0_hi_hi_hi_lo_9 = {regroupV0_hi_18[431:430], regroupV0_hi_18[399:398]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_9 = {regroupV0_hi_18[495:494], regroupV0_hi_18[463:462]};
  wire [7:0]        regroupV0_hi_hi_hi_26 = {regroupV0_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_9};
  wire [15:0]       regroupV0_hi_hi_26 = {regroupV0_hi_hi_hi_26, regroupV0_hi_hi_lo_26};
  wire [31:0]       regroupV0_hi_26 = {regroupV0_hi_hi_26, regroupV0_hi_lo_26};
  wire [3:0]        regroupV0_lo_lo_lo_lo_10 = {regroupV0_lo_18[49:48], regroupV0_lo_18[17:16]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_10 = {regroupV0_lo_18[113:112], regroupV0_lo_18[81:80]};
  wire [7:0]        regroupV0_lo_lo_lo_27 = {regroupV0_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_10};
  wire [3:0]        regroupV0_lo_lo_hi_lo_10 = {regroupV0_lo_18[177:176], regroupV0_lo_18[145:144]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_10 = {regroupV0_lo_18[241:240], regroupV0_lo_18[209:208]};
  wire [7:0]        regroupV0_lo_lo_hi_27 = {regroupV0_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_10};
  wire [15:0]       regroupV0_lo_lo_27 = {regroupV0_lo_lo_hi_27, regroupV0_lo_lo_lo_27};
  wire [3:0]        regroupV0_lo_hi_lo_lo_10 = {regroupV0_lo_18[305:304], regroupV0_lo_18[273:272]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_10 = {regroupV0_lo_18[369:368], regroupV0_lo_18[337:336]};
  wire [7:0]        regroupV0_lo_hi_lo_27 = {regroupV0_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_10};
  wire [3:0]        regroupV0_lo_hi_hi_lo_10 = {regroupV0_lo_18[433:432], regroupV0_lo_18[401:400]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_10 = {regroupV0_lo_18[497:496], regroupV0_lo_18[465:464]};
  wire [7:0]        regroupV0_lo_hi_hi_27 = {regroupV0_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_10};
  wire [15:0]       regroupV0_lo_hi_27 = {regroupV0_lo_hi_hi_27, regroupV0_lo_hi_lo_27};
  wire [31:0]       regroupV0_lo_27 = {regroupV0_lo_hi_27, regroupV0_lo_lo_27};
  wire [3:0]        regroupV0_hi_lo_lo_lo_10 = {regroupV0_hi_18[49:48], regroupV0_hi_18[17:16]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_10 = {regroupV0_hi_18[113:112], regroupV0_hi_18[81:80]};
  wire [7:0]        regroupV0_hi_lo_lo_27 = {regroupV0_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_10};
  wire [3:0]        regroupV0_hi_lo_hi_lo_10 = {regroupV0_hi_18[177:176], regroupV0_hi_18[145:144]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_10 = {regroupV0_hi_18[241:240], regroupV0_hi_18[209:208]};
  wire [7:0]        regroupV0_hi_lo_hi_27 = {regroupV0_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_10};
  wire [15:0]       regroupV0_hi_lo_27 = {regroupV0_hi_lo_hi_27, regroupV0_hi_lo_lo_27};
  wire [3:0]        regroupV0_hi_hi_lo_lo_10 = {regroupV0_hi_18[305:304], regroupV0_hi_18[273:272]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_10 = {regroupV0_hi_18[369:368], regroupV0_hi_18[337:336]};
  wire [7:0]        regroupV0_hi_hi_lo_27 = {regroupV0_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_10};
  wire [3:0]        regroupV0_hi_hi_hi_lo_10 = {regroupV0_hi_18[433:432], regroupV0_hi_18[401:400]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_10 = {regroupV0_hi_18[497:496], regroupV0_hi_18[465:464]};
  wire [7:0]        regroupV0_hi_hi_hi_27 = {regroupV0_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_10};
  wire [15:0]       regroupV0_hi_hi_27 = {regroupV0_hi_hi_hi_27, regroupV0_hi_hi_lo_27};
  wire [31:0]       regroupV0_hi_27 = {regroupV0_hi_hi_27, regroupV0_hi_lo_27};
  wire [3:0]        regroupV0_lo_lo_lo_lo_11 = {regroupV0_lo_18[51:50], regroupV0_lo_18[19:18]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_11 = {regroupV0_lo_18[115:114], regroupV0_lo_18[83:82]};
  wire [7:0]        regroupV0_lo_lo_lo_28 = {regroupV0_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_11};
  wire [3:0]        regroupV0_lo_lo_hi_lo_11 = {regroupV0_lo_18[179:178], regroupV0_lo_18[147:146]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_11 = {regroupV0_lo_18[243:242], regroupV0_lo_18[211:210]};
  wire [7:0]        regroupV0_lo_lo_hi_28 = {regroupV0_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_11};
  wire [15:0]       regroupV0_lo_lo_28 = {regroupV0_lo_lo_hi_28, regroupV0_lo_lo_lo_28};
  wire [3:0]        regroupV0_lo_hi_lo_lo_11 = {regroupV0_lo_18[307:306], regroupV0_lo_18[275:274]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_11 = {regroupV0_lo_18[371:370], regroupV0_lo_18[339:338]};
  wire [7:0]        regroupV0_lo_hi_lo_28 = {regroupV0_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_11};
  wire [3:0]        regroupV0_lo_hi_hi_lo_11 = {regroupV0_lo_18[435:434], regroupV0_lo_18[403:402]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_11 = {regroupV0_lo_18[499:498], regroupV0_lo_18[467:466]};
  wire [7:0]        regroupV0_lo_hi_hi_28 = {regroupV0_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_11};
  wire [15:0]       regroupV0_lo_hi_28 = {regroupV0_lo_hi_hi_28, regroupV0_lo_hi_lo_28};
  wire [31:0]       regroupV0_lo_28 = {regroupV0_lo_hi_28, regroupV0_lo_lo_28};
  wire [3:0]        regroupV0_hi_lo_lo_lo_11 = {regroupV0_hi_18[51:50], regroupV0_hi_18[19:18]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_11 = {regroupV0_hi_18[115:114], regroupV0_hi_18[83:82]};
  wire [7:0]        regroupV0_hi_lo_lo_28 = {regroupV0_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_11};
  wire [3:0]        regroupV0_hi_lo_hi_lo_11 = {regroupV0_hi_18[179:178], regroupV0_hi_18[147:146]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_11 = {regroupV0_hi_18[243:242], regroupV0_hi_18[211:210]};
  wire [7:0]        regroupV0_hi_lo_hi_28 = {regroupV0_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_11};
  wire [15:0]       regroupV0_hi_lo_28 = {regroupV0_hi_lo_hi_28, regroupV0_hi_lo_lo_28};
  wire [3:0]        regroupV0_hi_hi_lo_lo_11 = {regroupV0_hi_18[307:306], regroupV0_hi_18[275:274]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_11 = {regroupV0_hi_18[371:370], regroupV0_hi_18[339:338]};
  wire [7:0]        regroupV0_hi_hi_lo_28 = {regroupV0_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_11};
  wire [3:0]        regroupV0_hi_hi_hi_lo_11 = {regroupV0_hi_18[435:434], regroupV0_hi_18[403:402]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_11 = {regroupV0_hi_18[499:498], regroupV0_hi_18[467:466]};
  wire [7:0]        regroupV0_hi_hi_hi_28 = {regroupV0_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_11};
  wire [15:0]       regroupV0_hi_hi_28 = {regroupV0_hi_hi_hi_28, regroupV0_hi_hi_lo_28};
  wire [31:0]       regroupV0_hi_28 = {regroupV0_hi_hi_28, regroupV0_hi_lo_28};
  wire [3:0]        regroupV0_lo_lo_lo_lo_12 = {regroupV0_lo_18[53:52], regroupV0_lo_18[21:20]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_12 = {regroupV0_lo_18[117:116], regroupV0_lo_18[85:84]};
  wire [7:0]        regroupV0_lo_lo_lo_29 = {regroupV0_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_12};
  wire [3:0]        regroupV0_lo_lo_hi_lo_12 = {regroupV0_lo_18[181:180], regroupV0_lo_18[149:148]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_12 = {regroupV0_lo_18[245:244], regroupV0_lo_18[213:212]};
  wire [7:0]        regroupV0_lo_lo_hi_29 = {regroupV0_lo_lo_hi_hi_12, regroupV0_lo_lo_hi_lo_12};
  wire [15:0]       regroupV0_lo_lo_29 = {regroupV0_lo_lo_hi_29, regroupV0_lo_lo_lo_29};
  wire [3:0]        regroupV0_lo_hi_lo_lo_12 = {regroupV0_lo_18[309:308], regroupV0_lo_18[277:276]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_12 = {regroupV0_lo_18[373:372], regroupV0_lo_18[341:340]};
  wire [7:0]        regroupV0_lo_hi_lo_29 = {regroupV0_lo_hi_lo_hi_12, regroupV0_lo_hi_lo_lo_12};
  wire [3:0]        regroupV0_lo_hi_hi_lo_12 = {regroupV0_lo_18[437:436], regroupV0_lo_18[405:404]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_12 = {regroupV0_lo_18[501:500], regroupV0_lo_18[469:468]};
  wire [7:0]        regroupV0_lo_hi_hi_29 = {regroupV0_lo_hi_hi_hi_12, regroupV0_lo_hi_hi_lo_12};
  wire [15:0]       regroupV0_lo_hi_29 = {regroupV0_lo_hi_hi_29, regroupV0_lo_hi_lo_29};
  wire [31:0]       regroupV0_lo_29 = {regroupV0_lo_hi_29, regroupV0_lo_lo_29};
  wire [3:0]        regroupV0_hi_lo_lo_lo_12 = {regroupV0_hi_18[53:52], regroupV0_hi_18[21:20]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_12 = {regroupV0_hi_18[117:116], regroupV0_hi_18[85:84]};
  wire [7:0]        regroupV0_hi_lo_lo_29 = {regroupV0_hi_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_12};
  wire [3:0]        regroupV0_hi_lo_hi_lo_12 = {regroupV0_hi_18[181:180], regroupV0_hi_18[149:148]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_12 = {regroupV0_hi_18[245:244], regroupV0_hi_18[213:212]};
  wire [7:0]        regroupV0_hi_lo_hi_29 = {regroupV0_hi_lo_hi_hi_12, regroupV0_hi_lo_hi_lo_12};
  wire [15:0]       regroupV0_hi_lo_29 = {regroupV0_hi_lo_hi_29, regroupV0_hi_lo_lo_29};
  wire [3:0]        regroupV0_hi_hi_lo_lo_12 = {regroupV0_hi_18[309:308], regroupV0_hi_18[277:276]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_12 = {regroupV0_hi_18[373:372], regroupV0_hi_18[341:340]};
  wire [7:0]        regroupV0_hi_hi_lo_29 = {regroupV0_hi_hi_lo_hi_12, regroupV0_hi_hi_lo_lo_12};
  wire [3:0]        regroupV0_hi_hi_hi_lo_12 = {regroupV0_hi_18[437:436], regroupV0_hi_18[405:404]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_12 = {regroupV0_hi_18[501:500], regroupV0_hi_18[469:468]};
  wire [7:0]        regroupV0_hi_hi_hi_29 = {regroupV0_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_lo_12};
  wire [15:0]       regroupV0_hi_hi_29 = {regroupV0_hi_hi_hi_29, regroupV0_hi_hi_lo_29};
  wire [31:0]       regroupV0_hi_29 = {regroupV0_hi_hi_29, regroupV0_hi_lo_29};
  wire [3:0]        regroupV0_lo_lo_lo_lo_13 = {regroupV0_lo_18[55:54], regroupV0_lo_18[23:22]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_13 = {regroupV0_lo_18[119:118], regroupV0_lo_18[87:86]};
  wire [7:0]        regroupV0_lo_lo_lo_30 = {regroupV0_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_13};
  wire [3:0]        regroupV0_lo_lo_hi_lo_13 = {regroupV0_lo_18[183:182], regroupV0_lo_18[151:150]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_13 = {regroupV0_lo_18[247:246], regroupV0_lo_18[215:214]};
  wire [7:0]        regroupV0_lo_lo_hi_30 = {regroupV0_lo_lo_hi_hi_13, regroupV0_lo_lo_hi_lo_13};
  wire [15:0]       regroupV0_lo_lo_30 = {regroupV0_lo_lo_hi_30, regroupV0_lo_lo_lo_30};
  wire [3:0]        regroupV0_lo_hi_lo_lo_13 = {regroupV0_lo_18[311:310], regroupV0_lo_18[279:278]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_13 = {regroupV0_lo_18[375:374], regroupV0_lo_18[343:342]};
  wire [7:0]        regroupV0_lo_hi_lo_30 = {regroupV0_lo_hi_lo_hi_13, regroupV0_lo_hi_lo_lo_13};
  wire [3:0]        regroupV0_lo_hi_hi_lo_13 = {regroupV0_lo_18[439:438], regroupV0_lo_18[407:406]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_13 = {regroupV0_lo_18[503:502], regroupV0_lo_18[471:470]};
  wire [7:0]        regroupV0_lo_hi_hi_30 = {regroupV0_lo_hi_hi_hi_13, regroupV0_lo_hi_hi_lo_13};
  wire [15:0]       regroupV0_lo_hi_30 = {regroupV0_lo_hi_hi_30, regroupV0_lo_hi_lo_30};
  wire [31:0]       regroupV0_lo_30 = {regroupV0_lo_hi_30, regroupV0_lo_lo_30};
  wire [3:0]        regroupV0_hi_lo_lo_lo_13 = {regroupV0_hi_18[55:54], regroupV0_hi_18[23:22]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_13 = {regroupV0_hi_18[119:118], regroupV0_hi_18[87:86]};
  wire [7:0]        regroupV0_hi_lo_lo_30 = {regroupV0_hi_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_13};
  wire [3:0]        regroupV0_hi_lo_hi_lo_13 = {regroupV0_hi_18[183:182], regroupV0_hi_18[151:150]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_13 = {regroupV0_hi_18[247:246], regroupV0_hi_18[215:214]};
  wire [7:0]        regroupV0_hi_lo_hi_30 = {regroupV0_hi_lo_hi_hi_13, regroupV0_hi_lo_hi_lo_13};
  wire [15:0]       regroupV0_hi_lo_30 = {regroupV0_hi_lo_hi_30, regroupV0_hi_lo_lo_30};
  wire [3:0]        regroupV0_hi_hi_lo_lo_13 = {regroupV0_hi_18[311:310], regroupV0_hi_18[279:278]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_13 = {regroupV0_hi_18[375:374], regroupV0_hi_18[343:342]};
  wire [7:0]        regroupV0_hi_hi_lo_30 = {regroupV0_hi_hi_lo_hi_13, regroupV0_hi_hi_lo_lo_13};
  wire [3:0]        regroupV0_hi_hi_hi_lo_13 = {regroupV0_hi_18[439:438], regroupV0_hi_18[407:406]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_13 = {regroupV0_hi_18[503:502], regroupV0_hi_18[471:470]};
  wire [7:0]        regroupV0_hi_hi_hi_30 = {regroupV0_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_lo_13};
  wire [15:0]       regroupV0_hi_hi_30 = {regroupV0_hi_hi_hi_30, regroupV0_hi_hi_lo_30};
  wire [31:0]       regroupV0_hi_30 = {regroupV0_hi_hi_30, regroupV0_hi_lo_30};
  wire [3:0]        regroupV0_lo_lo_lo_lo_14 = {regroupV0_lo_18[57:56], regroupV0_lo_18[25:24]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_14 = {regroupV0_lo_18[121:120], regroupV0_lo_18[89:88]};
  wire [7:0]        regroupV0_lo_lo_lo_31 = {regroupV0_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_14};
  wire [3:0]        regroupV0_lo_lo_hi_lo_14 = {regroupV0_lo_18[185:184], regroupV0_lo_18[153:152]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_14 = {regroupV0_lo_18[249:248], regroupV0_lo_18[217:216]};
  wire [7:0]        regroupV0_lo_lo_hi_31 = {regroupV0_lo_lo_hi_hi_14, regroupV0_lo_lo_hi_lo_14};
  wire [15:0]       regroupV0_lo_lo_31 = {regroupV0_lo_lo_hi_31, regroupV0_lo_lo_lo_31};
  wire [3:0]        regroupV0_lo_hi_lo_lo_14 = {regroupV0_lo_18[313:312], regroupV0_lo_18[281:280]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_14 = {regroupV0_lo_18[377:376], regroupV0_lo_18[345:344]};
  wire [7:0]        regroupV0_lo_hi_lo_31 = {regroupV0_lo_hi_lo_hi_14, regroupV0_lo_hi_lo_lo_14};
  wire [3:0]        regroupV0_lo_hi_hi_lo_14 = {regroupV0_lo_18[441:440], regroupV0_lo_18[409:408]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_14 = {regroupV0_lo_18[505:504], regroupV0_lo_18[473:472]};
  wire [7:0]        regroupV0_lo_hi_hi_31 = {regroupV0_lo_hi_hi_hi_14, regroupV0_lo_hi_hi_lo_14};
  wire [15:0]       regroupV0_lo_hi_31 = {regroupV0_lo_hi_hi_31, regroupV0_lo_hi_lo_31};
  wire [31:0]       regroupV0_lo_31 = {regroupV0_lo_hi_31, regroupV0_lo_lo_31};
  wire [3:0]        regroupV0_hi_lo_lo_lo_14 = {regroupV0_hi_18[57:56], regroupV0_hi_18[25:24]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_14 = {regroupV0_hi_18[121:120], regroupV0_hi_18[89:88]};
  wire [7:0]        regroupV0_hi_lo_lo_31 = {regroupV0_hi_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_14};
  wire [3:0]        regroupV0_hi_lo_hi_lo_14 = {regroupV0_hi_18[185:184], regroupV0_hi_18[153:152]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_14 = {regroupV0_hi_18[249:248], regroupV0_hi_18[217:216]};
  wire [7:0]        regroupV0_hi_lo_hi_31 = {regroupV0_hi_lo_hi_hi_14, regroupV0_hi_lo_hi_lo_14};
  wire [15:0]       regroupV0_hi_lo_31 = {regroupV0_hi_lo_hi_31, regroupV0_hi_lo_lo_31};
  wire [3:0]        regroupV0_hi_hi_lo_lo_14 = {regroupV0_hi_18[313:312], regroupV0_hi_18[281:280]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_14 = {regroupV0_hi_18[377:376], regroupV0_hi_18[345:344]};
  wire [7:0]        regroupV0_hi_hi_lo_31 = {regroupV0_hi_hi_lo_hi_14, regroupV0_hi_hi_lo_lo_14};
  wire [3:0]        regroupV0_hi_hi_hi_lo_14 = {regroupV0_hi_18[441:440], regroupV0_hi_18[409:408]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_14 = {regroupV0_hi_18[505:504], regroupV0_hi_18[473:472]};
  wire [7:0]        regroupV0_hi_hi_hi_31 = {regroupV0_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_lo_14};
  wire [15:0]       regroupV0_hi_hi_31 = {regroupV0_hi_hi_hi_31, regroupV0_hi_hi_lo_31};
  wire [31:0]       regroupV0_hi_31 = {regroupV0_hi_hi_31, regroupV0_hi_lo_31};
  wire [3:0]        regroupV0_lo_lo_lo_lo_15 = {regroupV0_lo_18[59:58], regroupV0_lo_18[27:26]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_15 = {regroupV0_lo_18[123:122], regroupV0_lo_18[91:90]};
  wire [7:0]        regroupV0_lo_lo_lo_32 = {regroupV0_lo_lo_lo_hi_15, regroupV0_lo_lo_lo_lo_15};
  wire [3:0]        regroupV0_lo_lo_hi_lo_15 = {regroupV0_lo_18[187:186], regroupV0_lo_18[155:154]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_15 = {regroupV0_lo_18[251:250], regroupV0_lo_18[219:218]};
  wire [7:0]        regroupV0_lo_lo_hi_32 = {regroupV0_lo_lo_hi_hi_15, regroupV0_lo_lo_hi_lo_15};
  wire [15:0]       regroupV0_lo_lo_32 = {regroupV0_lo_lo_hi_32, regroupV0_lo_lo_lo_32};
  wire [3:0]        regroupV0_lo_hi_lo_lo_15 = {regroupV0_lo_18[315:314], regroupV0_lo_18[283:282]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_15 = {regroupV0_lo_18[379:378], regroupV0_lo_18[347:346]};
  wire [7:0]        regroupV0_lo_hi_lo_32 = {regroupV0_lo_hi_lo_hi_15, regroupV0_lo_hi_lo_lo_15};
  wire [3:0]        regroupV0_lo_hi_hi_lo_15 = {regroupV0_lo_18[443:442], regroupV0_lo_18[411:410]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_15 = {regroupV0_lo_18[507:506], regroupV0_lo_18[475:474]};
  wire [7:0]        regroupV0_lo_hi_hi_32 = {regroupV0_lo_hi_hi_hi_15, regroupV0_lo_hi_hi_lo_15};
  wire [15:0]       regroupV0_lo_hi_32 = {regroupV0_lo_hi_hi_32, regroupV0_lo_hi_lo_32};
  wire [31:0]       regroupV0_lo_32 = {regroupV0_lo_hi_32, regroupV0_lo_lo_32};
  wire [3:0]        regroupV0_hi_lo_lo_lo_15 = {regroupV0_hi_18[59:58], regroupV0_hi_18[27:26]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_15 = {regroupV0_hi_18[123:122], regroupV0_hi_18[91:90]};
  wire [7:0]        regroupV0_hi_lo_lo_32 = {regroupV0_hi_lo_lo_hi_15, regroupV0_hi_lo_lo_lo_15};
  wire [3:0]        regroupV0_hi_lo_hi_lo_15 = {regroupV0_hi_18[187:186], regroupV0_hi_18[155:154]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_15 = {regroupV0_hi_18[251:250], regroupV0_hi_18[219:218]};
  wire [7:0]        regroupV0_hi_lo_hi_32 = {regroupV0_hi_lo_hi_hi_15, regroupV0_hi_lo_hi_lo_15};
  wire [15:0]       regroupV0_hi_lo_32 = {regroupV0_hi_lo_hi_32, regroupV0_hi_lo_lo_32};
  wire [3:0]        regroupV0_hi_hi_lo_lo_15 = {regroupV0_hi_18[315:314], regroupV0_hi_18[283:282]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_15 = {regroupV0_hi_18[379:378], regroupV0_hi_18[347:346]};
  wire [7:0]        regroupV0_hi_hi_lo_32 = {regroupV0_hi_hi_lo_hi_15, regroupV0_hi_hi_lo_lo_15};
  wire [3:0]        regroupV0_hi_hi_hi_lo_15 = {regroupV0_hi_18[443:442], regroupV0_hi_18[411:410]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_15 = {regroupV0_hi_18[507:506], regroupV0_hi_18[475:474]};
  wire [7:0]        regroupV0_hi_hi_hi_32 = {regroupV0_hi_hi_hi_hi_15, regroupV0_hi_hi_hi_lo_15};
  wire [15:0]       regroupV0_hi_hi_32 = {regroupV0_hi_hi_hi_32, regroupV0_hi_hi_lo_32};
  wire [31:0]       regroupV0_hi_32 = {regroupV0_hi_hi_32, regroupV0_hi_lo_32};
  wire [3:0]        regroupV0_lo_lo_lo_lo_16 = {regroupV0_lo_18[61:60], regroupV0_lo_18[29:28]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_16 = {regroupV0_lo_18[125:124], regroupV0_lo_18[93:92]};
  wire [7:0]        regroupV0_lo_lo_lo_33 = {regroupV0_lo_lo_lo_hi_16, regroupV0_lo_lo_lo_lo_16};
  wire [3:0]        regroupV0_lo_lo_hi_lo_16 = {regroupV0_lo_18[189:188], regroupV0_lo_18[157:156]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_16 = {regroupV0_lo_18[253:252], regroupV0_lo_18[221:220]};
  wire [7:0]        regroupV0_lo_lo_hi_33 = {regroupV0_lo_lo_hi_hi_16, regroupV0_lo_lo_hi_lo_16};
  wire [15:0]       regroupV0_lo_lo_33 = {regroupV0_lo_lo_hi_33, regroupV0_lo_lo_lo_33};
  wire [3:0]        regroupV0_lo_hi_lo_lo_16 = {regroupV0_lo_18[317:316], regroupV0_lo_18[285:284]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_16 = {regroupV0_lo_18[381:380], regroupV0_lo_18[349:348]};
  wire [7:0]        regroupV0_lo_hi_lo_33 = {regroupV0_lo_hi_lo_hi_16, regroupV0_lo_hi_lo_lo_16};
  wire [3:0]        regroupV0_lo_hi_hi_lo_16 = {regroupV0_lo_18[445:444], regroupV0_lo_18[413:412]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_16 = {regroupV0_lo_18[509:508], regroupV0_lo_18[477:476]};
  wire [7:0]        regroupV0_lo_hi_hi_33 = {regroupV0_lo_hi_hi_hi_16, regroupV0_lo_hi_hi_lo_16};
  wire [15:0]       regroupV0_lo_hi_33 = {regroupV0_lo_hi_hi_33, regroupV0_lo_hi_lo_33};
  wire [31:0]       regroupV0_lo_33 = {regroupV0_lo_hi_33, regroupV0_lo_lo_33};
  wire [3:0]        regroupV0_hi_lo_lo_lo_16 = {regroupV0_hi_18[61:60], regroupV0_hi_18[29:28]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_16 = {regroupV0_hi_18[125:124], regroupV0_hi_18[93:92]};
  wire [7:0]        regroupV0_hi_lo_lo_33 = {regroupV0_hi_lo_lo_hi_16, regroupV0_hi_lo_lo_lo_16};
  wire [3:0]        regroupV0_hi_lo_hi_lo_16 = {regroupV0_hi_18[189:188], regroupV0_hi_18[157:156]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_16 = {regroupV0_hi_18[253:252], regroupV0_hi_18[221:220]};
  wire [7:0]        regroupV0_hi_lo_hi_33 = {regroupV0_hi_lo_hi_hi_16, regroupV0_hi_lo_hi_lo_16};
  wire [15:0]       regroupV0_hi_lo_33 = {regroupV0_hi_lo_hi_33, regroupV0_hi_lo_lo_33};
  wire [3:0]        regroupV0_hi_hi_lo_lo_16 = {regroupV0_hi_18[317:316], regroupV0_hi_18[285:284]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_16 = {regroupV0_hi_18[381:380], regroupV0_hi_18[349:348]};
  wire [7:0]        regroupV0_hi_hi_lo_33 = {regroupV0_hi_hi_lo_hi_16, regroupV0_hi_hi_lo_lo_16};
  wire [3:0]        regroupV0_hi_hi_hi_lo_16 = {regroupV0_hi_18[445:444], regroupV0_hi_18[413:412]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_16 = {regroupV0_hi_18[509:508], regroupV0_hi_18[477:476]};
  wire [7:0]        regroupV0_hi_hi_hi_33 = {regroupV0_hi_hi_hi_hi_16, regroupV0_hi_hi_hi_lo_16};
  wire [15:0]       regroupV0_hi_hi_33 = {regroupV0_hi_hi_hi_33, regroupV0_hi_hi_lo_33};
  wire [31:0]       regroupV0_hi_33 = {regroupV0_hi_hi_33, regroupV0_hi_lo_33};
  wire [3:0]        regroupV0_lo_lo_lo_lo_17 = {regroupV0_lo_18[63:62], regroupV0_lo_18[31:30]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_17 = {regroupV0_lo_18[127:126], regroupV0_lo_18[95:94]};
  wire [7:0]        regroupV0_lo_lo_lo_34 = {regroupV0_lo_lo_lo_hi_17, regroupV0_lo_lo_lo_lo_17};
  wire [3:0]        regroupV0_lo_lo_hi_lo_17 = {regroupV0_lo_18[191:190], regroupV0_lo_18[159:158]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_17 = {regroupV0_lo_18[255:254], regroupV0_lo_18[223:222]};
  wire [7:0]        regroupV0_lo_lo_hi_34 = {regroupV0_lo_lo_hi_hi_17, regroupV0_lo_lo_hi_lo_17};
  wire [15:0]       regroupV0_lo_lo_34 = {regroupV0_lo_lo_hi_34, regroupV0_lo_lo_lo_34};
  wire [3:0]        regroupV0_lo_hi_lo_lo_17 = {regroupV0_lo_18[319:318], regroupV0_lo_18[287:286]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_17 = {regroupV0_lo_18[383:382], regroupV0_lo_18[351:350]};
  wire [7:0]        regroupV0_lo_hi_lo_34 = {regroupV0_lo_hi_lo_hi_17, regroupV0_lo_hi_lo_lo_17};
  wire [3:0]        regroupV0_lo_hi_hi_lo_17 = {regroupV0_lo_18[447:446], regroupV0_lo_18[415:414]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_17 = {regroupV0_lo_18[511:510], regroupV0_lo_18[479:478]};
  wire [7:0]        regroupV0_lo_hi_hi_34 = {regroupV0_lo_hi_hi_hi_17, regroupV0_lo_hi_hi_lo_17};
  wire [15:0]       regroupV0_lo_hi_34 = {regroupV0_lo_hi_hi_34, regroupV0_lo_hi_lo_34};
  wire [31:0]       regroupV0_lo_34 = {regroupV0_lo_hi_34, regroupV0_lo_lo_34};
  wire [3:0]        regroupV0_hi_lo_lo_lo_17 = {regroupV0_hi_18[63:62], regroupV0_hi_18[31:30]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_17 = {regroupV0_hi_18[127:126], regroupV0_hi_18[95:94]};
  wire [7:0]        regroupV0_hi_lo_lo_34 = {regroupV0_hi_lo_lo_hi_17, regroupV0_hi_lo_lo_lo_17};
  wire [3:0]        regroupV0_hi_lo_hi_lo_17 = {regroupV0_hi_18[191:190], regroupV0_hi_18[159:158]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_17 = {regroupV0_hi_18[255:254], regroupV0_hi_18[223:222]};
  wire [7:0]        regroupV0_hi_lo_hi_34 = {regroupV0_hi_lo_hi_hi_17, regroupV0_hi_lo_hi_lo_17};
  wire [15:0]       regroupV0_hi_lo_34 = {regroupV0_hi_lo_hi_34, regroupV0_hi_lo_lo_34};
  wire [3:0]        regroupV0_hi_hi_lo_lo_17 = {regroupV0_hi_18[319:318], regroupV0_hi_18[287:286]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_17 = {regroupV0_hi_18[383:382], regroupV0_hi_18[351:350]};
  wire [7:0]        regroupV0_hi_hi_lo_34 = {regroupV0_hi_hi_lo_hi_17, regroupV0_hi_hi_lo_lo_17};
  wire [3:0]        regroupV0_hi_hi_hi_lo_17 = {regroupV0_hi_18[447:446], regroupV0_hi_18[415:414]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_17 = {regroupV0_hi_18[511:510], regroupV0_hi_18[479:478]};
  wire [7:0]        regroupV0_hi_hi_hi_34 = {regroupV0_hi_hi_hi_hi_17, regroupV0_hi_hi_hi_lo_17};
  wire [15:0]       regroupV0_hi_hi_34 = {regroupV0_hi_hi_hi_34, regroupV0_hi_hi_lo_34};
  wire [31:0]       regroupV0_hi_34 = {regroupV0_hi_hi_34, regroupV0_hi_lo_34};
  wire [127:0]      regroupV0_lo_lo_lo_35 = {regroupV0_hi_20, regroupV0_lo_20, regroupV0_hi_19, regroupV0_lo_19};
  wire [127:0]      regroupV0_lo_lo_hi_35 = {regroupV0_hi_22, regroupV0_lo_22, regroupV0_hi_21, regroupV0_lo_21};
  wire [255:0]      regroupV0_lo_lo_35 = {regroupV0_lo_lo_hi_35, regroupV0_lo_lo_lo_35};
  wire [127:0]      regroupV0_lo_hi_lo_35 = {regroupV0_hi_24, regroupV0_lo_24, regroupV0_hi_23, regroupV0_lo_23};
  wire [127:0]      regroupV0_lo_hi_hi_35 = {regroupV0_hi_26, regroupV0_lo_26, regroupV0_hi_25, regroupV0_lo_25};
  wire [255:0]      regroupV0_lo_hi_35 = {regroupV0_lo_hi_hi_35, regroupV0_lo_hi_lo_35};
  wire [511:0]      regroupV0_lo_35 = {regroupV0_lo_hi_35, regroupV0_lo_lo_35};
  wire [127:0]      regroupV0_hi_lo_lo_35 = {regroupV0_hi_28, regroupV0_lo_28, regroupV0_hi_27, regroupV0_lo_27};
  wire [127:0]      regroupV0_hi_lo_hi_35 = {regroupV0_hi_30, regroupV0_lo_30, regroupV0_hi_29, regroupV0_lo_29};
  wire [255:0]      regroupV0_hi_lo_35 = {regroupV0_hi_lo_hi_35, regroupV0_hi_lo_lo_35};
  wire [127:0]      regroupV0_hi_hi_lo_35 = {regroupV0_hi_32, regroupV0_lo_32, regroupV0_hi_31, regroupV0_lo_31};
  wire [127:0]      regroupV0_hi_hi_hi_35 = {regroupV0_hi_34, regroupV0_lo_34, regroupV0_hi_33, regroupV0_lo_33};
  wire [255:0]      regroupV0_hi_hi_35 = {regroupV0_hi_hi_hi_35, regroupV0_hi_hi_lo_35};
  wire [511:0]      regroupV0_hi_35 = {regroupV0_hi_hi_35, regroupV0_hi_lo_35};
  wire [1023:0]     regroupV0_1 = {regroupV0_hi_35, regroupV0_lo_35};
  wire [127:0]      regroupV0_lo_lo_lo_36 = {regroupV0_lo_lo_lo_hi_18, regroupV0_lo_lo_lo_lo_18};
  wire [127:0]      regroupV0_lo_lo_hi_36 = {regroupV0_lo_lo_hi_hi_18, regroupV0_lo_lo_hi_lo_18};
  wire [255:0]      regroupV0_lo_lo_36 = {regroupV0_lo_lo_hi_36, regroupV0_lo_lo_lo_36};
  wire [127:0]      regroupV0_lo_hi_lo_36 = {regroupV0_lo_hi_lo_hi_18, regroupV0_lo_hi_lo_lo_18};
  wire [127:0]      regroupV0_lo_hi_hi_36 = {regroupV0_lo_hi_hi_hi_18, regroupV0_lo_hi_hi_lo_18};
  wire [255:0]      regroupV0_lo_hi_36 = {regroupV0_lo_hi_hi_36, regroupV0_lo_hi_lo_36};
  wire [511:0]      regroupV0_lo_36 = {regroupV0_lo_hi_36, regroupV0_lo_lo_36};
  wire [127:0]      regroupV0_hi_lo_lo_36 = {regroupV0_hi_lo_lo_hi_18, regroupV0_hi_lo_lo_lo_18};
  wire [127:0]      regroupV0_hi_lo_hi_36 = {regroupV0_hi_lo_hi_hi_18, regroupV0_hi_lo_hi_lo_18};
  wire [255:0]      regroupV0_hi_lo_36 = {regroupV0_hi_lo_hi_36, regroupV0_hi_lo_lo_36};
  wire [127:0]      regroupV0_hi_hi_lo_36 = {regroupV0_hi_hi_lo_hi_18, regroupV0_hi_hi_lo_lo_18};
  wire [127:0]      regroupV0_hi_hi_hi_36 = {regroupV0_hi_hi_hi_hi_18, regroupV0_hi_hi_hi_lo_18};
  wire [255:0]      regroupV0_hi_hi_36 = {regroupV0_hi_hi_hi_36, regroupV0_hi_hi_lo_36};
  wire [511:0]      regroupV0_hi_36 = {regroupV0_hi_hi_36, regroupV0_hi_lo_36};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo = {regroupV0_lo_36[16], regroupV0_lo_36[0]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi = {regroupV0_lo_36[48], regroupV0_lo_36[32]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_19 = {regroupV0_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo = {regroupV0_lo_36[80], regroupV0_lo_36[64]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi = {regroupV0_lo_36[112], regroupV0_lo_36[96]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_19 = {regroupV0_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo};
  wire [7:0]        regroupV0_lo_lo_lo_37 = {regroupV0_lo_lo_lo_hi_19, regroupV0_lo_lo_lo_lo_19};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo = {regroupV0_lo_36[144], regroupV0_lo_36[128]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi = {regroupV0_lo_36[176], regroupV0_lo_36[160]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_19 = {regroupV0_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo = {regroupV0_lo_36[208], regroupV0_lo_36[192]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi = {regroupV0_lo_36[240], regroupV0_lo_36[224]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_19 = {regroupV0_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo};
  wire [7:0]        regroupV0_lo_lo_hi_37 = {regroupV0_lo_lo_hi_hi_19, regroupV0_lo_lo_hi_lo_19};
  wire [15:0]       regroupV0_lo_lo_37 = {regroupV0_lo_lo_hi_37, regroupV0_lo_lo_lo_37};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo = {regroupV0_lo_36[272], regroupV0_lo_36[256]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi = {regroupV0_lo_36[304], regroupV0_lo_36[288]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_19 = {regroupV0_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo = {regroupV0_lo_36[336], regroupV0_lo_36[320]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi = {regroupV0_lo_36[368], regroupV0_lo_36[352]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_19 = {regroupV0_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo};
  wire [7:0]        regroupV0_lo_hi_lo_37 = {regroupV0_lo_hi_lo_hi_19, regroupV0_lo_hi_lo_lo_19};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo = {regroupV0_lo_36[400], regroupV0_lo_36[384]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi = {regroupV0_lo_36[432], regroupV0_lo_36[416]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_19 = {regroupV0_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo = {regroupV0_lo_36[464], regroupV0_lo_36[448]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi = {regroupV0_lo_36[496], regroupV0_lo_36[480]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_19 = {regroupV0_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo};
  wire [7:0]        regroupV0_lo_hi_hi_37 = {regroupV0_lo_hi_hi_hi_19, regroupV0_lo_hi_hi_lo_19};
  wire [15:0]       regroupV0_lo_hi_37 = {regroupV0_lo_hi_hi_37, regroupV0_lo_hi_lo_37};
  wire [31:0]       regroupV0_lo_37 = {regroupV0_lo_hi_37, regroupV0_lo_lo_37};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo = {regroupV0_hi_36[16], regroupV0_hi_36[0]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi = {regroupV0_hi_36[48], regroupV0_hi_36[32]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_19 = {regroupV0_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo = {regroupV0_hi_36[80], regroupV0_hi_36[64]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi = {regroupV0_hi_36[112], regroupV0_hi_36[96]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_19 = {regroupV0_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo};
  wire [7:0]        regroupV0_hi_lo_lo_37 = {regroupV0_hi_lo_lo_hi_19, regroupV0_hi_lo_lo_lo_19};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo = {regroupV0_hi_36[144], regroupV0_hi_36[128]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi = {regroupV0_hi_36[176], regroupV0_hi_36[160]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_19 = {regroupV0_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo = {regroupV0_hi_36[208], regroupV0_hi_36[192]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi = {regroupV0_hi_36[240], regroupV0_hi_36[224]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_19 = {regroupV0_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo};
  wire [7:0]        regroupV0_hi_lo_hi_37 = {regroupV0_hi_lo_hi_hi_19, regroupV0_hi_lo_hi_lo_19};
  wire [15:0]       regroupV0_hi_lo_37 = {regroupV0_hi_lo_hi_37, regroupV0_hi_lo_lo_37};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo = {regroupV0_hi_36[272], regroupV0_hi_36[256]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi = {regroupV0_hi_36[304], regroupV0_hi_36[288]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_19 = {regroupV0_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo = {regroupV0_hi_36[336], regroupV0_hi_36[320]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi = {regroupV0_hi_36[368], regroupV0_hi_36[352]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_19 = {regroupV0_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo};
  wire [7:0]        regroupV0_hi_hi_lo_37 = {regroupV0_hi_hi_lo_hi_19, regroupV0_hi_hi_lo_lo_19};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo = {regroupV0_hi_36[400], regroupV0_hi_36[384]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi = {regroupV0_hi_36[432], regroupV0_hi_36[416]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_19 = {regroupV0_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo = {regroupV0_hi_36[464], regroupV0_hi_36[448]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi = {regroupV0_hi_36[496], regroupV0_hi_36[480]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_19 = {regroupV0_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo};
  wire [7:0]        regroupV0_hi_hi_hi_37 = {regroupV0_hi_hi_hi_hi_19, regroupV0_hi_hi_hi_lo_19};
  wire [15:0]       regroupV0_hi_hi_37 = {regroupV0_hi_hi_hi_37, regroupV0_hi_hi_lo_37};
  wire [31:0]       regroupV0_hi_37 = {regroupV0_hi_hi_37, regroupV0_hi_lo_37};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_1 = {regroupV0_lo_36[17], regroupV0_lo_36[1]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_1 = {regroupV0_lo_36[49], regroupV0_lo_36[33]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_20 = {regroupV0_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_1 = {regroupV0_lo_36[81], regroupV0_lo_36[65]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_1 = {regroupV0_lo_36[113], regroupV0_lo_36[97]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_20 = {regroupV0_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_lo_38 = {regroupV0_lo_lo_lo_hi_20, regroupV0_lo_lo_lo_lo_20};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_1 = {regroupV0_lo_36[145], regroupV0_lo_36[129]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_1 = {regroupV0_lo_36[177], regroupV0_lo_36[161]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_20 = {regroupV0_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_1 = {regroupV0_lo_36[209], regroupV0_lo_36[193]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_1 = {regroupV0_lo_36[241], regroupV0_lo_36[225]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_20 = {regroupV0_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_lo_hi_38 = {regroupV0_lo_lo_hi_hi_20, regroupV0_lo_lo_hi_lo_20};
  wire [15:0]       regroupV0_lo_lo_38 = {regroupV0_lo_lo_hi_38, regroupV0_lo_lo_lo_38};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_1 = {regroupV0_lo_36[273], regroupV0_lo_36[257]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_1 = {regroupV0_lo_36[305], regroupV0_lo_36[289]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_20 = {regroupV0_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_1 = {regroupV0_lo_36[337], regroupV0_lo_36[321]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_1 = {regroupV0_lo_36[369], regroupV0_lo_36[353]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_20 = {regroupV0_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_lo_38 = {regroupV0_lo_hi_lo_hi_20, regroupV0_lo_hi_lo_lo_20};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_1 = {regroupV0_lo_36[401], regroupV0_lo_36[385]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_1 = {regroupV0_lo_36[433], regroupV0_lo_36[417]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_20 = {regroupV0_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_1 = {regroupV0_lo_36[465], regroupV0_lo_36[449]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_1 = {regroupV0_lo_36[497], regroupV0_lo_36[481]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_20 = {regroupV0_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_lo_hi_hi_38 = {regroupV0_lo_hi_hi_hi_20, regroupV0_lo_hi_hi_lo_20};
  wire [15:0]       regroupV0_lo_hi_38 = {regroupV0_lo_hi_hi_38, regroupV0_lo_hi_lo_38};
  wire [31:0]       regroupV0_lo_38 = {regroupV0_lo_hi_38, regroupV0_lo_lo_38};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_1 = {regroupV0_hi_36[17], regroupV0_hi_36[1]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_1 = {regroupV0_hi_36[49], regroupV0_hi_36[33]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_20 = {regroupV0_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_1 = {regroupV0_hi_36[81], regroupV0_hi_36[65]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_1 = {regroupV0_hi_36[113], regroupV0_hi_36[97]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_20 = {regroupV0_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_lo_38 = {regroupV0_hi_lo_lo_hi_20, regroupV0_hi_lo_lo_lo_20};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_1 = {regroupV0_hi_36[145], regroupV0_hi_36[129]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_1 = {regroupV0_hi_36[177], regroupV0_hi_36[161]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_20 = {regroupV0_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_1 = {regroupV0_hi_36[209], regroupV0_hi_36[193]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_1 = {regroupV0_hi_36[241], regroupV0_hi_36[225]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_20 = {regroupV0_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_lo_hi_38 = {regroupV0_hi_lo_hi_hi_20, regroupV0_hi_lo_hi_lo_20};
  wire [15:0]       regroupV0_hi_lo_38 = {regroupV0_hi_lo_hi_38, regroupV0_hi_lo_lo_38};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_1 = {regroupV0_hi_36[273], regroupV0_hi_36[257]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_1 = {regroupV0_hi_36[305], regroupV0_hi_36[289]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_20 = {regroupV0_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_1 = {regroupV0_hi_36[337], regroupV0_hi_36[321]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_1 = {regroupV0_hi_36[369], regroupV0_hi_36[353]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_20 = {regroupV0_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_lo_38 = {regroupV0_hi_hi_lo_hi_20, regroupV0_hi_hi_lo_lo_20};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_1 = {regroupV0_hi_36[401], regroupV0_hi_36[385]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_1 = {regroupV0_hi_36[433], regroupV0_hi_36[417]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_20 = {regroupV0_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_1};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_1 = {regroupV0_hi_36[465], regroupV0_hi_36[449]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_1 = {regroupV0_hi_36[497], regroupV0_hi_36[481]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_20 = {regroupV0_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_1};
  wire [7:0]        regroupV0_hi_hi_hi_38 = {regroupV0_hi_hi_hi_hi_20, regroupV0_hi_hi_hi_lo_20};
  wire [15:0]       regroupV0_hi_hi_38 = {regroupV0_hi_hi_hi_38, regroupV0_hi_hi_lo_38};
  wire [31:0]       regroupV0_hi_38 = {regroupV0_hi_hi_38, regroupV0_hi_lo_38};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_2 = {regroupV0_lo_36[18], regroupV0_lo_36[2]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_2 = {regroupV0_lo_36[50], regroupV0_lo_36[34]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_21 = {regroupV0_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_2 = {regroupV0_lo_36[82], regroupV0_lo_36[66]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_2 = {regroupV0_lo_36[114], regroupV0_lo_36[98]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_21 = {regroupV0_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_lo_39 = {regroupV0_lo_lo_lo_hi_21, regroupV0_lo_lo_lo_lo_21};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_2 = {regroupV0_lo_36[146], regroupV0_lo_36[130]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_2 = {regroupV0_lo_36[178], regroupV0_lo_36[162]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_21 = {regroupV0_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_2 = {regroupV0_lo_36[210], regroupV0_lo_36[194]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_2 = {regroupV0_lo_36[242], regroupV0_lo_36[226]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_21 = {regroupV0_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_lo_hi_39 = {regroupV0_lo_lo_hi_hi_21, regroupV0_lo_lo_hi_lo_21};
  wire [15:0]       regroupV0_lo_lo_39 = {regroupV0_lo_lo_hi_39, regroupV0_lo_lo_lo_39};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_2 = {regroupV0_lo_36[274], regroupV0_lo_36[258]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_2 = {regroupV0_lo_36[306], regroupV0_lo_36[290]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_21 = {regroupV0_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_2 = {regroupV0_lo_36[338], regroupV0_lo_36[322]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_2 = {regroupV0_lo_36[370], regroupV0_lo_36[354]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_21 = {regroupV0_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_lo_39 = {regroupV0_lo_hi_lo_hi_21, regroupV0_lo_hi_lo_lo_21};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_2 = {regroupV0_lo_36[402], regroupV0_lo_36[386]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_2 = {regroupV0_lo_36[434], regroupV0_lo_36[418]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_21 = {regroupV0_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_2 = {regroupV0_lo_36[466], regroupV0_lo_36[450]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_2 = {regroupV0_lo_36[498], regroupV0_lo_36[482]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_21 = {regroupV0_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_lo_hi_hi_39 = {regroupV0_lo_hi_hi_hi_21, regroupV0_lo_hi_hi_lo_21};
  wire [15:0]       regroupV0_lo_hi_39 = {regroupV0_lo_hi_hi_39, regroupV0_lo_hi_lo_39};
  wire [31:0]       regroupV0_lo_39 = {regroupV0_lo_hi_39, regroupV0_lo_lo_39};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_2 = {regroupV0_hi_36[18], regroupV0_hi_36[2]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_2 = {regroupV0_hi_36[50], regroupV0_hi_36[34]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_21 = {regroupV0_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_2 = {regroupV0_hi_36[82], regroupV0_hi_36[66]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_2 = {regroupV0_hi_36[114], regroupV0_hi_36[98]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_21 = {regroupV0_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_lo_39 = {regroupV0_hi_lo_lo_hi_21, regroupV0_hi_lo_lo_lo_21};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_2 = {regroupV0_hi_36[146], regroupV0_hi_36[130]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_2 = {regroupV0_hi_36[178], regroupV0_hi_36[162]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_21 = {regroupV0_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_2 = {regroupV0_hi_36[210], regroupV0_hi_36[194]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_2 = {regroupV0_hi_36[242], regroupV0_hi_36[226]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_21 = {regroupV0_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_lo_hi_39 = {regroupV0_hi_lo_hi_hi_21, regroupV0_hi_lo_hi_lo_21};
  wire [15:0]       regroupV0_hi_lo_39 = {regroupV0_hi_lo_hi_39, regroupV0_hi_lo_lo_39};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_2 = {regroupV0_hi_36[274], regroupV0_hi_36[258]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_2 = {regroupV0_hi_36[306], regroupV0_hi_36[290]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_21 = {regroupV0_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_2 = {regroupV0_hi_36[338], regroupV0_hi_36[322]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_2 = {regroupV0_hi_36[370], regroupV0_hi_36[354]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_21 = {regroupV0_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_lo_39 = {regroupV0_hi_hi_lo_hi_21, regroupV0_hi_hi_lo_lo_21};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_2 = {regroupV0_hi_36[402], regroupV0_hi_36[386]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_2 = {regroupV0_hi_36[434], regroupV0_hi_36[418]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_21 = {regroupV0_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_2};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_2 = {regroupV0_hi_36[466], regroupV0_hi_36[450]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_2 = {regroupV0_hi_36[498], regroupV0_hi_36[482]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_21 = {regroupV0_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_2};
  wire [7:0]        regroupV0_hi_hi_hi_39 = {regroupV0_hi_hi_hi_hi_21, regroupV0_hi_hi_hi_lo_21};
  wire [15:0]       regroupV0_hi_hi_39 = {regroupV0_hi_hi_hi_39, regroupV0_hi_hi_lo_39};
  wire [31:0]       regroupV0_hi_39 = {regroupV0_hi_hi_39, regroupV0_hi_lo_39};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_3 = {regroupV0_lo_36[19], regroupV0_lo_36[3]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_3 = {regroupV0_lo_36[51], regroupV0_lo_36[35]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_22 = {regroupV0_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_3 = {regroupV0_lo_36[83], regroupV0_lo_36[67]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_3 = {regroupV0_lo_36[115], regroupV0_lo_36[99]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_22 = {regroupV0_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_lo_40 = {regroupV0_lo_lo_lo_hi_22, regroupV0_lo_lo_lo_lo_22};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_3 = {regroupV0_lo_36[147], regroupV0_lo_36[131]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_3 = {regroupV0_lo_36[179], regroupV0_lo_36[163]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_22 = {regroupV0_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_3 = {regroupV0_lo_36[211], regroupV0_lo_36[195]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_3 = {regroupV0_lo_36[243], regroupV0_lo_36[227]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_22 = {regroupV0_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_lo_hi_40 = {regroupV0_lo_lo_hi_hi_22, regroupV0_lo_lo_hi_lo_22};
  wire [15:0]       regroupV0_lo_lo_40 = {regroupV0_lo_lo_hi_40, regroupV0_lo_lo_lo_40};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_3 = {regroupV0_lo_36[275], regroupV0_lo_36[259]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_3 = {regroupV0_lo_36[307], regroupV0_lo_36[291]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_22 = {regroupV0_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_3 = {regroupV0_lo_36[339], regroupV0_lo_36[323]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_3 = {regroupV0_lo_36[371], regroupV0_lo_36[355]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_22 = {regroupV0_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_lo_40 = {regroupV0_lo_hi_lo_hi_22, regroupV0_lo_hi_lo_lo_22};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_3 = {regroupV0_lo_36[403], regroupV0_lo_36[387]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_3 = {regroupV0_lo_36[435], regroupV0_lo_36[419]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_22 = {regroupV0_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_3 = {regroupV0_lo_36[467], regroupV0_lo_36[451]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_3 = {regroupV0_lo_36[499], regroupV0_lo_36[483]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_22 = {regroupV0_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_lo_hi_hi_40 = {regroupV0_lo_hi_hi_hi_22, regroupV0_lo_hi_hi_lo_22};
  wire [15:0]       regroupV0_lo_hi_40 = {regroupV0_lo_hi_hi_40, regroupV0_lo_hi_lo_40};
  wire [31:0]       regroupV0_lo_40 = {regroupV0_lo_hi_40, regroupV0_lo_lo_40};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_3 = {regroupV0_hi_36[19], regroupV0_hi_36[3]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_3 = {regroupV0_hi_36[51], regroupV0_hi_36[35]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_22 = {regroupV0_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_3 = {regroupV0_hi_36[83], regroupV0_hi_36[67]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_3 = {regroupV0_hi_36[115], regroupV0_hi_36[99]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_22 = {regroupV0_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_lo_40 = {regroupV0_hi_lo_lo_hi_22, regroupV0_hi_lo_lo_lo_22};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_3 = {regroupV0_hi_36[147], regroupV0_hi_36[131]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_3 = {regroupV0_hi_36[179], regroupV0_hi_36[163]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_22 = {regroupV0_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_3 = {regroupV0_hi_36[211], regroupV0_hi_36[195]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_3 = {regroupV0_hi_36[243], regroupV0_hi_36[227]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_22 = {regroupV0_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_lo_hi_40 = {regroupV0_hi_lo_hi_hi_22, regroupV0_hi_lo_hi_lo_22};
  wire [15:0]       regroupV0_hi_lo_40 = {regroupV0_hi_lo_hi_40, regroupV0_hi_lo_lo_40};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_3 = {regroupV0_hi_36[275], regroupV0_hi_36[259]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_3 = {regroupV0_hi_36[307], regroupV0_hi_36[291]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_22 = {regroupV0_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_3 = {regroupV0_hi_36[339], regroupV0_hi_36[323]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_3 = {regroupV0_hi_36[371], regroupV0_hi_36[355]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_22 = {regroupV0_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_lo_40 = {regroupV0_hi_hi_lo_hi_22, regroupV0_hi_hi_lo_lo_22};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_3 = {regroupV0_hi_36[403], regroupV0_hi_36[387]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_3 = {regroupV0_hi_36[435], regroupV0_hi_36[419]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_22 = {regroupV0_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_3};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_3 = {regroupV0_hi_36[467], regroupV0_hi_36[451]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_3 = {regroupV0_hi_36[499], regroupV0_hi_36[483]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_22 = {regroupV0_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_3};
  wire [7:0]        regroupV0_hi_hi_hi_40 = {regroupV0_hi_hi_hi_hi_22, regroupV0_hi_hi_hi_lo_22};
  wire [15:0]       regroupV0_hi_hi_40 = {regroupV0_hi_hi_hi_40, regroupV0_hi_hi_lo_40};
  wire [31:0]       regroupV0_hi_40 = {regroupV0_hi_hi_40, regroupV0_hi_lo_40};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_4 = {regroupV0_lo_36[20], regroupV0_lo_36[4]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_4 = {regroupV0_lo_36[52], regroupV0_lo_36[36]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_23 = {regroupV0_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_4};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_4 = {regroupV0_lo_36[84], regroupV0_lo_36[68]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_4 = {regroupV0_lo_36[116], regroupV0_lo_36[100]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_23 = {regroupV0_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_lo_41 = {regroupV0_lo_lo_lo_hi_23, regroupV0_lo_lo_lo_lo_23};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_4 = {regroupV0_lo_36[148], regroupV0_lo_36[132]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_4 = {regroupV0_lo_36[180], regroupV0_lo_36[164]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_23 = {regroupV0_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_4};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_4 = {regroupV0_lo_36[212], regroupV0_lo_36[196]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_4 = {regroupV0_lo_36[244], regroupV0_lo_36[228]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_23 = {regroupV0_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_4};
  wire [7:0]        regroupV0_lo_lo_hi_41 = {regroupV0_lo_lo_hi_hi_23, regroupV0_lo_lo_hi_lo_23};
  wire [15:0]       regroupV0_lo_lo_41 = {regroupV0_lo_lo_hi_41, regroupV0_lo_lo_lo_41};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_4 = {regroupV0_lo_36[276], regroupV0_lo_36[260]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_4 = {regroupV0_lo_36[308], regroupV0_lo_36[292]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_23 = {regroupV0_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_4};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_4 = {regroupV0_lo_36[340], regroupV0_lo_36[324]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_4 = {regroupV0_lo_36[372], regroupV0_lo_36[356]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_23 = {regroupV0_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_4};
  wire [7:0]        regroupV0_lo_hi_lo_41 = {regroupV0_lo_hi_lo_hi_23, regroupV0_lo_hi_lo_lo_23};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_4 = {regroupV0_lo_36[404], regroupV0_lo_36[388]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_4 = {regroupV0_lo_36[436], regroupV0_lo_36[420]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_23 = {regroupV0_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_4};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_4 = {regroupV0_lo_36[468], regroupV0_lo_36[452]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_4 = {regroupV0_lo_36[500], regroupV0_lo_36[484]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_23 = {regroupV0_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_4};
  wire [7:0]        regroupV0_lo_hi_hi_41 = {regroupV0_lo_hi_hi_hi_23, regroupV0_lo_hi_hi_lo_23};
  wire [15:0]       regroupV0_lo_hi_41 = {regroupV0_lo_hi_hi_41, regroupV0_lo_hi_lo_41};
  wire [31:0]       regroupV0_lo_41 = {regroupV0_lo_hi_41, regroupV0_lo_lo_41};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_4 = {regroupV0_hi_36[20], regroupV0_hi_36[4]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_4 = {regroupV0_hi_36[52], regroupV0_hi_36[36]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_23 = {regroupV0_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_4};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_4 = {regroupV0_hi_36[84], regroupV0_hi_36[68]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_4 = {regroupV0_hi_36[116], regroupV0_hi_36[100]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_23 = {regroupV0_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_4};
  wire [7:0]        regroupV0_hi_lo_lo_41 = {regroupV0_hi_lo_lo_hi_23, regroupV0_hi_lo_lo_lo_23};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_4 = {regroupV0_hi_36[148], regroupV0_hi_36[132]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_4 = {regroupV0_hi_36[180], regroupV0_hi_36[164]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_23 = {regroupV0_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_4};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_4 = {regroupV0_hi_36[212], regroupV0_hi_36[196]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_4 = {regroupV0_hi_36[244], regroupV0_hi_36[228]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_23 = {regroupV0_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_4};
  wire [7:0]        regroupV0_hi_lo_hi_41 = {regroupV0_hi_lo_hi_hi_23, regroupV0_hi_lo_hi_lo_23};
  wire [15:0]       regroupV0_hi_lo_41 = {regroupV0_hi_lo_hi_41, regroupV0_hi_lo_lo_41};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_4 = {regroupV0_hi_36[276], regroupV0_hi_36[260]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_4 = {regroupV0_hi_36[308], regroupV0_hi_36[292]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_23 = {regroupV0_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_4};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_4 = {regroupV0_hi_36[340], regroupV0_hi_36[324]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_4 = {regroupV0_hi_36[372], regroupV0_hi_36[356]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_23 = {regroupV0_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_4};
  wire [7:0]        regroupV0_hi_hi_lo_41 = {regroupV0_hi_hi_lo_hi_23, regroupV0_hi_hi_lo_lo_23};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_4 = {regroupV0_hi_36[404], regroupV0_hi_36[388]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_4 = {regroupV0_hi_36[436], regroupV0_hi_36[420]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_23 = {regroupV0_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_4};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_4 = {regroupV0_hi_36[468], regroupV0_hi_36[452]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_4 = {regroupV0_hi_36[500], regroupV0_hi_36[484]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_23 = {regroupV0_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_4};
  wire [7:0]        regroupV0_hi_hi_hi_41 = {regroupV0_hi_hi_hi_hi_23, regroupV0_hi_hi_hi_lo_23};
  wire [15:0]       regroupV0_hi_hi_41 = {regroupV0_hi_hi_hi_41, regroupV0_hi_hi_lo_41};
  wire [31:0]       regroupV0_hi_41 = {regroupV0_hi_hi_41, regroupV0_hi_lo_41};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_5 = {regroupV0_lo_36[21], regroupV0_lo_36[5]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_5 = {regroupV0_lo_36[53], regroupV0_lo_36[37]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_24 = {regroupV0_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_5};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_5 = {regroupV0_lo_36[85], regroupV0_lo_36[69]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_5 = {regroupV0_lo_36[117], regroupV0_lo_36[101]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_24 = {regroupV0_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_lo_42 = {regroupV0_lo_lo_lo_hi_24, regroupV0_lo_lo_lo_lo_24};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_5 = {regroupV0_lo_36[149], regroupV0_lo_36[133]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_5 = {regroupV0_lo_36[181], regroupV0_lo_36[165]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_24 = {regroupV0_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_5};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_5 = {regroupV0_lo_36[213], regroupV0_lo_36[197]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_5 = {regroupV0_lo_36[245], regroupV0_lo_36[229]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_24 = {regroupV0_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_5};
  wire [7:0]        regroupV0_lo_lo_hi_42 = {regroupV0_lo_lo_hi_hi_24, regroupV0_lo_lo_hi_lo_24};
  wire [15:0]       regroupV0_lo_lo_42 = {regroupV0_lo_lo_hi_42, regroupV0_lo_lo_lo_42};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_5 = {regroupV0_lo_36[277], regroupV0_lo_36[261]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_5 = {regroupV0_lo_36[309], regroupV0_lo_36[293]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_24 = {regroupV0_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_5};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_5 = {regroupV0_lo_36[341], regroupV0_lo_36[325]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_5 = {regroupV0_lo_36[373], regroupV0_lo_36[357]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_24 = {regroupV0_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_5};
  wire [7:0]        regroupV0_lo_hi_lo_42 = {regroupV0_lo_hi_lo_hi_24, regroupV0_lo_hi_lo_lo_24};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_5 = {regroupV0_lo_36[405], regroupV0_lo_36[389]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_5 = {regroupV0_lo_36[437], regroupV0_lo_36[421]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_24 = {regroupV0_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_5};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_5 = {regroupV0_lo_36[469], regroupV0_lo_36[453]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_5 = {regroupV0_lo_36[501], regroupV0_lo_36[485]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_24 = {regroupV0_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_5};
  wire [7:0]        regroupV0_lo_hi_hi_42 = {regroupV0_lo_hi_hi_hi_24, regroupV0_lo_hi_hi_lo_24};
  wire [15:0]       regroupV0_lo_hi_42 = {regroupV0_lo_hi_hi_42, regroupV0_lo_hi_lo_42};
  wire [31:0]       regroupV0_lo_42 = {regroupV0_lo_hi_42, regroupV0_lo_lo_42};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_5 = {regroupV0_hi_36[21], regroupV0_hi_36[5]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_5 = {regroupV0_hi_36[53], regroupV0_hi_36[37]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_24 = {regroupV0_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_5};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_5 = {regroupV0_hi_36[85], regroupV0_hi_36[69]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_5 = {regroupV0_hi_36[117], regroupV0_hi_36[101]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_24 = {regroupV0_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_5};
  wire [7:0]        regroupV0_hi_lo_lo_42 = {regroupV0_hi_lo_lo_hi_24, regroupV0_hi_lo_lo_lo_24};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_5 = {regroupV0_hi_36[149], regroupV0_hi_36[133]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_5 = {regroupV0_hi_36[181], regroupV0_hi_36[165]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_24 = {regroupV0_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_5};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_5 = {regroupV0_hi_36[213], regroupV0_hi_36[197]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_5 = {regroupV0_hi_36[245], regroupV0_hi_36[229]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_24 = {regroupV0_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_5};
  wire [7:0]        regroupV0_hi_lo_hi_42 = {regroupV0_hi_lo_hi_hi_24, regroupV0_hi_lo_hi_lo_24};
  wire [15:0]       regroupV0_hi_lo_42 = {regroupV0_hi_lo_hi_42, regroupV0_hi_lo_lo_42};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_5 = {regroupV0_hi_36[277], regroupV0_hi_36[261]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_5 = {regroupV0_hi_36[309], regroupV0_hi_36[293]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_24 = {regroupV0_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_5};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_5 = {regroupV0_hi_36[341], regroupV0_hi_36[325]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_5 = {regroupV0_hi_36[373], regroupV0_hi_36[357]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_24 = {regroupV0_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_5};
  wire [7:0]        regroupV0_hi_hi_lo_42 = {regroupV0_hi_hi_lo_hi_24, regroupV0_hi_hi_lo_lo_24};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_5 = {regroupV0_hi_36[405], regroupV0_hi_36[389]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_5 = {regroupV0_hi_36[437], regroupV0_hi_36[421]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_24 = {regroupV0_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_5};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_5 = {regroupV0_hi_36[469], regroupV0_hi_36[453]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_5 = {regroupV0_hi_36[501], regroupV0_hi_36[485]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_24 = {regroupV0_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_5};
  wire [7:0]        regroupV0_hi_hi_hi_42 = {regroupV0_hi_hi_hi_hi_24, regroupV0_hi_hi_hi_lo_24};
  wire [15:0]       regroupV0_hi_hi_42 = {regroupV0_hi_hi_hi_42, regroupV0_hi_hi_lo_42};
  wire [31:0]       regroupV0_hi_42 = {regroupV0_hi_hi_42, regroupV0_hi_lo_42};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_6 = {regroupV0_lo_36[22], regroupV0_lo_36[6]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_6 = {regroupV0_lo_36[54], regroupV0_lo_36[38]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_25 = {regroupV0_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_6};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_6 = {regroupV0_lo_36[86], regroupV0_lo_36[70]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_6 = {regroupV0_lo_36[118], regroupV0_lo_36[102]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_25 = {regroupV0_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_lo_43 = {regroupV0_lo_lo_lo_hi_25, regroupV0_lo_lo_lo_lo_25};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_6 = {regroupV0_lo_36[150], regroupV0_lo_36[134]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_6 = {regroupV0_lo_36[182], regroupV0_lo_36[166]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_25 = {regroupV0_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_6};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_6 = {regroupV0_lo_36[214], regroupV0_lo_36[198]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_6 = {regroupV0_lo_36[246], regroupV0_lo_36[230]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_25 = {regroupV0_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_6};
  wire [7:0]        regroupV0_lo_lo_hi_43 = {regroupV0_lo_lo_hi_hi_25, regroupV0_lo_lo_hi_lo_25};
  wire [15:0]       regroupV0_lo_lo_43 = {regroupV0_lo_lo_hi_43, regroupV0_lo_lo_lo_43};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_6 = {regroupV0_lo_36[278], regroupV0_lo_36[262]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_6 = {regroupV0_lo_36[310], regroupV0_lo_36[294]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_25 = {regroupV0_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_6};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_6 = {regroupV0_lo_36[342], regroupV0_lo_36[326]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_6 = {regroupV0_lo_36[374], regroupV0_lo_36[358]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_25 = {regroupV0_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_6};
  wire [7:0]        regroupV0_lo_hi_lo_43 = {regroupV0_lo_hi_lo_hi_25, regroupV0_lo_hi_lo_lo_25};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_6 = {regroupV0_lo_36[406], regroupV0_lo_36[390]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_6 = {regroupV0_lo_36[438], regroupV0_lo_36[422]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_25 = {regroupV0_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_6};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_6 = {regroupV0_lo_36[470], regroupV0_lo_36[454]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_6 = {regroupV0_lo_36[502], regroupV0_lo_36[486]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_25 = {regroupV0_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_6};
  wire [7:0]        regroupV0_lo_hi_hi_43 = {regroupV0_lo_hi_hi_hi_25, regroupV0_lo_hi_hi_lo_25};
  wire [15:0]       regroupV0_lo_hi_43 = {regroupV0_lo_hi_hi_43, regroupV0_lo_hi_lo_43};
  wire [31:0]       regroupV0_lo_43 = {regroupV0_lo_hi_43, regroupV0_lo_lo_43};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_6 = {regroupV0_hi_36[22], regroupV0_hi_36[6]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_6 = {regroupV0_hi_36[54], regroupV0_hi_36[38]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_25 = {regroupV0_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_6};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_6 = {regroupV0_hi_36[86], regroupV0_hi_36[70]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_6 = {regroupV0_hi_36[118], regroupV0_hi_36[102]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_25 = {regroupV0_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_6};
  wire [7:0]        regroupV0_hi_lo_lo_43 = {regroupV0_hi_lo_lo_hi_25, regroupV0_hi_lo_lo_lo_25};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_6 = {regroupV0_hi_36[150], regroupV0_hi_36[134]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_6 = {regroupV0_hi_36[182], regroupV0_hi_36[166]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_25 = {regroupV0_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_6};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_6 = {regroupV0_hi_36[214], regroupV0_hi_36[198]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_6 = {regroupV0_hi_36[246], regroupV0_hi_36[230]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_25 = {regroupV0_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_6};
  wire [7:0]        regroupV0_hi_lo_hi_43 = {regroupV0_hi_lo_hi_hi_25, regroupV0_hi_lo_hi_lo_25};
  wire [15:0]       regroupV0_hi_lo_43 = {regroupV0_hi_lo_hi_43, regroupV0_hi_lo_lo_43};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_6 = {regroupV0_hi_36[278], regroupV0_hi_36[262]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_6 = {regroupV0_hi_36[310], regroupV0_hi_36[294]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_25 = {regroupV0_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_6};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_6 = {regroupV0_hi_36[342], regroupV0_hi_36[326]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_6 = {regroupV0_hi_36[374], regroupV0_hi_36[358]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_25 = {regroupV0_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_6};
  wire [7:0]        regroupV0_hi_hi_lo_43 = {regroupV0_hi_hi_lo_hi_25, regroupV0_hi_hi_lo_lo_25};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_6 = {regroupV0_hi_36[406], regroupV0_hi_36[390]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_6 = {regroupV0_hi_36[438], regroupV0_hi_36[422]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_25 = {regroupV0_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_6};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_6 = {regroupV0_hi_36[470], regroupV0_hi_36[454]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_6 = {regroupV0_hi_36[502], regroupV0_hi_36[486]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_25 = {regroupV0_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_6};
  wire [7:0]        regroupV0_hi_hi_hi_43 = {regroupV0_hi_hi_hi_hi_25, regroupV0_hi_hi_hi_lo_25};
  wire [15:0]       regroupV0_hi_hi_43 = {regroupV0_hi_hi_hi_43, regroupV0_hi_hi_lo_43};
  wire [31:0]       regroupV0_hi_43 = {regroupV0_hi_hi_43, regroupV0_hi_lo_43};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_7 = {regroupV0_lo_36[23], regroupV0_lo_36[7]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_7 = {regroupV0_lo_36[55], regroupV0_lo_36[39]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_26 = {regroupV0_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_7};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_7 = {regroupV0_lo_36[87], regroupV0_lo_36[71]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_7 = {regroupV0_lo_36[119], regroupV0_lo_36[103]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_26 = {regroupV0_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_lo_44 = {regroupV0_lo_lo_lo_hi_26, regroupV0_lo_lo_lo_lo_26};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_7 = {regroupV0_lo_36[151], regroupV0_lo_36[135]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_7 = {regroupV0_lo_36[183], regroupV0_lo_36[167]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_26 = {regroupV0_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_7};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_7 = {regroupV0_lo_36[215], regroupV0_lo_36[199]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_7 = {regroupV0_lo_36[247], regroupV0_lo_36[231]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_26 = {regroupV0_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_7};
  wire [7:0]        regroupV0_lo_lo_hi_44 = {regroupV0_lo_lo_hi_hi_26, regroupV0_lo_lo_hi_lo_26};
  wire [15:0]       regroupV0_lo_lo_44 = {regroupV0_lo_lo_hi_44, regroupV0_lo_lo_lo_44};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_7 = {regroupV0_lo_36[279], regroupV0_lo_36[263]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_7 = {regroupV0_lo_36[311], regroupV0_lo_36[295]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_26 = {regroupV0_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_7};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_7 = {regroupV0_lo_36[343], regroupV0_lo_36[327]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_7 = {regroupV0_lo_36[375], regroupV0_lo_36[359]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_26 = {regroupV0_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_7};
  wire [7:0]        regroupV0_lo_hi_lo_44 = {regroupV0_lo_hi_lo_hi_26, regroupV0_lo_hi_lo_lo_26};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_7 = {regroupV0_lo_36[407], regroupV0_lo_36[391]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_7 = {regroupV0_lo_36[439], regroupV0_lo_36[423]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_26 = {regroupV0_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_7};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_7 = {regroupV0_lo_36[471], regroupV0_lo_36[455]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_7 = {regroupV0_lo_36[503], regroupV0_lo_36[487]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_26 = {regroupV0_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_7};
  wire [7:0]        regroupV0_lo_hi_hi_44 = {regroupV0_lo_hi_hi_hi_26, regroupV0_lo_hi_hi_lo_26};
  wire [15:0]       regroupV0_lo_hi_44 = {regroupV0_lo_hi_hi_44, regroupV0_lo_hi_lo_44};
  wire [31:0]       regroupV0_lo_44 = {regroupV0_lo_hi_44, regroupV0_lo_lo_44};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_7 = {regroupV0_hi_36[23], regroupV0_hi_36[7]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_7 = {regroupV0_hi_36[55], regroupV0_hi_36[39]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_26 = {regroupV0_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_7};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_7 = {regroupV0_hi_36[87], regroupV0_hi_36[71]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_7 = {regroupV0_hi_36[119], regroupV0_hi_36[103]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_26 = {regroupV0_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_7};
  wire [7:0]        regroupV0_hi_lo_lo_44 = {regroupV0_hi_lo_lo_hi_26, regroupV0_hi_lo_lo_lo_26};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_7 = {regroupV0_hi_36[151], regroupV0_hi_36[135]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_7 = {regroupV0_hi_36[183], regroupV0_hi_36[167]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_26 = {regroupV0_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_7};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_7 = {regroupV0_hi_36[215], regroupV0_hi_36[199]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_7 = {regroupV0_hi_36[247], regroupV0_hi_36[231]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_26 = {regroupV0_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_7};
  wire [7:0]        regroupV0_hi_lo_hi_44 = {regroupV0_hi_lo_hi_hi_26, regroupV0_hi_lo_hi_lo_26};
  wire [15:0]       regroupV0_hi_lo_44 = {regroupV0_hi_lo_hi_44, regroupV0_hi_lo_lo_44};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_7 = {regroupV0_hi_36[279], regroupV0_hi_36[263]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_7 = {regroupV0_hi_36[311], regroupV0_hi_36[295]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_26 = {regroupV0_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_7};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_7 = {regroupV0_hi_36[343], regroupV0_hi_36[327]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_7 = {regroupV0_hi_36[375], regroupV0_hi_36[359]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_26 = {regroupV0_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_7};
  wire [7:0]        regroupV0_hi_hi_lo_44 = {regroupV0_hi_hi_lo_hi_26, regroupV0_hi_hi_lo_lo_26};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_7 = {regroupV0_hi_36[407], regroupV0_hi_36[391]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_7 = {regroupV0_hi_36[439], regroupV0_hi_36[423]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_26 = {regroupV0_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_7};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_7 = {regroupV0_hi_36[471], regroupV0_hi_36[455]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_7 = {regroupV0_hi_36[503], regroupV0_hi_36[487]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_26 = {regroupV0_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_7};
  wire [7:0]        regroupV0_hi_hi_hi_44 = {regroupV0_hi_hi_hi_hi_26, regroupV0_hi_hi_hi_lo_26};
  wire [15:0]       regroupV0_hi_hi_44 = {regroupV0_hi_hi_hi_44, regroupV0_hi_hi_lo_44};
  wire [31:0]       regroupV0_hi_44 = {regroupV0_hi_hi_44, regroupV0_hi_lo_44};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_8 = {regroupV0_lo_36[24], regroupV0_lo_36[8]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_8 = {regroupV0_lo_36[56], regroupV0_lo_36[40]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_27 = {regroupV0_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_8};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_8 = {regroupV0_lo_36[88], regroupV0_lo_36[72]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_8 = {regroupV0_lo_36[120], regroupV0_lo_36[104]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_27 = {regroupV0_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_8};
  wire [7:0]        regroupV0_lo_lo_lo_45 = {regroupV0_lo_lo_lo_hi_27, regroupV0_lo_lo_lo_lo_27};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_8 = {regroupV0_lo_36[152], regroupV0_lo_36[136]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_8 = {regroupV0_lo_36[184], regroupV0_lo_36[168]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_27 = {regroupV0_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_8};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_8 = {regroupV0_lo_36[216], regroupV0_lo_36[200]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_8 = {regroupV0_lo_36[248], regroupV0_lo_36[232]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_27 = {regroupV0_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_8};
  wire [7:0]        regroupV0_lo_lo_hi_45 = {regroupV0_lo_lo_hi_hi_27, regroupV0_lo_lo_hi_lo_27};
  wire [15:0]       regroupV0_lo_lo_45 = {regroupV0_lo_lo_hi_45, regroupV0_lo_lo_lo_45};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_8 = {regroupV0_lo_36[280], regroupV0_lo_36[264]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_8 = {regroupV0_lo_36[312], regroupV0_lo_36[296]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_27 = {regroupV0_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_8};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_8 = {regroupV0_lo_36[344], regroupV0_lo_36[328]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_8 = {regroupV0_lo_36[376], regroupV0_lo_36[360]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_27 = {regroupV0_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_8};
  wire [7:0]        regroupV0_lo_hi_lo_45 = {regroupV0_lo_hi_lo_hi_27, regroupV0_lo_hi_lo_lo_27};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_8 = {regroupV0_lo_36[408], regroupV0_lo_36[392]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_8 = {regroupV0_lo_36[440], regroupV0_lo_36[424]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_27 = {regroupV0_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_8};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_8 = {regroupV0_lo_36[472], regroupV0_lo_36[456]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_8 = {regroupV0_lo_36[504], regroupV0_lo_36[488]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_27 = {regroupV0_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_8};
  wire [7:0]        regroupV0_lo_hi_hi_45 = {regroupV0_lo_hi_hi_hi_27, regroupV0_lo_hi_hi_lo_27};
  wire [15:0]       regroupV0_lo_hi_45 = {regroupV0_lo_hi_hi_45, regroupV0_lo_hi_lo_45};
  wire [31:0]       regroupV0_lo_45 = {regroupV0_lo_hi_45, regroupV0_lo_lo_45};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_8 = {regroupV0_hi_36[24], regroupV0_hi_36[8]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_8 = {regroupV0_hi_36[56], regroupV0_hi_36[40]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_27 = {regroupV0_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_8};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_8 = {regroupV0_hi_36[88], regroupV0_hi_36[72]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_8 = {regroupV0_hi_36[120], regroupV0_hi_36[104]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_27 = {regroupV0_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_8};
  wire [7:0]        regroupV0_hi_lo_lo_45 = {regroupV0_hi_lo_lo_hi_27, regroupV0_hi_lo_lo_lo_27};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_8 = {regroupV0_hi_36[152], regroupV0_hi_36[136]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_8 = {regroupV0_hi_36[184], regroupV0_hi_36[168]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_27 = {regroupV0_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_8};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_8 = {regroupV0_hi_36[216], regroupV0_hi_36[200]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_8 = {regroupV0_hi_36[248], regroupV0_hi_36[232]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_27 = {regroupV0_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_8};
  wire [7:0]        regroupV0_hi_lo_hi_45 = {regroupV0_hi_lo_hi_hi_27, regroupV0_hi_lo_hi_lo_27};
  wire [15:0]       regroupV0_hi_lo_45 = {regroupV0_hi_lo_hi_45, regroupV0_hi_lo_lo_45};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_8 = {regroupV0_hi_36[280], regroupV0_hi_36[264]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_8 = {regroupV0_hi_36[312], regroupV0_hi_36[296]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_27 = {regroupV0_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_8};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_8 = {regroupV0_hi_36[344], regroupV0_hi_36[328]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_8 = {regroupV0_hi_36[376], regroupV0_hi_36[360]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_27 = {regroupV0_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_8};
  wire [7:0]        regroupV0_hi_hi_lo_45 = {regroupV0_hi_hi_lo_hi_27, regroupV0_hi_hi_lo_lo_27};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_8 = {regroupV0_hi_36[408], regroupV0_hi_36[392]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_8 = {regroupV0_hi_36[440], regroupV0_hi_36[424]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_27 = {regroupV0_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_8};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_8 = {regroupV0_hi_36[472], regroupV0_hi_36[456]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_8 = {regroupV0_hi_36[504], regroupV0_hi_36[488]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_27 = {regroupV0_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_8};
  wire [7:0]        regroupV0_hi_hi_hi_45 = {regroupV0_hi_hi_hi_hi_27, regroupV0_hi_hi_hi_lo_27};
  wire [15:0]       regroupV0_hi_hi_45 = {regroupV0_hi_hi_hi_45, regroupV0_hi_hi_lo_45};
  wire [31:0]       regroupV0_hi_45 = {regroupV0_hi_hi_45, regroupV0_hi_lo_45};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_9 = {regroupV0_lo_36[25], regroupV0_lo_36[9]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_9 = {regroupV0_lo_36[57], regroupV0_lo_36[41]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_28 = {regroupV0_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_9};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_9 = {regroupV0_lo_36[89], regroupV0_lo_36[73]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_9 = {regroupV0_lo_36[121], regroupV0_lo_36[105]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_28 = {regroupV0_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_9};
  wire [7:0]        regroupV0_lo_lo_lo_46 = {regroupV0_lo_lo_lo_hi_28, regroupV0_lo_lo_lo_lo_28};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_9 = {regroupV0_lo_36[153], regroupV0_lo_36[137]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_9 = {regroupV0_lo_36[185], regroupV0_lo_36[169]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_28 = {regroupV0_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_9};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_9 = {regroupV0_lo_36[217], regroupV0_lo_36[201]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_9 = {regroupV0_lo_36[249], regroupV0_lo_36[233]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_28 = {regroupV0_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_9};
  wire [7:0]        regroupV0_lo_lo_hi_46 = {regroupV0_lo_lo_hi_hi_28, regroupV0_lo_lo_hi_lo_28};
  wire [15:0]       regroupV0_lo_lo_46 = {regroupV0_lo_lo_hi_46, regroupV0_lo_lo_lo_46};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_9 = {regroupV0_lo_36[281], regroupV0_lo_36[265]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_9 = {regroupV0_lo_36[313], regroupV0_lo_36[297]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_28 = {regroupV0_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_9};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_9 = {regroupV0_lo_36[345], regroupV0_lo_36[329]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_9 = {regroupV0_lo_36[377], regroupV0_lo_36[361]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_28 = {regroupV0_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_9};
  wire [7:0]        regroupV0_lo_hi_lo_46 = {regroupV0_lo_hi_lo_hi_28, regroupV0_lo_hi_lo_lo_28};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_9 = {regroupV0_lo_36[409], regroupV0_lo_36[393]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_9 = {regroupV0_lo_36[441], regroupV0_lo_36[425]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_28 = {regroupV0_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_9};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_9 = {regroupV0_lo_36[473], regroupV0_lo_36[457]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_9 = {regroupV0_lo_36[505], regroupV0_lo_36[489]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_28 = {regroupV0_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_9};
  wire [7:0]        regroupV0_lo_hi_hi_46 = {regroupV0_lo_hi_hi_hi_28, regroupV0_lo_hi_hi_lo_28};
  wire [15:0]       regroupV0_lo_hi_46 = {regroupV0_lo_hi_hi_46, regroupV0_lo_hi_lo_46};
  wire [31:0]       regroupV0_lo_46 = {regroupV0_lo_hi_46, regroupV0_lo_lo_46};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_9 = {regroupV0_hi_36[25], regroupV0_hi_36[9]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_9 = {regroupV0_hi_36[57], regroupV0_hi_36[41]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_28 = {regroupV0_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_9};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_9 = {regroupV0_hi_36[89], regroupV0_hi_36[73]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_9 = {regroupV0_hi_36[121], regroupV0_hi_36[105]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_28 = {regroupV0_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_9};
  wire [7:0]        regroupV0_hi_lo_lo_46 = {regroupV0_hi_lo_lo_hi_28, regroupV0_hi_lo_lo_lo_28};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_9 = {regroupV0_hi_36[153], regroupV0_hi_36[137]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_9 = {regroupV0_hi_36[185], regroupV0_hi_36[169]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_28 = {regroupV0_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_9};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_9 = {regroupV0_hi_36[217], regroupV0_hi_36[201]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_9 = {regroupV0_hi_36[249], regroupV0_hi_36[233]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_28 = {regroupV0_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_9};
  wire [7:0]        regroupV0_hi_lo_hi_46 = {regroupV0_hi_lo_hi_hi_28, regroupV0_hi_lo_hi_lo_28};
  wire [15:0]       regroupV0_hi_lo_46 = {regroupV0_hi_lo_hi_46, regroupV0_hi_lo_lo_46};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_9 = {regroupV0_hi_36[281], regroupV0_hi_36[265]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_9 = {regroupV0_hi_36[313], regroupV0_hi_36[297]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_28 = {regroupV0_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_9};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_9 = {regroupV0_hi_36[345], regroupV0_hi_36[329]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_9 = {regroupV0_hi_36[377], regroupV0_hi_36[361]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_28 = {regroupV0_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_9};
  wire [7:0]        regroupV0_hi_hi_lo_46 = {regroupV0_hi_hi_lo_hi_28, regroupV0_hi_hi_lo_lo_28};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_9 = {regroupV0_hi_36[409], regroupV0_hi_36[393]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_9 = {regroupV0_hi_36[441], regroupV0_hi_36[425]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_28 = {regroupV0_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_9};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_9 = {regroupV0_hi_36[473], regroupV0_hi_36[457]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_9 = {regroupV0_hi_36[505], regroupV0_hi_36[489]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_28 = {regroupV0_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_9};
  wire [7:0]        regroupV0_hi_hi_hi_46 = {regroupV0_hi_hi_hi_hi_28, regroupV0_hi_hi_hi_lo_28};
  wire [15:0]       regroupV0_hi_hi_46 = {regroupV0_hi_hi_hi_46, regroupV0_hi_hi_lo_46};
  wire [31:0]       regroupV0_hi_46 = {regroupV0_hi_hi_46, regroupV0_hi_lo_46};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_10 = {regroupV0_lo_36[26], regroupV0_lo_36[10]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_10 = {regroupV0_lo_36[58], regroupV0_lo_36[42]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_29 = {regroupV0_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_10};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_10 = {regroupV0_lo_36[90], regroupV0_lo_36[74]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_10 = {regroupV0_lo_36[122], regroupV0_lo_36[106]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_29 = {regroupV0_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_10};
  wire [7:0]        regroupV0_lo_lo_lo_47 = {regroupV0_lo_lo_lo_hi_29, regroupV0_lo_lo_lo_lo_29};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_10 = {regroupV0_lo_36[154], regroupV0_lo_36[138]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_10 = {regroupV0_lo_36[186], regroupV0_lo_36[170]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_29 = {regroupV0_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_10};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_10 = {regroupV0_lo_36[218], regroupV0_lo_36[202]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_10 = {regroupV0_lo_36[250], regroupV0_lo_36[234]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_29 = {regroupV0_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_10};
  wire [7:0]        regroupV0_lo_lo_hi_47 = {regroupV0_lo_lo_hi_hi_29, regroupV0_lo_lo_hi_lo_29};
  wire [15:0]       regroupV0_lo_lo_47 = {regroupV0_lo_lo_hi_47, regroupV0_lo_lo_lo_47};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_10 = {regroupV0_lo_36[282], regroupV0_lo_36[266]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_10 = {regroupV0_lo_36[314], regroupV0_lo_36[298]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_29 = {regroupV0_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_10};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_10 = {regroupV0_lo_36[346], regroupV0_lo_36[330]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_10 = {regroupV0_lo_36[378], regroupV0_lo_36[362]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_29 = {regroupV0_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_10};
  wire [7:0]        regroupV0_lo_hi_lo_47 = {regroupV0_lo_hi_lo_hi_29, regroupV0_lo_hi_lo_lo_29};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_10 = {regroupV0_lo_36[410], regroupV0_lo_36[394]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_10 = {regroupV0_lo_36[442], regroupV0_lo_36[426]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_29 = {regroupV0_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_10};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_10 = {regroupV0_lo_36[474], regroupV0_lo_36[458]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_10 = {regroupV0_lo_36[506], regroupV0_lo_36[490]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_29 = {regroupV0_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_10};
  wire [7:0]        regroupV0_lo_hi_hi_47 = {regroupV0_lo_hi_hi_hi_29, regroupV0_lo_hi_hi_lo_29};
  wire [15:0]       regroupV0_lo_hi_47 = {regroupV0_lo_hi_hi_47, regroupV0_lo_hi_lo_47};
  wire [31:0]       regroupV0_lo_47 = {regroupV0_lo_hi_47, regroupV0_lo_lo_47};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_10 = {regroupV0_hi_36[26], regroupV0_hi_36[10]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_10 = {regroupV0_hi_36[58], regroupV0_hi_36[42]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_29 = {regroupV0_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_10};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_10 = {regroupV0_hi_36[90], regroupV0_hi_36[74]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_10 = {regroupV0_hi_36[122], regroupV0_hi_36[106]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_29 = {regroupV0_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_10};
  wire [7:0]        regroupV0_hi_lo_lo_47 = {regroupV0_hi_lo_lo_hi_29, regroupV0_hi_lo_lo_lo_29};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_10 = {regroupV0_hi_36[154], regroupV0_hi_36[138]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_10 = {regroupV0_hi_36[186], regroupV0_hi_36[170]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_29 = {regroupV0_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_10};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_10 = {regroupV0_hi_36[218], regroupV0_hi_36[202]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_10 = {regroupV0_hi_36[250], regroupV0_hi_36[234]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_29 = {regroupV0_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_10};
  wire [7:0]        regroupV0_hi_lo_hi_47 = {regroupV0_hi_lo_hi_hi_29, regroupV0_hi_lo_hi_lo_29};
  wire [15:0]       regroupV0_hi_lo_47 = {regroupV0_hi_lo_hi_47, regroupV0_hi_lo_lo_47};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_10 = {regroupV0_hi_36[282], regroupV0_hi_36[266]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_10 = {regroupV0_hi_36[314], regroupV0_hi_36[298]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_29 = {regroupV0_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_10};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_10 = {regroupV0_hi_36[346], regroupV0_hi_36[330]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_10 = {regroupV0_hi_36[378], regroupV0_hi_36[362]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_29 = {regroupV0_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_10};
  wire [7:0]        regroupV0_hi_hi_lo_47 = {regroupV0_hi_hi_lo_hi_29, regroupV0_hi_hi_lo_lo_29};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_10 = {regroupV0_hi_36[410], regroupV0_hi_36[394]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_10 = {regroupV0_hi_36[442], regroupV0_hi_36[426]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_29 = {regroupV0_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_10};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_10 = {regroupV0_hi_36[474], regroupV0_hi_36[458]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_10 = {regroupV0_hi_36[506], regroupV0_hi_36[490]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_29 = {regroupV0_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_10};
  wire [7:0]        regroupV0_hi_hi_hi_47 = {regroupV0_hi_hi_hi_hi_29, regroupV0_hi_hi_hi_lo_29};
  wire [15:0]       regroupV0_hi_hi_47 = {regroupV0_hi_hi_hi_47, regroupV0_hi_hi_lo_47};
  wire [31:0]       regroupV0_hi_47 = {regroupV0_hi_hi_47, regroupV0_hi_lo_47};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_11 = {regroupV0_lo_36[27], regroupV0_lo_36[11]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_11 = {regroupV0_lo_36[59], regroupV0_lo_36[43]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_30 = {regroupV0_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_11};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_11 = {regroupV0_lo_36[91], regroupV0_lo_36[75]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_11 = {regroupV0_lo_36[123], regroupV0_lo_36[107]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_30 = {regroupV0_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_11};
  wire [7:0]        regroupV0_lo_lo_lo_48 = {regroupV0_lo_lo_lo_hi_30, regroupV0_lo_lo_lo_lo_30};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_11 = {regroupV0_lo_36[155], regroupV0_lo_36[139]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_11 = {regroupV0_lo_36[187], regroupV0_lo_36[171]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_30 = {regroupV0_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_11};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_11 = {regroupV0_lo_36[219], regroupV0_lo_36[203]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_11 = {regroupV0_lo_36[251], regroupV0_lo_36[235]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_30 = {regroupV0_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_11};
  wire [7:0]        regroupV0_lo_lo_hi_48 = {regroupV0_lo_lo_hi_hi_30, regroupV0_lo_lo_hi_lo_30};
  wire [15:0]       regroupV0_lo_lo_48 = {regroupV0_lo_lo_hi_48, regroupV0_lo_lo_lo_48};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_11 = {regroupV0_lo_36[283], regroupV0_lo_36[267]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_11 = {regroupV0_lo_36[315], regroupV0_lo_36[299]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_30 = {regroupV0_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_11};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_11 = {regroupV0_lo_36[347], regroupV0_lo_36[331]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_11 = {regroupV0_lo_36[379], regroupV0_lo_36[363]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_30 = {regroupV0_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_11};
  wire [7:0]        regroupV0_lo_hi_lo_48 = {regroupV0_lo_hi_lo_hi_30, regroupV0_lo_hi_lo_lo_30};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_11 = {regroupV0_lo_36[411], regroupV0_lo_36[395]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_11 = {regroupV0_lo_36[443], regroupV0_lo_36[427]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_30 = {regroupV0_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_11};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_11 = {regroupV0_lo_36[475], regroupV0_lo_36[459]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_11 = {regroupV0_lo_36[507], regroupV0_lo_36[491]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_30 = {regroupV0_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_11};
  wire [7:0]        regroupV0_lo_hi_hi_48 = {regroupV0_lo_hi_hi_hi_30, regroupV0_lo_hi_hi_lo_30};
  wire [15:0]       regroupV0_lo_hi_48 = {regroupV0_lo_hi_hi_48, regroupV0_lo_hi_lo_48};
  wire [31:0]       regroupV0_lo_48 = {regroupV0_lo_hi_48, regroupV0_lo_lo_48};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_11 = {regroupV0_hi_36[27], regroupV0_hi_36[11]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_11 = {regroupV0_hi_36[59], regroupV0_hi_36[43]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_30 = {regroupV0_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_11};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_11 = {regroupV0_hi_36[91], regroupV0_hi_36[75]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_11 = {regroupV0_hi_36[123], regroupV0_hi_36[107]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_30 = {regroupV0_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_11};
  wire [7:0]        regroupV0_hi_lo_lo_48 = {regroupV0_hi_lo_lo_hi_30, regroupV0_hi_lo_lo_lo_30};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_11 = {regroupV0_hi_36[155], regroupV0_hi_36[139]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_11 = {regroupV0_hi_36[187], regroupV0_hi_36[171]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_30 = {regroupV0_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_11};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_11 = {regroupV0_hi_36[219], regroupV0_hi_36[203]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_11 = {regroupV0_hi_36[251], regroupV0_hi_36[235]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_30 = {regroupV0_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_11};
  wire [7:0]        regroupV0_hi_lo_hi_48 = {regroupV0_hi_lo_hi_hi_30, regroupV0_hi_lo_hi_lo_30};
  wire [15:0]       regroupV0_hi_lo_48 = {regroupV0_hi_lo_hi_48, regroupV0_hi_lo_lo_48};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_11 = {regroupV0_hi_36[283], regroupV0_hi_36[267]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_11 = {regroupV0_hi_36[315], regroupV0_hi_36[299]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_30 = {regroupV0_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_11};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_11 = {regroupV0_hi_36[347], regroupV0_hi_36[331]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_11 = {regroupV0_hi_36[379], regroupV0_hi_36[363]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_30 = {regroupV0_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_11};
  wire [7:0]        regroupV0_hi_hi_lo_48 = {regroupV0_hi_hi_lo_hi_30, regroupV0_hi_hi_lo_lo_30};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_11 = {regroupV0_hi_36[411], regroupV0_hi_36[395]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_11 = {regroupV0_hi_36[443], regroupV0_hi_36[427]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_30 = {regroupV0_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_11};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_11 = {regroupV0_hi_36[475], regroupV0_hi_36[459]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_11 = {regroupV0_hi_36[507], regroupV0_hi_36[491]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_30 = {regroupV0_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_11};
  wire [7:0]        regroupV0_hi_hi_hi_48 = {regroupV0_hi_hi_hi_hi_30, regroupV0_hi_hi_hi_lo_30};
  wire [15:0]       regroupV0_hi_hi_48 = {regroupV0_hi_hi_hi_48, regroupV0_hi_hi_lo_48};
  wire [31:0]       regroupV0_hi_48 = {regroupV0_hi_hi_48, regroupV0_hi_lo_48};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_12 = {regroupV0_lo_36[28], regroupV0_lo_36[12]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_12 = {regroupV0_lo_36[60], regroupV0_lo_36[44]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_31 = {regroupV0_lo_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_lo_12};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_12 = {regroupV0_lo_36[92], regroupV0_lo_36[76]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_12 = {regroupV0_lo_36[124], regroupV0_lo_36[108]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_31 = {regroupV0_lo_lo_lo_hi_hi_12, regroupV0_lo_lo_lo_hi_lo_12};
  wire [7:0]        regroupV0_lo_lo_lo_49 = {regroupV0_lo_lo_lo_hi_31, regroupV0_lo_lo_lo_lo_31};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_12 = {regroupV0_lo_36[156], regroupV0_lo_36[140]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_12 = {regroupV0_lo_36[188], regroupV0_lo_36[172]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_31 = {regroupV0_lo_lo_hi_lo_hi_12, regroupV0_lo_lo_hi_lo_lo_12};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_12 = {regroupV0_lo_36[220], regroupV0_lo_36[204]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_12 = {regroupV0_lo_36[252], regroupV0_lo_36[236]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_31 = {regroupV0_lo_lo_hi_hi_hi_12, regroupV0_lo_lo_hi_hi_lo_12};
  wire [7:0]        regroupV0_lo_lo_hi_49 = {regroupV0_lo_lo_hi_hi_31, regroupV0_lo_lo_hi_lo_31};
  wire [15:0]       regroupV0_lo_lo_49 = {regroupV0_lo_lo_hi_49, regroupV0_lo_lo_lo_49};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_12 = {regroupV0_lo_36[284], regroupV0_lo_36[268]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_12 = {regroupV0_lo_36[316], regroupV0_lo_36[300]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_31 = {regroupV0_lo_hi_lo_lo_hi_12, regroupV0_lo_hi_lo_lo_lo_12};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_12 = {regroupV0_lo_36[348], regroupV0_lo_36[332]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_12 = {regroupV0_lo_36[380], regroupV0_lo_36[364]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_31 = {regroupV0_lo_hi_lo_hi_hi_12, regroupV0_lo_hi_lo_hi_lo_12};
  wire [7:0]        regroupV0_lo_hi_lo_49 = {regroupV0_lo_hi_lo_hi_31, regroupV0_lo_hi_lo_lo_31};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_12 = {regroupV0_lo_36[412], regroupV0_lo_36[396]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_12 = {regroupV0_lo_36[444], regroupV0_lo_36[428]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_31 = {regroupV0_lo_hi_hi_lo_hi_12, regroupV0_lo_hi_hi_lo_lo_12};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_12 = {regroupV0_lo_36[476], regroupV0_lo_36[460]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_12 = {regroupV0_lo_36[508], regroupV0_lo_36[492]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_31 = {regroupV0_lo_hi_hi_hi_hi_12, regroupV0_lo_hi_hi_hi_lo_12};
  wire [7:0]        regroupV0_lo_hi_hi_49 = {regroupV0_lo_hi_hi_hi_31, regroupV0_lo_hi_hi_lo_31};
  wire [15:0]       regroupV0_lo_hi_49 = {regroupV0_lo_hi_hi_49, regroupV0_lo_hi_lo_49};
  wire [31:0]       regroupV0_lo_49 = {regroupV0_lo_hi_49, regroupV0_lo_lo_49};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_12 = {regroupV0_hi_36[28], regroupV0_hi_36[12]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_12 = {regroupV0_hi_36[60], regroupV0_hi_36[44]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_31 = {regroupV0_hi_lo_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_lo_12};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_12 = {regroupV0_hi_36[92], regroupV0_hi_36[76]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_12 = {regroupV0_hi_36[124], regroupV0_hi_36[108]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_31 = {regroupV0_hi_lo_lo_hi_hi_12, regroupV0_hi_lo_lo_hi_lo_12};
  wire [7:0]        regroupV0_hi_lo_lo_49 = {regroupV0_hi_lo_lo_hi_31, regroupV0_hi_lo_lo_lo_31};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_12 = {regroupV0_hi_36[156], regroupV0_hi_36[140]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_12 = {regroupV0_hi_36[188], regroupV0_hi_36[172]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_31 = {regroupV0_hi_lo_hi_lo_hi_12, regroupV0_hi_lo_hi_lo_lo_12};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_12 = {regroupV0_hi_36[220], regroupV0_hi_36[204]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_12 = {regroupV0_hi_36[252], regroupV0_hi_36[236]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_31 = {regroupV0_hi_lo_hi_hi_hi_12, regroupV0_hi_lo_hi_hi_lo_12};
  wire [7:0]        regroupV0_hi_lo_hi_49 = {regroupV0_hi_lo_hi_hi_31, regroupV0_hi_lo_hi_lo_31};
  wire [15:0]       regroupV0_hi_lo_49 = {regroupV0_hi_lo_hi_49, regroupV0_hi_lo_lo_49};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_12 = {regroupV0_hi_36[284], regroupV0_hi_36[268]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_12 = {regroupV0_hi_36[316], regroupV0_hi_36[300]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_31 = {regroupV0_hi_hi_lo_lo_hi_12, regroupV0_hi_hi_lo_lo_lo_12};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_12 = {regroupV0_hi_36[348], regroupV0_hi_36[332]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_12 = {regroupV0_hi_36[380], regroupV0_hi_36[364]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_31 = {regroupV0_hi_hi_lo_hi_hi_12, regroupV0_hi_hi_lo_hi_lo_12};
  wire [7:0]        regroupV0_hi_hi_lo_49 = {regroupV0_hi_hi_lo_hi_31, regroupV0_hi_hi_lo_lo_31};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_12 = {regroupV0_hi_36[412], regroupV0_hi_36[396]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_12 = {regroupV0_hi_36[444], regroupV0_hi_36[428]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_31 = {regroupV0_hi_hi_hi_lo_hi_12, regroupV0_hi_hi_hi_lo_lo_12};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_12 = {regroupV0_hi_36[476], regroupV0_hi_36[460]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_12 = {regroupV0_hi_36[508], regroupV0_hi_36[492]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_31 = {regroupV0_hi_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_hi_lo_12};
  wire [7:0]        regroupV0_hi_hi_hi_49 = {regroupV0_hi_hi_hi_hi_31, regroupV0_hi_hi_hi_lo_31};
  wire [15:0]       regroupV0_hi_hi_49 = {regroupV0_hi_hi_hi_49, regroupV0_hi_hi_lo_49};
  wire [31:0]       regroupV0_hi_49 = {regroupV0_hi_hi_49, regroupV0_hi_lo_49};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_13 = {regroupV0_lo_36[29], regroupV0_lo_36[13]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_13 = {regroupV0_lo_36[61], regroupV0_lo_36[45]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_32 = {regroupV0_lo_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_lo_13};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_13 = {regroupV0_lo_36[93], regroupV0_lo_36[77]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_13 = {regroupV0_lo_36[125], regroupV0_lo_36[109]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_32 = {regroupV0_lo_lo_lo_hi_hi_13, regroupV0_lo_lo_lo_hi_lo_13};
  wire [7:0]        regroupV0_lo_lo_lo_50 = {regroupV0_lo_lo_lo_hi_32, regroupV0_lo_lo_lo_lo_32};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_13 = {regroupV0_lo_36[157], regroupV0_lo_36[141]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_13 = {regroupV0_lo_36[189], regroupV0_lo_36[173]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_32 = {regroupV0_lo_lo_hi_lo_hi_13, regroupV0_lo_lo_hi_lo_lo_13};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_13 = {regroupV0_lo_36[221], regroupV0_lo_36[205]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_13 = {regroupV0_lo_36[253], regroupV0_lo_36[237]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_32 = {regroupV0_lo_lo_hi_hi_hi_13, regroupV0_lo_lo_hi_hi_lo_13};
  wire [7:0]        regroupV0_lo_lo_hi_50 = {regroupV0_lo_lo_hi_hi_32, regroupV0_lo_lo_hi_lo_32};
  wire [15:0]       regroupV0_lo_lo_50 = {regroupV0_lo_lo_hi_50, regroupV0_lo_lo_lo_50};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_13 = {regroupV0_lo_36[285], regroupV0_lo_36[269]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_13 = {regroupV0_lo_36[317], regroupV0_lo_36[301]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_32 = {regroupV0_lo_hi_lo_lo_hi_13, regroupV0_lo_hi_lo_lo_lo_13};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_13 = {regroupV0_lo_36[349], regroupV0_lo_36[333]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_13 = {regroupV0_lo_36[381], regroupV0_lo_36[365]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_32 = {regroupV0_lo_hi_lo_hi_hi_13, regroupV0_lo_hi_lo_hi_lo_13};
  wire [7:0]        regroupV0_lo_hi_lo_50 = {regroupV0_lo_hi_lo_hi_32, regroupV0_lo_hi_lo_lo_32};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_13 = {regroupV0_lo_36[413], regroupV0_lo_36[397]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_13 = {regroupV0_lo_36[445], regroupV0_lo_36[429]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_32 = {regroupV0_lo_hi_hi_lo_hi_13, regroupV0_lo_hi_hi_lo_lo_13};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_13 = {regroupV0_lo_36[477], regroupV0_lo_36[461]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_13 = {regroupV0_lo_36[509], regroupV0_lo_36[493]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_32 = {regroupV0_lo_hi_hi_hi_hi_13, regroupV0_lo_hi_hi_hi_lo_13};
  wire [7:0]        regroupV0_lo_hi_hi_50 = {regroupV0_lo_hi_hi_hi_32, regroupV0_lo_hi_hi_lo_32};
  wire [15:0]       regroupV0_lo_hi_50 = {regroupV0_lo_hi_hi_50, regroupV0_lo_hi_lo_50};
  wire [31:0]       regroupV0_lo_50 = {regroupV0_lo_hi_50, regroupV0_lo_lo_50};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_13 = {regroupV0_hi_36[29], regroupV0_hi_36[13]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_13 = {regroupV0_hi_36[61], regroupV0_hi_36[45]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_32 = {regroupV0_hi_lo_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_lo_13};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_13 = {regroupV0_hi_36[93], regroupV0_hi_36[77]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_13 = {regroupV0_hi_36[125], regroupV0_hi_36[109]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_32 = {regroupV0_hi_lo_lo_hi_hi_13, regroupV0_hi_lo_lo_hi_lo_13};
  wire [7:0]        regroupV0_hi_lo_lo_50 = {regroupV0_hi_lo_lo_hi_32, regroupV0_hi_lo_lo_lo_32};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_13 = {regroupV0_hi_36[157], regroupV0_hi_36[141]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_13 = {regroupV0_hi_36[189], regroupV0_hi_36[173]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_32 = {regroupV0_hi_lo_hi_lo_hi_13, regroupV0_hi_lo_hi_lo_lo_13};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_13 = {regroupV0_hi_36[221], regroupV0_hi_36[205]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_13 = {regroupV0_hi_36[253], regroupV0_hi_36[237]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_32 = {regroupV0_hi_lo_hi_hi_hi_13, regroupV0_hi_lo_hi_hi_lo_13};
  wire [7:0]        regroupV0_hi_lo_hi_50 = {regroupV0_hi_lo_hi_hi_32, regroupV0_hi_lo_hi_lo_32};
  wire [15:0]       regroupV0_hi_lo_50 = {regroupV0_hi_lo_hi_50, regroupV0_hi_lo_lo_50};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_13 = {regroupV0_hi_36[285], regroupV0_hi_36[269]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_13 = {regroupV0_hi_36[317], regroupV0_hi_36[301]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_32 = {regroupV0_hi_hi_lo_lo_hi_13, regroupV0_hi_hi_lo_lo_lo_13};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_13 = {regroupV0_hi_36[349], regroupV0_hi_36[333]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_13 = {regroupV0_hi_36[381], regroupV0_hi_36[365]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_32 = {regroupV0_hi_hi_lo_hi_hi_13, regroupV0_hi_hi_lo_hi_lo_13};
  wire [7:0]        regroupV0_hi_hi_lo_50 = {regroupV0_hi_hi_lo_hi_32, regroupV0_hi_hi_lo_lo_32};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_13 = {regroupV0_hi_36[413], regroupV0_hi_36[397]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_13 = {regroupV0_hi_36[445], regroupV0_hi_36[429]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_32 = {regroupV0_hi_hi_hi_lo_hi_13, regroupV0_hi_hi_hi_lo_lo_13};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_13 = {regroupV0_hi_36[477], regroupV0_hi_36[461]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_13 = {regroupV0_hi_36[509], regroupV0_hi_36[493]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_32 = {regroupV0_hi_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_hi_lo_13};
  wire [7:0]        regroupV0_hi_hi_hi_50 = {regroupV0_hi_hi_hi_hi_32, regroupV0_hi_hi_hi_lo_32};
  wire [15:0]       regroupV0_hi_hi_50 = {regroupV0_hi_hi_hi_50, regroupV0_hi_hi_lo_50};
  wire [31:0]       regroupV0_hi_50 = {regroupV0_hi_hi_50, regroupV0_hi_lo_50};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_14 = {regroupV0_lo_36[30], regroupV0_lo_36[14]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_14 = {regroupV0_lo_36[62], regroupV0_lo_36[46]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_33 = {regroupV0_lo_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_lo_14};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_14 = {regroupV0_lo_36[94], regroupV0_lo_36[78]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_14 = {regroupV0_lo_36[126], regroupV0_lo_36[110]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_33 = {regroupV0_lo_lo_lo_hi_hi_14, regroupV0_lo_lo_lo_hi_lo_14};
  wire [7:0]        regroupV0_lo_lo_lo_51 = {regroupV0_lo_lo_lo_hi_33, regroupV0_lo_lo_lo_lo_33};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_14 = {regroupV0_lo_36[158], regroupV0_lo_36[142]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_14 = {regroupV0_lo_36[190], regroupV0_lo_36[174]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_33 = {regroupV0_lo_lo_hi_lo_hi_14, regroupV0_lo_lo_hi_lo_lo_14};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_14 = {regroupV0_lo_36[222], regroupV0_lo_36[206]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_14 = {regroupV0_lo_36[254], regroupV0_lo_36[238]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_33 = {regroupV0_lo_lo_hi_hi_hi_14, regroupV0_lo_lo_hi_hi_lo_14};
  wire [7:0]        regroupV0_lo_lo_hi_51 = {regroupV0_lo_lo_hi_hi_33, regroupV0_lo_lo_hi_lo_33};
  wire [15:0]       regroupV0_lo_lo_51 = {regroupV0_lo_lo_hi_51, regroupV0_lo_lo_lo_51};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_14 = {regroupV0_lo_36[286], regroupV0_lo_36[270]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_14 = {regroupV0_lo_36[318], regroupV0_lo_36[302]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_33 = {regroupV0_lo_hi_lo_lo_hi_14, regroupV0_lo_hi_lo_lo_lo_14};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_14 = {regroupV0_lo_36[350], regroupV0_lo_36[334]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_14 = {regroupV0_lo_36[382], regroupV0_lo_36[366]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_33 = {regroupV0_lo_hi_lo_hi_hi_14, regroupV0_lo_hi_lo_hi_lo_14};
  wire [7:0]        regroupV0_lo_hi_lo_51 = {regroupV0_lo_hi_lo_hi_33, regroupV0_lo_hi_lo_lo_33};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_14 = {regroupV0_lo_36[414], regroupV0_lo_36[398]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_14 = {regroupV0_lo_36[446], regroupV0_lo_36[430]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_33 = {regroupV0_lo_hi_hi_lo_hi_14, regroupV0_lo_hi_hi_lo_lo_14};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_14 = {regroupV0_lo_36[478], regroupV0_lo_36[462]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_14 = {regroupV0_lo_36[510], regroupV0_lo_36[494]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_33 = {regroupV0_lo_hi_hi_hi_hi_14, regroupV0_lo_hi_hi_hi_lo_14};
  wire [7:0]        regroupV0_lo_hi_hi_51 = {regroupV0_lo_hi_hi_hi_33, regroupV0_lo_hi_hi_lo_33};
  wire [15:0]       regroupV0_lo_hi_51 = {regroupV0_lo_hi_hi_51, regroupV0_lo_hi_lo_51};
  wire [31:0]       regroupV0_lo_51 = {regroupV0_lo_hi_51, regroupV0_lo_lo_51};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_14 = {regroupV0_hi_36[30], regroupV0_hi_36[14]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_14 = {regroupV0_hi_36[62], regroupV0_hi_36[46]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_33 = {regroupV0_hi_lo_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_lo_14};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_14 = {regroupV0_hi_36[94], regroupV0_hi_36[78]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_14 = {regroupV0_hi_36[126], regroupV0_hi_36[110]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_33 = {regroupV0_hi_lo_lo_hi_hi_14, regroupV0_hi_lo_lo_hi_lo_14};
  wire [7:0]        regroupV0_hi_lo_lo_51 = {regroupV0_hi_lo_lo_hi_33, regroupV0_hi_lo_lo_lo_33};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_14 = {regroupV0_hi_36[158], regroupV0_hi_36[142]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_14 = {regroupV0_hi_36[190], regroupV0_hi_36[174]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_33 = {regroupV0_hi_lo_hi_lo_hi_14, regroupV0_hi_lo_hi_lo_lo_14};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_14 = {regroupV0_hi_36[222], regroupV0_hi_36[206]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_14 = {regroupV0_hi_36[254], regroupV0_hi_36[238]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_33 = {regroupV0_hi_lo_hi_hi_hi_14, regroupV0_hi_lo_hi_hi_lo_14};
  wire [7:0]        regroupV0_hi_lo_hi_51 = {regroupV0_hi_lo_hi_hi_33, regroupV0_hi_lo_hi_lo_33};
  wire [15:0]       regroupV0_hi_lo_51 = {regroupV0_hi_lo_hi_51, regroupV0_hi_lo_lo_51};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_14 = {regroupV0_hi_36[286], regroupV0_hi_36[270]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_14 = {regroupV0_hi_36[318], regroupV0_hi_36[302]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_33 = {regroupV0_hi_hi_lo_lo_hi_14, regroupV0_hi_hi_lo_lo_lo_14};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_14 = {regroupV0_hi_36[350], regroupV0_hi_36[334]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_14 = {regroupV0_hi_36[382], regroupV0_hi_36[366]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_33 = {regroupV0_hi_hi_lo_hi_hi_14, regroupV0_hi_hi_lo_hi_lo_14};
  wire [7:0]        regroupV0_hi_hi_lo_51 = {regroupV0_hi_hi_lo_hi_33, regroupV0_hi_hi_lo_lo_33};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_14 = {regroupV0_hi_36[414], regroupV0_hi_36[398]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_14 = {regroupV0_hi_36[446], regroupV0_hi_36[430]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_33 = {regroupV0_hi_hi_hi_lo_hi_14, regroupV0_hi_hi_hi_lo_lo_14};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_14 = {regroupV0_hi_36[478], regroupV0_hi_36[462]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_14 = {regroupV0_hi_36[510], regroupV0_hi_36[494]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_33 = {regroupV0_hi_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_hi_lo_14};
  wire [7:0]        regroupV0_hi_hi_hi_51 = {regroupV0_hi_hi_hi_hi_33, regroupV0_hi_hi_hi_lo_33};
  wire [15:0]       regroupV0_hi_hi_51 = {regroupV0_hi_hi_hi_51, regroupV0_hi_hi_lo_51};
  wire [31:0]       regroupV0_hi_51 = {regroupV0_hi_hi_51, regroupV0_hi_lo_51};
  wire [1:0]        regroupV0_lo_lo_lo_lo_lo_15 = {regroupV0_lo_36[31], regroupV0_lo_36[15]};
  wire [1:0]        regroupV0_lo_lo_lo_lo_hi_15 = {regroupV0_lo_36[63], regroupV0_lo_36[47]};
  wire [3:0]        regroupV0_lo_lo_lo_lo_34 = {regroupV0_lo_lo_lo_lo_hi_15, regroupV0_lo_lo_lo_lo_lo_15};
  wire [1:0]        regroupV0_lo_lo_lo_hi_lo_15 = {regroupV0_lo_36[95], regroupV0_lo_36[79]};
  wire [1:0]        regroupV0_lo_lo_lo_hi_hi_15 = {regroupV0_lo_36[127], regroupV0_lo_36[111]};
  wire [3:0]        regroupV0_lo_lo_lo_hi_34 = {regroupV0_lo_lo_lo_hi_hi_15, regroupV0_lo_lo_lo_hi_lo_15};
  wire [7:0]        regroupV0_lo_lo_lo_52 = {regroupV0_lo_lo_lo_hi_34, regroupV0_lo_lo_lo_lo_34};
  wire [1:0]        regroupV0_lo_lo_hi_lo_lo_15 = {regroupV0_lo_36[159], regroupV0_lo_36[143]};
  wire [1:0]        regroupV0_lo_lo_hi_lo_hi_15 = {regroupV0_lo_36[191], regroupV0_lo_36[175]};
  wire [3:0]        regroupV0_lo_lo_hi_lo_34 = {regroupV0_lo_lo_hi_lo_hi_15, regroupV0_lo_lo_hi_lo_lo_15};
  wire [1:0]        regroupV0_lo_lo_hi_hi_lo_15 = {regroupV0_lo_36[223], regroupV0_lo_36[207]};
  wire [1:0]        regroupV0_lo_lo_hi_hi_hi_15 = {regroupV0_lo_36[255], regroupV0_lo_36[239]};
  wire [3:0]        regroupV0_lo_lo_hi_hi_34 = {regroupV0_lo_lo_hi_hi_hi_15, regroupV0_lo_lo_hi_hi_lo_15};
  wire [7:0]        regroupV0_lo_lo_hi_52 = {regroupV0_lo_lo_hi_hi_34, regroupV0_lo_lo_hi_lo_34};
  wire [15:0]       regroupV0_lo_lo_52 = {regroupV0_lo_lo_hi_52, regroupV0_lo_lo_lo_52};
  wire [1:0]        regroupV0_lo_hi_lo_lo_lo_15 = {regroupV0_lo_36[287], regroupV0_lo_36[271]};
  wire [1:0]        regroupV0_lo_hi_lo_lo_hi_15 = {regroupV0_lo_36[319], regroupV0_lo_36[303]};
  wire [3:0]        regroupV0_lo_hi_lo_lo_34 = {regroupV0_lo_hi_lo_lo_hi_15, regroupV0_lo_hi_lo_lo_lo_15};
  wire [1:0]        regroupV0_lo_hi_lo_hi_lo_15 = {regroupV0_lo_36[351], regroupV0_lo_36[335]};
  wire [1:0]        regroupV0_lo_hi_lo_hi_hi_15 = {regroupV0_lo_36[383], regroupV0_lo_36[367]};
  wire [3:0]        regroupV0_lo_hi_lo_hi_34 = {regroupV0_lo_hi_lo_hi_hi_15, regroupV0_lo_hi_lo_hi_lo_15};
  wire [7:0]        regroupV0_lo_hi_lo_52 = {regroupV0_lo_hi_lo_hi_34, regroupV0_lo_hi_lo_lo_34};
  wire [1:0]        regroupV0_lo_hi_hi_lo_lo_15 = {regroupV0_lo_36[415], regroupV0_lo_36[399]};
  wire [1:0]        regroupV0_lo_hi_hi_lo_hi_15 = {regroupV0_lo_36[447], regroupV0_lo_36[431]};
  wire [3:0]        regroupV0_lo_hi_hi_lo_34 = {regroupV0_lo_hi_hi_lo_hi_15, regroupV0_lo_hi_hi_lo_lo_15};
  wire [1:0]        regroupV0_lo_hi_hi_hi_lo_15 = {regroupV0_lo_36[479], regroupV0_lo_36[463]};
  wire [1:0]        regroupV0_lo_hi_hi_hi_hi_15 = {regroupV0_lo_36[511], regroupV0_lo_36[495]};
  wire [3:0]        regroupV0_lo_hi_hi_hi_34 = {regroupV0_lo_hi_hi_hi_hi_15, regroupV0_lo_hi_hi_hi_lo_15};
  wire [7:0]        regroupV0_lo_hi_hi_52 = {regroupV0_lo_hi_hi_hi_34, regroupV0_lo_hi_hi_lo_34};
  wire [15:0]       regroupV0_lo_hi_52 = {regroupV0_lo_hi_hi_52, regroupV0_lo_hi_lo_52};
  wire [31:0]       regroupV0_lo_52 = {regroupV0_lo_hi_52, regroupV0_lo_lo_52};
  wire [1:0]        regroupV0_hi_lo_lo_lo_lo_15 = {regroupV0_hi_36[31], regroupV0_hi_36[15]};
  wire [1:0]        regroupV0_hi_lo_lo_lo_hi_15 = {regroupV0_hi_36[63], regroupV0_hi_36[47]};
  wire [3:0]        regroupV0_hi_lo_lo_lo_34 = {regroupV0_hi_lo_lo_lo_hi_15, regroupV0_hi_lo_lo_lo_lo_15};
  wire [1:0]        regroupV0_hi_lo_lo_hi_lo_15 = {regroupV0_hi_36[95], regroupV0_hi_36[79]};
  wire [1:0]        regroupV0_hi_lo_lo_hi_hi_15 = {regroupV0_hi_36[127], regroupV0_hi_36[111]};
  wire [3:0]        regroupV0_hi_lo_lo_hi_34 = {regroupV0_hi_lo_lo_hi_hi_15, regroupV0_hi_lo_lo_hi_lo_15};
  wire [7:0]        regroupV0_hi_lo_lo_52 = {regroupV0_hi_lo_lo_hi_34, regroupV0_hi_lo_lo_lo_34};
  wire [1:0]        regroupV0_hi_lo_hi_lo_lo_15 = {regroupV0_hi_36[159], regroupV0_hi_36[143]};
  wire [1:0]        regroupV0_hi_lo_hi_lo_hi_15 = {regroupV0_hi_36[191], regroupV0_hi_36[175]};
  wire [3:0]        regroupV0_hi_lo_hi_lo_34 = {regroupV0_hi_lo_hi_lo_hi_15, regroupV0_hi_lo_hi_lo_lo_15};
  wire [1:0]        regroupV0_hi_lo_hi_hi_lo_15 = {regroupV0_hi_36[223], regroupV0_hi_36[207]};
  wire [1:0]        regroupV0_hi_lo_hi_hi_hi_15 = {regroupV0_hi_36[255], regroupV0_hi_36[239]};
  wire [3:0]        regroupV0_hi_lo_hi_hi_34 = {regroupV0_hi_lo_hi_hi_hi_15, regroupV0_hi_lo_hi_hi_lo_15};
  wire [7:0]        regroupV0_hi_lo_hi_52 = {regroupV0_hi_lo_hi_hi_34, regroupV0_hi_lo_hi_lo_34};
  wire [15:0]       regroupV0_hi_lo_52 = {regroupV0_hi_lo_hi_52, regroupV0_hi_lo_lo_52};
  wire [1:0]        regroupV0_hi_hi_lo_lo_lo_15 = {regroupV0_hi_36[287], regroupV0_hi_36[271]};
  wire [1:0]        regroupV0_hi_hi_lo_lo_hi_15 = {regroupV0_hi_36[319], regroupV0_hi_36[303]};
  wire [3:0]        regroupV0_hi_hi_lo_lo_34 = {regroupV0_hi_hi_lo_lo_hi_15, regroupV0_hi_hi_lo_lo_lo_15};
  wire [1:0]        regroupV0_hi_hi_lo_hi_lo_15 = {regroupV0_hi_36[351], regroupV0_hi_36[335]};
  wire [1:0]        regroupV0_hi_hi_lo_hi_hi_15 = {regroupV0_hi_36[383], regroupV0_hi_36[367]};
  wire [3:0]        regroupV0_hi_hi_lo_hi_34 = {regroupV0_hi_hi_lo_hi_hi_15, regroupV0_hi_hi_lo_hi_lo_15};
  wire [7:0]        regroupV0_hi_hi_lo_52 = {regroupV0_hi_hi_lo_hi_34, regroupV0_hi_hi_lo_lo_34};
  wire [1:0]        regroupV0_hi_hi_hi_lo_lo_15 = {regroupV0_hi_36[415], regroupV0_hi_36[399]};
  wire [1:0]        regroupV0_hi_hi_hi_lo_hi_15 = {regroupV0_hi_36[447], regroupV0_hi_36[431]};
  wire [3:0]        regroupV0_hi_hi_hi_lo_34 = {regroupV0_hi_hi_hi_lo_hi_15, regroupV0_hi_hi_hi_lo_lo_15};
  wire [1:0]        regroupV0_hi_hi_hi_hi_lo_15 = {regroupV0_hi_36[479], regroupV0_hi_36[463]};
  wire [1:0]        regroupV0_hi_hi_hi_hi_hi_15 = {regroupV0_hi_36[511], regroupV0_hi_36[495]};
  wire [3:0]        regroupV0_hi_hi_hi_hi_34 = {regroupV0_hi_hi_hi_hi_hi_15, regroupV0_hi_hi_hi_hi_lo_15};
  wire [7:0]        regroupV0_hi_hi_hi_52 = {regroupV0_hi_hi_hi_hi_34, regroupV0_hi_hi_hi_lo_34};
  wire [15:0]       regroupV0_hi_hi_52 = {regroupV0_hi_hi_hi_52, regroupV0_hi_hi_lo_52};
  wire [31:0]       regroupV0_hi_52 = {regroupV0_hi_hi_52, regroupV0_hi_lo_52};
  wire [127:0]      regroupV0_lo_lo_lo_53 = {regroupV0_hi_38, regroupV0_lo_38, regroupV0_hi_37, regroupV0_lo_37};
  wire [127:0]      regroupV0_lo_lo_hi_53 = {regroupV0_hi_40, regroupV0_lo_40, regroupV0_hi_39, regroupV0_lo_39};
  wire [255:0]      regroupV0_lo_lo_53 = {regroupV0_lo_lo_hi_53, regroupV0_lo_lo_lo_53};
  wire [127:0]      regroupV0_lo_hi_lo_53 = {regroupV0_hi_42, regroupV0_lo_42, regroupV0_hi_41, regroupV0_lo_41};
  wire [127:0]      regroupV0_lo_hi_hi_53 = {regroupV0_hi_44, regroupV0_lo_44, regroupV0_hi_43, regroupV0_lo_43};
  wire [255:0]      regroupV0_lo_hi_53 = {regroupV0_lo_hi_hi_53, regroupV0_lo_hi_lo_53};
  wire [511:0]      regroupV0_lo_53 = {regroupV0_lo_hi_53, regroupV0_lo_lo_53};
  wire [127:0]      regroupV0_hi_lo_lo_53 = {regroupV0_hi_46, regroupV0_lo_46, regroupV0_hi_45, regroupV0_lo_45};
  wire [127:0]      regroupV0_hi_lo_hi_53 = {regroupV0_hi_48, regroupV0_lo_48, regroupV0_hi_47, regroupV0_lo_47};
  wire [255:0]      regroupV0_hi_lo_53 = {regroupV0_hi_lo_hi_53, regroupV0_hi_lo_lo_53};
  wire [127:0]      regroupV0_hi_hi_lo_53 = {regroupV0_hi_50, regroupV0_lo_50, regroupV0_hi_49, regroupV0_lo_49};
  wire [127:0]      regroupV0_hi_hi_hi_53 = {regroupV0_hi_52, regroupV0_lo_52, regroupV0_hi_51, regroupV0_lo_51};
  wire [255:0]      regroupV0_hi_hi_53 = {regroupV0_hi_hi_hi_53, regroupV0_hi_hi_lo_53};
  wire [511:0]      regroupV0_hi_53 = {regroupV0_hi_hi_53, regroupV0_hi_lo_53};
  wire [1023:0]     regroupV0_2 = {regroupV0_hi_53, regroupV0_lo_53};
  wire [3:0]        _v0SelectBySew_T = 4'h1 << laneMaskSewSelect_0;
  wire [63:0]       v0SelectBySew = (_v0SelectBySew_T[0] ? regroupV0_0[63:0] : 64'h0) | (_v0SelectBySew_T[1] ? regroupV0_1[63:0] : 64'h0) | (_v0SelectBySew_T[2] ? regroupV0_2[63:0] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_9 = 4'h1 << laneMaskSewSelect_1;
  wire [63:0]       v0SelectBySew_1 = (_v0SelectBySew_T_9[0] ? regroupV0_0[127:64] : 64'h0) | (_v0SelectBySew_T_9[1] ? regroupV0_1[127:64] : 64'h0) | (_v0SelectBySew_T_9[2] ? regroupV0_2[127:64] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_18 = 4'h1 << laneMaskSewSelect_2;
  wire [63:0]       v0SelectBySew_2 = (_v0SelectBySew_T_18[0] ? regroupV0_0[191:128] : 64'h0) | (_v0SelectBySew_T_18[1] ? regroupV0_1[191:128] : 64'h0) | (_v0SelectBySew_T_18[2] ? regroupV0_2[191:128] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_27 = 4'h1 << laneMaskSewSelect_3;
  wire [63:0]       v0SelectBySew_3 = (_v0SelectBySew_T_27[0] ? regroupV0_0[255:192] : 64'h0) | (_v0SelectBySew_T_27[1] ? regroupV0_1[255:192] : 64'h0) | (_v0SelectBySew_T_27[2] ? regroupV0_2[255:192] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_36 = 4'h1 << laneMaskSewSelect_4;
  wire [63:0]       v0SelectBySew_4 = (_v0SelectBySew_T_36[0] ? regroupV0_0[319:256] : 64'h0) | (_v0SelectBySew_T_36[1] ? regroupV0_1[319:256] : 64'h0) | (_v0SelectBySew_T_36[2] ? regroupV0_2[319:256] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_45 = 4'h1 << laneMaskSewSelect_5;
  wire [63:0]       v0SelectBySew_5 = (_v0SelectBySew_T_45[0] ? regroupV0_0[383:320] : 64'h0) | (_v0SelectBySew_T_45[1] ? regroupV0_1[383:320] : 64'h0) | (_v0SelectBySew_T_45[2] ? regroupV0_2[383:320] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_54 = 4'h1 << laneMaskSewSelect_6;
  wire [63:0]       v0SelectBySew_6 = (_v0SelectBySew_T_54[0] ? regroupV0_0[447:384] : 64'h0) | (_v0SelectBySew_T_54[1] ? regroupV0_1[447:384] : 64'h0) | (_v0SelectBySew_T_54[2] ? regroupV0_2[447:384] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_63 = 4'h1 << laneMaskSewSelect_7;
  wire [63:0]       v0SelectBySew_7 = (_v0SelectBySew_T_63[0] ? regroupV0_0[511:448] : 64'h0) | (_v0SelectBySew_T_63[1] ? regroupV0_1[511:448] : 64'h0) | (_v0SelectBySew_T_63[2] ? regroupV0_2[511:448] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_72 = 4'h1 << laneMaskSewSelect_8;
  wire [63:0]       v0SelectBySew_8 = (_v0SelectBySew_T_72[0] ? regroupV0_0[575:512] : 64'h0) | (_v0SelectBySew_T_72[1] ? regroupV0_1[575:512] : 64'h0) | (_v0SelectBySew_T_72[2] ? regroupV0_2[575:512] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_81 = 4'h1 << laneMaskSewSelect_9;
  wire [63:0]       v0SelectBySew_9 = (_v0SelectBySew_T_81[0] ? regroupV0_0[639:576] : 64'h0) | (_v0SelectBySew_T_81[1] ? regroupV0_1[639:576] : 64'h0) | (_v0SelectBySew_T_81[2] ? regroupV0_2[639:576] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_90 = 4'h1 << laneMaskSewSelect_10;
  wire [63:0]       v0SelectBySew_10 = (_v0SelectBySew_T_90[0] ? regroupV0_0[703:640] : 64'h0) | (_v0SelectBySew_T_90[1] ? regroupV0_1[703:640] : 64'h0) | (_v0SelectBySew_T_90[2] ? regroupV0_2[703:640] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_99 = 4'h1 << laneMaskSewSelect_11;
  wire [63:0]       v0SelectBySew_11 = (_v0SelectBySew_T_99[0] ? regroupV0_0[767:704] : 64'h0) | (_v0SelectBySew_T_99[1] ? regroupV0_1[767:704] : 64'h0) | (_v0SelectBySew_T_99[2] ? regroupV0_2[767:704] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_108 = 4'h1 << laneMaskSewSelect_12;
  wire [63:0]       v0SelectBySew_12 = (_v0SelectBySew_T_108[0] ? regroupV0_0[831:768] : 64'h0) | (_v0SelectBySew_T_108[1] ? regroupV0_1[831:768] : 64'h0) | (_v0SelectBySew_T_108[2] ? regroupV0_2[831:768] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_117 = 4'h1 << laneMaskSewSelect_13;
  wire [63:0]       v0SelectBySew_13 = (_v0SelectBySew_T_117[0] ? regroupV0_0[895:832] : 64'h0) | (_v0SelectBySew_T_117[1] ? regroupV0_1[895:832] : 64'h0) | (_v0SelectBySew_T_117[2] ? regroupV0_2[895:832] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_126 = 4'h1 << laneMaskSewSelect_14;
  wire [63:0]       v0SelectBySew_14 = (_v0SelectBySew_T_126[0] ? regroupV0_0[959:896] : 64'h0) | (_v0SelectBySew_T_126[1] ? regroupV0_1[959:896] : 64'h0) | (_v0SelectBySew_T_126[2] ? regroupV0_2[959:896] : 64'h0);
  wire [3:0]        _v0SelectBySew_T_135 = 4'h1 << laneMaskSewSelect_15;
  wire [63:0]       v0SelectBySew_15 = (_v0SelectBySew_T_135[0] ? regroupV0_0[1023:960] : 64'h0) | (_v0SelectBySew_T_135[1] ? regroupV0_1[1023:960] : 64'h0) | (_v0SelectBySew_T_135[2] ? regroupV0_2[1023:960] : 64'h0);
  wire [3:0]        intLMULInput = 4'h1 << instReq_bits_vlmul[1:0];
  wire [12:0]       _dataPosition_T_1 = {3'h0, instReq_bits_readFromScala[9:0]} << instReq_bits_sew;
  wire [9:0]        dataPosition = _dataPosition_T_1[9:0];
  wire [3:0]        _sewOHInput_T = 4'h1 << instReq_bits_sew;
  wire [2:0]        sewOHInput = _sewOHInput_T[2:0];
  wire [1:0]        dataOffset = {dataPosition[1] & (|(sewOHInput[1:0])), dataPosition[0] & sewOHInput[0]};
  wire [3:0]        accessLane = dataPosition[5:2];
  wire [3:0]        dataGroup = dataPosition[9:6];
  wire              offset = dataGroup[0];
  wire [2:0]        accessRegGrowth = dataGroup[3:1];
  wire [2:0]        reallyGrowth = accessRegGrowth;
  wire [4:0]        decimalProportion = {offset, accessLane};
  wire [2:0]        decimal = decimalProportion[4:2];
  wire              notNeedRead = |{instReq_bits_vlmul[2] & decimal >= intLMULInput[3:1] | ~(instReq_bits_vlmul[2]) & {1'h0, accessRegGrowth} >= intLMULInput, instReq_bits_readFromScala[31:10]};
  reg  [1:0]        gatherReadState;
  wire              gatherSRead = gatherReadState == 2'h1;
  wire              gatherWaiteRead = gatherReadState == 2'h2;
  assign gatherResponse = &gatherReadState;
  wire              gatherData_valid_0 = gatherResponse;
  reg  [1:0]        gatherDatOffset;
  reg  [3:0]        gatherLane;
  reg               gatherOffset;
  reg  [2:0]        gatherGrowth;
  reg  [2:0]        instReg_instructionIndex;
  wire [2:0]        exeResp_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_4_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_5_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_6_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_7_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_8_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_9_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_10_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_11_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_12_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_13_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_14_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        exeResp_15_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_4_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_5_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_6_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_7_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_8_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_9_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_10_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_11_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_12_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_13_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_14_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        readChannel_15_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]        writeRequest_0_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_1_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_2_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_3_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_4_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_5_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_6_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_7_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_8_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_9_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_10_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_11_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_12_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_13_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_14_index = instReg_instructionIndex;
  wire [2:0]        writeRequest_15_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_0_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_1_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_2_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_3_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_4_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_5_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_6_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_7_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_8_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_9_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_10_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_11_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_12_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_13_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_14_enq_bits_index = instReg_instructionIndex;
  wire [2:0]        writeQueue_15_enq_bits_index = instReg_instructionIndex;
  reg               instReg_decodeResult_orderReduce;
  reg               instReg_decodeResult_floatMul;
  reg  [1:0]        instReg_decodeResult_fpExecutionType;
  reg               instReg_decodeResult_float;
  reg               instReg_decodeResult_specialSlot;
  reg  [4:0]        instReg_decodeResult_topUop;
  reg               instReg_decodeResult_popCount;
  reg               instReg_decodeResult_ffo;
  reg               instReg_decodeResult_average;
  reg               instReg_decodeResult_reverse;
  reg               instReg_decodeResult_dontNeedExecuteInLane;
  reg               instReg_decodeResult_scheduler;
  reg               instReg_decodeResult_sReadVD;
  reg               instReg_decodeResult_vtype;
  reg               instReg_decodeResult_sWrite;
  reg               instReg_decodeResult_crossRead;
  reg               instReg_decodeResult_crossWrite;
  reg               instReg_decodeResult_maskUnit;
  reg               instReg_decodeResult_special;
  reg               instReg_decodeResult_saturate;
  reg               instReg_decodeResult_vwmacc;
  reg               instReg_decodeResult_readOnly;
  reg               instReg_decodeResult_maskSource;
  reg               instReg_decodeResult_maskDestination;
  reg               instReg_decodeResult_maskLogic;
  reg  [3:0]        instReg_decodeResult_uop;
  reg               instReg_decodeResult_iota;
  reg               instReg_decodeResult_mv;
  reg               instReg_decodeResult_extend;
  reg               instReg_decodeResult_unOrderWrite;
  reg               instReg_decodeResult_compress;
  reg               instReg_decodeResult_gather16;
  reg               instReg_decodeResult_gather;
  reg               instReg_decodeResult_slid;
  reg               instReg_decodeResult_targetRd;
  reg               instReg_decodeResult_widenReduce;
  reg               instReg_decodeResult_red;
  reg               instReg_decodeResult_nr;
  reg               instReg_decodeResult_itype;
  reg               instReg_decodeResult_unsigned1;
  reg               instReg_decodeResult_unsigned0;
  reg               instReg_decodeResult_other;
  reg               instReg_decodeResult_multiCycle;
  reg               instReg_decodeResult_divider;
  reg               instReg_decodeResult_multiplier;
  reg               instReg_decodeResult_shift;
  reg               instReg_decodeResult_adder;
  reg               instReg_decodeResult_logic;
  reg  [31:0]       instReg_readFromScala;
  reg  [1:0]        instReg_sew;
  reg  [2:0]        instReg_vlmul;
  reg               instReg_maskType;
  reg  [2:0]        instReg_vxrm;
  reg  [4:0]        instReg_vs2;
  reg  [4:0]        instReg_vs1;
  reg  [4:0]        instReg_vd;
  wire [4:0]        writeRequest_0_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_1_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_2_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_3_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_4_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_5_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_6_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_7_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_8_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_9_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_10_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_11_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_12_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_13_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_14_writeData_vd = instReg_vd;
  wire [4:0]        writeRequest_15_writeData_vd = instReg_vd;
  reg  [10:0]       instReg_vl;
  wire [10:0]       reduceLastDataNeed_byteForVl = instReg_vl;
  wire              enqMvRD = instReq_bits_decodeResult_topUop == 5'hB;
  reg               instVlValid;
  wire              gatherRequestFire = gatherReadState == 2'h0 & gatherRead & ~instVlValid;
  wire              viotaReq = instReq_bits_decodeResult_topUop == 5'h8;
  reg               readVS1Reg_dataValid;
  reg               readVS1Reg_requestSend;
  reg               readVS1Reg_sendToExecution;
  reg  [31:0]       readVS1Reg_data;
  reg  [3:0]        readVS1Reg_readIndex;
  wire [3:0]        _sew1H_T = 4'h1 << instReg_sew;
  wire [2:0]        sew1H = _sew1H_T[2:0];
  wire [3:0]        unitType = 4'h1 << instReg_decodeResult_topUop[4:3];
  wire [3:0]        subType = 4'h1 << instReg_decodeResult_topUop[2:1];
  wire              readType = unitType[0];
  wire              gather16 = instReg_decodeResult_topUop == 5'h5;
  wire              maskDestinationType = instReg_decodeResult_topUop == 5'h18;
  wire              compress = instReg_decodeResult_topUop[4:1] == 4'h4;
  wire              viota = instReg_decodeResult_topUop == 5'h8;
  wire              mv = instReg_decodeResult_topUop[4:1] == 4'h5;
  wire              mvRd = instReg_decodeResult_topUop == 5'hB;
  wire              mvVd = instReg_decodeResult_topUop == 5'hA;
  wire              orderReduce = {instReg_decodeResult_topUop[4:2], instReg_decodeResult_topUop[0]} == 4'hB;
  wire              ffo = instReg_decodeResult_topUop[4:1] == 4'h7;
  wire              extendType = unitType[3] & (subType[2] | subType[1]);
  wire              readValid = readType & instVlValid;
  wire              noSource = mv | viota;
  wire              allGroupExecute = maskDestinationType | unitType[2] | compress | ffo;
  wire              useDefaultSew = readType & ~gather16;
  wire [1:0]        _dataSplitSew_T_11 = useDefaultSew ? instReg_sew : 2'h0;
  wire [1:0]        dataSplitSew = {_dataSplitSew_T_11[1], _dataSplitSew_T_11[0] | unitType[3] & subType[1] | gather16} | {allGroupExecute, 1'h0};
  wire              sourceDataUseDefaultSew = ~(unitType[3] | gather16);
  wire [1:0]        _sourceDataEEW_T_6 = (sourceDataUseDefaultSew ? instReg_sew : 2'h0) | (unitType[3] ? instReg_sew >> subType[2:1] : 2'h0);
  wire [1:0]        sourceDataEEW = {_sourceDataEEW_T_6[1], _sourceDataEEW_T_6[0] | gather16};
  wire [3:0]        executeIndexGrowth = 4'h1 << dataSplitSew;
  wire [1:0]        lastExecuteIndex = {2{executeIndexGrowth[0]}} | {executeIndexGrowth[1], 1'h0};
  wire [3:0]        _sourceDataEEW1H_T = 4'h1 << sourceDataEEW;
  wire [2:0]        sourceDataEEW1H = _sourceDataEEW1H_T[2:0];
  wire [9:0]        lastElementIndex = instReg_vl[9:0] - {9'h0, |instReg_vl};
  wire [9:0]        processingVl_lastByteIndex = lastElementIndex;
  wire              maskFormatSource = ffo | maskDestinationType;
  wire [5:0]        processingVl_lastGroupRemaining = processingVl_lastByteIndex[5:0];
  wire [3:0]        processingVl_0_1 = processingVl_lastByteIndex[9:6];
  wire [3:0]        processingVl_lastLaneIndex = processingVl_lastGroupRemaining[5:2];
  wire [15:0]       _processingVl_lastGroupDataNeed_T = 16'h1 << processingVl_lastLaneIndex;
  wire [14:0]       _GEN_15 = _processingVl_lastGroupDataNeed_T[14:0] | _processingVl_lastGroupDataNeed_T[15:1];
  wire [13:0]       _GEN_16 = _GEN_15[13:0] | {_processingVl_lastGroupDataNeed_T[15], _GEN_15[14:2]};
  wire [11:0]       _GEN_17 = _GEN_16[11:0] | {_processingVl_lastGroupDataNeed_T[15], _GEN_15[14], _GEN_16[13:4]};
  wire [15:0]       processingVl_0_2 = {_processingVl_lastGroupDataNeed_T[15], _GEN_15[14], _GEN_16[13:12], _GEN_17[11:8], _GEN_17[7:0] | {_processingVl_lastGroupDataNeed_T[15], _GEN_15[14], _GEN_16[13:12], _GEN_17[11:8]}};
  wire [10:0]       processingVl_lastByteIndex_1 = {lastElementIndex, 1'h0};
  wire [5:0]        processingVl_lastGroupRemaining_1 = processingVl_lastByteIndex_1[5:0];
  wire [4:0]        processingVl_1_1 = processingVl_lastByteIndex_1[10:6];
  wire [3:0]        processingVl_lastLaneIndex_1 = processingVl_lastGroupRemaining_1[5:2];
  wire [15:0]       _processingVl_lastGroupDataNeed_T_9 = 16'h1 << processingVl_lastLaneIndex_1;
  wire [14:0]       _GEN_18 = _processingVl_lastGroupDataNeed_T_9[14:0] | _processingVl_lastGroupDataNeed_T_9[15:1];
  wire [13:0]       _GEN_19 = _GEN_18[13:0] | {_processingVl_lastGroupDataNeed_T_9[15], _GEN_18[14:2]};
  wire [11:0]       _GEN_20 = _GEN_19[11:0] | {_processingVl_lastGroupDataNeed_T_9[15], _GEN_18[14], _GEN_19[13:4]};
  wire [15:0]       processingVl_1_2 = {_processingVl_lastGroupDataNeed_T_9[15], _GEN_18[14], _GEN_19[13:12], _GEN_20[11:8], _GEN_20[7:0] | {_processingVl_lastGroupDataNeed_T_9[15], _GEN_18[14], _GEN_19[13:12], _GEN_20[11:8]}};
  wire [11:0]       processingVl_lastByteIndex_2 = {lastElementIndex, 2'h0};
  wire [5:0]        processingVl_lastGroupRemaining_2 = processingVl_lastByteIndex_2[5:0];
  wire [5:0]        processingVl_2_1 = processingVl_lastByteIndex_2[11:6];
  wire [3:0]        processingVl_lastLaneIndex_2 = processingVl_lastGroupRemaining_2[5:2];
  wire [15:0]       _processingVl_lastGroupDataNeed_T_18 = 16'h1 << processingVl_lastLaneIndex_2;
  wire [14:0]       _GEN_21 = _processingVl_lastGroupDataNeed_T_18[14:0] | _processingVl_lastGroupDataNeed_T_18[15:1];
  wire [13:0]       _GEN_22 = _GEN_21[13:0] | {_processingVl_lastGroupDataNeed_T_18[15], _GEN_21[14:2]};
  wire [11:0]       _GEN_23 = _GEN_22[11:0] | {_processingVl_lastGroupDataNeed_T_18[15], _GEN_21[14], _GEN_22[13:4]};
  wire [15:0]       processingVl_2_2 = {_processingVl_lastGroupDataNeed_T_18[15], _GEN_21[14], _GEN_22[13:12], _GEN_23[11:8], _GEN_23[7:0] | {_processingVl_lastGroupDataNeed_T_18[15], _GEN_21[14], _GEN_22[13:12], _GEN_23[11:8]}};
  wire [8:0]        processingMaskVl_lastGroupRemaining = lastElementIndex[8:0];
  wire [8:0]        elementTailForMaskDestination = lastElementIndex[8:0];
  wire              processingMaskVl_lastGroupMisAlign = |processingMaskVl_lastGroupRemaining;
  wire              processingMaskVl_0_1 = lastElementIndex[9];
  wire [3:0]        processingMaskVl_lastLaneIndex = processingMaskVl_lastGroupRemaining[8:5] - {3'h0, processingMaskVl_lastGroupRemaining[4:0] == 5'h0};
  wire [15:0]       _processingMaskVl_dataNeedForPL_T = 16'h1 << processingMaskVl_lastLaneIndex;
  wire [14:0]       _GEN_24 = _processingMaskVl_dataNeedForPL_T[14:0] | _processingMaskVl_dataNeedForPL_T[15:1];
  wire [13:0]       _GEN_25 = _GEN_24[13:0] | {_processingMaskVl_dataNeedForPL_T[15], _GEN_24[14:2]};
  wire [11:0]       _GEN_26 = _GEN_25[11:0] | {_processingMaskVl_dataNeedForPL_T[15], _GEN_24[14], _GEN_25[13:4]};
  wire [15:0]       processingMaskVl_dataNeedForPL = {_processingMaskVl_dataNeedForPL_T[15], _GEN_24[14], _GEN_25[13:12], _GEN_26[11:8], _GEN_26[7:0] | {_processingMaskVl_dataNeedForPL_T[15], _GEN_24[14], _GEN_25[13:12], _GEN_26[11:8]}};
  wire              processingMaskVl_dataNeedForNPL_misAlign = |(processingMaskVl_lastGroupRemaining[1:0]);
  wire [7:0]        processingMaskVl_dataNeedForNPL_datapathSize = {1'h0, processingMaskVl_lastGroupRemaining[8:2]} + {7'h0, processingMaskVl_dataNeedForNPL_misAlign};
  wire              processingMaskVl_dataNeedForNPL_allNeed = |(processingMaskVl_dataNeedForNPL_datapathSize[7:4]);
  wire [3:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex = processingMaskVl_dataNeedForNPL_datapathSize[3:0];
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T = 16'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex;
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_3 = _processingMaskVl_dataNeedForNPL_dataNeed_T | {_processingMaskVl_dataNeedForNPL_dataNeed_T[14:0], 1'h0};
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_6 = _processingMaskVl_dataNeedForNPL_dataNeed_T_3 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_3[13:0], 2'h0};
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_9 = _processingMaskVl_dataNeedForNPL_dataNeed_T_6 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_6[11:0], 4'h0};
  wire [15:0]       processingMaskVl_dataNeedForNPL_dataNeed = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_9 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_9[7:0], 8'h0}) | {16{processingMaskVl_dataNeedForNPL_allNeed}};
  wire              processingMaskVl_dataNeedForNPL_misAlign_1 = processingMaskVl_lastGroupRemaining[0];
  wire [8:0]        processingMaskVl_dataNeedForNPL_datapathSize_1 = {1'h0, processingMaskVl_lastGroupRemaining[8:1]} + {8'h0, processingMaskVl_dataNeedForNPL_misAlign_1};
  wire              processingMaskVl_dataNeedForNPL_allNeed_1 = |(processingMaskVl_dataNeedForNPL_datapathSize_1[8:4]);
  wire [3:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex_1 = processingMaskVl_dataNeedForNPL_datapathSize_1[3:0];
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_16 = 16'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_1;
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_19 = _processingMaskVl_dataNeedForNPL_dataNeed_T_16 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_16[14:0], 1'h0};
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_22 = _processingMaskVl_dataNeedForNPL_dataNeed_T_19 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_19[13:0], 2'h0};
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_25 = _processingMaskVl_dataNeedForNPL_dataNeed_T_22 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_22[11:0], 4'h0};
  wire [15:0]       processingMaskVl_dataNeedForNPL_dataNeed_1 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_25 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_25[7:0], 8'h0}) | {16{processingMaskVl_dataNeedForNPL_allNeed_1}};
  wire [9:0]        processingMaskVl_dataNeedForNPL_datapathSize_2 = {1'h0, processingMaskVl_lastGroupRemaining};
  wire              processingMaskVl_dataNeedForNPL_allNeed_2 = |(processingMaskVl_dataNeedForNPL_datapathSize_2[9:4]);
  wire [3:0]        processingMaskVl_dataNeedForNPL_lastLaneIndex_2 = processingMaskVl_dataNeedForNPL_datapathSize_2[3:0];
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_32 = 16'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_2;
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_35 = _processingMaskVl_dataNeedForNPL_dataNeed_T_32 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_32[14:0], 1'h0};
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_38 = _processingMaskVl_dataNeedForNPL_dataNeed_T_35 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_35[13:0], 2'h0};
  wire [15:0]       _processingMaskVl_dataNeedForNPL_dataNeed_T_41 = _processingMaskVl_dataNeedForNPL_dataNeed_T_38 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_38[11:0], 4'h0};
  wire [15:0]       processingMaskVl_dataNeedForNPL_dataNeed_2 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_41 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_41[7:0], 8'h0}) | {16{processingMaskVl_dataNeedForNPL_allNeed_2}};
  wire [15:0]       processingMaskVl_dataNeedForNPL =
    (sew1H[0] ? processingMaskVl_dataNeedForNPL_dataNeed : 16'h0) | (sew1H[1] ? processingMaskVl_dataNeedForNPL_dataNeed_1 : 16'h0) | (sew1H[2] ? processingMaskVl_dataNeedForNPL_dataNeed_2 : 16'h0);
  wire [15:0]       processingMaskVl_0_2 = ffo ? processingMaskVl_dataNeedForPL : processingMaskVl_dataNeedForNPL;
  wire              reduceLastDataNeed_vlMSB = |(reduceLastDataNeed_byteForVl[10:6]);
  wire [5:0]        reduceLastDataNeed_vlLSB = instReg_vl[5:0];
  wire [5:0]        reduceLastDataNeed_vlLSB_1 = instReg_vl[5:0];
  wire [5:0]        reduceLastDataNeed_vlLSB_2 = instReg_vl[5:0];
  wire [3:0]        reduceLastDataNeed_lsbDSize = reduceLastDataNeed_vlLSB[5:2] - {3'h0, reduceLastDataNeed_vlLSB[1:0] == 2'h0};
  wire [15:0]       _reduceLastDataNeed_T = 16'h1 << reduceLastDataNeed_lsbDSize;
  wire [14:0]       _GEN_27 = _reduceLastDataNeed_T[14:0] | _reduceLastDataNeed_T[15:1];
  wire [13:0]       _GEN_28 = _GEN_27[13:0] | {_reduceLastDataNeed_T[15], _GEN_27[14:2]};
  wire [11:0]       _GEN_29 = _GEN_28[11:0] | {_reduceLastDataNeed_T[15], _GEN_27[14], _GEN_28[13:4]};
  wire [11:0]       reduceLastDataNeed_byteForVl_1 = {instReg_vl, 1'h0};
  wire              reduceLastDataNeed_vlMSB_1 = |(reduceLastDataNeed_byteForVl_1[11:6]);
  wire [3:0]        reduceLastDataNeed_lsbDSize_1 = reduceLastDataNeed_vlLSB_1[5:2] - {3'h0, reduceLastDataNeed_vlLSB_1[1:0] == 2'h0};
  wire [15:0]       _reduceLastDataNeed_T_12 = 16'h1 << reduceLastDataNeed_lsbDSize_1;
  wire [14:0]       _GEN_30 = _reduceLastDataNeed_T_12[14:0] | _reduceLastDataNeed_T_12[15:1];
  wire [13:0]       _GEN_31 = _GEN_30[13:0] | {_reduceLastDataNeed_T_12[15], _GEN_30[14:2]};
  wire [11:0]       _GEN_32 = _GEN_31[11:0] | {_reduceLastDataNeed_T_12[15], _GEN_30[14], _GEN_31[13:4]};
  wire [12:0]       reduceLastDataNeed_byteForVl_2 = {instReg_vl, 2'h0};
  wire              reduceLastDataNeed_vlMSB_2 = |(reduceLastDataNeed_byteForVl_2[12:6]);
  wire [3:0]        reduceLastDataNeed_lsbDSize_2 = reduceLastDataNeed_vlLSB_2[5:2] - {3'h0, reduceLastDataNeed_vlLSB_2[1:0] == 2'h0};
  wire [15:0]       _reduceLastDataNeed_T_24 = 16'h1 << reduceLastDataNeed_lsbDSize_2;
  wire [14:0]       _GEN_33 = _reduceLastDataNeed_T_24[14:0] | _reduceLastDataNeed_T_24[15:1];
  wire [13:0]       _GEN_34 = _GEN_33[13:0] | {_reduceLastDataNeed_T_24[15], _GEN_33[14:2]};
  wire [11:0]       _GEN_35 = _GEN_34[11:0] | {_reduceLastDataNeed_T_24[15], _GEN_33[14], _GEN_34[13:4]};
  wire [15:0]       reduceLastDataNeed =
    (sew1H[0] ? {_reduceLastDataNeed_T[15], _GEN_27[14], _GEN_28[13:12], _GEN_29[11:8], _GEN_29[7:0] | {_reduceLastDataNeed_T[15], _GEN_27[14], _GEN_28[13:12], _GEN_29[11:8]}} | {16{reduceLastDataNeed_vlMSB}} : 16'h0)
    | (sew1H[1] ? {_reduceLastDataNeed_T_12[15], _GEN_30[14], _GEN_31[13:12], _GEN_32[11:8], _GEN_32[7:0] | {_reduceLastDataNeed_T_12[15], _GEN_30[14], _GEN_31[13:12], _GEN_32[11:8]}} | {16{reduceLastDataNeed_vlMSB_1}} : 16'h0)
    | (sew1H[2] ? {_reduceLastDataNeed_T_24[15], _GEN_33[14], _GEN_34[13:12], _GEN_35[11:8], _GEN_35[7:0] | {_reduceLastDataNeed_T_24[15], _GEN_33[14], _GEN_34[13:12], _GEN_35[11:8]}} | {16{reduceLastDataNeed_vlMSB_2}} : 16'h0);
  wire [1:0]        dataSourceSew = unitType[3] ? instReg_sew - instReg_decodeResult_topUop[2:1] : gather16 ? 2'h1 : instReg_sew;
  wire [3:0]        _dataSourceSew1H_T = 4'h1 << dataSourceSew;
  wire [2:0]        dataSourceSew1H = _dataSourceSew1H_T[2:0];
  wire              unorderReduce = ~orderReduce & unitType[2];
  wire              normalFormat = ~maskFormatSource & ~unorderReduce & ~mv;
  wire [5:0]        lastGroupForInstruction =
    {1'h0, {1'h0, {3'h0, maskFormatSource & processingMaskVl_0_1} | (normalFormat & dataSourceSew1H[0] ? processingVl_0_1 : 4'h0)} | (normalFormat & dataSourceSew1H[1] ? processingVl_1_1 : 5'h0)}
    | (normalFormat & dataSourceSew1H[2] ? processingVl_2_1 : 6'h0);
  wire [4:0]        popDataNeed_dataPathGroups = lastElementIndex[9:5];
  wire [3:0]        popDataNeed_lastLaneIndex = popDataNeed_dataPathGroups[3:0];
  wire              popDataNeed_lagerThanDLen = popDataNeed_dataPathGroups[4];
  wire [15:0]       _popDataNeed_T = 16'h1 << popDataNeed_lastLaneIndex;
  wire [14:0]       _GEN_36 = _popDataNeed_T[14:0] | _popDataNeed_T[15:1];
  wire [13:0]       _GEN_37 = _GEN_36[13:0] | {_popDataNeed_T[15], _GEN_36[14:2]};
  wire [11:0]       _GEN_38 = _GEN_37[11:0] | {_popDataNeed_T[15], _GEN_36[14], _GEN_37[13:4]};
  wire [15:0]       popDataNeed = {_popDataNeed_T[15], _GEN_36[14], _GEN_37[13:12], _GEN_38[11:8], _GEN_38[7:0] | {_popDataNeed_T[15], _GEN_36[14], _GEN_37[13:12], _GEN_38[11:8]}} | {16{popDataNeed_lagerThanDLen}};
  wire [15:0]       lastGroupDataNeed =
    (unorderReduce & instReg_decodeResult_popCount ? popDataNeed : 16'h0) | (unorderReduce & ~instReg_decodeResult_popCount ? reduceLastDataNeed : 16'h0) | (maskFormatSource ? processingMaskVl_0_2 : 16'h0)
    | (normalFormat & dataSourceSew1H[0] ? processingVl_0_2 : 16'h0) | (normalFormat & dataSourceSew1H[1] ? processingVl_1_2 : 16'h0) | (normalFormat & dataSourceSew1H[2] ? processingVl_2_2 : 16'h0);
  wire [1:0]        exeRequestQueue_queue_dataIn_lo = {exeRequestQueue_0_enq_bits_ffo, exeRequestQueue_0_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi = {exeRequestQueue_0_enq_bits_source1, exeRequestQueue_0_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi = {exeRequestQueue_queue_dataIn_hi_hi, exeRequestQueue_0_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn = {exeRequestQueue_queue_dataIn_hi, exeRequestQueue_queue_dataIn_lo};
  wire              exeRequestQueue_queue_dataOut_fpReduceValid = _exeRequestQueue_queue_fifo_data_out[0];
  wire              exeRequestQueue_queue_dataOut_ffo = _exeRequestQueue_queue_fifo_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_index = _exeRequestQueue_queue_fifo_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_source2 = _exeRequestQueue_queue_fifo_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_source1 = _exeRequestQueue_queue_fifo_data_out[68:37];
  wire              exeRequestQueue_0_enq_ready = ~_exeRequestQueue_queue_fifo_full;
  wire              exeRequestQueue_0_deq_ready;
  wire              exeRequestQueue_0_deq_valid = ~_exeRequestQueue_queue_fifo_empty | exeRequestQueue_0_enq_valid;
  wire [31:0]       exeRequestQueue_0_deq_bits_source1 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source1 : exeRequestQueue_queue_dataOut_source1;
  wire [31:0]       exeRequestQueue_0_deq_bits_source2 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source2 : exeRequestQueue_queue_dataOut_source2;
  wire [2:0]        exeRequestQueue_0_deq_bits_index = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_index : exeRequestQueue_queue_dataOut_index;
  wire              exeRequestQueue_0_deq_bits_ffo = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_ffo : exeRequestQueue_queue_dataOut_ffo;
  wire              exeRequestQueue_0_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_fpReduceValid;
  wire              tokenIO_0_maskRequestRelease_0 = exeRequestQueue_0_deq_ready & exeRequestQueue_0_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_1 = {exeRequestQueue_1_enq_bits_ffo, exeRequestQueue_1_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_1 = {exeRequestQueue_1_enq_bits_source1, exeRequestQueue_1_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_1 = {exeRequestQueue_queue_dataIn_hi_hi_1, exeRequestQueue_1_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_1 = {exeRequestQueue_queue_dataIn_hi_1, exeRequestQueue_queue_dataIn_lo_1};
  wire              exeRequestQueue_queue_dataOut_1_fpReduceValid = _exeRequestQueue_queue_fifo_1_data_out[0];
  wire              exeRequestQueue_queue_dataOut_1_ffo = _exeRequestQueue_queue_fifo_1_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_1_index = _exeRequestQueue_queue_fifo_1_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_1_source2 = _exeRequestQueue_queue_fifo_1_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_1_source1 = _exeRequestQueue_queue_fifo_1_data_out[68:37];
  wire              exeRequestQueue_1_enq_ready = ~_exeRequestQueue_queue_fifo_1_full;
  wire              exeRequestQueue_1_deq_ready;
  wire              exeRequestQueue_1_deq_valid = ~_exeRequestQueue_queue_fifo_1_empty | exeRequestQueue_1_enq_valid;
  wire [31:0]       exeRequestQueue_1_deq_bits_source1 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source1 : exeRequestQueue_queue_dataOut_1_source1;
  wire [31:0]       exeRequestQueue_1_deq_bits_source2 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source2 : exeRequestQueue_queue_dataOut_1_source2;
  wire [2:0]        exeRequestQueue_1_deq_bits_index = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_index : exeRequestQueue_queue_dataOut_1_index;
  wire              exeRequestQueue_1_deq_bits_ffo = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_ffo : exeRequestQueue_queue_dataOut_1_ffo;
  wire              exeRequestQueue_1_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_1_fpReduceValid;
  wire              tokenIO_1_maskRequestRelease_0 = exeRequestQueue_1_deq_ready & exeRequestQueue_1_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_2 = {exeRequestQueue_2_enq_bits_ffo, exeRequestQueue_2_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_2 = {exeRequestQueue_2_enq_bits_source1, exeRequestQueue_2_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_2 = {exeRequestQueue_queue_dataIn_hi_hi_2, exeRequestQueue_2_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_2 = {exeRequestQueue_queue_dataIn_hi_2, exeRequestQueue_queue_dataIn_lo_2};
  wire              exeRequestQueue_queue_dataOut_2_fpReduceValid = _exeRequestQueue_queue_fifo_2_data_out[0];
  wire              exeRequestQueue_queue_dataOut_2_ffo = _exeRequestQueue_queue_fifo_2_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_2_index = _exeRequestQueue_queue_fifo_2_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_2_source2 = _exeRequestQueue_queue_fifo_2_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_2_source1 = _exeRequestQueue_queue_fifo_2_data_out[68:37];
  wire              exeRequestQueue_2_enq_ready = ~_exeRequestQueue_queue_fifo_2_full;
  wire              exeRequestQueue_2_deq_ready;
  wire              exeRequestQueue_2_deq_valid = ~_exeRequestQueue_queue_fifo_2_empty | exeRequestQueue_2_enq_valid;
  wire [31:0]       exeRequestQueue_2_deq_bits_source1 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source1 : exeRequestQueue_queue_dataOut_2_source1;
  wire [31:0]       exeRequestQueue_2_deq_bits_source2 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source2 : exeRequestQueue_queue_dataOut_2_source2;
  wire [2:0]        exeRequestQueue_2_deq_bits_index = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_index : exeRequestQueue_queue_dataOut_2_index;
  wire              exeRequestQueue_2_deq_bits_ffo = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_ffo : exeRequestQueue_queue_dataOut_2_ffo;
  wire              exeRequestQueue_2_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_2_fpReduceValid;
  wire              tokenIO_2_maskRequestRelease_0 = exeRequestQueue_2_deq_ready & exeRequestQueue_2_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_3 = {exeRequestQueue_3_enq_bits_ffo, exeRequestQueue_3_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_3 = {exeRequestQueue_3_enq_bits_source1, exeRequestQueue_3_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_3 = {exeRequestQueue_queue_dataIn_hi_hi_3, exeRequestQueue_3_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_3 = {exeRequestQueue_queue_dataIn_hi_3, exeRequestQueue_queue_dataIn_lo_3};
  wire              exeRequestQueue_queue_dataOut_3_fpReduceValid = _exeRequestQueue_queue_fifo_3_data_out[0];
  wire              exeRequestQueue_queue_dataOut_3_ffo = _exeRequestQueue_queue_fifo_3_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_3_index = _exeRequestQueue_queue_fifo_3_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_3_source2 = _exeRequestQueue_queue_fifo_3_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_3_source1 = _exeRequestQueue_queue_fifo_3_data_out[68:37];
  wire              exeRequestQueue_3_enq_ready = ~_exeRequestQueue_queue_fifo_3_full;
  wire              exeRequestQueue_3_deq_ready;
  wire              exeRequestQueue_3_deq_valid = ~_exeRequestQueue_queue_fifo_3_empty | exeRequestQueue_3_enq_valid;
  wire [31:0]       exeRequestQueue_3_deq_bits_source1 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source1 : exeRequestQueue_queue_dataOut_3_source1;
  wire [31:0]       exeRequestQueue_3_deq_bits_source2 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source2 : exeRequestQueue_queue_dataOut_3_source2;
  wire [2:0]        exeRequestQueue_3_deq_bits_index = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_index : exeRequestQueue_queue_dataOut_3_index;
  wire              exeRequestQueue_3_deq_bits_ffo = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_ffo : exeRequestQueue_queue_dataOut_3_ffo;
  wire              exeRequestQueue_3_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_3_fpReduceValid;
  wire              tokenIO_3_maskRequestRelease_0 = exeRequestQueue_3_deq_ready & exeRequestQueue_3_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_4 = {exeRequestQueue_4_enq_bits_ffo, exeRequestQueue_4_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_4 = {exeRequestQueue_4_enq_bits_source1, exeRequestQueue_4_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_4 = {exeRequestQueue_queue_dataIn_hi_hi_4, exeRequestQueue_4_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_4 = {exeRequestQueue_queue_dataIn_hi_4, exeRequestQueue_queue_dataIn_lo_4};
  wire              exeRequestQueue_queue_dataOut_4_fpReduceValid = _exeRequestQueue_queue_fifo_4_data_out[0];
  wire              exeRequestQueue_queue_dataOut_4_ffo = _exeRequestQueue_queue_fifo_4_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_4_index = _exeRequestQueue_queue_fifo_4_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_4_source2 = _exeRequestQueue_queue_fifo_4_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_4_source1 = _exeRequestQueue_queue_fifo_4_data_out[68:37];
  wire              exeRequestQueue_4_enq_ready = ~_exeRequestQueue_queue_fifo_4_full;
  wire              exeRequestQueue_4_deq_ready;
  wire              exeRequestQueue_4_deq_valid = ~_exeRequestQueue_queue_fifo_4_empty | exeRequestQueue_4_enq_valid;
  wire [31:0]       exeRequestQueue_4_deq_bits_source1 = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_source1 : exeRequestQueue_queue_dataOut_4_source1;
  wire [31:0]       exeRequestQueue_4_deq_bits_source2 = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_source2 : exeRequestQueue_queue_dataOut_4_source2;
  wire [2:0]        exeRequestQueue_4_deq_bits_index = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_index : exeRequestQueue_queue_dataOut_4_index;
  wire              exeRequestQueue_4_deq_bits_ffo = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_ffo : exeRequestQueue_queue_dataOut_4_ffo;
  wire              exeRequestQueue_4_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_4_empty ? exeRequestQueue_4_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_4_fpReduceValid;
  wire              tokenIO_4_maskRequestRelease_0 = exeRequestQueue_4_deq_ready & exeRequestQueue_4_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_5 = {exeRequestQueue_5_enq_bits_ffo, exeRequestQueue_5_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_5 = {exeRequestQueue_5_enq_bits_source1, exeRequestQueue_5_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_5 = {exeRequestQueue_queue_dataIn_hi_hi_5, exeRequestQueue_5_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_5 = {exeRequestQueue_queue_dataIn_hi_5, exeRequestQueue_queue_dataIn_lo_5};
  wire              exeRequestQueue_queue_dataOut_5_fpReduceValid = _exeRequestQueue_queue_fifo_5_data_out[0];
  wire              exeRequestQueue_queue_dataOut_5_ffo = _exeRequestQueue_queue_fifo_5_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_5_index = _exeRequestQueue_queue_fifo_5_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_5_source2 = _exeRequestQueue_queue_fifo_5_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_5_source1 = _exeRequestQueue_queue_fifo_5_data_out[68:37];
  wire              exeRequestQueue_5_enq_ready = ~_exeRequestQueue_queue_fifo_5_full;
  wire              exeRequestQueue_5_deq_ready;
  wire              exeRequestQueue_5_deq_valid = ~_exeRequestQueue_queue_fifo_5_empty | exeRequestQueue_5_enq_valid;
  wire [31:0]       exeRequestQueue_5_deq_bits_source1 = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_source1 : exeRequestQueue_queue_dataOut_5_source1;
  wire [31:0]       exeRequestQueue_5_deq_bits_source2 = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_source2 : exeRequestQueue_queue_dataOut_5_source2;
  wire [2:0]        exeRequestQueue_5_deq_bits_index = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_index : exeRequestQueue_queue_dataOut_5_index;
  wire              exeRequestQueue_5_deq_bits_ffo = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_ffo : exeRequestQueue_queue_dataOut_5_ffo;
  wire              exeRequestQueue_5_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_5_empty ? exeRequestQueue_5_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_5_fpReduceValid;
  wire              tokenIO_5_maskRequestRelease_0 = exeRequestQueue_5_deq_ready & exeRequestQueue_5_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_6 = {exeRequestQueue_6_enq_bits_ffo, exeRequestQueue_6_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_6 = {exeRequestQueue_6_enq_bits_source1, exeRequestQueue_6_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_6 = {exeRequestQueue_queue_dataIn_hi_hi_6, exeRequestQueue_6_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_6 = {exeRequestQueue_queue_dataIn_hi_6, exeRequestQueue_queue_dataIn_lo_6};
  wire              exeRequestQueue_queue_dataOut_6_fpReduceValid = _exeRequestQueue_queue_fifo_6_data_out[0];
  wire              exeRequestQueue_queue_dataOut_6_ffo = _exeRequestQueue_queue_fifo_6_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_6_index = _exeRequestQueue_queue_fifo_6_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_6_source2 = _exeRequestQueue_queue_fifo_6_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_6_source1 = _exeRequestQueue_queue_fifo_6_data_out[68:37];
  wire              exeRequestQueue_6_enq_ready = ~_exeRequestQueue_queue_fifo_6_full;
  wire              exeRequestQueue_6_deq_ready;
  wire              exeRequestQueue_6_deq_valid = ~_exeRequestQueue_queue_fifo_6_empty | exeRequestQueue_6_enq_valid;
  wire [31:0]       exeRequestQueue_6_deq_bits_source1 = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_source1 : exeRequestQueue_queue_dataOut_6_source1;
  wire [31:0]       exeRequestQueue_6_deq_bits_source2 = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_source2 : exeRequestQueue_queue_dataOut_6_source2;
  wire [2:0]        exeRequestQueue_6_deq_bits_index = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_index : exeRequestQueue_queue_dataOut_6_index;
  wire              exeRequestQueue_6_deq_bits_ffo = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_ffo : exeRequestQueue_queue_dataOut_6_ffo;
  wire              exeRequestQueue_6_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_6_empty ? exeRequestQueue_6_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_6_fpReduceValid;
  wire              tokenIO_6_maskRequestRelease_0 = exeRequestQueue_6_deq_ready & exeRequestQueue_6_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_7 = {exeRequestQueue_7_enq_bits_ffo, exeRequestQueue_7_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_7 = {exeRequestQueue_7_enq_bits_source1, exeRequestQueue_7_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_7 = {exeRequestQueue_queue_dataIn_hi_hi_7, exeRequestQueue_7_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_7 = {exeRequestQueue_queue_dataIn_hi_7, exeRequestQueue_queue_dataIn_lo_7};
  wire              exeRequestQueue_queue_dataOut_7_fpReduceValid = _exeRequestQueue_queue_fifo_7_data_out[0];
  wire              exeRequestQueue_queue_dataOut_7_ffo = _exeRequestQueue_queue_fifo_7_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_7_index = _exeRequestQueue_queue_fifo_7_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_7_source2 = _exeRequestQueue_queue_fifo_7_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_7_source1 = _exeRequestQueue_queue_fifo_7_data_out[68:37];
  wire              exeRequestQueue_7_enq_ready = ~_exeRequestQueue_queue_fifo_7_full;
  wire              exeRequestQueue_7_deq_ready;
  wire              exeRequestQueue_7_deq_valid = ~_exeRequestQueue_queue_fifo_7_empty | exeRequestQueue_7_enq_valid;
  wire [31:0]       exeRequestQueue_7_deq_bits_source1 = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_source1 : exeRequestQueue_queue_dataOut_7_source1;
  wire [31:0]       exeRequestQueue_7_deq_bits_source2 = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_source2 : exeRequestQueue_queue_dataOut_7_source2;
  wire [2:0]        exeRequestQueue_7_deq_bits_index = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_index : exeRequestQueue_queue_dataOut_7_index;
  wire              exeRequestQueue_7_deq_bits_ffo = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_ffo : exeRequestQueue_queue_dataOut_7_ffo;
  wire              exeRequestQueue_7_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_7_empty ? exeRequestQueue_7_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_7_fpReduceValid;
  wire              tokenIO_7_maskRequestRelease_0 = exeRequestQueue_7_deq_ready & exeRequestQueue_7_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_8 = {exeRequestQueue_8_enq_bits_ffo, exeRequestQueue_8_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_8 = {exeRequestQueue_8_enq_bits_source1, exeRequestQueue_8_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_8 = {exeRequestQueue_queue_dataIn_hi_hi_8, exeRequestQueue_8_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_8 = {exeRequestQueue_queue_dataIn_hi_8, exeRequestQueue_queue_dataIn_lo_8};
  wire              exeRequestQueue_queue_dataOut_8_fpReduceValid = _exeRequestQueue_queue_fifo_8_data_out[0];
  wire              exeRequestQueue_queue_dataOut_8_ffo = _exeRequestQueue_queue_fifo_8_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_8_index = _exeRequestQueue_queue_fifo_8_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_8_source2 = _exeRequestQueue_queue_fifo_8_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_8_source1 = _exeRequestQueue_queue_fifo_8_data_out[68:37];
  wire              exeRequestQueue_8_enq_ready = ~_exeRequestQueue_queue_fifo_8_full;
  wire              exeRequestQueue_8_deq_ready;
  wire              exeRequestQueue_8_deq_valid = ~_exeRequestQueue_queue_fifo_8_empty | exeRequestQueue_8_enq_valid;
  wire [31:0]       exeRequestQueue_8_deq_bits_source1 = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_source1 : exeRequestQueue_queue_dataOut_8_source1;
  wire [31:0]       exeRequestQueue_8_deq_bits_source2 = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_source2 : exeRequestQueue_queue_dataOut_8_source2;
  wire [2:0]        exeRequestQueue_8_deq_bits_index = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_index : exeRequestQueue_queue_dataOut_8_index;
  wire              exeRequestQueue_8_deq_bits_ffo = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_ffo : exeRequestQueue_queue_dataOut_8_ffo;
  wire              exeRequestQueue_8_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_8_empty ? exeRequestQueue_8_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_8_fpReduceValid;
  wire              tokenIO_8_maskRequestRelease_0 = exeRequestQueue_8_deq_ready & exeRequestQueue_8_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_9 = {exeRequestQueue_9_enq_bits_ffo, exeRequestQueue_9_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_9 = {exeRequestQueue_9_enq_bits_source1, exeRequestQueue_9_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_9 = {exeRequestQueue_queue_dataIn_hi_hi_9, exeRequestQueue_9_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_9 = {exeRequestQueue_queue_dataIn_hi_9, exeRequestQueue_queue_dataIn_lo_9};
  wire              exeRequestQueue_queue_dataOut_9_fpReduceValid = _exeRequestQueue_queue_fifo_9_data_out[0];
  wire              exeRequestQueue_queue_dataOut_9_ffo = _exeRequestQueue_queue_fifo_9_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_9_index = _exeRequestQueue_queue_fifo_9_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_9_source2 = _exeRequestQueue_queue_fifo_9_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_9_source1 = _exeRequestQueue_queue_fifo_9_data_out[68:37];
  wire              exeRequestQueue_9_enq_ready = ~_exeRequestQueue_queue_fifo_9_full;
  wire              exeRequestQueue_9_deq_ready;
  wire              exeRequestQueue_9_deq_valid = ~_exeRequestQueue_queue_fifo_9_empty | exeRequestQueue_9_enq_valid;
  wire [31:0]       exeRequestQueue_9_deq_bits_source1 = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_source1 : exeRequestQueue_queue_dataOut_9_source1;
  wire [31:0]       exeRequestQueue_9_deq_bits_source2 = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_source2 : exeRequestQueue_queue_dataOut_9_source2;
  wire [2:0]        exeRequestQueue_9_deq_bits_index = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_index : exeRequestQueue_queue_dataOut_9_index;
  wire              exeRequestQueue_9_deq_bits_ffo = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_ffo : exeRequestQueue_queue_dataOut_9_ffo;
  wire              exeRequestQueue_9_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_9_empty ? exeRequestQueue_9_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_9_fpReduceValid;
  wire              tokenIO_9_maskRequestRelease_0 = exeRequestQueue_9_deq_ready & exeRequestQueue_9_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_10 = {exeRequestQueue_10_enq_bits_ffo, exeRequestQueue_10_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_10 = {exeRequestQueue_10_enq_bits_source1, exeRequestQueue_10_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_10 = {exeRequestQueue_queue_dataIn_hi_hi_10, exeRequestQueue_10_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_10 = {exeRequestQueue_queue_dataIn_hi_10, exeRequestQueue_queue_dataIn_lo_10};
  wire              exeRequestQueue_queue_dataOut_10_fpReduceValid = _exeRequestQueue_queue_fifo_10_data_out[0];
  wire              exeRequestQueue_queue_dataOut_10_ffo = _exeRequestQueue_queue_fifo_10_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_10_index = _exeRequestQueue_queue_fifo_10_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_10_source2 = _exeRequestQueue_queue_fifo_10_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_10_source1 = _exeRequestQueue_queue_fifo_10_data_out[68:37];
  wire              exeRequestQueue_10_enq_ready = ~_exeRequestQueue_queue_fifo_10_full;
  wire              exeRequestQueue_10_deq_ready;
  wire              exeRequestQueue_10_deq_valid = ~_exeRequestQueue_queue_fifo_10_empty | exeRequestQueue_10_enq_valid;
  wire [31:0]       exeRequestQueue_10_deq_bits_source1 = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_source1 : exeRequestQueue_queue_dataOut_10_source1;
  wire [31:0]       exeRequestQueue_10_deq_bits_source2 = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_source2 : exeRequestQueue_queue_dataOut_10_source2;
  wire [2:0]        exeRequestQueue_10_deq_bits_index = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_index : exeRequestQueue_queue_dataOut_10_index;
  wire              exeRequestQueue_10_deq_bits_ffo = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_ffo : exeRequestQueue_queue_dataOut_10_ffo;
  wire              exeRequestQueue_10_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_10_empty ? exeRequestQueue_10_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_10_fpReduceValid;
  wire              tokenIO_10_maskRequestRelease_0 = exeRequestQueue_10_deq_ready & exeRequestQueue_10_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_11 = {exeRequestQueue_11_enq_bits_ffo, exeRequestQueue_11_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_11 = {exeRequestQueue_11_enq_bits_source1, exeRequestQueue_11_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_11 = {exeRequestQueue_queue_dataIn_hi_hi_11, exeRequestQueue_11_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_11 = {exeRequestQueue_queue_dataIn_hi_11, exeRequestQueue_queue_dataIn_lo_11};
  wire              exeRequestQueue_queue_dataOut_11_fpReduceValid = _exeRequestQueue_queue_fifo_11_data_out[0];
  wire              exeRequestQueue_queue_dataOut_11_ffo = _exeRequestQueue_queue_fifo_11_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_11_index = _exeRequestQueue_queue_fifo_11_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_11_source2 = _exeRequestQueue_queue_fifo_11_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_11_source1 = _exeRequestQueue_queue_fifo_11_data_out[68:37];
  wire              exeRequestQueue_11_enq_ready = ~_exeRequestQueue_queue_fifo_11_full;
  wire              exeRequestQueue_11_deq_ready;
  wire              exeRequestQueue_11_deq_valid = ~_exeRequestQueue_queue_fifo_11_empty | exeRequestQueue_11_enq_valid;
  wire [31:0]       exeRequestQueue_11_deq_bits_source1 = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_source1 : exeRequestQueue_queue_dataOut_11_source1;
  wire [31:0]       exeRequestQueue_11_deq_bits_source2 = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_source2 : exeRequestQueue_queue_dataOut_11_source2;
  wire [2:0]        exeRequestQueue_11_deq_bits_index = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_index : exeRequestQueue_queue_dataOut_11_index;
  wire              exeRequestQueue_11_deq_bits_ffo = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_ffo : exeRequestQueue_queue_dataOut_11_ffo;
  wire              exeRequestQueue_11_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_11_empty ? exeRequestQueue_11_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_11_fpReduceValid;
  wire              tokenIO_11_maskRequestRelease_0 = exeRequestQueue_11_deq_ready & exeRequestQueue_11_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_12 = {exeRequestQueue_12_enq_bits_ffo, exeRequestQueue_12_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_12 = {exeRequestQueue_12_enq_bits_source1, exeRequestQueue_12_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_12 = {exeRequestQueue_queue_dataIn_hi_hi_12, exeRequestQueue_12_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_12 = {exeRequestQueue_queue_dataIn_hi_12, exeRequestQueue_queue_dataIn_lo_12};
  wire              exeRequestQueue_queue_dataOut_12_fpReduceValid = _exeRequestQueue_queue_fifo_12_data_out[0];
  wire              exeRequestQueue_queue_dataOut_12_ffo = _exeRequestQueue_queue_fifo_12_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_12_index = _exeRequestQueue_queue_fifo_12_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_12_source2 = _exeRequestQueue_queue_fifo_12_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_12_source1 = _exeRequestQueue_queue_fifo_12_data_out[68:37];
  wire              exeRequestQueue_12_enq_ready = ~_exeRequestQueue_queue_fifo_12_full;
  wire              exeRequestQueue_12_deq_ready;
  wire              exeRequestQueue_12_deq_valid = ~_exeRequestQueue_queue_fifo_12_empty | exeRequestQueue_12_enq_valid;
  wire [31:0]       exeRequestQueue_12_deq_bits_source1 = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_source1 : exeRequestQueue_queue_dataOut_12_source1;
  wire [31:0]       exeRequestQueue_12_deq_bits_source2 = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_source2 : exeRequestQueue_queue_dataOut_12_source2;
  wire [2:0]        exeRequestQueue_12_deq_bits_index = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_index : exeRequestQueue_queue_dataOut_12_index;
  wire              exeRequestQueue_12_deq_bits_ffo = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_ffo : exeRequestQueue_queue_dataOut_12_ffo;
  wire              exeRequestQueue_12_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_12_empty ? exeRequestQueue_12_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_12_fpReduceValid;
  wire              tokenIO_12_maskRequestRelease_0 = exeRequestQueue_12_deq_ready & exeRequestQueue_12_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_13 = {exeRequestQueue_13_enq_bits_ffo, exeRequestQueue_13_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_13 = {exeRequestQueue_13_enq_bits_source1, exeRequestQueue_13_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_13 = {exeRequestQueue_queue_dataIn_hi_hi_13, exeRequestQueue_13_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_13 = {exeRequestQueue_queue_dataIn_hi_13, exeRequestQueue_queue_dataIn_lo_13};
  wire              exeRequestQueue_queue_dataOut_13_fpReduceValid = _exeRequestQueue_queue_fifo_13_data_out[0];
  wire              exeRequestQueue_queue_dataOut_13_ffo = _exeRequestQueue_queue_fifo_13_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_13_index = _exeRequestQueue_queue_fifo_13_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_13_source2 = _exeRequestQueue_queue_fifo_13_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_13_source1 = _exeRequestQueue_queue_fifo_13_data_out[68:37];
  wire              exeRequestQueue_13_enq_ready = ~_exeRequestQueue_queue_fifo_13_full;
  wire              exeRequestQueue_13_deq_ready;
  wire              exeRequestQueue_13_deq_valid = ~_exeRequestQueue_queue_fifo_13_empty | exeRequestQueue_13_enq_valid;
  wire [31:0]       exeRequestQueue_13_deq_bits_source1 = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_source1 : exeRequestQueue_queue_dataOut_13_source1;
  wire [31:0]       exeRequestQueue_13_deq_bits_source2 = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_source2 : exeRequestQueue_queue_dataOut_13_source2;
  wire [2:0]        exeRequestQueue_13_deq_bits_index = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_index : exeRequestQueue_queue_dataOut_13_index;
  wire              exeRequestQueue_13_deq_bits_ffo = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_ffo : exeRequestQueue_queue_dataOut_13_ffo;
  wire              exeRequestQueue_13_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_13_empty ? exeRequestQueue_13_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_13_fpReduceValid;
  wire              tokenIO_13_maskRequestRelease_0 = exeRequestQueue_13_deq_ready & exeRequestQueue_13_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_14 = {exeRequestQueue_14_enq_bits_ffo, exeRequestQueue_14_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_14 = {exeRequestQueue_14_enq_bits_source1, exeRequestQueue_14_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_14 = {exeRequestQueue_queue_dataIn_hi_hi_14, exeRequestQueue_14_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_14 = {exeRequestQueue_queue_dataIn_hi_14, exeRequestQueue_queue_dataIn_lo_14};
  wire              exeRequestQueue_queue_dataOut_14_fpReduceValid = _exeRequestQueue_queue_fifo_14_data_out[0];
  wire              exeRequestQueue_queue_dataOut_14_ffo = _exeRequestQueue_queue_fifo_14_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_14_index = _exeRequestQueue_queue_fifo_14_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_14_source2 = _exeRequestQueue_queue_fifo_14_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_14_source1 = _exeRequestQueue_queue_fifo_14_data_out[68:37];
  wire              exeRequestQueue_14_enq_ready = ~_exeRequestQueue_queue_fifo_14_full;
  wire              exeRequestQueue_14_deq_ready;
  wire              exeRequestQueue_14_deq_valid = ~_exeRequestQueue_queue_fifo_14_empty | exeRequestQueue_14_enq_valid;
  wire [31:0]       exeRequestQueue_14_deq_bits_source1 = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_source1 : exeRequestQueue_queue_dataOut_14_source1;
  wire [31:0]       exeRequestQueue_14_deq_bits_source2 = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_source2 : exeRequestQueue_queue_dataOut_14_source2;
  wire [2:0]        exeRequestQueue_14_deq_bits_index = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_index : exeRequestQueue_queue_dataOut_14_index;
  wire              exeRequestQueue_14_deq_bits_ffo = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_ffo : exeRequestQueue_queue_dataOut_14_ffo;
  wire              exeRequestQueue_14_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_14_empty ? exeRequestQueue_14_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_14_fpReduceValid;
  wire              tokenIO_14_maskRequestRelease_0 = exeRequestQueue_14_deq_ready & exeRequestQueue_14_deq_valid;
  wire [1:0]        exeRequestQueue_queue_dataIn_lo_15 = {exeRequestQueue_15_enq_bits_ffo, exeRequestQueue_15_enq_bits_fpReduceValid};
  wire [63:0]       exeRequestQueue_queue_dataIn_hi_hi_15 = {exeRequestQueue_15_enq_bits_source1, exeRequestQueue_15_enq_bits_source2};
  wire [66:0]       exeRequestQueue_queue_dataIn_hi_15 = {exeRequestQueue_queue_dataIn_hi_hi_15, exeRequestQueue_15_enq_bits_index};
  wire [68:0]       exeRequestQueue_queue_dataIn_15 = {exeRequestQueue_queue_dataIn_hi_15, exeRequestQueue_queue_dataIn_lo_15};
  wire              exeRequestQueue_queue_dataOut_15_fpReduceValid = _exeRequestQueue_queue_fifo_15_data_out[0];
  wire              exeRequestQueue_queue_dataOut_15_ffo = _exeRequestQueue_queue_fifo_15_data_out[1];
  wire [2:0]        exeRequestQueue_queue_dataOut_15_index = _exeRequestQueue_queue_fifo_15_data_out[4:2];
  wire [31:0]       exeRequestQueue_queue_dataOut_15_source2 = _exeRequestQueue_queue_fifo_15_data_out[36:5];
  wire [31:0]       exeRequestQueue_queue_dataOut_15_source1 = _exeRequestQueue_queue_fifo_15_data_out[68:37];
  wire              exeRequestQueue_15_enq_ready = ~_exeRequestQueue_queue_fifo_15_full;
  wire              exeRequestQueue_15_deq_ready;
  wire              exeRequestQueue_15_deq_valid = ~_exeRequestQueue_queue_fifo_15_empty | exeRequestQueue_15_enq_valid;
  wire [31:0]       exeRequestQueue_15_deq_bits_source1 = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_source1 : exeRequestQueue_queue_dataOut_15_source1;
  wire [31:0]       exeRequestQueue_15_deq_bits_source2 = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_source2 : exeRequestQueue_queue_dataOut_15_source2;
  wire [2:0]        exeRequestQueue_15_deq_bits_index = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_index : exeRequestQueue_queue_dataOut_15_index;
  wire              exeRequestQueue_15_deq_bits_ffo = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_ffo : exeRequestQueue_queue_dataOut_15_ffo;
  wire              exeRequestQueue_15_deq_bits_fpReduceValid = _exeRequestQueue_queue_fifo_15_empty ? exeRequestQueue_15_enq_bits_fpReduceValid : exeRequestQueue_queue_dataOut_15_fpReduceValid;
  wire              tokenIO_15_maskRequestRelease_0 = exeRequestQueue_15_deq_ready & exeRequestQueue_15_deq_valid;
  reg               exeReqReg_0_valid;
  reg  [31:0]       exeReqReg_0_bits_source1;
  reg  [31:0]       exeReqReg_0_bits_source2;
  reg  [2:0]        exeReqReg_0_bits_index;
  reg               exeReqReg_0_bits_ffo;
  reg               exeReqReg_0_bits_fpReduceValid;
  reg               exeReqReg_1_valid;
  reg  [31:0]       exeReqReg_1_bits_source1;
  reg  [31:0]       exeReqReg_1_bits_source2;
  reg  [2:0]        exeReqReg_1_bits_index;
  reg               exeReqReg_1_bits_ffo;
  reg               exeReqReg_1_bits_fpReduceValid;
  reg               exeReqReg_2_valid;
  reg  [31:0]       exeReqReg_2_bits_source1;
  reg  [31:0]       exeReqReg_2_bits_source2;
  reg  [2:0]        exeReqReg_2_bits_index;
  reg               exeReqReg_2_bits_ffo;
  reg               exeReqReg_2_bits_fpReduceValid;
  reg               exeReqReg_3_valid;
  reg  [31:0]       exeReqReg_3_bits_source1;
  reg  [31:0]       exeReqReg_3_bits_source2;
  reg  [2:0]        exeReqReg_3_bits_index;
  reg               exeReqReg_3_bits_ffo;
  reg               exeReqReg_3_bits_fpReduceValid;
  reg               exeReqReg_4_valid;
  reg  [31:0]       exeReqReg_4_bits_source1;
  reg  [31:0]       exeReqReg_4_bits_source2;
  reg  [2:0]        exeReqReg_4_bits_index;
  reg               exeReqReg_4_bits_ffo;
  reg               exeReqReg_4_bits_fpReduceValid;
  reg               exeReqReg_5_valid;
  reg  [31:0]       exeReqReg_5_bits_source1;
  reg  [31:0]       exeReqReg_5_bits_source2;
  reg  [2:0]        exeReqReg_5_bits_index;
  reg               exeReqReg_5_bits_ffo;
  reg               exeReqReg_5_bits_fpReduceValid;
  reg               exeReqReg_6_valid;
  reg  [31:0]       exeReqReg_6_bits_source1;
  reg  [31:0]       exeReqReg_6_bits_source2;
  reg  [2:0]        exeReqReg_6_bits_index;
  reg               exeReqReg_6_bits_ffo;
  reg               exeReqReg_6_bits_fpReduceValid;
  reg               exeReqReg_7_valid;
  reg  [31:0]       exeReqReg_7_bits_source1;
  reg  [31:0]       exeReqReg_7_bits_source2;
  reg  [2:0]        exeReqReg_7_bits_index;
  reg               exeReqReg_7_bits_ffo;
  reg               exeReqReg_7_bits_fpReduceValid;
  reg               exeReqReg_8_valid;
  reg  [31:0]       exeReqReg_8_bits_source1;
  reg  [31:0]       exeReqReg_8_bits_source2;
  reg  [2:0]        exeReqReg_8_bits_index;
  reg               exeReqReg_8_bits_ffo;
  reg               exeReqReg_8_bits_fpReduceValid;
  reg               exeReqReg_9_valid;
  reg  [31:0]       exeReqReg_9_bits_source1;
  reg  [31:0]       exeReqReg_9_bits_source2;
  reg  [2:0]        exeReqReg_9_bits_index;
  reg               exeReqReg_9_bits_ffo;
  reg               exeReqReg_9_bits_fpReduceValid;
  reg               exeReqReg_10_valid;
  reg  [31:0]       exeReqReg_10_bits_source1;
  reg  [31:0]       exeReqReg_10_bits_source2;
  reg  [2:0]        exeReqReg_10_bits_index;
  reg               exeReqReg_10_bits_ffo;
  reg               exeReqReg_10_bits_fpReduceValid;
  reg               exeReqReg_11_valid;
  reg  [31:0]       exeReqReg_11_bits_source1;
  reg  [31:0]       exeReqReg_11_bits_source2;
  reg  [2:0]        exeReqReg_11_bits_index;
  reg               exeReqReg_11_bits_ffo;
  reg               exeReqReg_11_bits_fpReduceValid;
  reg               exeReqReg_12_valid;
  reg  [31:0]       exeReqReg_12_bits_source1;
  reg  [31:0]       exeReqReg_12_bits_source2;
  reg  [2:0]        exeReqReg_12_bits_index;
  reg               exeReqReg_12_bits_ffo;
  reg               exeReqReg_12_bits_fpReduceValid;
  reg               exeReqReg_13_valid;
  reg  [31:0]       exeReqReg_13_bits_source1;
  reg  [31:0]       exeReqReg_13_bits_source2;
  reg  [2:0]        exeReqReg_13_bits_index;
  reg               exeReqReg_13_bits_ffo;
  reg               exeReqReg_13_bits_fpReduceValid;
  reg               exeReqReg_14_valid;
  reg  [31:0]       exeReqReg_14_bits_source1;
  reg  [31:0]       exeReqReg_14_bits_source2;
  reg  [2:0]        exeReqReg_14_bits_index;
  reg               exeReqReg_14_bits_ffo;
  reg               exeReqReg_14_bits_fpReduceValid;
  reg               exeReqReg_15_valid;
  reg  [31:0]       exeReqReg_15_bits_source1;
  reg  [31:0]       exeReqReg_15_bits_source2;
  reg  [2:0]        exeReqReg_15_bits_index;
  reg               exeReqReg_15_bits_ffo;
  reg               exeReqReg_15_bits_fpReduceValid;
  reg  [4:0]        requestCounter;
  wire [5:0]        _GEN_39 = {1'h0, requestCounter};
  wire              counterValid = _GEN_39 <= lastGroupForInstruction;
  wire              lastGroup = _GEN_39 == lastGroupForInstruction | ~orderReduce & unitType[2] | mv;
  wire [127:0]      slideAddressGen_slideMaskInput_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo};
  wire [511:0]      slideAddressGen_slideMaskInput_lo = {slideAddressGen_slideMaskInput_lo_hi, slideAddressGen_slideMaskInput_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo};
  wire [127:0]      slideAddressGen_slideMaskInput_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo};
  wire [255:0]      slideAddressGen_slideMaskInput_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo};
  wire [511:0]      slideAddressGen_slideMaskInput_hi = {slideAddressGen_slideMaskInput_hi_hi, slideAddressGen_slideMaskInput_hi_lo};
  wire [63:0][15:0] _GEN_40 =
    {{slideAddressGen_slideMaskInput_hi[511:496]},
     {slideAddressGen_slideMaskInput_hi[495:480]},
     {slideAddressGen_slideMaskInput_hi[479:464]},
     {slideAddressGen_slideMaskInput_hi[463:448]},
     {slideAddressGen_slideMaskInput_hi[447:432]},
     {slideAddressGen_slideMaskInput_hi[431:416]},
     {slideAddressGen_slideMaskInput_hi[415:400]},
     {slideAddressGen_slideMaskInput_hi[399:384]},
     {slideAddressGen_slideMaskInput_hi[383:368]},
     {slideAddressGen_slideMaskInput_hi[367:352]},
     {slideAddressGen_slideMaskInput_hi[351:336]},
     {slideAddressGen_slideMaskInput_hi[335:320]},
     {slideAddressGen_slideMaskInput_hi[319:304]},
     {slideAddressGen_slideMaskInput_hi[303:288]},
     {slideAddressGen_slideMaskInput_hi[287:272]},
     {slideAddressGen_slideMaskInput_hi[271:256]},
     {slideAddressGen_slideMaskInput_hi[255:240]},
     {slideAddressGen_slideMaskInput_hi[239:224]},
     {slideAddressGen_slideMaskInput_hi[223:208]},
     {slideAddressGen_slideMaskInput_hi[207:192]},
     {slideAddressGen_slideMaskInput_hi[191:176]},
     {slideAddressGen_slideMaskInput_hi[175:160]},
     {slideAddressGen_slideMaskInput_hi[159:144]},
     {slideAddressGen_slideMaskInput_hi[143:128]},
     {slideAddressGen_slideMaskInput_hi[127:112]},
     {slideAddressGen_slideMaskInput_hi[111:96]},
     {slideAddressGen_slideMaskInput_hi[95:80]},
     {slideAddressGen_slideMaskInput_hi[79:64]},
     {slideAddressGen_slideMaskInput_hi[63:48]},
     {slideAddressGen_slideMaskInput_hi[47:32]},
     {slideAddressGen_slideMaskInput_hi[31:16]},
     {slideAddressGen_slideMaskInput_hi[15:0]},
     {slideAddressGen_slideMaskInput_lo[511:496]},
     {slideAddressGen_slideMaskInput_lo[495:480]},
     {slideAddressGen_slideMaskInput_lo[479:464]},
     {slideAddressGen_slideMaskInput_lo[463:448]},
     {slideAddressGen_slideMaskInput_lo[447:432]},
     {slideAddressGen_slideMaskInput_lo[431:416]},
     {slideAddressGen_slideMaskInput_lo[415:400]},
     {slideAddressGen_slideMaskInput_lo[399:384]},
     {slideAddressGen_slideMaskInput_lo[383:368]},
     {slideAddressGen_slideMaskInput_lo[367:352]},
     {slideAddressGen_slideMaskInput_lo[351:336]},
     {slideAddressGen_slideMaskInput_lo[335:320]},
     {slideAddressGen_slideMaskInput_lo[319:304]},
     {slideAddressGen_slideMaskInput_lo[303:288]},
     {slideAddressGen_slideMaskInput_lo[287:272]},
     {slideAddressGen_slideMaskInput_lo[271:256]},
     {slideAddressGen_slideMaskInput_lo[255:240]},
     {slideAddressGen_slideMaskInput_lo[239:224]},
     {slideAddressGen_slideMaskInput_lo[223:208]},
     {slideAddressGen_slideMaskInput_lo[207:192]},
     {slideAddressGen_slideMaskInput_lo[191:176]},
     {slideAddressGen_slideMaskInput_lo[175:160]},
     {slideAddressGen_slideMaskInput_lo[159:144]},
     {slideAddressGen_slideMaskInput_lo[143:128]},
     {slideAddressGen_slideMaskInput_lo[127:112]},
     {slideAddressGen_slideMaskInput_lo[111:96]},
     {slideAddressGen_slideMaskInput_lo[95:80]},
     {slideAddressGen_slideMaskInput_lo[79:64]},
     {slideAddressGen_slideMaskInput_lo[63:48]},
     {slideAddressGen_slideMaskInput_lo[47:32]},
     {slideAddressGen_slideMaskInput_lo[31:16]},
     {slideAddressGen_slideMaskInput_lo[15:0]}};
  wire              lastExecuteGroupDeq;
  wire              viotaCounterAdd;
  wire              groupCounterAdd = noSource ? viotaCounterAdd : lastExecuteGroupDeq;
  wire [15:0]       groupDataNeed = lastGroup ? lastGroupDataNeed : 16'hFFFF;
  reg  [1:0]        executeIndex;
  reg  [15:0]       readIssueStageState_groupReadState;
  reg  [15:0]       readIssueStageState_needRead;
  wire [15:0]       readWaitQueue_enq_bits_needRead = readIssueStageState_needRead;
  reg  [15:0]       readIssueStageState_elementValid;
  wire [15:0]       readWaitQueue_enq_bits_sourceValid = readIssueStageState_elementValid;
  reg  [15:0]       readIssueStageState_replaceVs1;
  wire [15:0]       readWaitQueue_enq_bits_replaceVs1 = readIssueStageState_replaceVs1;
  reg  [15:0]       readIssueStageState_readOffset;
  reg  [3:0]        readIssueStageState_accessLane_0;
  reg  [3:0]        readIssueStageState_accessLane_1;
  wire [3:0]        selectExecuteReq_1_bits_readLane = readIssueStageState_accessLane_1;
  reg  [3:0]        readIssueStageState_accessLane_2;
  wire [3:0]        selectExecuteReq_2_bits_readLane = readIssueStageState_accessLane_2;
  reg  [3:0]        readIssueStageState_accessLane_3;
  wire [3:0]        selectExecuteReq_3_bits_readLane = readIssueStageState_accessLane_3;
  reg  [3:0]        readIssueStageState_accessLane_4;
  wire [3:0]        selectExecuteReq_4_bits_readLane = readIssueStageState_accessLane_4;
  reg  [3:0]        readIssueStageState_accessLane_5;
  wire [3:0]        selectExecuteReq_5_bits_readLane = readIssueStageState_accessLane_5;
  reg  [3:0]        readIssueStageState_accessLane_6;
  wire [3:0]        selectExecuteReq_6_bits_readLane = readIssueStageState_accessLane_6;
  reg  [3:0]        readIssueStageState_accessLane_7;
  wire [3:0]        selectExecuteReq_7_bits_readLane = readIssueStageState_accessLane_7;
  reg  [3:0]        readIssueStageState_accessLane_8;
  wire [3:0]        selectExecuteReq_8_bits_readLane = readIssueStageState_accessLane_8;
  reg  [3:0]        readIssueStageState_accessLane_9;
  wire [3:0]        selectExecuteReq_9_bits_readLane = readIssueStageState_accessLane_9;
  reg  [3:0]        readIssueStageState_accessLane_10;
  wire [3:0]        selectExecuteReq_10_bits_readLane = readIssueStageState_accessLane_10;
  reg  [3:0]        readIssueStageState_accessLane_11;
  wire [3:0]        selectExecuteReq_11_bits_readLane = readIssueStageState_accessLane_11;
  reg  [3:0]        readIssueStageState_accessLane_12;
  wire [3:0]        selectExecuteReq_12_bits_readLane = readIssueStageState_accessLane_12;
  reg  [3:0]        readIssueStageState_accessLane_13;
  wire [3:0]        selectExecuteReq_13_bits_readLane = readIssueStageState_accessLane_13;
  reg  [3:0]        readIssueStageState_accessLane_14;
  wire [3:0]        selectExecuteReq_14_bits_readLane = readIssueStageState_accessLane_14;
  reg  [3:0]        readIssueStageState_accessLane_15;
  wire [3:0]        selectExecuteReq_15_bits_readLane = readIssueStageState_accessLane_15;
  reg  [2:0]        readIssueStageState_vsGrowth_0;
  reg  [2:0]        readIssueStageState_vsGrowth_1;
  reg  [2:0]        readIssueStageState_vsGrowth_2;
  reg  [2:0]        readIssueStageState_vsGrowth_3;
  reg  [2:0]        readIssueStageState_vsGrowth_4;
  reg  [2:0]        readIssueStageState_vsGrowth_5;
  reg  [2:0]        readIssueStageState_vsGrowth_6;
  reg  [2:0]        readIssueStageState_vsGrowth_7;
  reg  [2:0]        readIssueStageState_vsGrowth_8;
  reg  [2:0]        readIssueStageState_vsGrowth_9;
  reg  [2:0]        readIssueStageState_vsGrowth_10;
  reg  [2:0]        readIssueStageState_vsGrowth_11;
  reg  [2:0]        readIssueStageState_vsGrowth_12;
  reg  [2:0]        readIssueStageState_vsGrowth_13;
  reg  [2:0]        readIssueStageState_vsGrowth_14;
  reg  [2:0]        readIssueStageState_vsGrowth_15;
  reg  [6:0]        readIssueStageState_executeGroup;
  wire [6:0]        readWaitQueue_enq_bits_executeGroup = readIssueStageState_executeGroup;
  reg  [31:0]       readIssueStageState_readDataOffset;
  reg               readIssueStageState_last;
  wire              readWaitQueue_enq_bits_last = readIssueStageState_last;
  reg               readIssueStageValid;
  wire [4:0]        accessCountQueue_enq_bits_0 = accessCountEnq_0;
  wire [4:0]        accessCountQueue_enq_bits_1 = accessCountEnq_1;
  wire [4:0]        accessCountQueue_enq_bits_2 = accessCountEnq_2;
  wire [4:0]        accessCountQueue_enq_bits_3 = accessCountEnq_3;
  wire [4:0]        accessCountQueue_enq_bits_4 = accessCountEnq_4;
  wire [4:0]        accessCountQueue_enq_bits_5 = accessCountEnq_5;
  wire [4:0]        accessCountQueue_enq_bits_6 = accessCountEnq_6;
  wire [4:0]        accessCountQueue_enq_bits_7 = accessCountEnq_7;
  wire [4:0]        accessCountQueue_enq_bits_8 = accessCountEnq_8;
  wire [4:0]        accessCountQueue_enq_bits_9 = accessCountEnq_9;
  wire [4:0]        accessCountQueue_enq_bits_10 = accessCountEnq_10;
  wire [4:0]        accessCountQueue_enq_bits_11 = accessCountEnq_11;
  wire [4:0]        accessCountQueue_enq_bits_12 = accessCountEnq_12;
  wire [4:0]        accessCountQueue_enq_bits_13 = accessCountEnq_13;
  wire [4:0]        accessCountQueue_enq_bits_14 = accessCountEnq_14;
  wire [4:0]        accessCountQueue_enq_bits_15 = accessCountEnq_15;
  wire              readIssueStageEnq;
  wire              accessCountQueue_deq_valid;
  assign accessCountQueue_deq_valid = ~_accessCountQueue_fifo_empty;
  wire [4:0]        accessCountQueue_dataOut_0;
  wire [4:0]        accessCountQueue_dataOut_1;
  wire [4:0]        accessCountQueue_dataOut_2;
  wire [4:0]        accessCountQueue_dataOut_3;
  wire [4:0]        accessCountQueue_dataOut_4;
  wire [4:0]        accessCountQueue_dataOut_5;
  wire [4:0]        accessCountQueue_dataOut_6;
  wire [4:0]        accessCountQueue_dataOut_7;
  wire [4:0]        accessCountQueue_dataOut_8;
  wire [4:0]        accessCountQueue_dataOut_9;
  wire [4:0]        accessCountQueue_dataOut_10;
  wire [4:0]        accessCountQueue_dataOut_11;
  wire [4:0]        accessCountQueue_dataOut_12;
  wire [4:0]        accessCountQueue_dataOut_13;
  wire [4:0]        accessCountQueue_dataOut_14;
  wire [4:0]        accessCountQueue_dataOut_15;
  wire [9:0]        accessCountQueue_dataIn_lo_lo_lo = {accessCountQueue_enq_bits_1, accessCountQueue_enq_bits_0};
  wire [9:0]        accessCountQueue_dataIn_lo_lo_hi = {accessCountQueue_enq_bits_3, accessCountQueue_enq_bits_2};
  wire [19:0]       accessCountQueue_dataIn_lo_lo = {accessCountQueue_dataIn_lo_lo_hi, accessCountQueue_dataIn_lo_lo_lo};
  wire [9:0]        accessCountQueue_dataIn_lo_hi_lo = {accessCountQueue_enq_bits_5, accessCountQueue_enq_bits_4};
  wire [9:0]        accessCountQueue_dataIn_lo_hi_hi = {accessCountQueue_enq_bits_7, accessCountQueue_enq_bits_6};
  wire [19:0]       accessCountQueue_dataIn_lo_hi = {accessCountQueue_dataIn_lo_hi_hi, accessCountQueue_dataIn_lo_hi_lo};
  wire [39:0]       accessCountQueue_dataIn_lo = {accessCountQueue_dataIn_lo_hi, accessCountQueue_dataIn_lo_lo};
  wire [9:0]        accessCountQueue_dataIn_hi_lo_lo = {accessCountQueue_enq_bits_9, accessCountQueue_enq_bits_8};
  wire [9:0]        accessCountQueue_dataIn_hi_lo_hi = {accessCountQueue_enq_bits_11, accessCountQueue_enq_bits_10};
  wire [19:0]       accessCountQueue_dataIn_hi_lo = {accessCountQueue_dataIn_hi_lo_hi, accessCountQueue_dataIn_hi_lo_lo};
  wire [9:0]        accessCountQueue_dataIn_hi_hi_lo = {accessCountQueue_enq_bits_13, accessCountQueue_enq_bits_12};
  wire [9:0]        accessCountQueue_dataIn_hi_hi_hi = {accessCountQueue_enq_bits_15, accessCountQueue_enq_bits_14};
  wire [19:0]       accessCountQueue_dataIn_hi_hi = {accessCountQueue_dataIn_hi_hi_hi, accessCountQueue_dataIn_hi_hi_lo};
  wire [39:0]       accessCountQueue_dataIn_hi = {accessCountQueue_dataIn_hi_hi, accessCountQueue_dataIn_hi_lo};
  wire [79:0]       accessCountQueue_dataIn = {accessCountQueue_dataIn_hi, accessCountQueue_dataIn_lo};
  assign accessCountQueue_dataOut_0 = _accessCountQueue_fifo_data_out[4:0];
  assign accessCountQueue_dataOut_1 = _accessCountQueue_fifo_data_out[9:5];
  assign accessCountQueue_dataOut_2 = _accessCountQueue_fifo_data_out[14:10];
  assign accessCountQueue_dataOut_3 = _accessCountQueue_fifo_data_out[19:15];
  assign accessCountQueue_dataOut_4 = _accessCountQueue_fifo_data_out[24:20];
  assign accessCountQueue_dataOut_5 = _accessCountQueue_fifo_data_out[29:25];
  assign accessCountQueue_dataOut_6 = _accessCountQueue_fifo_data_out[34:30];
  assign accessCountQueue_dataOut_7 = _accessCountQueue_fifo_data_out[39:35];
  assign accessCountQueue_dataOut_8 = _accessCountQueue_fifo_data_out[44:40];
  assign accessCountQueue_dataOut_9 = _accessCountQueue_fifo_data_out[49:45];
  assign accessCountQueue_dataOut_10 = _accessCountQueue_fifo_data_out[54:50];
  assign accessCountQueue_dataOut_11 = _accessCountQueue_fifo_data_out[59:55];
  assign accessCountQueue_dataOut_12 = _accessCountQueue_fifo_data_out[64:60];
  assign accessCountQueue_dataOut_13 = _accessCountQueue_fifo_data_out[69:65];
  assign accessCountQueue_dataOut_14 = _accessCountQueue_fifo_data_out[74:70];
  assign accessCountQueue_dataOut_15 = _accessCountQueue_fifo_data_out[79:75];
  wire [4:0]        accessCountQueue_deq_bits_0 = accessCountQueue_dataOut_0;
  wire [4:0]        accessCountQueue_deq_bits_1 = accessCountQueue_dataOut_1;
  wire [4:0]        accessCountQueue_deq_bits_2 = accessCountQueue_dataOut_2;
  wire [4:0]        accessCountQueue_deq_bits_3 = accessCountQueue_dataOut_3;
  wire [4:0]        accessCountQueue_deq_bits_4 = accessCountQueue_dataOut_4;
  wire [4:0]        accessCountQueue_deq_bits_5 = accessCountQueue_dataOut_5;
  wire [4:0]        accessCountQueue_deq_bits_6 = accessCountQueue_dataOut_6;
  wire [4:0]        accessCountQueue_deq_bits_7 = accessCountQueue_dataOut_7;
  wire [4:0]        accessCountQueue_deq_bits_8 = accessCountQueue_dataOut_8;
  wire [4:0]        accessCountQueue_deq_bits_9 = accessCountQueue_dataOut_9;
  wire [4:0]        accessCountQueue_deq_bits_10 = accessCountQueue_dataOut_10;
  wire [4:0]        accessCountQueue_deq_bits_11 = accessCountQueue_dataOut_11;
  wire [4:0]        accessCountQueue_deq_bits_12 = accessCountQueue_dataOut_12;
  wire [4:0]        accessCountQueue_deq_bits_13 = accessCountQueue_dataOut_13;
  wire [4:0]        accessCountQueue_deq_bits_14 = accessCountQueue_dataOut_14;
  wire [4:0]        accessCountQueue_deq_bits_15 = accessCountQueue_dataOut_15;
  wire              accessCountQueue_enq_ready = ~_accessCountQueue_fifo_full;
  wire              accessCountQueue_enq_valid;
  wire              accessCountQueue_deq_ready;
  wire [6:0]        _extendGroupCount_T_1 = {requestCounter, executeIndex};
  wire [6:0]        _executeGroup_T_8 = executeIndexGrowth[0] ? _extendGroupCount_T_1 : 7'h0;
  wire [5:0]        _GEN_41 = _executeGroup_T_8[5:0] | (executeIndexGrowth[1] ? {requestCounter, executeIndex[1]} : 6'h0);
  wire [6:0]        executeGroup = {_executeGroup_T_8[6], _GEN_41[5], _GEN_41[4:0] | (executeIndexGrowth[2] ? requestCounter : 5'h0)};
  wire              vlMisAlign;
  assign vlMisAlign = |(instReg_vl[3:0]);
  wire [6:0]        lastexecuteGroup = instReg_vl[10:4] - {6'h0, ~vlMisAlign};
  wire              isVlBoundary = executeGroup == lastexecuteGroup;
  wire              validExecuteGroup = executeGroup <= lastexecuteGroup;
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_49 = 16'h1 << instReg_vl[3:0];
  wire [15:0]       _vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_49 | {_maskSplit_vlBoundaryCorrection_T_49[14:0], 1'h0};
  wire [15:0]       _vlBoundaryCorrection_T_8 = _vlBoundaryCorrection_T_5 | {_vlBoundaryCorrection_T_5[13:0], 2'h0};
  wire [15:0]       _vlBoundaryCorrection_T_11 = _vlBoundaryCorrection_T_8 | {_vlBoundaryCorrection_T_8[11:0], 4'h0};
  wire [15:0]       vlBoundaryCorrection = ~({16{vlMisAlign & isVlBoundary}} & (_vlBoundaryCorrection_T_11 | {_vlBoundaryCorrection_T_11[7:0], 8'h0})) & {16{validExecuteGroup}};
  wire [127:0]      selectReadStageMask_lo_lo_lo = {selectReadStageMask_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo};
  wire [127:0]      selectReadStageMask_lo_lo_hi = {selectReadStageMask_lo_lo_hi_hi, selectReadStageMask_lo_lo_hi_lo};
  wire [255:0]      selectReadStageMask_lo_lo = {selectReadStageMask_lo_lo_hi, selectReadStageMask_lo_lo_lo};
  wire [127:0]      selectReadStageMask_lo_hi_lo = {selectReadStageMask_lo_hi_lo_hi, selectReadStageMask_lo_hi_lo_lo};
  wire [127:0]      selectReadStageMask_lo_hi_hi = {selectReadStageMask_lo_hi_hi_hi, selectReadStageMask_lo_hi_hi_lo};
  wire [255:0]      selectReadStageMask_lo_hi = {selectReadStageMask_lo_hi_hi, selectReadStageMask_lo_hi_lo};
  wire [511:0]      selectReadStageMask_lo = {selectReadStageMask_lo_hi, selectReadStageMask_lo_lo};
  wire [127:0]      selectReadStageMask_hi_lo_lo = {selectReadStageMask_hi_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo};
  wire [127:0]      selectReadStageMask_hi_lo_hi = {selectReadStageMask_hi_lo_hi_hi, selectReadStageMask_hi_lo_hi_lo};
  wire [255:0]      selectReadStageMask_hi_lo = {selectReadStageMask_hi_lo_hi, selectReadStageMask_hi_lo_lo};
  wire [127:0]      selectReadStageMask_hi_hi_lo = {selectReadStageMask_hi_hi_lo_hi, selectReadStageMask_hi_hi_lo_lo};
  wire [127:0]      selectReadStageMask_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_lo};
  wire [255:0]      selectReadStageMask_hi_hi = {selectReadStageMask_hi_hi_hi, selectReadStageMask_hi_hi_lo};
  wire [511:0]      selectReadStageMask_hi = {selectReadStageMask_hi_hi, selectReadStageMask_hi_lo};
  wire [63:0][15:0] _GEN_42 =
    {{selectReadStageMask_hi[511:496]},
     {selectReadStageMask_hi[495:480]},
     {selectReadStageMask_hi[479:464]},
     {selectReadStageMask_hi[463:448]},
     {selectReadStageMask_hi[447:432]},
     {selectReadStageMask_hi[431:416]},
     {selectReadStageMask_hi[415:400]},
     {selectReadStageMask_hi[399:384]},
     {selectReadStageMask_hi[383:368]},
     {selectReadStageMask_hi[367:352]},
     {selectReadStageMask_hi[351:336]},
     {selectReadStageMask_hi[335:320]},
     {selectReadStageMask_hi[319:304]},
     {selectReadStageMask_hi[303:288]},
     {selectReadStageMask_hi[287:272]},
     {selectReadStageMask_hi[271:256]},
     {selectReadStageMask_hi[255:240]},
     {selectReadStageMask_hi[239:224]},
     {selectReadStageMask_hi[223:208]},
     {selectReadStageMask_hi[207:192]},
     {selectReadStageMask_hi[191:176]},
     {selectReadStageMask_hi[175:160]},
     {selectReadStageMask_hi[159:144]},
     {selectReadStageMask_hi[143:128]},
     {selectReadStageMask_hi[127:112]},
     {selectReadStageMask_hi[111:96]},
     {selectReadStageMask_hi[95:80]},
     {selectReadStageMask_hi[79:64]},
     {selectReadStageMask_hi[63:48]},
     {selectReadStageMask_hi[47:32]},
     {selectReadStageMask_hi[31:16]},
     {selectReadStageMask_hi[15:0]},
     {selectReadStageMask_lo[511:496]},
     {selectReadStageMask_lo[495:480]},
     {selectReadStageMask_lo[479:464]},
     {selectReadStageMask_lo[463:448]},
     {selectReadStageMask_lo[447:432]},
     {selectReadStageMask_lo[431:416]},
     {selectReadStageMask_lo[415:400]},
     {selectReadStageMask_lo[399:384]},
     {selectReadStageMask_lo[383:368]},
     {selectReadStageMask_lo[367:352]},
     {selectReadStageMask_lo[351:336]},
     {selectReadStageMask_lo[335:320]},
     {selectReadStageMask_lo[319:304]},
     {selectReadStageMask_lo[303:288]},
     {selectReadStageMask_lo[287:272]},
     {selectReadStageMask_lo[271:256]},
     {selectReadStageMask_lo[255:240]},
     {selectReadStageMask_lo[239:224]},
     {selectReadStageMask_lo[223:208]},
     {selectReadStageMask_lo[207:192]},
     {selectReadStageMask_lo[191:176]},
     {selectReadStageMask_lo[175:160]},
     {selectReadStageMask_lo[159:144]},
     {selectReadStageMask_lo[143:128]},
     {selectReadStageMask_lo[127:112]},
     {selectReadStageMask_lo[111:96]},
     {selectReadStageMask_lo[95:80]},
     {selectReadStageMask_lo[79:64]},
     {selectReadStageMask_lo[63:48]},
     {selectReadStageMask_lo[47:32]},
     {selectReadStageMask_lo[31:16]},
     {selectReadStageMask_lo[15:0]}};
  wire [15:0]       readMaskCorrection = (instReg_maskType ? _GEN_42[executeGroup[5:0]] : 16'hFFFF) & vlBoundaryCorrection;
  wire [127:0]      maskSplit_maskSelect_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo};
  wire [127:0]      maskSplit_maskSelect_lo_lo_hi = {maskSplit_maskSelect_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo};
  wire [255:0]      maskSplit_maskSelect_lo_lo = {maskSplit_maskSelect_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo};
  wire [127:0]      maskSplit_maskSelect_lo_hi_lo = {maskSplit_maskSelect_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo};
  wire [127:0]      maskSplit_maskSelect_lo_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo};
  wire [255:0]      maskSplit_maskSelect_lo_hi = {maskSplit_maskSelect_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo};
  wire [511:0]      maskSplit_maskSelect_lo = {maskSplit_maskSelect_lo_hi, maskSplit_maskSelect_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_lo_lo = {maskSplit_maskSelect_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_lo_hi = {maskSplit_maskSelect_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo};
  wire [255:0]      maskSplit_maskSelect_hi_lo = {maskSplit_maskSelect_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_hi_lo = {maskSplit_maskSelect_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo};
  wire [127:0]      maskSplit_maskSelect_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo};
  wire [255:0]      maskSplit_maskSelect_hi_hi = {maskSplit_maskSelect_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo};
  wire [511:0]      maskSplit_maskSelect_hi = {maskSplit_maskSelect_hi_hi, maskSplit_maskSelect_hi_lo};
  wire [4:0]        executeGroupCounter;
  wire              maskSplit_vlMisAlign = |(instReg_vl[5:0]);
  wire [4:0]        maskSplit_lastexecuteGroup = instReg_vl[10:6] - {4'h0, ~maskSplit_vlMisAlign};
  wire              maskSplit_isVlBoundary = executeGroupCounter == maskSplit_lastexecuteGroup;
  wire              maskSplit_validExecuteGroup = executeGroupCounter <= maskSplit_lastexecuteGroup;
  wire [63:0]       _maskSplit_vlBoundaryCorrection_T_2 = 64'h1 << instReg_vl[5:0];
  wire [63:0]       _maskSplit_vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_2 | {_maskSplit_vlBoundaryCorrection_T_2[62:0], 1'h0};
  wire [63:0]       _maskSplit_vlBoundaryCorrection_T_8 = _maskSplit_vlBoundaryCorrection_T_5 | {_maskSplit_vlBoundaryCorrection_T_5[61:0], 2'h0};
  wire [63:0]       _maskSplit_vlBoundaryCorrection_T_11 = _maskSplit_vlBoundaryCorrection_T_8 | {_maskSplit_vlBoundaryCorrection_T_8[59:0], 4'h0};
  wire [63:0]       _maskSplit_vlBoundaryCorrection_T_14 = _maskSplit_vlBoundaryCorrection_T_11 | {_maskSplit_vlBoundaryCorrection_T_11[55:0], 8'h0};
  wire [63:0]       _maskSplit_vlBoundaryCorrection_T_17 = _maskSplit_vlBoundaryCorrection_T_14 | {_maskSplit_vlBoundaryCorrection_T_14[47:0], 16'h0};
  wire [63:0]       maskSplit_vlBoundaryCorrection = ~({64{maskSplit_vlMisAlign & maskSplit_isVlBoundary}} & (_maskSplit_vlBoundaryCorrection_T_17 | {_maskSplit_vlBoundaryCorrection_T_17[31:0], 32'h0})) & {64{maskSplit_validExecuteGroup}};
  wire [15:0][63:0] _GEN_43 =
    {{maskSplit_maskSelect_hi[511:448]},
     {maskSplit_maskSelect_hi[447:384]},
     {maskSplit_maskSelect_hi[383:320]},
     {maskSplit_maskSelect_hi[319:256]},
     {maskSplit_maskSelect_hi[255:192]},
     {maskSplit_maskSelect_hi[191:128]},
     {maskSplit_maskSelect_hi[127:64]},
     {maskSplit_maskSelect_hi[63:0]},
     {maskSplit_maskSelect_lo[511:448]},
     {maskSplit_maskSelect_lo[447:384]},
     {maskSplit_maskSelect_lo[383:320]},
     {maskSplit_maskSelect_lo[319:256]},
     {maskSplit_maskSelect_lo[255:192]},
     {maskSplit_maskSelect_lo[191:128]},
     {maskSplit_maskSelect_lo[127:64]},
     {maskSplit_maskSelect_lo[63:0]}};
  wire [63:0]       maskSplit_0_2 = (instReg_maskType ? _GEN_43[executeGroupCounter[3:0]] : 64'hFFFFFFFFFFFFFFFF) & maskSplit_vlBoundaryCorrection;
  wire [1:0]        maskSplit_byteMask_lo_lo_lo_lo_lo = maskSplit_0_2[1:0];
  wire [1:0]        maskSplit_byteMask_lo_lo_lo_lo_hi = maskSplit_0_2[3:2];
  wire [3:0]        maskSplit_byteMask_lo_lo_lo_lo = {maskSplit_byteMask_lo_lo_lo_lo_hi, maskSplit_byteMask_lo_lo_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_lo_lo_hi_lo = maskSplit_0_2[5:4];
  wire [1:0]        maskSplit_byteMask_lo_lo_lo_hi_hi = maskSplit_0_2[7:6];
  wire [3:0]        maskSplit_byteMask_lo_lo_lo_hi = {maskSplit_byteMask_lo_lo_lo_hi_hi, maskSplit_byteMask_lo_lo_lo_hi_lo};
  wire [7:0]        maskSplit_byteMask_lo_lo_lo = {maskSplit_byteMask_lo_lo_lo_hi, maskSplit_byteMask_lo_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_lo_hi_lo_lo = maskSplit_0_2[9:8];
  wire [1:0]        maskSplit_byteMask_lo_lo_hi_lo_hi = maskSplit_0_2[11:10];
  wire [3:0]        maskSplit_byteMask_lo_lo_hi_lo = {maskSplit_byteMask_lo_lo_hi_lo_hi, maskSplit_byteMask_lo_lo_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_lo_hi_hi_lo = maskSplit_0_2[13:12];
  wire [1:0]        maskSplit_byteMask_lo_lo_hi_hi_hi = maskSplit_0_2[15:14];
  wire [3:0]        maskSplit_byteMask_lo_lo_hi_hi = {maskSplit_byteMask_lo_lo_hi_hi_hi, maskSplit_byteMask_lo_lo_hi_hi_lo};
  wire [7:0]        maskSplit_byteMask_lo_lo_hi = {maskSplit_byteMask_lo_lo_hi_hi, maskSplit_byteMask_lo_lo_hi_lo};
  wire [15:0]       maskSplit_byteMask_lo_lo = {maskSplit_byteMask_lo_lo_hi, maskSplit_byteMask_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_hi_lo_lo_lo = maskSplit_0_2[17:16];
  wire [1:0]        maskSplit_byteMask_lo_hi_lo_lo_hi = maskSplit_0_2[19:18];
  wire [3:0]        maskSplit_byteMask_lo_hi_lo_lo = {maskSplit_byteMask_lo_hi_lo_lo_hi, maskSplit_byteMask_lo_hi_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_hi_lo_hi_lo = maskSplit_0_2[21:20];
  wire [1:0]        maskSplit_byteMask_lo_hi_lo_hi_hi = maskSplit_0_2[23:22];
  wire [3:0]        maskSplit_byteMask_lo_hi_lo_hi = {maskSplit_byteMask_lo_hi_lo_hi_hi, maskSplit_byteMask_lo_hi_lo_hi_lo};
  wire [7:0]        maskSplit_byteMask_lo_hi_lo = {maskSplit_byteMask_lo_hi_lo_hi, maskSplit_byteMask_lo_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_hi_hi_lo_lo = maskSplit_0_2[25:24];
  wire [1:0]        maskSplit_byteMask_lo_hi_hi_lo_hi = maskSplit_0_2[27:26];
  wire [3:0]        maskSplit_byteMask_lo_hi_hi_lo = {maskSplit_byteMask_lo_hi_hi_lo_hi, maskSplit_byteMask_lo_hi_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_lo_hi_hi_hi_lo = maskSplit_0_2[29:28];
  wire [1:0]        maskSplit_byteMask_lo_hi_hi_hi_hi = maskSplit_0_2[31:30];
  wire [3:0]        maskSplit_byteMask_lo_hi_hi_hi = {maskSplit_byteMask_lo_hi_hi_hi_hi, maskSplit_byteMask_lo_hi_hi_hi_lo};
  wire [7:0]        maskSplit_byteMask_lo_hi_hi = {maskSplit_byteMask_lo_hi_hi_hi, maskSplit_byteMask_lo_hi_hi_lo};
  wire [15:0]       maskSplit_byteMask_lo_hi = {maskSplit_byteMask_lo_hi_hi, maskSplit_byteMask_lo_hi_lo};
  wire [31:0]       maskSplit_byteMask_lo = {maskSplit_byteMask_lo_hi, maskSplit_byteMask_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_lo_lo_lo_lo = maskSplit_0_2[33:32];
  wire [1:0]        maskSplit_byteMask_hi_lo_lo_lo_hi = maskSplit_0_2[35:34];
  wire [3:0]        maskSplit_byteMask_hi_lo_lo_lo = {maskSplit_byteMask_hi_lo_lo_lo_hi, maskSplit_byteMask_hi_lo_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_lo_lo_hi_lo = maskSplit_0_2[37:36];
  wire [1:0]        maskSplit_byteMask_hi_lo_lo_hi_hi = maskSplit_0_2[39:38];
  wire [3:0]        maskSplit_byteMask_hi_lo_lo_hi = {maskSplit_byteMask_hi_lo_lo_hi_hi, maskSplit_byteMask_hi_lo_lo_hi_lo};
  wire [7:0]        maskSplit_byteMask_hi_lo_lo = {maskSplit_byteMask_hi_lo_lo_hi, maskSplit_byteMask_hi_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_lo_hi_lo_lo = maskSplit_0_2[41:40];
  wire [1:0]        maskSplit_byteMask_hi_lo_hi_lo_hi = maskSplit_0_2[43:42];
  wire [3:0]        maskSplit_byteMask_hi_lo_hi_lo = {maskSplit_byteMask_hi_lo_hi_lo_hi, maskSplit_byteMask_hi_lo_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_lo_hi_hi_lo = maskSplit_0_2[45:44];
  wire [1:0]        maskSplit_byteMask_hi_lo_hi_hi_hi = maskSplit_0_2[47:46];
  wire [3:0]        maskSplit_byteMask_hi_lo_hi_hi = {maskSplit_byteMask_hi_lo_hi_hi_hi, maskSplit_byteMask_hi_lo_hi_hi_lo};
  wire [7:0]        maskSplit_byteMask_hi_lo_hi = {maskSplit_byteMask_hi_lo_hi_hi, maskSplit_byteMask_hi_lo_hi_lo};
  wire [15:0]       maskSplit_byteMask_hi_lo = {maskSplit_byteMask_hi_lo_hi, maskSplit_byteMask_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_hi_lo_lo_lo = maskSplit_0_2[49:48];
  wire [1:0]        maskSplit_byteMask_hi_hi_lo_lo_hi = maskSplit_0_2[51:50];
  wire [3:0]        maskSplit_byteMask_hi_hi_lo_lo = {maskSplit_byteMask_hi_hi_lo_lo_hi, maskSplit_byteMask_hi_hi_lo_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_hi_lo_hi_lo = maskSplit_0_2[53:52];
  wire [1:0]        maskSplit_byteMask_hi_hi_lo_hi_hi = maskSplit_0_2[55:54];
  wire [3:0]        maskSplit_byteMask_hi_hi_lo_hi = {maskSplit_byteMask_hi_hi_lo_hi_hi, maskSplit_byteMask_hi_hi_lo_hi_lo};
  wire [7:0]        maskSplit_byteMask_hi_hi_lo = {maskSplit_byteMask_hi_hi_lo_hi, maskSplit_byteMask_hi_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_hi_hi_lo_lo = maskSplit_0_2[57:56];
  wire [1:0]        maskSplit_byteMask_hi_hi_hi_lo_hi = maskSplit_0_2[59:58];
  wire [3:0]        maskSplit_byteMask_hi_hi_hi_lo = {maskSplit_byteMask_hi_hi_hi_lo_hi, maskSplit_byteMask_hi_hi_hi_lo_lo};
  wire [1:0]        maskSplit_byteMask_hi_hi_hi_hi_lo = maskSplit_0_2[61:60];
  wire [1:0]        maskSplit_byteMask_hi_hi_hi_hi_hi = maskSplit_0_2[63:62];
  wire [3:0]        maskSplit_byteMask_hi_hi_hi_hi = {maskSplit_byteMask_hi_hi_hi_hi_hi, maskSplit_byteMask_hi_hi_hi_hi_lo};
  wire [7:0]        maskSplit_byteMask_hi_hi_hi = {maskSplit_byteMask_hi_hi_hi_hi, maskSplit_byteMask_hi_hi_hi_lo};
  wire [15:0]       maskSplit_byteMask_hi_hi = {maskSplit_byteMask_hi_hi_hi, maskSplit_byteMask_hi_hi_lo};
  wire [31:0]       maskSplit_byteMask_hi = {maskSplit_byteMask_hi_hi, maskSplit_byteMask_hi_lo};
  wire [63:0]       maskSplit_0_1 = {maskSplit_byteMask_hi, maskSplit_byteMask_lo};
  wire [127:0]      maskSplit_maskSelect_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_1};
  wire [511:0]      maskSplit_maskSelect_lo_1 = {maskSplit_maskSelect_lo_hi_1, maskSplit_maskSelect_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_1};
  wire [127:0]      maskSplit_maskSelect_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_1};
  wire [255:0]      maskSplit_maskSelect_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_1};
  wire [511:0]      maskSplit_maskSelect_hi_1 = {maskSplit_maskSelect_hi_hi_1, maskSplit_maskSelect_hi_lo_1};
  wire              maskSplit_vlMisAlign_1 = |(instReg_vl[4:0]);
  wire [5:0]        maskSplit_lastexecuteGroup_1 = instReg_vl[10:5] - {5'h0, ~maskSplit_vlMisAlign_1};
  wire [5:0]        _GEN_44 = {1'h0, executeGroupCounter};
  wire              maskSplit_isVlBoundary_1 = _GEN_44 == maskSplit_lastexecuteGroup_1;
  wire              maskSplit_validExecuteGroup_1 = _GEN_44 <= maskSplit_lastexecuteGroup_1;
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_27 = 32'h1 << instReg_vl[4:0];
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_30 = _maskSplit_vlBoundaryCorrection_T_27 | {_maskSplit_vlBoundaryCorrection_T_27[30:0], 1'h0};
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_33 = _maskSplit_vlBoundaryCorrection_T_30 | {_maskSplit_vlBoundaryCorrection_T_30[29:0], 2'h0};
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_36 = _maskSplit_vlBoundaryCorrection_T_33 | {_maskSplit_vlBoundaryCorrection_T_33[27:0], 4'h0};
  wire [31:0]       _maskSplit_vlBoundaryCorrection_T_39 = _maskSplit_vlBoundaryCorrection_T_36 | {_maskSplit_vlBoundaryCorrection_T_36[23:0], 8'h0};
  wire [31:0]       maskSplit_vlBoundaryCorrection_1 =
    ~({32{maskSplit_vlMisAlign_1 & maskSplit_isVlBoundary_1}} & (_maskSplit_vlBoundaryCorrection_T_39 | {_maskSplit_vlBoundaryCorrection_T_39[15:0], 16'h0})) & {32{maskSplit_validExecuteGroup_1}};
  wire [31:0][31:0] _GEN_45 =
    {{maskSplit_maskSelect_hi_1[511:480]},
     {maskSplit_maskSelect_hi_1[479:448]},
     {maskSplit_maskSelect_hi_1[447:416]},
     {maskSplit_maskSelect_hi_1[415:384]},
     {maskSplit_maskSelect_hi_1[383:352]},
     {maskSplit_maskSelect_hi_1[351:320]},
     {maskSplit_maskSelect_hi_1[319:288]},
     {maskSplit_maskSelect_hi_1[287:256]},
     {maskSplit_maskSelect_hi_1[255:224]},
     {maskSplit_maskSelect_hi_1[223:192]},
     {maskSplit_maskSelect_hi_1[191:160]},
     {maskSplit_maskSelect_hi_1[159:128]},
     {maskSplit_maskSelect_hi_1[127:96]},
     {maskSplit_maskSelect_hi_1[95:64]},
     {maskSplit_maskSelect_hi_1[63:32]},
     {maskSplit_maskSelect_hi_1[31:0]},
     {maskSplit_maskSelect_lo_1[511:480]},
     {maskSplit_maskSelect_lo_1[479:448]},
     {maskSplit_maskSelect_lo_1[447:416]},
     {maskSplit_maskSelect_lo_1[415:384]},
     {maskSplit_maskSelect_lo_1[383:352]},
     {maskSplit_maskSelect_lo_1[351:320]},
     {maskSplit_maskSelect_lo_1[319:288]},
     {maskSplit_maskSelect_lo_1[287:256]},
     {maskSplit_maskSelect_lo_1[255:224]},
     {maskSplit_maskSelect_lo_1[223:192]},
     {maskSplit_maskSelect_lo_1[191:160]},
     {maskSplit_maskSelect_lo_1[159:128]},
     {maskSplit_maskSelect_lo_1[127:96]},
     {maskSplit_maskSelect_lo_1[95:64]},
     {maskSplit_maskSelect_lo_1[63:32]},
     {maskSplit_maskSelect_lo_1[31:0]}};
  wire [31:0]       maskSplit_1_2 = (instReg_maskType ? _GEN_45[executeGroupCounter] : 32'hFFFFFFFF) & maskSplit_vlBoundaryCorrection_1;
  wire [3:0]        maskSplit_byteMask_lo_lo_lo_lo_1 = {{2{maskSplit_1_2[1]}}, {2{maskSplit_1_2[0]}}};
  wire [3:0]        maskSplit_byteMask_lo_lo_lo_hi_1 = {{2{maskSplit_1_2[3]}}, {2{maskSplit_1_2[2]}}};
  wire [7:0]        maskSplit_byteMask_lo_lo_lo_1 = {maskSplit_byteMask_lo_lo_lo_hi_1, maskSplit_byteMask_lo_lo_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_lo_lo_hi_lo_1 = {{2{maskSplit_1_2[5]}}, {2{maskSplit_1_2[4]}}};
  wire [3:0]        maskSplit_byteMask_lo_lo_hi_hi_1 = {{2{maskSplit_1_2[7]}}, {2{maskSplit_1_2[6]}}};
  wire [7:0]        maskSplit_byteMask_lo_lo_hi_1 = {maskSplit_byteMask_lo_lo_hi_hi_1, maskSplit_byteMask_lo_lo_hi_lo_1};
  wire [15:0]       maskSplit_byteMask_lo_lo_1 = {maskSplit_byteMask_lo_lo_hi_1, maskSplit_byteMask_lo_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_lo_hi_lo_lo_1 = {{2{maskSplit_1_2[9]}}, {2{maskSplit_1_2[8]}}};
  wire [3:0]        maskSplit_byteMask_lo_hi_lo_hi_1 = {{2{maskSplit_1_2[11]}}, {2{maskSplit_1_2[10]}}};
  wire [7:0]        maskSplit_byteMask_lo_hi_lo_1 = {maskSplit_byteMask_lo_hi_lo_hi_1, maskSplit_byteMask_lo_hi_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_lo_hi_hi_lo_1 = {{2{maskSplit_1_2[13]}}, {2{maskSplit_1_2[12]}}};
  wire [3:0]        maskSplit_byteMask_lo_hi_hi_hi_1 = {{2{maskSplit_1_2[15]}}, {2{maskSplit_1_2[14]}}};
  wire [7:0]        maskSplit_byteMask_lo_hi_hi_1 = {maskSplit_byteMask_lo_hi_hi_hi_1, maskSplit_byteMask_lo_hi_hi_lo_1};
  wire [15:0]       maskSplit_byteMask_lo_hi_1 = {maskSplit_byteMask_lo_hi_hi_1, maskSplit_byteMask_lo_hi_lo_1};
  wire [31:0]       maskSplit_byteMask_lo_1 = {maskSplit_byteMask_lo_hi_1, maskSplit_byteMask_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_hi_lo_lo_lo_1 = {{2{maskSplit_1_2[17]}}, {2{maskSplit_1_2[16]}}};
  wire [3:0]        maskSplit_byteMask_hi_lo_lo_hi_1 = {{2{maskSplit_1_2[19]}}, {2{maskSplit_1_2[18]}}};
  wire [7:0]        maskSplit_byteMask_hi_lo_lo_1 = {maskSplit_byteMask_hi_lo_lo_hi_1, maskSplit_byteMask_hi_lo_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_hi_lo_hi_lo_1 = {{2{maskSplit_1_2[21]}}, {2{maskSplit_1_2[20]}}};
  wire [3:0]        maskSplit_byteMask_hi_lo_hi_hi_1 = {{2{maskSplit_1_2[23]}}, {2{maskSplit_1_2[22]}}};
  wire [7:0]        maskSplit_byteMask_hi_lo_hi_1 = {maskSplit_byteMask_hi_lo_hi_hi_1, maskSplit_byteMask_hi_lo_hi_lo_1};
  wire [15:0]       maskSplit_byteMask_hi_lo_1 = {maskSplit_byteMask_hi_lo_hi_1, maskSplit_byteMask_hi_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_hi_hi_lo_lo_1 = {{2{maskSplit_1_2[25]}}, {2{maskSplit_1_2[24]}}};
  wire [3:0]        maskSplit_byteMask_hi_hi_lo_hi_1 = {{2{maskSplit_1_2[27]}}, {2{maskSplit_1_2[26]}}};
  wire [7:0]        maskSplit_byteMask_hi_hi_lo_1 = {maskSplit_byteMask_hi_hi_lo_hi_1, maskSplit_byteMask_hi_hi_lo_lo_1};
  wire [3:0]        maskSplit_byteMask_hi_hi_hi_lo_1 = {{2{maskSplit_1_2[29]}}, {2{maskSplit_1_2[28]}}};
  wire [3:0]        maskSplit_byteMask_hi_hi_hi_hi_1 = {{2{maskSplit_1_2[31]}}, {2{maskSplit_1_2[30]}}};
  wire [7:0]        maskSplit_byteMask_hi_hi_hi_1 = {maskSplit_byteMask_hi_hi_hi_hi_1, maskSplit_byteMask_hi_hi_hi_lo_1};
  wire [15:0]       maskSplit_byteMask_hi_hi_1 = {maskSplit_byteMask_hi_hi_hi_1, maskSplit_byteMask_hi_hi_lo_1};
  wire [31:0]       maskSplit_byteMask_hi_1 = {maskSplit_byteMask_hi_hi_1, maskSplit_byteMask_hi_lo_1};
  wire [63:0]       maskSplit_1_1 = {maskSplit_byteMask_hi_1, maskSplit_byteMask_lo_1};
  wire [127:0]      maskSplit_maskSelect_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_2};
  wire [511:0]      maskSplit_maskSelect_lo_2 = {maskSplit_maskSelect_lo_hi_2, maskSplit_maskSelect_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_2};
  wire [127:0]      maskSplit_maskSelect_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_2};
  wire [255:0]      maskSplit_maskSelect_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_2};
  wire [511:0]      maskSplit_maskSelect_hi_2 = {maskSplit_maskSelect_hi_hi_2, maskSplit_maskSelect_hi_lo_2};
  wire              maskSplit_vlMisAlign_2;
  assign maskSplit_vlMisAlign_2 = |(instReg_vl[3:0]);
  wire [6:0]        maskSplit_lastexecuteGroup_2 = instReg_vl[10:4] - {6'h0, ~maskSplit_vlMisAlign_2};
  wire [6:0]        _GEN_46 = {2'h0, executeGroupCounter};
  wire              maskSplit_isVlBoundary_2 = _GEN_46 == maskSplit_lastexecuteGroup_2;
  wire              maskSplit_validExecuteGroup_2 = _GEN_46 <= maskSplit_lastexecuteGroup_2;
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_52 = _maskSplit_vlBoundaryCorrection_T_49 | {_maskSplit_vlBoundaryCorrection_T_49[14:0], 1'h0};
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_55 = _maskSplit_vlBoundaryCorrection_T_52 | {_maskSplit_vlBoundaryCorrection_T_52[13:0], 2'h0};
  wire [15:0]       _maskSplit_vlBoundaryCorrection_T_58 = _maskSplit_vlBoundaryCorrection_T_55 | {_maskSplit_vlBoundaryCorrection_T_55[11:0], 4'h0};
  wire [15:0]       maskSplit_vlBoundaryCorrection_2 =
    ~({16{maskSplit_vlMisAlign_2 & maskSplit_isVlBoundary_2}} & (_maskSplit_vlBoundaryCorrection_T_58 | {_maskSplit_vlBoundaryCorrection_T_58[7:0], 8'h0})) & {16{maskSplit_validExecuteGroup_2}};
  wire [31:0][15:0] _GEN_47 =
    {{maskSplit_maskSelect_lo_2[511:496]},
     {maskSplit_maskSelect_lo_2[495:480]},
     {maskSplit_maskSelect_lo_2[479:464]},
     {maskSplit_maskSelect_lo_2[463:448]},
     {maskSplit_maskSelect_lo_2[447:432]},
     {maskSplit_maskSelect_lo_2[431:416]},
     {maskSplit_maskSelect_lo_2[415:400]},
     {maskSplit_maskSelect_lo_2[399:384]},
     {maskSplit_maskSelect_lo_2[383:368]},
     {maskSplit_maskSelect_lo_2[367:352]},
     {maskSplit_maskSelect_lo_2[351:336]},
     {maskSplit_maskSelect_lo_2[335:320]},
     {maskSplit_maskSelect_lo_2[319:304]},
     {maskSplit_maskSelect_lo_2[303:288]},
     {maskSplit_maskSelect_lo_2[287:272]},
     {maskSplit_maskSelect_lo_2[271:256]},
     {maskSplit_maskSelect_lo_2[255:240]},
     {maskSplit_maskSelect_lo_2[239:224]},
     {maskSplit_maskSelect_lo_2[223:208]},
     {maskSplit_maskSelect_lo_2[207:192]},
     {maskSplit_maskSelect_lo_2[191:176]},
     {maskSplit_maskSelect_lo_2[175:160]},
     {maskSplit_maskSelect_lo_2[159:144]},
     {maskSplit_maskSelect_lo_2[143:128]},
     {maskSplit_maskSelect_lo_2[127:112]},
     {maskSplit_maskSelect_lo_2[111:96]},
     {maskSplit_maskSelect_lo_2[95:80]},
     {maskSplit_maskSelect_lo_2[79:64]},
     {maskSplit_maskSelect_lo_2[63:48]},
     {maskSplit_maskSelect_lo_2[47:32]},
     {maskSplit_maskSelect_lo_2[31:16]},
     {maskSplit_maskSelect_lo_2[15:0]}};
  wire [15:0]       maskSplit_2_2 = (instReg_maskType ? _GEN_47[executeGroupCounter] : 16'hFFFF) & maskSplit_vlBoundaryCorrection_2;
  wire [7:0]        maskSplit_byteMask_lo_lo_lo_2 = {{4{maskSplit_2_2[1]}}, {4{maskSplit_2_2[0]}}};
  wire [7:0]        maskSplit_byteMask_lo_lo_hi_2 = {{4{maskSplit_2_2[3]}}, {4{maskSplit_2_2[2]}}};
  wire [15:0]       maskSplit_byteMask_lo_lo_2 = {maskSplit_byteMask_lo_lo_hi_2, maskSplit_byteMask_lo_lo_lo_2};
  wire [7:0]        maskSplit_byteMask_lo_hi_lo_2 = {{4{maskSplit_2_2[5]}}, {4{maskSplit_2_2[4]}}};
  wire [7:0]        maskSplit_byteMask_lo_hi_hi_2 = {{4{maskSplit_2_2[7]}}, {4{maskSplit_2_2[6]}}};
  wire [15:0]       maskSplit_byteMask_lo_hi_2 = {maskSplit_byteMask_lo_hi_hi_2, maskSplit_byteMask_lo_hi_lo_2};
  wire [31:0]       maskSplit_byteMask_lo_2 = {maskSplit_byteMask_lo_hi_2, maskSplit_byteMask_lo_lo_2};
  wire [7:0]        maskSplit_byteMask_hi_lo_lo_2 = {{4{maskSplit_2_2[9]}}, {4{maskSplit_2_2[8]}}};
  wire [7:0]        maskSplit_byteMask_hi_lo_hi_2 = {{4{maskSplit_2_2[11]}}, {4{maskSplit_2_2[10]}}};
  wire [15:0]       maskSplit_byteMask_hi_lo_2 = {maskSplit_byteMask_hi_lo_hi_2, maskSplit_byteMask_hi_lo_lo_2};
  wire [7:0]        maskSplit_byteMask_hi_hi_lo_2 = {{4{maskSplit_2_2[13]}}, {4{maskSplit_2_2[12]}}};
  wire [7:0]        maskSplit_byteMask_hi_hi_hi_2 = {{4{maskSplit_2_2[15]}}, {4{maskSplit_2_2[14]}}};
  wire [15:0]       maskSplit_byteMask_hi_hi_2 = {maskSplit_byteMask_hi_hi_hi_2, maskSplit_byteMask_hi_hi_lo_2};
  wire [31:0]       maskSplit_byteMask_hi_2 = {maskSplit_byteMask_hi_hi_2, maskSplit_byteMask_hi_lo_2};
  wire [63:0]       maskSplit_2_1 = {maskSplit_byteMask_hi_2, maskSplit_byteMask_lo_2};
  wire [63:0]       executeByteMask = (sew1H[0] ? maskSplit_0_1 : 64'h0) | (sew1H[1] ? maskSplit_1_1 : 64'h0) | (sew1H[2] ? maskSplit_2_1 : 64'h0);
  wire [63:0]       _executeElementMask_T_3 = sew1H[0] ? maskSplit_0_2 : 64'h0;
  wire [31:0]       _GEN_48 = _executeElementMask_T_3[31:0] | (sew1H[1] ? maskSplit_1_2 : 32'h0);
  wire [63:0]       executeElementMask = {_executeElementMask_T_3[63:32], _GEN_48[31:16], _GEN_48[15:0] | (sew1H[2] ? maskSplit_2_2 : 16'h0)};
  wire [127:0]      maskForDestination_lo_lo_lo = {maskForDestination_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo};
  wire [127:0]      maskForDestination_lo_lo_hi = {maskForDestination_lo_lo_hi_hi, maskForDestination_lo_lo_hi_lo};
  wire [255:0]      maskForDestination_lo_lo = {maskForDestination_lo_lo_hi, maskForDestination_lo_lo_lo};
  wire [127:0]      maskForDestination_lo_hi_lo = {maskForDestination_lo_hi_lo_hi, maskForDestination_lo_hi_lo_lo};
  wire [127:0]      maskForDestination_lo_hi_hi = {maskForDestination_lo_hi_hi_hi, maskForDestination_lo_hi_hi_lo};
  wire [255:0]      maskForDestination_lo_hi = {maskForDestination_lo_hi_hi, maskForDestination_lo_hi_lo};
  wire [511:0]      maskForDestination_lo = {maskForDestination_lo_hi, maskForDestination_lo_lo};
  wire [127:0]      maskForDestination_hi_lo_lo = {maskForDestination_hi_lo_lo_hi, maskForDestination_hi_lo_lo_lo};
  wire [127:0]      maskForDestination_hi_lo_hi = {maskForDestination_hi_lo_hi_hi, maskForDestination_hi_lo_hi_lo};
  wire [255:0]      maskForDestination_hi_lo = {maskForDestination_hi_lo_hi, maskForDestination_hi_lo_lo};
  wire [127:0]      maskForDestination_hi_hi_lo = {maskForDestination_hi_hi_lo_hi, maskForDestination_hi_hi_lo_lo};
  wire [127:0]      maskForDestination_hi_hi_hi = {maskForDestination_hi_hi_hi_hi, maskForDestination_hi_hi_hi_lo};
  wire [255:0]      maskForDestination_hi_hi = {maskForDestination_hi_hi_hi, maskForDestination_hi_hi_lo};
  wire [511:0]      maskForDestination_hi = {maskForDestination_hi_hi, maskForDestination_hi_lo};
  wire              vs1Split_vs1SetIndex = requestCounter[0];
  wire [511:0]      _lastGroupMask_T = 512'h1 << elementTailForMaskDestination;
  wire [510:0]      _GEN_49 = _lastGroupMask_T[510:0] | _lastGroupMask_T[511:1];
  wire [509:0]      _GEN_50 = _GEN_49[509:0] | {_lastGroupMask_T[511], _GEN_49[510:2]};
  wire [507:0]      _GEN_51 = _GEN_50[507:0] | {_lastGroupMask_T[511], _GEN_49[510], _GEN_50[509:4]};
  wire [503:0]      _GEN_52 = _GEN_51[503:0] | {_lastGroupMask_T[511], _GEN_49[510], _GEN_50[509:508], _GEN_51[507:8]};
  wire [495:0]      _GEN_53 = _GEN_52[495:0] | {_lastGroupMask_T[511], _GEN_49[510], _GEN_50[509:508], _GEN_51[507:504], _GEN_52[503:16]};
  wire [479:0]      _GEN_54 = _GEN_53[479:0] | {_lastGroupMask_T[511], _GEN_49[510], _GEN_50[509:508], _GEN_51[507:504], _GEN_52[503:496], _GEN_53[495:32]};
  wire [447:0]      _GEN_55 = _GEN_54[447:0] | {_lastGroupMask_T[511], _GEN_49[510], _GEN_50[509:508], _GEN_51[507:504], _GEN_52[503:496], _GEN_53[495:480], _GEN_54[479:64]};
  wire [383:0]      _GEN_56 = _GEN_55[383:0] | {_lastGroupMask_T[511], _GEN_49[510], _GEN_50[509:508], _GEN_51[507:504], _GEN_52[503:496], _GEN_53[495:480], _GEN_54[479:448], _GEN_55[447:128]};
  wire [511:0]      lastGroupMask =
    {_lastGroupMask_T[511],
     _GEN_49[510],
     _GEN_50[509:508],
     _GEN_51[507:504],
     _GEN_52[503:496],
     _GEN_53[495:480],
     _GEN_54[479:448],
     _GEN_55[447:384],
     _GEN_56[383:256],
     _GEN_56[255:0] | {_lastGroupMask_T[511], _GEN_49[510], _GEN_50[509:508], _GEN_51[507:504], _GEN_52[503:496], _GEN_53[495:480], _GEN_54[479:448], _GEN_55[447:384], _GEN_56[383:256]}};
  wire [511:0]      currentMaskGroupForDestination =
    (lastGroup ? lastGroupMask : 512'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
    & (instReg_maskType & ~instReg_decodeResult_maskSource
         ? (vs1Split_vs1SetIndex ? maskForDestination_hi : maskForDestination_lo)
         : 512'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF);
  wire [63:0]       _GEN_57 = {exeReqReg_1_bits_source1, exeReqReg_0_bits_source1};
  wire [63:0]       groupSourceData_lo_lo_lo;
  assign groupSourceData_lo_lo_lo = _GEN_57;
  wire [63:0]       source1_lo_lo_lo;
  assign source1_lo_lo_lo = _GEN_57;
  wire [63:0]       _GEN_58 = {exeReqReg_3_bits_source1, exeReqReg_2_bits_source1};
  wire [63:0]       groupSourceData_lo_lo_hi;
  assign groupSourceData_lo_lo_hi = _GEN_58;
  wire [63:0]       source1_lo_lo_hi;
  assign source1_lo_lo_hi = _GEN_58;
  wire [127:0]      groupSourceData_lo_lo = {groupSourceData_lo_lo_hi, groupSourceData_lo_lo_lo};
  wire [63:0]       _GEN_59 = {exeReqReg_5_bits_source1, exeReqReg_4_bits_source1};
  wire [63:0]       groupSourceData_lo_hi_lo;
  assign groupSourceData_lo_hi_lo = _GEN_59;
  wire [63:0]       source1_lo_hi_lo;
  assign source1_lo_hi_lo = _GEN_59;
  wire [63:0]       _GEN_60 = {exeReqReg_7_bits_source1, exeReqReg_6_bits_source1};
  wire [63:0]       groupSourceData_lo_hi_hi;
  assign groupSourceData_lo_hi_hi = _GEN_60;
  wire [63:0]       source1_lo_hi_hi;
  assign source1_lo_hi_hi = _GEN_60;
  wire [127:0]      groupSourceData_lo_hi = {groupSourceData_lo_hi_hi, groupSourceData_lo_hi_lo};
  wire [255:0]      groupSourceData_lo = {groupSourceData_lo_hi, groupSourceData_lo_lo};
  wire [63:0]       _GEN_61 = {exeReqReg_9_bits_source1, exeReqReg_8_bits_source1};
  wire [63:0]       groupSourceData_hi_lo_lo;
  assign groupSourceData_hi_lo_lo = _GEN_61;
  wire [63:0]       source1_hi_lo_lo;
  assign source1_hi_lo_lo = _GEN_61;
  wire [63:0]       _GEN_62 = {exeReqReg_11_bits_source1, exeReqReg_10_bits_source1};
  wire [63:0]       groupSourceData_hi_lo_hi;
  assign groupSourceData_hi_lo_hi = _GEN_62;
  wire [63:0]       source1_hi_lo_hi;
  assign source1_hi_lo_hi = _GEN_62;
  wire [127:0]      groupSourceData_hi_lo = {groupSourceData_hi_lo_hi, groupSourceData_hi_lo_lo};
  wire [63:0]       _GEN_63 = {exeReqReg_13_bits_source1, exeReqReg_12_bits_source1};
  wire [63:0]       groupSourceData_hi_hi_lo;
  assign groupSourceData_hi_hi_lo = _GEN_63;
  wire [63:0]       source1_hi_hi_lo;
  assign source1_hi_hi_lo = _GEN_63;
  wire [63:0]       _GEN_64 = {exeReqReg_15_bits_source1, exeReqReg_14_bits_source1};
  wire [63:0]       groupSourceData_hi_hi_hi;
  assign groupSourceData_hi_hi_hi = _GEN_64;
  wire [63:0]       source1_hi_hi_hi;
  assign source1_hi_hi_hi = _GEN_64;
  wire [127:0]      groupSourceData_hi_hi = {groupSourceData_hi_hi_hi, groupSourceData_hi_hi_lo};
  wire [255:0]      groupSourceData_hi = {groupSourceData_hi_hi, groupSourceData_hi_lo};
  wire [511:0]      groupSourceData = {groupSourceData_hi, groupSourceData_lo};
  wire [1:0]        _GEN_65 = {exeReqReg_1_valid, exeReqReg_0_valid};
  wire [1:0]        groupSourceValid_lo_lo_lo;
  assign groupSourceValid_lo_lo_lo = _GEN_65;
  wire [1:0]        view__in_bits_validInput_lo_lo_lo;
  assign view__in_bits_validInput_lo_lo_lo = _GEN_65;
  wire [1:0]        view__in_bits_sourceValid_lo_lo_lo;
  assign view__in_bits_sourceValid_lo_lo_lo = _GEN_65;
  wire [1:0]        _GEN_66 = {exeReqReg_3_valid, exeReqReg_2_valid};
  wire [1:0]        groupSourceValid_lo_lo_hi;
  assign groupSourceValid_lo_lo_hi = _GEN_66;
  wire [1:0]        view__in_bits_validInput_lo_lo_hi;
  assign view__in_bits_validInput_lo_lo_hi = _GEN_66;
  wire [1:0]        view__in_bits_sourceValid_lo_lo_hi;
  assign view__in_bits_sourceValid_lo_lo_hi = _GEN_66;
  wire [3:0]        groupSourceValid_lo_lo = {groupSourceValid_lo_lo_hi, groupSourceValid_lo_lo_lo};
  wire [1:0]        _GEN_67 = {exeReqReg_5_valid, exeReqReg_4_valid};
  wire [1:0]        groupSourceValid_lo_hi_lo;
  assign groupSourceValid_lo_hi_lo = _GEN_67;
  wire [1:0]        view__in_bits_validInput_lo_hi_lo;
  assign view__in_bits_validInput_lo_hi_lo = _GEN_67;
  wire [1:0]        view__in_bits_sourceValid_lo_hi_lo;
  assign view__in_bits_sourceValid_lo_hi_lo = _GEN_67;
  wire [1:0]        _GEN_68 = {exeReqReg_7_valid, exeReqReg_6_valid};
  wire [1:0]        groupSourceValid_lo_hi_hi;
  assign groupSourceValid_lo_hi_hi = _GEN_68;
  wire [1:0]        view__in_bits_validInput_lo_hi_hi;
  assign view__in_bits_validInput_lo_hi_hi = _GEN_68;
  wire [1:0]        view__in_bits_sourceValid_lo_hi_hi;
  assign view__in_bits_sourceValid_lo_hi_hi = _GEN_68;
  wire [3:0]        groupSourceValid_lo_hi = {groupSourceValid_lo_hi_hi, groupSourceValid_lo_hi_lo};
  wire [7:0]        groupSourceValid_lo = {groupSourceValid_lo_hi, groupSourceValid_lo_lo};
  wire [1:0]        _GEN_69 = {exeReqReg_9_valid, exeReqReg_8_valid};
  wire [1:0]        groupSourceValid_hi_lo_lo;
  assign groupSourceValid_hi_lo_lo = _GEN_69;
  wire [1:0]        view__in_bits_validInput_hi_lo_lo;
  assign view__in_bits_validInput_hi_lo_lo = _GEN_69;
  wire [1:0]        view__in_bits_sourceValid_hi_lo_lo;
  assign view__in_bits_sourceValid_hi_lo_lo = _GEN_69;
  wire [1:0]        _GEN_70 = {exeReqReg_11_valid, exeReqReg_10_valid};
  wire [1:0]        groupSourceValid_hi_lo_hi;
  assign groupSourceValid_hi_lo_hi = _GEN_70;
  wire [1:0]        view__in_bits_validInput_hi_lo_hi;
  assign view__in_bits_validInput_hi_lo_hi = _GEN_70;
  wire [1:0]        view__in_bits_sourceValid_hi_lo_hi;
  assign view__in_bits_sourceValid_hi_lo_hi = _GEN_70;
  wire [3:0]        groupSourceValid_hi_lo = {groupSourceValid_hi_lo_hi, groupSourceValid_hi_lo_lo};
  wire [1:0]        _GEN_71 = {exeReqReg_13_valid, exeReqReg_12_valid};
  wire [1:0]        groupSourceValid_hi_hi_lo;
  assign groupSourceValid_hi_hi_lo = _GEN_71;
  wire [1:0]        view__in_bits_validInput_hi_hi_lo;
  assign view__in_bits_validInput_hi_hi_lo = _GEN_71;
  wire [1:0]        view__in_bits_sourceValid_hi_hi_lo;
  assign view__in_bits_sourceValid_hi_hi_lo = _GEN_71;
  wire [1:0]        _GEN_72 = {exeReqReg_15_valid, exeReqReg_14_valid};
  wire [1:0]        groupSourceValid_hi_hi_hi;
  assign groupSourceValid_hi_hi_hi = _GEN_72;
  wire [1:0]        view__in_bits_validInput_hi_hi_hi;
  assign view__in_bits_validInput_hi_hi_hi = _GEN_72;
  wire [1:0]        view__in_bits_sourceValid_hi_hi_hi;
  assign view__in_bits_sourceValid_hi_hi_hi = _GEN_72;
  wire [3:0]        groupSourceValid_hi_hi = {groupSourceValid_hi_hi_hi, groupSourceValid_hi_hi_lo};
  wire [7:0]        groupSourceValid_hi = {groupSourceValid_hi_hi, groupSourceValid_hi_lo};
  wire [15:0]       groupSourceValid = {groupSourceValid_hi, groupSourceValid_lo};
  wire [1:0]        shifterSize = (sourceDataEEW1H[0] ? executeIndex : 2'h0) | (sourceDataEEW1H[1] ? {executeIndex[1], 1'h0} : 2'h0);
  wire [3:0]        _shifterSource_T = 4'h1 << shifterSize;
  wire [511:0]      _shifterSource_T_8 = _shifterSource_T[0] ? groupSourceData : 512'h0;
  wire [383:0]      _GEN_73 = _shifterSource_T_8[383:0] | (_shifterSource_T[1] ? groupSourceData[511:128] : 384'h0);
  wire [255:0]      _GEN_74 = _GEN_73[255:0] | (_shifterSource_T[2] ? groupSourceData[511:256] : 256'h0);
  wire [511:0]      shifterSource = {_shifterSource_T_8[511:384], _GEN_73[383:256], _GEN_74[255:128], _GEN_74[127:0] | (_shifterSource_T[3] ? groupSourceData[511:384] : 128'h0)};
  wire [7:0]        selectValid_lo_lo_lo = {{4{groupSourceValid[1]}}, {4{groupSourceValid[0]}}};
  wire [7:0]        selectValid_lo_lo_hi = {{4{groupSourceValid[3]}}, {4{groupSourceValid[2]}}};
  wire [15:0]       selectValid_lo_lo = {selectValid_lo_lo_hi, selectValid_lo_lo_lo};
  wire [7:0]        selectValid_lo_hi_lo = {{4{groupSourceValid[5]}}, {4{groupSourceValid[4]}}};
  wire [7:0]        selectValid_lo_hi_hi = {{4{groupSourceValid[7]}}, {4{groupSourceValid[6]}}};
  wire [15:0]       selectValid_lo_hi = {selectValid_lo_hi_hi, selectValid_lo_hi_lo};
  wire [31:0]       selectValid_lo = {selectValid_lo_hi, selectValid_lo_lo};
  wire [7:0]        selectValid_hi_lo_lo = {{4{groupSourceValid[9]}}, {4{groupSourceValid[8]}}};
  wire [7:0]        selectValid_hi_lo_hi = {{4{groupSourceValid[11]}}, {4{groupSourceValid[10]}}};
  wire [15:0]       selectValid_hi_lo = {selectValid_hi_lo_hi, selectValid_hi_lo_lo};
  wire [7:0]        selectValid_hi_hi_lo = {{4{groupSourceValid[13]}}, {4{groupSourceValid[12]}}};
  wire [7:0]        selectValid_hi_hi_hi = {{4{groupSourceValid[15]}}, {4{groupSourceValid[14]}}};
  wire [15:0]       selectValid_hi_hi = {selectValid_hi_hi_hi, selectValid_hi_hi_lo};
  wire [31:0]       selectValid_hi = {selectValid_hi_hi, selectValid_hi_lo};
  wire [3:0]        selectValid_lo_lo_lo_1 = {{2{groupSourceValid[1]}}, {2{groupSourceValid[0]}}};
  wire [3:0]        selectValid_lo_lo_hi_1 = {{2{groupSourceValid[3]}}, {2{groupSourceValid[2]}}};
  wire [7:0]        selectValid_lo_lo_1 = {selectValid_lo_lo_hi_1, selectValid_lo_lo_lo_1};
  wire [3:0]        selectValid_lo_hi_lo_1 = {{2{groupSourceValid[5]}}, {2{groupSourceValid[4]}}};
  wire [3:0]        selectValid_lo_hi_hi_1 = {{2{groupSourceValid[7]}}, {2{groupSourceValid[6]}}};
  wire [7:0]        selectValid_lo_hi_1 = {selectValid_lo_hi_hi_1, selectValid_lo_hi_lo_1};
  wire [15:0]       selectValid_lo_1 = {selectValid_lo_hi_1, selectValid_lo_lo_1};
  wire [3:0]        selectValid_hi_lo_lo_1 = {{2{groupSourceValid[9]}}, {2{groupSourceValid[8]}}};
  wire [3:0]        selectValid_hi_lo_hi_1 = {{2{groupSourceValid[11]}}, {2{groupSourceValid[10]}}};
  wire [7:0]        selectValid_hi_lo_1 = {selectValid_hi_lo_hi_1, selectValid_hi_lo_lo_1};
  wire [3:0]        selectValid_hi_hi_lo_1 = {{2{groupSourceValid[13]}}, {2{groupSourceValid[12]}}};
  wire [3:0]        selectValid_hi_hi_hi_1 = {{2{groupSourceValid[15]}}, {2{groupSourceValid[14]}}};
  wire [7:0]        selectValid_hi_hi_1 = {selectValid_hi_hi_hi_1, selectValid_hi_hi_lo_1};
  wire [15:0]       selectValid_hi_1 = {selectValid_hi_hi_1, selectValid_hi_lo_1};
  wire [3:0][15:0]  _GEN_75 = {{selectValid_hi[31:16]}, {selectValid_hi[15:0]}, {selectValid_lo[31:16]}, {selectValid_lo[15:0]}};
  wire [15:0]       selectValid = (sourceDataEEW1H[0] ? _GEN_75[executeIndex] : 16'h0) | (sourceDataEEW1H[1] ? (executeIndex[1] ? selectValid_hi_1 : selectValid_lo_1) : 16'h0) | (sourceDataEEW1H[2] ? groupSourceValid : 16'h0);
  wire [31:0]       source_0 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[7:0] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[15:0] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[31:0] : 32'h0);
  wire [31:0]       source_1 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[15:8] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[31:16] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[63:32] : 32'h0);
  wire [31:0]       source_2 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[23:16] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[47:32] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[95:64] : 32'h0);
  wire [31:0]       source_3 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[31:24] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[63:48] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[127:96] : 32'h0);
  wire [31:0]       source_4 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[39:32] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[79:64] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[159:128] : 32'h0);
  wire [31:0]       source_5 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[47:40] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[95:80] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[191:160] : 32'h0);
  wire [31:0]       source_6 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[55:48] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[111:96] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[223:192] : 32'h0);
  wire [31:0]       source_7 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[63:56] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[127:112] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[255:224] : 32'h0);
  wire [31:0]       source_8 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[71:64] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[143:128] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[287:256] : 32'h0);
  wire [31:0]       source_9 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[79:72] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[159:144] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[319:288] : 32'h0);
  wire [31:0]       source_10 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[87:80] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[175:160] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[351:320] : 32'h0);
  wire [31:0]       source_11 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[95:88] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[191:176] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[383:352] : 32'h0);
  wire [31:0]       source_12 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[103:96] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[207:192] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[415:384] : 32'h0);
  wire [31:0]       source_13 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[111:104] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[223:208] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[447:416] : 32'h0);
  wire [31:0]       source_14 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[119:112] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[239:224] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[479:448] : 32'h0);
  wire [31:0]       source_15 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[127:120] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[255:240] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[511:480] : 32'h0);
  wire [15:0]       _GEN_76 = selectValid & readMaskCorrection;
  wire [15:0]       checkVec_validVec;
  assign checkVec_validVec = _GEN_76;
  wire [15:0]       checkVec_validVec_1;
  assign checkVec_validVec_1 = _GEN_76;
  wire [15:0]       checkVec_validVec_2;
  assign checkVec_validVec_2 = _GEN_76;
  wire              checkVec_checkResultVec_0_6 = checkVec_validVec[0];
  wire [3:0]        _GEN_77 = 4'h1 << instReg_vlmul[1:0];
  wire [3:0]        checkVec_checkResultVec_intLMULInput;
  assign checkVec_checkResultVec_intLMULInput = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_1;
  assign checkVec_checkResultVec_intLMULInput_1 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_2;
  assign checkVec_checkResultVec_intLMULInput_2 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_3;
  assign checkVec_checkResultVec_intLMULInput_3 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_4;
  assign checkVec_checkResultVec_intLMULInput_4 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_5;
  assign checkVec_checkResultVec_intLMULInput_5 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_6;
  assign checkVec_checkResultVec_intLMULInput_6 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_7;
  assign checkVec_checkResultVec_intLMULInput_7 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_8;
  assign checkVec_checkResultVec_intLMULInput_8 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_9;
  assign checkVec_checkResultVec_intLMULInput_9 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_10;
  assign checkVec_checkResultVec_intLMULInput_10 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_11;
  assign checkVec_checkResultVec_intLMULInput_11 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_12;
  assign checkVec_checkResultVec_intLMULInput_12 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_13;
  assign checkVec_checkResultVec_intLMULInput_13 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_14;
  assign checkVec_checkResultVec_intLMULInput_14 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_15;
  assign checkVec_checkResultVec_intLMULInput_15 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_16;
  assign checkVec_checkResultVec_intLMULInput_16 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_17;
  assign checkVec_checkResultVec_intLMULInput_17 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_18;
  assign checkVec_checkResultVec_intLMULInput_18 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_19;
  assign checkVec_checkResultVec_intLMULInput_19 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_20;
  assign checkVec_checkResultVec_intLMULInput_20 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_21;
  assign checkVec_checkResultVec_intLMULInput_21 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_22;
  assign checkVec_checkResultVec_intLMULInput_22 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_23;
  assign checkVec_checkResultVec_intLMULInput_23 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_24;
  assign checkVec_checkResultVec_intLMULInput_24 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_25;
  assign checkVec_checkResultVec_intLMULInput_25 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_26;
  assign checkVec_checkResultVec_intLMULInput_26 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_27;
  assign checkVec_checkResultVec_intLMULInput_27 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_28;
  assign checkVec_checkResultVec_intLMULInput_28 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_29;
  assign checkVec_checkResultVec_intLMULInput_29 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_30;
  assign checkVec_checkResultVec_intLMULInput_30 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_31;
  assign checkVec_checkResultVec_intLMULInput_31 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_32;
  assign checkVec_checkResultVec_intLMULInput_32 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_33;
  assign checkVec_checkResultVec_intLMULInput_33 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_34;
  assign checkVec_checkResultVec_intLMULInput_34 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_35;
  assign checkVec_checkResultVec_intLMULInput_35 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_36;
  assign checkVec_checkResultVec_intLMULInput_36 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_37;
  assign checkVec_checkResultVec_intLMULInput_37 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_38;
  assign checkVec_checkResultVec_intLMULInput_38 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_39;
  assign checkVec_checkResultVec_intLMULInput_39 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_40;
  assign checkVec_checkResultVec_intLMULInput_40 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_41;
  assign checkVec_checkResultVec_intLMULInput_41 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_42;
  assign checkVec_checkResultVec_intLMULInput_42 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_43;
  assign checkVec_checkResultVec_intLMULInput_43 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_44;
  assign checkVec_checkResultVec_intLMULInput_44 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_45;
  assign checkVec_checkResultVec_intLMULInput_45 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_46;
  assign checkVec_checkResultVec_intLMULInput_46 = _GEN_77;
  wire [3:0]        checkVec_checkResultVec_intLMULInput_47;
  assign checkVec_checkResultVec_intLMULInput_47 = _GEN_77;
  wire [9:0]        checkVec_checkResultVec_dataPosition = source_0[9:0];
  wire [3:0]        checkVec_checkResultVec_0_0 = 4'h1 << checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]        checkVec_checkResultVec_0_1 = checkVec_checkResultVec_dataPosition[1:0];
  wire [3:0]        checkVec_checkResultVec_0_2 = checkVec_checkResultVec_dataPosition[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup = checkVec_checkResultVec_dataPosition[9:6];
  wire              checkVec_checkResultVec_0_3 = checkVec_checkResultVec_dataGroup[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth = checkVec_checkResultVec_dataGroup[3:1];
  wire [2:0]        checkVec_checkResultVec_0_4 = checkVec_checkResultVec_accessRegGrowth;
  wire [4:0]        checkVec_checkResultVec_decimalProportion = {checkVec_checkResultVec_0_3, checkVec_checkResultVec_0_2};
  wire [2:0]        checkVec_checkResultVec_decimal = checkVec_checkResultVec_decimalProportion[4:2];
  wire              checkVec_checkResultVec_overlap =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal >= checkVec_checkResultVec_intLMULInput[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth} >= checkVec_checkResultVec_intLMULInput, source_0[31:10]};
  wire              checkVec_checkResultVec_0_5 = checkVec_checkResultVec_overlap | ~checkVec_checkResultVec_0_6;
  wire              checkVec_checkResultVec_1_6 = checkVec_validVec[1];
  wire [9:0]        checkVec_checkResultVec_dataPosition_1 = source_1[9:0];
  wire [3:0]        checkVec_checkResultVec_1_0 = 4'h1 << checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]        checkVec_checkResultVec_1_1 = checkVec_checkResultVec_dataPosition_1[1:0];
  wire [3:0]        checkVec_checkResultVec_1_2 = checkVec_checkResultVec_dataPosition_1[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_1 = checkVec_checkResultVec_dataPosition_1[9:6];
  wire              checkVec_checkResultVec_1_3 = checkVec_checkResultVec_dataGroup_1[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_1 = checkVec_checkResultVec_dataGroup_1[3:1];
  wire [2:0]        checkVec_checkResultVec_1_4 = checkVec_checkResultVec_accessRegGrowth_1;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_1 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_1_2};
  wire [2:0]        checkVec_checkResultVec_decimal_1 = checkVec_checkResultVec_decimalProportion_1[4:2];
  wire              checkVec_checkResultVec_overlap_1 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_1 >= checkVec_checkResultVec_intLMULInput_1[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_1} >= checkVec_checkResultVec_intLMULInput_1, source_1[31:10]};
  wire              checkVec_checkResultVec_1_5 = checkVec_checkResultVec_overlap_1 | ~checkVec_checkResultVec_1_6;
  wire              checkVec_checkResultVec_2_6 = checkVec_validVec[2];
  wire [9:0]        checkVec_checkResultVec_dataPosition_2 = source_2[9:0];
  wire [3:0]        checkVec_checkResultVec_2_0 = 4'h1 << checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]        checkVec_checkResultVec_2_1 = checkVec_checkResultVec_dataPosition_2[1:0];
  wire [3:0]        checkVec_checkResultVec_2_2 = checkVec_checkResultVec_dataPosition_2[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_2 = checkVec_checkResultVec_dataPosition_2[9:6];
  wire              checkVec_checkResultVec_2_3 = checkVec_checkResultVec_dataGroup_2[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_2 = checkVec_checkResultVec_dataGroup_2[3:1];
  wire [2:0]        checkVec_checkResultVec_2_4 = checkVec_checkResultVec_accessRegGrowth_2;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_2 = {checkVec_checkResultVec_2_3, checkVec_checkResultVec_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_2 = checkVec_checkResultVec_decimalProportion_2[4:2];
  wire              checkVec_checkResultVec_overlap_2 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_2 >= checkVec_checkResultVec_intLMULInput_2[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_2} >= checkVec_checkResultVec_intLMULInput_2, source_2[31:10]};
  wire              checkVec_checkResultVec_2_5 = checkVec_checkResultVec_overlap_2 | ~checkVec_checkResultVec_2_6;
  wire              checkVec_checkResultVec_3_6 = checkVec_validVec[3];
  wire [9:0]        checkVec_checkResultVec_dataPosition_3 = source_3[9:0];
  wire [3:0]        checkVec_checkResultVec_3_0 = 4'h1 << checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]        checkVec_checkResultVec_3_1 = checkVec_checkResultVec_dataPosition_3[1:0];
  wire [3:0]        checkVec_checkResultVec_3_2 = checkVec_checkResultVec_dataPosition_3[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_3 = checkVec_checkResultVec_dataPosition_3[9:6];
  wire              checkVec_checkResultVec_3_3 = checkVec_checkResultVec_dataGroup_3[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_3 = checkVec_checkResultVec_dataGroup_3[3:1];
  wire [2:0]        checkVec_checkResultVec_3_4 = checkVec_checkResultVec_accessRegGrowth_3;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_3_2};
  wire [2:0]        checkVec_checkResultVec_decimal_3 = checkVec_checkResultVec_decimalProportion_3[4:2];
  wire              checkVec_checkResultVec_overlap_3 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_3 >= checkVec_checkResultVec_intLMULInput_3[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_3} >= checkVec_checkResultVec_intLMULInput_3, source_3[31:10]};
  wire              checkVec_checkResultVec_3_5 = checkVec_checkResultVec_overlap_3 | ~checkVec_checkResultVec_3_6;
  wire              checkVec_checkResultVec_4_6 = checkVec_validVec[4];
  wire [9:0]        checkVec_checkResultVec_dataPosition_4 = source_4[9:0];
  wire [3:0]        checkVec_checkResultVec_4_0 = 4'h1 << checkVec_checkResultVec_dataPosition_4[1:0];
  wire [1:0]        checkVec_checkResultVec_4_1 = checkVec_checkResultVec_dataPosition_4[1:0];
  wire [3:0]        checkVec_checkResultVec_4_2 = checkVec_checkResultVec_dataPosition_4[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_4 = checkVec_checkResultVec_dataPosition_4[9:6];
  wire              checkVec_checkResultVec_4_3 = checkVec_checkResultVec_dataGroup_4[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_4 = checkVec_checkResultVec_dataGroup_4[3:1];
  wire [2:0]        checkVec_checkResultVec_4_4 = checkVec_checkResultVec_accessRegGrowth_4;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_4 = {checkVec_checkResultVec_4_3, checkVec_checkResultVec_4_2};
  wire [2:0]        checkVec_checkResultVec_decimal_4 = checkVec_checkResultVec_decimalProportion_4[4:2];
  wire              checkVec_checkResultVec_overlap_4 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_4 >= checkVec_checkResultVec_intLMULInput_4[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_4} >= checkVec_checkResultVec_intLMULInput_4, source_4[31:10]};
  wire              checkVec_checkResultVec_4_5 = checkVec_checkResultVec_overlap_4 | ~checkVec_checkResultVec_4_6;
  wire              checkVec_checkResultVec_5_6 = checkVec_validVec[5];
  wire [9:0]        checkVec_checkResultVec_dataPosition_5 = source_5[9:0];
  wire [3:0]        checkVec_checkResultVec_5_0 = 4'h1 << checkVec_checkResultVec_dataPosition_5[1:0];
  wire [1:0]        checkVec_checkResultVec_5_1 = checkVec_checkResultVec_dataPosition_5[1:0];
  wire [3:0]        checkVec_checkResultVec_5_2 = checkVec_checkResultVec_dataPosition_5[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_5 = checkVec_checkResultVec_dataPosition_5[9:6];
  wire              checkVec_checkResultVec_5_3 = checkVec_checkResultVec_dataGroup_5[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_5 = checkVec_checkResultVec_dataGroup_5[3:1];
  wire [2:0]        checkVec_checkResultVec_5_4 = checkVec_checkResultVec_accessRegGrowth_5;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_5 = {checkVec_checkResultVec_5_3, checkVec_checkResultVec_5_2};
  wire [2:0]        checkVec_checkResultVec_decimal_5 = checkVec_checkResultVec_decimalProportion_5[4:2];
  wire              checkVec_checkResultVec_overlap_5 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_5 >= checkVec_checkResultVec_intLMULInput_5[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_5} >= checkVec_checkResultVec_intLMULInput_5, source_5[31:10]};
  wire              checkVec_checkResultVec_5_5 = checkVec_checkResultVec_overlap_5 | ~checkVec_checkResultVec_5_6;
  wire              checkVec_checkResultVec_6_6 = checkVec_validVec[6];
  wire [9:0]        checkVec_checkResultVec_dataPosition_6 = source_6[9:0];
  wire [3:0]        checkVec_checkResultVec_6_0 = 4'h1 << checkVec_checkResultVec_dataPosition_6[1:0];
  wire [1:0]        checkVec_checkResultVec_6_1 = checkVec_checkResultVec_dataPosition_6[1:0];
  wire [3:0]        checkVec_checkResultVec_6_2 = checkVec_checkResultVec_dataPosition_6[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_6 = checkVec_checkResultVec_dataPosition_6[9:6];
  wire              checkVec_checkResultVec_6_3 = checkVec_checkResultVec_dataGroup_6[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_6 = checkVec_checkResultVec_dataGroup_6[3:1];
  wire [2:0]        checkVec_checkResultVec_6_4 = checkVec_checkResultVec_accessRegGrowth_6;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_6 = {checkVec_checkResultVec_6_3, checkVec_checkResultVec_6_2};
  wire [2:0]        checkVec_checkResultVec_decimal_6 = checkVec_checkResultVec_decimalProportion_6[4:2];
  wire              checkVec_checkResultVec_overlap_6 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_6 >= checkVec_checkResultVec_intLMULInput_6[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_6} >= checkVec_checkResultVec_intLMULInput_6, source_6[31:10]};
  wire              checkVec_checkResultVec_6_5 = checkVec_checkResultVec_overlap_6 | ~checkVec_checkResultVec_6_6;
  wire              checkVec_checkResultVec_7_6 = checkVec_validVec[7];
  wire [9:0]        checkVec_checkResultVec_dataPosition_7 = source_7[9:0];
  wire [3:0]        checkVec_checkResultVec_7_0 = 4'h1 << checkVec_checkResultVec_dataPosition_7[1:0];
  wire [1:0]        checkVec_checkResultVec_7_1 = checkVec_checkResultVec_dataPosition_7[1:0];
  wire [3:0]        checkVec_checkResultVec_7_2 = checkVec_checkResultVec_dataPosition_7[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_7 = checkVec_checkResultVec_dataPosition_7[9:6];
  wire              checkVec_checkResultVec_7_3 = checkVec_checkResultVec_dataGroup_7[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_7 = checkVec_checkResultVec_dataGroup_7[3:1];
  wire [2:0]        checkVec_checkResultVec_7_4 = checkVec_checkResultVec_accessRegGrowth_7;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_7 = {checkVec_checkResultVec_7_3, checkVec_checkResultVec_7_2};
  wire [2:0]        checkVec_checkResultVec_decimal_7 = checkVec_checkResultVec_decimalProportion_7[4:2];
  wire              checkVec_checkResultVec_overlap_7 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_7 >= checkVec_checkResultVec_intLMULInput_7[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_7} >= checkVec_checkResultVec_intLMULInput_7, source_7[31:10]};
  wire              checkVec_checkResultVec_7_5 = checkVec_checkResultVec_overlap_7 | ~checkVec_checkResultVec_7_6;
  wire              checkVec_checkResultVec_8_6 = checkVec_validVec[8];
  wire [9:0]        checkVec_checkResultVec_dataPosition_8 = source_8[9:0];
  wire [3:0]        checkVec_checkResultVec_8_0 = 4'h1 << checkVec_checkResultVec_dataPosition_8[1:0];
  wire [1:0]        checkVec_checkResultVec_8_1 = checkVec_checkResultVec_dataPosition_8[1:0];
  wire [3:0]        checkVec_checkResultVec_8_2 = checkVec_checkResultVec_dataPosition_8[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_8 = checkVec_checkResultVec_dataPosition_8[9:6];
  wire              checkVec_checkResultVec_8_3 = checkVec_checkResultVec_dataGroup_8[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_8 = checkVec_checkResultVec_dataGroup_8[3:1];
  wire [2:0]        checkVec_checkResultVec_8_4 = checkVec_checkResultVec_accessRegGrowth_8;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_8 = {checkVec_checkResultVec_8_3, checkVec_checkResultVec_8_2};
  wire [2:0]        checkVec_checkResultVec_decimal_8 = checkVec_checkResultVec_decimalProportion_8[4:2];
  wire              checkVec_checkResultVec_overlap_8 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_8 >= checkVec_checkResultVec_intLMULInput_8[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_8} >= checkVec_checkResultVec_intLMULInput_8, source_8[31:10]};
  wire              checkVec_checkResultVec_8_5 = checkVec_checkResultVec_overlap_8 | ~checkVec_checkResultVec_8_6;
  wire              checkVec_checkResultVec_9_6 = checkVec_validVec[9];
  wire [9:0]        checkVec_checkResultVec_dataPosition_9 = source_9[9:0];
  wire [3:0]        checkVec_checkResultVec_9_0 = 4'h1 << checkVec_checkResultVec_dataPosition_9[1:0];
  wire [1:0]        checkVec_checkResultVec_9_1 = checkVec_checkResultVec_dataPosition_9[1:0];
  wire [3:0]        checkVec_checkResultVec_9_2 = checkVec_checkResultVec_dataPosition_9[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_9 = checkVec_checkResultVec_dataPosition_9[9:6];
  wire              checkVec_checkResultVec_9_3 = checkVec_checkResultVec_dataGroup_9[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_9 = checkVec_checkResultVec_dataGroup_9[3:1];
  wire [2:0]        checkVec_checkResultVec_9_4 = checkVec_checkResultVec_accessRegGrowth_9;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_9 = {checkVec_checkResultVec_9_3, checkVec_checkResultVec_9_2};
  wire [2:0]        checkVec_checkResultVec_decimal_9 = checkVec_checkResultVec_decimalProportion_9[4:2];
  wire              checkVec_checkResultVec_overlap_9 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_9 >= checkVec_checkResultVec_intLMULInput_9[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_9} >= checkVec_checkResultVec_intLMULInput_9, source_9[31:10]};
  wire              checkVec_checkResultVec_9_5 = checkVec_checkResultVec_overlap_9 | ~checkVec_checkResultVec_9_6;
  wire              checkVec_checkResultVec_10_6 = checkVec_validVec[10];
  wire [9:0]        checkVec_checkResultVec_dataPosition_10 = source_10[9:0];
  wire [3:0]        checkVec_checkResultVec_10_0 = 4'h1 << checkVec_checkResultVec_dataPosition_10[1:0];
  wire [1:0]        checkVec_checkResultVec_10_1 = checkVec_checkResultVec_dataPosition_10[1:0];
  wire [3:0]        checkVec_checkResultVec_10_2 = checkVec_checkResultVec_dataPosition_10[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_10 = checkVec_checkResultVec_dataPosition_10[9:6];
  wire              checkVec_checkResultVec_10_3 = checkVec_checkResultVec_dataGroup_10[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_10 = checkVec_checkResultVec_dataGroup_10[3:1];
  wire [2:0]        checkVec_checkResultVec_10_4 = checkVec_checkResultVec_accessRegGrowth_10;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_10 = {checkVec_checkResultVec_10_3, checkVec_checkResultVec_10_2};
  wire [2:0]        checkVec_checkResultVec_decimal_10 = checkVec_checkResultVec_decimalProportion_10[4:2];
  wire              checkVec_checkResultVec_overlap_10 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_10 >= checkVec_checkResultVec_intLMULInput_10[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_10} >= checkVec_checkResultVec_intLMULInput_10,
      source_10[31:10]};
  wire              checkVec_checkResultVec_10_5 = checkVec_checkResultVec_overlap_10 | ~checkVec_checkResultVec_10_6;
  wire              checkVec_checkResultVec_11_6 = checkVec_validVec[11];
  wire [9:0]        checkVec_checkResultVec_dataPosition_11 = source_11[9:0];
  wire [3:0]        checkVec_checkResultVec_11_0 = 4'h1 << checkVec_checkResultVec_dataPosition_11[1:0];
  wire [1:0]        checkVec_checkResultVec_11_1 = checkVec_checkResultVec_dataPosition_11[1:0];
  wire [3:0]        checkVec_checkResultVec_11_2 = checkVec_checkResultVec_dataPosition_11[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_11 = checkVec_checkResultVec_dataPosition_11[9:6];
  wire              checkVec_checkResultVec_11_3 = checkVec_checkResultVec_dataGroup_11[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_11 = checkVec_checkResultVec_dataGroup_11[3:1];
  wire [2:0]        checkVec_checkResultVec_11_4 = checkVec_checkResultVec_accessRegGrowth_11;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_11 = {checkVec_checkResultVec_11_3, checkVec_checkResultVec_11_2};
  wire [2:0]        checkVec_checkResultVec_decimal_11 = checkVec_checkResultVec_decimalProportion_11[4:2];
  wire              checkVec_checkResultVec_overlap_11 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_11 >= checkVec_checkResultVec_intLMULInput_11[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_11} >= checkVec_checkResultVec_intLMULInput_11,
      source_11[31:10]};
  wire              checkVec_checkResultVec_11_5 = checkVec_checkResultVec_overlap_11 | ~checkVec_checkResultVec_11_6;
  wire              checkVec_checkResultVec_12_6 = checkVec_validVec[12];
  wire [9:0]        checkVec_checkResultVec_dataPosition_12 = source_12[9:0];
  wire [3:0]        checkVec_checkResultVec_12_0 = 4'h1 << checkVec_checkResultVec_dataPosition_12[1:0];
  wire [1:0]        checkVec_checkResultVec_12_1 = checkVec_checkResultVec_dataPosition_12[1:0];
  wire [3:0]        checkVec_checkResultVec_12_2 = checkVec_checkResultVec_dataPosition_12[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_12 = checkVec_checkResultVec_dataPosition_12[9:6];
  wire              checkVec_checkResultVec_12_3 = checkVec_checkResultVec_dataGroup_12[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_12 = checkVec_checkResultVec_dataGroup_12[3:1];
  wire [2:0]        checkVec_checkResultVec_12_4 = checkVec_checkResultVec_accessRegGrowth_12;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_12 = {checkVec_checkResultVec_12_3, checkVec_checkResultVec_12_2};
  wire [2:0]        checkVec_checkResultVec_decimal_12 = checkVec_checkResultVec_decimalProportion_12[4:2];
  wire              checkVec_checkResultVec_overlap_12 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_12 >= checkVec_checkResultVec_intLMULInput_12[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_12} >= checkVec_checkResultVec_intLMULInput_12,
      source_12[31:10]};
  wire              checkVec_checkResultVec_12_5 = checkVec_checkResultVec_overlap_12 | ~checkVec_checkResultVec_12_6;
  wire              checkVec_checkResultVec_13_6 = checkVec_validVec[13];
  wire [9:0]        checkVec_checkResultVec_dataPosition_13 = source_13[9:0];
  wire [3:0]        checkVec_checkResultVec_13_0 = 4'h1 << checkVec_checkResultVec_dataPosition_13[1:0];
  wire [1:0]        checkVec_checkResultVec_13_1 = checkVec_checkResultVec_dataPosition_13[1:0];
  wire [3:0]        checkVec_checkResultVec_13_2 = checkVec_checkResultVec_dataPosition_13[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_13 = checkVec_checkResultVec_dataPosition_13[9:6];
  wire              checkVec_checkResultVec_13_3 = checkVec_checkResultVec_dataGroup_13[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_13 = checkVec_checkResultVec_dataGroup_13[3:1];
  wire [2:0]        checkVec_checkResultVec_13_4 = checkVec_checkResultVec_accessRegGrowth_13;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_13 = {checkVec_checkResultVec_13_3, checkVec_checkResultVec_13_2};
  wire [2:0]        checkVec_checkResultVec_decimal_13 = checkVec_checkResultVec_decimalProportion_13[4:2];
  wire              checkVec_checkResultVec_overlap_13 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_13 >= checkVec_checkResultVec_intLMULInput_13[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_13} >= checkVec_checkResultVec_intLMULInput_13,
      source_13[31:10]};
  wire              checkVec_checkResultVec_13_5 = checkVec_checkResultVec_overlap_13 | ~checkVec_checkResultVec_13_6;
  wire              checkVec_checkResultVec_14_6 = checkVec_validVec[14];
  wire [9:0]        checkVec_checkResultVec_dataPosition_14 = source_14[9:0];
  wire [3:0]        checkVec_checkResultVec_14_0 = 4'h1 << checkVec_checkResultVec_dataPosition_14[1:0];
  wire [1:0]        checkVec_checkResultVec_14_1 = checkVec_checkResultVec_dataPosition_14[1:0];
  wire [3:0]        checkVec_checkResultVec_14_2 = checkVec_checkResultVec_dataPosition_14[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_14 = checkVec_checkResultVec_dataPosition_14[9:6];
  wire              checkVec_checkResultVec_14_3 = checkVec_checkResultVec_dataGroup_14[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_14 = checkVec_checkResultVec_dataGroup_14[3:1];
  wire [2:0]        checkVec_checkResultVec_14_4 = checkVec_checkResultVec_accessRegGrowth_14;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_14 = {checkVec_checkResultVec_14_3, checkVec_checkResultVec_14_2};
  wire [2:0]        checkVec_checkResultVec_decimal_14 = checkVec_checkResultVec_decimalProportion_14[4:2];
  wire              checkVec_checkResultVec_overlap_14 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_14 >= checkVec_checkResultVec_intLMULInput_14[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_14} >= checkVec_checkResultVec_intLMULInput_14,
      source_14[31:10]};
  wire              checkVec_checkResultVec_14_5 = checkVec_checkResultVec_overlap_14 | ~checkVec_checkResultVec_14_6;
  wire              checkVec_checkResultVec_15_6 = checkVec_validVec[15];
  wire [9:0]        checkVec_checkResultVec_dataPosition_15 = source_15[9:0];
  wire [3:0]        checkVec_checkResultVec_15_0 = 4'h1 << checkVec_checkResultVec_dataPosition_15[1:0];
  wire [1:0]        checkVec_checkResultVec_15_1 = checkVec_checkResultVec_dataPosition_15[1:0];
  wire [3:0]        checkVec_checkResultVec_15_2 = checkVec_checkResultVec_dataPosition_15[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_15 = checkVec_checkResultVec_dataPosition_15[9:6];
  wire              checkVec_checkResultVec_15_3 = checkVec_checkResultVec_dataGroup_15[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_15 = checkVec_checkResultVec_dataGroup_15[3:1];
  wire [2:0]        checkVec_checkResultVec_15_4 = checkVec_checkResultVec_accessRegGrowth_15;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_15 = {checkVec_checkResultVec_15_3, checkVec_checkResultVec_15_2};
  wire [2:0]        checkVec_checkResultVec_decimal_15 = checkVec_checkResultVec_decimalProportion_15[4:2];
  wire              checkVec_checkResultVec_overlap_15 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_15 >= checkVec_checkResultVec_intLMULInput_15[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_15} >= checkVec_checkResultVec_intLMULInput_15,
      source_15[31:10]};
  wire              checkVec_checkResultVec_15_5 = checkVec_checkResultVec_overlap_15 | ~checkVec_checkResultVec_15_6;
  wire [7:0]        checkVec_checkResult_lo_lo_lo = {checkVec_checkResultVec_1_0, checkVec_checkResultVec_0_0};
  wire [7:0]        checkVec_checkResult_lo_lo_hi = {checkVec_checkResultVec_3_0, checkVec_checkResultVec_2_0};
  wire [15:0]       checkVec_checkResult_lo_lo = {checkVec_checkResult_lo_lo_hi, checkVec_checkResult_lo_lo_lo};
  wire [7:0]        checkVec_checkResult_lo_hi_lo = {checkVec_checkResultVec_5_0, checkVec_checkResultVec_4_0};
  wire [7:0]        checkVec_checkResult_lo_hi_hi = {checkVec_checkResultVec_7_0, checkVec_checkResultVec_6_0};
  wire [15:0]       checkVec_checkResult_lo_hi = {checkVec_checkResult_lo_hi_hi, checkVec_checkResult_lo_hi_lo};
  wire [31:0]       checkVec_checkResult_lo = {checkVec_checkResult_lo_hi, checkVec_checkResult_lo_lo};
  wire [7:0]        checkVec_checkResult_hi_lo_lo = {checkVec_checkResultVec_9_0, checkVec_checkResultVec_8_0};
  wire [7:0]        checkVec_checkResult_hi_lo_hi = {checkVec_checkResultVec_11_0, checkVec_checkResultVec_10_0};
  wire [15:0]       checkVec_checkResult_hi_lo = {checkVec_checkResult_hi_lo_hi, checkVec_checkResult_hi_lo_lo};
  wire [7:0]        checkVec_checkResult_hi_hi_lo = {checkVec_checkResultVec_13_0, checkVec_checkResultVec_12_0};
  wire [7:0]        checkVec_checkResult_hi_hi_hi = {checkVec_checkResultVec_15_0, checkVec_checkResultVec_14_0};
  wire [15:0]       checkVec_checkResult_hi_hi = {checkVec_checkResult_hi_hi_hi, checkVec_checkResult_hi_hi_lo};
  wire [31:0]       checkVec_checkResult_hi = {checkVec_checkResult_hi_hi, checkVec_checkResult_hi_lo};
  wire [63:0]       checkVec_0_0 = {checkVec_checkResult_hi, checkVec_checkResult_lo};
  wire [3:0]        checkVec_checkResult_lo_lo_lo_1 = {checkVec_checkResultVec_1_1, checkVec_checkResultVec_0_1};
  wire [3:0]        checkVec_checkResult_lo_lo_hi_1 = {checkVec_checkResultVec_3_1, checkVec_checkResultVec_2_1};
  wire [7:0]        checkVec_checkResult_lo_lo_1 = {checkVec_checkResult_lo_lo_hi_1, checkVec_checkResult_lo_lo_lo_1};
  wire [3:0]        checkVec_checkResult_lo_hi_lo_1 = {checkVec_checkResultVec_5_1, checkVec_checkResultVec_4_1};
  wire [3:0]        checkVec_checkResult_lo_hi_hi_1 = {checkVec_checkResultVec_7_1, checkVec_checkResultVec_6_1};
  wire [7:0]        checkVec_checkResult_lo_hi_1 = {checkVec_checkResult_lo_hi_hi_1, checkVec_checkResult_lo_hi_lo_1};
  wire [15:0]       checkVec_checkResult_lo_1 = {checkVec_checkResult_lo_hi_1, checkVec_checkResult_lo_lo_1};
  wire [3:0]        checkVec_checkResult_hi_lo_lo_1 = {checkVec_checkResultVec_9_1, checkVec_checkResultVec_8_1};
  wire [3:0]        checkVec_checkResult_hi_lo_hi_1 = {checkVec_checkResultVec_11_1, checkVec_checkResultVec_10_1};
  wire [7:0]        checkVec_checkResult_hi_lo_1 = {checkVec_checkResult_hi_lo_hi_1, checkVec_checkResult_hi_lo_lo_1};
  wire [3:0]        checkVec_checkResult_hi_hi_lo_1 = {checkVec_checkResultVec_13_1, checkVec_checkResultVec_12_1};
  wire [3:0]        checkVec_checkResult_hi_hi_hi_1 = {checkVec_checkResultVec_15_1, checkVec_checkResultVec_14_1};
  wire [7:0]        checkVec_checkResult_hi_hi_1 = {checkVec_checkResult_hi_hi_hi_1, checkVec_checkResult_hi_hi_lo_1};
  wire [15:0]       checkVec_checkResult_hi_1 = {checkVec_checkResult_hi_hi_1, checkVec_checkResult_hi_lo_1};
  wire [31:0]       checkVec_0_1 = {checkVec_checkResult_hi_1, checkVec_checkResult_lo_1};
  wire [7:0]        checkVec_checkResult_lo_lo_lo_2 = {checkVec_checkResultVec_1_2, checkVec_checkResultVec_0_2};
  wire [7:0]        checkVec_checkResult_lo_lo_hi_2 = {checkVec_checkResultVec_3_2, checkVec_checkResultVec_2_2};
  wire [15:0]       checkVec_checkResult_lo_lo_2 = {checkVec_checkResult_lo_lo_hi_2, checkVec_checkResult_lo_lo_lo_2};
  wire [7:0]        checkVec_checkResult_lo_hi_lo_2 = {checkVec_checkResultVec_5_2, checkVec_checkResultVec_4_2};
  wire [7:0]        checkVec_checkResult_lo_hi_hi_2 = {checkVec_checkResultVec_7_2, checkVec_checkResultVec_6_2};
  wire [15:0]       checkVec_checkResult_lo_hi_2 = {checkVec_checkResult_lo_hi_hi_2, checkVec_checkResult_lo_hi_lo_2};
  wire [31:0]       checkVec_checkResult_lo_2 = {checkVec_checkResult_lo_hi_2, checkVec_checkResult_lo_lo_2};
  wire [7:0]        checkVec_checkResult_hi_lo_lo_2 = {checkVec_checkResultVec_9_2, checkVec_checkResultVec_8_2};
  wire [7:0]        checkVec_checkResult_hi_lo_hi_2 = {checkVec_checkResultVec_11_2, checkVec_checkResultVec_10_2};
  wire [15:0]       checkVec_checkResult_hi_lo_2 = {checkVec_checkResult_hi_lo_hi_2, checkVec_checkResult_hi_lo_lo_2};
  wire [7:0]        checkVec_checkResult_hi_hi_lo_2 = {checkVec_checkResultVec_13_2, checkVec_checkResultVec_12_2};
  wire [7:0]        checkVec_checkResult_hi_hi_hi_2 = {checkVec_checkResultVec_15_2, checkVec_checkResultVec_14_2};
  wire [15:0]       checkVec_checkResult_hi_hi_2 = {checkVec_checkResult_hi_hi_hi_2, checkVec_checkResult_hi_hi_lo_2};
  wire [31:0]       checkVec_checkResult_hi_2 = {checkVec_checkResult_hi_hi_2, checkVec_checkResult_hi_lo_2};
  wire [63:0]       checkVec_0_2 = {checkVec_checkResult_hi_2, checkVec_checkResult_lo_2};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_3 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_0_3};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_2_3};
  wire [3:0]        checkVec_checkResult_lo_lo_3 = {checkVec_checkResult_lo_lo_hi_3, checkVec_checkResult_lo_lo_lo_3};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_3 = {checkVec_checkResultVec_5_3, checkVec_checkResultVec_4_3};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_3 = {checkVec_checkResultVec_7_3, checkVec_checkResultVec_6_3};
  wire [3:0]        checkVec_checkResult_lo_hi_3 = {checkVec_checkResult_lo_hi_hi_3, checkVec_checkResult_lo_hi_lo_3};
  wire [7:0]        checkVec_checkResult_lo_3 = {checkVec_checkResult_lo_hi_3, checkVec_checkResult_lo_lo_3};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_3 = {checkVec_checkResultVec_9_3, checkVec_checkResultVec_8_3};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_3 = {checkVec_checkResultVec_11_3, checkVec_checkResultVec_10_3};
  wire [3:0]        checkVec_checkResult_hi_lo_3 = {checkVec_checkResult_hi_lo_hi_3, checkVec_checkResult_hi_lo_lo_3};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_3 = {checkVec_checkResultVec_13_3, checkVec_checkResultVec_12_3};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_3 = {checkVec_checkResultVec_15_3, checkVec_checkResultVec_14_3};
  wire [3:0]        checkVec_checkResult_hi_hi_3 = {checkVec_checkResult_hi_hi_hi_3, checkVec_checkResult_hi_hi_lo_3};
  wire [7:0]        checkVec_checkResult_hi_3 = {checkVec_checkResult_hi_hi_3, checkVec_checkResult_hi_lo_3};
  wire [15:0]       checkVec_0_3 = {checkVec_checkResult_hi_3, checkVec_checkResult_lo_3};
  wire [5:0]        checkVec_checkResult_lo_lo_lo_4 = {checkVec_checkResultVec_1_4, checkVec_checkResultVec_0_4};
  wire [5:0]        checkVec_checkResult_lo_lo_hi_4 = {checkVec_checkResultVec_3_4, checkVec_checkResultVec_2_4};
  wire [11:0]       checkVec_checkResult_lo_lo_4 = {checkVec_checkResult_lo_lo_hi_4, checkVec_checkResult_lo_lo_lo_4};
  wire [5:0]        checkVec_checkResult_lo_hi_lo_4 = {checkVec_checkResultVec_5_4, checkVec_checkResultVec_4_4};
  wire [5:0]        checkVec_checkResult_lo_hi_hi_4 = {checkVec_checkResultVec_7_4, checkVec_checkResultVec_6_4};
  wire [11:0]       checkVec_checkResult_lo_hi_4 = {checkVec_checkResult_lo_hi_hi_4, checkVec_checkResult_lo_hi_lo_4};
  wire [23:0]       checkVec_checkResult_lo_4 = {checkVec_checkResult_lo_hi_4, checkVec_checkResult_lo_lo_4};
  wire [5:0]        checkVec_checkResult_hi_lo_lo_4 = {checkVec_checkResultVec_9_4, checkVec_checkResultVec_8_4};
  wire [5:0]        checkVec_checkResult_hi_lo_hi_4 = {checkVec_checkResultVec_11_4, checkVec_checkResultVec_10_4};
  wire [11:0]       checkVec_checkResult_hi_lo_4 = {checkVec_checkResult_hi_lo_hi_4, checkVec_checkResult_hi_lo_lo_4};
  wire [5:0]        checkVec_checkResult_hi_hi_lo_4 = {checkVec_checkResultVec_13_4, checkVec_checkResultVec_12_4};
  wire [5:0]        checkVec_checkResult_hi_hi_hi_4 = {checkVec_checkResultVec_15_4, checkVec_checkResultVec_14_4};
  wire [11:0]       checkVec_checkResult_hi_hi_4 = {checkVec_checkResult_hi_hi_hi_4, checkVec_checkResult_hi_hi_lo_4};
  wire [23:0]       checkVec_checkResult_hi_4 = {checkVec_checkResult_hi_hi_4, checkVec_checkResult_hi_lo_4};
  wire [47:0]       checkVec_0_4 = {checkVec_checkResult_hi_4, checkVec_checkResult_lo_4};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_5 = {checkVec_checkResultVec_1_5, checkVec_checkResultVec_0_5};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_5 = {checkVec_checkResultVec_3_5, checkVec_checkResultVec_2_5};
  wire [3:0]        checkVec_checkResult_lo_lo_5 = {checkVec_checkResult_lo_lo_hi_5, checkVec_checkResult_lo_lo_lo_5};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_5 = {checkVec_checkResultVec_5_5, checkVec_checkResultVec_4_5};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_5 = {checkVec_checkResultVec_7_5, checkVec_checkResultVec_6_5};
  wire [3:0]        checkVec_checkResult_lo_hi_5 = {checkVec_checkResult_lo_hi_hi_5, checkVec_checkResult_lo_hi_lo_5};
  wire [7:0]        checkVec_checkResult_lo_5 = {checkVec_checkResult_lo_hi_5, checkVec_checkResult_lo_lo_5};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_5 = {checkVec_checkResultVec_9_5, checkVec_checkResultVec_8_5};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_5 = {checkVec_checkResultVec_11_5, checkVec_checkResultVec_10_5};
  wire [3:0]        checkVec_checkResult_hi_lo_5 = {checkVec_checkResult_hi_lo_hi_5, checkVec_checkResult_hi_lo_lo_5};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_5 = {checkVec_checkResultVec_13_5, checkVec_checkResultVec_12_5};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_5 = {checkVec_checkResultVec_15_5, checkVec_checkResultVec_14_5};
  wire [3:0]        checkVec_checkResult_hi_hi_5 = {checkVec_checkResult_hi_hi_hi_5, checkVec_checkResult_hi_hi_lo_5};
  wire [7:0]        checkVec_checkResult_hi_5 = {checkVec_checkResult_hi_hi_5, checkVec_checkResult_hi_lo_5};
  wire [15:0]       checkVec_0_5 = {checkVec_checkResult_hi_5, checkVec_checkResult_lo_5};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_6 = {checkVec_checkResultVec_1_6, checkVec_checkResultVec_0_6};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_6 = {checkVec_checkResultVec_3_6, checkVec_checkResultVec_2_6};
  wire [3:0]        checkVec_checkResult_lo_lo_6 = {checkVec_checkResult_lo_lo_hi_6, checkVec_checkResult_lo_lo_lo_6};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_6 = {checkVec_checkResultVec_5_6, checkVec_checkResultVec_4_6};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_6 = {checkVec_checkResultVec_7_6, checkVec_checkResultVec_6_6};
  wire [3:0]        checkVec_checkResult_lo_hi_6 = {checkVec_checkResult_lo_hi_hi_6, checkVec_checkResult_lo_hi_lo_6};
  wire [7:0]        checkVec_checkResult_lo_6 = {checkVec_checkResult_lo_hi_6, checkVec_checkResult_lo_lo_6};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_6 = {checkVec_checkResultVec_9_6, checkVec_checkResultVec_8_6};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_6 = {checkVec_checkResultVec_11_6, checkVec_checkResultVec_10_6};
  wire [3:0]        checkVec_checkResult_hi_lo_6 = {checkVec_checkResult_hi_lo_hi_6, checkVec_checkResult_hi_lo_lo_6};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_6 = {checkVec_checkResultVec_13_6, checkVec_checkResultVec_12_6};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_6 = {checkVec_checkResultVec_15_6, checkVec_checkResultVec_14_6};
  wire [3:0]        checkVec_checkResult_hi_hi_6 = {checkVec_checkResult_hi_hi_hi_6, checkVec_checkResult_hi_hi_lo_6};
  wire [7:0]        checkVec_checkResult_hi_6 = {checkVec_checkResult_hi_hi_6, checkVec_checkResult_hi_lo_6};
  wire [15:0]       checkVec_0_6 = {checkVec_checkResult_hi_6, checkVec_checkResult_lo_6};
  wire              checkVec_checkResultVec_0_6_1 = checkVec_validVec_1[0];
  wire [9:0]        checkVec_checkResultVec_dataPosition_16 = {source_0[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_131 = 2'h1 << checkVec_checkResultVec_dataPosition_16[1];
  wire [3:0]        checkVec_checkResultVec_0_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_131[1]}}, {2{_checkVec_checkResultVec_accessMask_T_131[0]}}};
  wire [1:0]        checkVec_checkResultVec_0_1_1 = {checkVec_checkResultVec_dataPosition_16[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_0_2_1 = checkVec_checkResultVec_dataPosition_16[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_16 = checkVec_checkResultVec_dataPosition_16[9:6];
  wire              checkVec_checkResultVec_0_3_1 = checkVec_checkResultVec_dataGroup_16[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_16 = checkVec_checkResultVec_dataGroup_16[3:1];
  wire [2:0]        checkVec_checkResultVec_0_4_1 = checkVec_checkResultVec_accessRegGrowth_16;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_16 = {checkVec_checkResultVec_0_3_1, checkVec_checkResultVec_0_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_16 = checkVec_checkResultVec_decimalProportion_16[4:2];
  wire              checkVec_checkResultVec_overlap_16 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_16 >= checkVec_checkResultVec_intLMULInput_16[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_16} >= checkVec_checkResultVec_intLMULInput_16,
      source_0[31:10]};
  wire              checkVec_checkResultVec_0_5_1 = checkVec_checkResultVec_overlap_16 | ~checkVec_checkResultVec_0_6_1;
  wire              checkVec_checkResultVec_1_6_1 = checkVec_validVec_1[1];
  wire [9:0]        checkVec_checkResultVec_dataPosition_17 = {source_1[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_139 = 2'h1 << checkVec_checkResultVec_dataPosition_17[1];
  wire [3:0]        checkVec_checkResultVec_1_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_139[1]}}, {2{_checkVec_checkResultVec_accessMask_T_139[0]}}};
  wire [1:0]        checkVec_checkResultVec_1_1_1 = {checkVec_checkResultVec_dataPosition_17[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_1_2_1 = checkVec_checkResultVec_dataPosition_17[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_17 = checkVec_checkResultVec_dataPosition_17[9:6];
  wire              checkVec_checkResultVec_1_3_1 = checkVec_checkResultVec_dataGroup_17[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_17 = checkVec_checkResultVec_dataGroup_17[3:1];
  wire [2:0]        checkVec_checkResultVec_1_4_1 = checkVec_checkResultVec_accessRegGrowth_17;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_17 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_1_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_17 = checkVec_checkResultVec_decimalProportion_17[4:2];
  wire              checkVec_checkResultVec_overlap_17 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_17 >= checkVec_checkResultVec_intLMULInput_17[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_17} >= checkVec_checkResultVec_intLMULInput_17,
      source_1[31:10]};
  wire              checkVec_checkResultVec_1_5_1 = checkVec_checkResultVec_overlap_17 | ~checkVec_checkResultVec_1_6_1;
  wire              checkVec_checkResultVec_2_6_1 = checkVec_validVec_1[2];
  wire [9:0]        checkVec_checkResultVec_dataPosition_18 = {source_2[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_147 = 2'h1 << checkVec_checkResultVec_dataPosition_18[1];
  wire [3:0]        checkVec_checkResultVec_2_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_147[1]}}, {2{_checkVec_checkResultVec_accessMask_T_147[0]}}};
  wire [1:0]        checkVec_checkResultVec_2_1_1 = {checkVec_checkResultVec_dataPosition_18[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_2_2_1 = checkVec_checkResultVec_dataPosition_18[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_18 = checkVec_checkResultVec_dataPosition_18[9:6];
  wire              checkVec_checkResultVec_2_3_1 = checkVec_checkResultVec_dataGroup_18[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_18 = checkVec_checkResultVec_dataGroup_18[3:1];
  wire [2:0]        checkVec_checkResultVec_2_4_1 = checkVec_checkResultVec_accessRegGrowth_18;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_18 = {checkVec_checkResultVec_2_3_1, checkVec_checkResultVec_2_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_18 = checkVec_checkResultVec_decimalProportion_18[4:2];
  wire              checkVec_checkResultVec_overlap_18 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_18 >= checkVec_checkResultVec_intLMULInput_18[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_18} >= checkVec_checkResultVec_intLMULInput_18,
      source_2[31:10]};
  wire              checkVec_checkResultVec_2_5_1 = checkVec_checkResultVec_overlap_18 | ~checkVec_checkResultVec_2_6_1;
  wire              checkVec_checkResultVec_3_6_1 = checkVec_validVec_1[3];
  wire [9:0]        checkVec_checkResultVec_dataPosition_19 = {source_3[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_155 = 2'h1 << checkVec_checkResultVec_dataPosition_19[1];
  wire [3:0]        checkVec_checkResultVec_3_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_155[1]}}, {2{_checkVec_checkResultVec_accessMask_T_155[0]}}};
  wire [1:0]        checkVec_checkResultVec_3_1_1 = {checkVec_checkResultVec_dataPosition_19[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_3_2_1 = checkVec_checkResultVec_dataPosition_19[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_19 = checkVec_checkResultVec_dataPosition_19[9:6];
  wire              checkVec_checkResultVec_3_3_1 = checkVec_checkResultVec_dataGroup_19[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_19 = checkVec_checkResultVec_dataGroup_19[3:1];
  wire [2:0]        checkVec_checkResultVec_3_4_1 = checkVec_checkResultVec_accessRegGrowth_19;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_19 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_3_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_19 = checkVec_checkResultVec_decimalProportion_19[4:2];
  wire              checkVec_checkResultVec_overlap_19 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_19 >= checkVec_checkResultVec_intLMULInput_19[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_19} >= checkVec_checkResultVec_intLMULInput_19,
      source_3[31:10]};
  wire              checkVec_checkResultVec_3_5_1 = checkVec_checkResultVec_overlap_19 | ~checkVec_checkResultVec_3_6_1;
  wire              checkVec_checkResultVec_4_6_1 = checkVec_validVec_1[4];
  wire [9:0]        checkVec_checkResultVec_dataPosition_20 = {source_4[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_163 = 2'h1 << checkVec_checkResultVec_dataPosition_20[1];
  wire [3:0]        checkVec_checkResultVec_4_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_163[1]}}, {2{_checkVec_checkResultVec_accessMask_T_163[0]}}};
  wire [1:0]        checkVec_checkResultVec_4_1_1 = {checkVec_checkResultVec_dataPosition_20[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_4_2_1 = checkVec_checkResultVec_dataPosition_20[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_20 = checkVec_checkResultVec_dataPosition_20[9:6];
  wire              checkVec_checkResultVec_4_3_1 = checkVec_checkResultVec_dataGroup_20[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_20 = checkVec_checkResultVec_dataGroup_20[3:1];
  wire [2:0]        checkVec_checkResultVec_4_4_1 = checkVec_checkResultVec_accessRegGrowth_20;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_20 = {checkVec_checkResultVec_4_3_1, checkVec_checkResultVec_4_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_20 = checkVec_checkResultVec_decimalProportion_20[4:2];
  wire              checkVec_checkResultVec_overlap_20 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_20 >= checkVec_checkResultVec_intLMULInput_20[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_20} >= checkVec_checkResultVec_intLMULInput_20,
      source_4[31:10]};
  wire              checkVec_checkResultVec_4_5_1 = checkVec_checkResultVec_overlap_20 | ~checkVec_checkResultVec_4_6_1;
  wire              checkVec_checkResultVec_5_6_1 = checkVec_validVec_1[5];
  wire [9:0]        checkVec_checkResultVec_dataPosition_21 = {source_5[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_171 = 2'h1 << checkVec_checkResultVec_dataPosition_21[1];
  wire [3:0]        checkVec_checkResultVec_5_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_171[1]}}, {2{_checkVec_checkResultVec_accessMask_T_171[0]}}};
  wire [1:0]        checkVec_checkResultVec_5_1_1 = {checkVec_checkResultVec_dataPosition_21[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_5_2_1 = checkVec_checkResultVec_dataPosition_21[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_21 = checkVec_checkResultVec_dataPosition_21[9:6];
  wire              checkVec_checkResultVec_5_3_1 = checkVec_checkResultVec_dataGroup_21[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_21 = checkVec_checkResultVec_dataGroup_21[3:1];
  wire [2:0]        checkVec_checkResultVec_5_4_1 = checkVec_checkResultVec_accessRegGrowth_21;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_21 = {checkVec_checkResultVec_5_3_1, checkVec_checkResultVec_5_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_21 = checkVec_checkResultVec_decimalProportion_21[4:2];
  wire              checkVec_checkResultVec_overlap_21 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_21 >= checkVec_checkResultVec_intLMULInput_21[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_21} >= checkVec_checkResultVec_intLMULInput_21,
      source_5[31:10]};
  wire              checkVec_checkResultVec_5_5_1 = checkVec_checkResultVec_overlap_21 | ~checkVec_checkResultVec_5_6_1;
  wire              checkVec_checkResultVec_6_6_1 = checkVec_validVec_1[6];
  wire [9:0]        checkVec_checkResultVec_dataPosition_22 = {source_6[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_179 = 2'h1 << checkVec_checkResultVec_dataPosition_22[1];
  wire [3:0]        checkVec_checkResultVec_6_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_179[1]}}, {2{_checkVec_checkResultVec_accessMask_T_179[0]}}};
  wire [1:0]        checkVec_checkResultVec_6_1_1 = {checkVec_checkResultVec_dataPosition_22[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_6_2_1 = checkVec_checkResultVec_dataPosition_22[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_22 = checkVec_checkResultVec_dataPosition_22[9:6];
  wire              checkVec_checkResultVec_6_3_1 = checkVec_checkResultVec_dataGroup_22[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_22 = checkVec_checkResultVec_dataGroup_22[3:1];
  wire [2:0]        checkVec_checkResultVec_6_4_1 = checkVec_checkResultVec_accessRegGrowth_22;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_22 = {checkVec_checkResultVec_6_3_1, checkVec_checkResultVec_6_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_22 = checkVec_checkResultVec_decimalProportion_22[4:2];
  wire              checkVec_checkResultVec_overlap_22 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_22 >= checkVec_checkResultVec_intLMULInput_22[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_22} >= checkVec_checkResultVec_intLMULInput_22,
      source_6[31:10]};
  wire              checkVec_checkResultVec_6_5_1 = checkVec_checkResultVec_overlap_22 | ~checkVec_checkResultVec_6_6_1;
  wire              checkVec_checkResultVec_7_6_1 = checkVec_validVec_1[7];
  wire [9:0]        checkVec_checkResultVec_dataPosition_23 = {source_7[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_187 = 2'h1 << checkVec_checkResultVec_dataPosition_23[1];
  wire [3:0]        checkVec_checkResultVec_7_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_187[1]}}, {2{_checkVec_checkResultVec_accessMask_T_187[0]}}};
  wire [1:0]        checkVec_checkResultVec_7_1_1 = {checkVec_checkResultVec_dataPosition_23[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_7_2_1 = checkVec_checkResultVec_dataPosition_23[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_23 = checkVec_checkResultVec_dataPosition_23[9:6];
  wire              checkVec_checkResultVec_7_3_1 = checkVec_checkResultVec_dataGroup_23[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_23 = checkVec_checkResultVec_dataGroup_23[3:1];
  wire [2:0]        checkVec_checkResultVec_7_4_1 = checkVec_checkResultVec_accessRegGrowth_23;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_23 = {checkVec_checkResultVec_7_3_1, checkVec_checkResultVec_7_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_23 = checkVec_checkResultVec_decimalProportion_23[4:2];
  wire              checkVec_checkResultVec_overlap_23 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_23 >= checkVec_checkResultVec_intLMULInput_23[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_23} >= checkVec_checkResultVec_intLMULInput_23,
      source_7[31:10]};
  wire              checkVec_checkResultVec_7_5_1 = checkVec_checkResultVec_overlap_23 | ~checkVec_checkResultVec_7_6_1;
  wire              checkVec_checkResultVec_8_6_1 = checkVec_validVec_1[8];
  wire [9:0]        checkVec_checkResultVec_dataPosition_24 = {source_8[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_195 = 2'h1 << checkVec_checkResultVec_dataPosition_24[1];
  wire [3:0]        checkVec_checkResultVec_8_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_195[1]}}, {2{_checkVec_checkResultVec_accessMask_T_195[0]}}};
  wire [1:0]        checkVec_checkResultVec_8_1_1 = {checkVec_checkResultVec_dataPosition_24[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_8_2_1 = checkVec_checkResultVec_dataPosition_24[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_24 = checkVec_checkResultVec_dataPosition_24[9:6];
  wire              checkVec_checkResultVec_8_3_1 = checkVec_checkResultVec_dataGroup_24[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_24 = checkVec_checkResultVec_dataGroup_24[3:1];
  wire [2:0]        checkVec_checkResultVec_8_4_1 = checkVec_checkResultVec_accessRegGrowth_24;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_24 = {checkVec_checkResultVec_8_3_1, checkVec_checkResultVec_8_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_24 = checkVec_checkResultVec_decimalProportion_24[4:2];
  wire              checkVec_checkResultVec_overlap_24 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_24 >= checkVec_checkResultVec_intLMULInput_24[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_24} >= checkVec_checkResultVec_intLMULInput_24,
      source_8[31:10]};
  wire              checkVec_checkResultVec_8_5_1 = checkVec_checkResultVec_overlap_24 | ~checkVec_checkResultVec_8_6_1;
  wire              checkVec_checkResultVec_9_6_1 = checkVec_validVec_1[9];
  wire [9:0]        checkVec_checkResultVec_dataPosition_25 = {source_9[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_203 = 2'h1 << checkVec_checkResultVec_dataPosition_25[1];
  wire [3:0]        checkVec_checkResultVec_9_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_203[1]}}, {2{_checkVec_checkResultVec_accessMask_T_203[0]}}};
  wire [1:0]        checkVec_checkResultVec_9_1_1 = {checkVec_checkResultVec_dataPosition_25[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_9_2_1 = checkVec_checkResultVec_dataPosition_25[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_25 = checkVec_checkResultVec_dataPosition_25[9:6];
  wire              checkVec_checkResultVec_9_3_1 = checkVec_checkResultVec_dataGroup_25[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_25 = checkVec_checkResultVec_dataGroup_25[3:1];
  wire [2:0]        checkVec_checkResultVec_9_4_1 = checkVec_checkResultVec_accessRegGrowth_25;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_25 = {checkVec_checkResultVec_9_3_1, checkVec_checkResultVec_9_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_25 = checkVec_checkResultVec_decimalProportion_25[4:2];
  wire              checkVec_checkResultVec_overlap_25 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_25 >= checkVec_checkResultVec_intLMULInput_25[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_25} >= checkVec_checkResultVec_intLMULInput_25,
      source_9[31:10]};
  wire              checkVec_checkResultVec_9_5_1 = checkVec_checkResultVec_overlap_25 | ~checkVec_checkResultVec_9_6_1;
  wire              checkVec_checkResultVec_10_6_1 = checkVec_validVec_1[10];
  wire [9:0]        checkVec_checkResultVec_dataPosition_26 = {source_10[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_211 = 2'h1 << checkVec_checkResultVec_dataPosition_26[1];
  wire [3:0]        checkVec_checkResultVec_10_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_211[1]}}, {2{_checkVec_checkResultVec_accessMask_T_211[0]}}};
  wire [1:0]        checkVec_checkResultVec_10_1_1 = {checkVec_checkResultVec_dataPosition_26[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_10_2_1 = checkVec_checkResultVec_dataPosition_26[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_26 = checkVec_checkResultVec_dataPosition_26[9:6];
  wire              checkVec_checkResultVec_10_3_1 = checkVec_checkResultVec_dataGroup_26[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_26 = checkVec_checkResultVec_dataGroup_26[3:1];
  wire [2:0]        checkVec_checkResultVec_10_4_1 = checkVec_checkResultVec_accessRegGrowth_26;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_26 = {checkVec_checkResultVec_10_3_1, checkVec_checkResultVec_10_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_26 = checkVec_checkResultVec_decimalProportion_26[4:2];
  wire              checkVec_checkResultVec_overlap_26 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_26 >= checkVec_checkResultVec_intLMULInput_26[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_26} >= checkVec_checkResultVec_intLMULInput_26,
      source_10[31:10]};
  wire              checkVec_checkResultVec_10_5_1 = checkVec_checkResultVec_overlap_26 | ~checkVec_checkResultVec_10_6_1;
  wire              checkVec_checkResultVec_11_6_1 = checkVec_validVec_1[11];
  wire [9:0]        checkVec_checkResultVec_dataPosition_27 = {source_11[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_219 = 2'h1 << checkVec_checkResultVec_dataPosition_27[1];
  wire [3:0]        checkVec_checkResultVec_11_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_219[1]}}, {2{_checkVec_checkResultVec_accessMask_T_219[0]}}};
  wire [1:0]        checkVec_checkResultVec_11_1_1 = {checkVec_checkResultVec_dataPosition_27[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_11_2_1 = checkVec_checkResultVec_dataPosition_27[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_27 = checkVec_checkResultVec_dataPosition_27[9:6];
  wire              checkVec_checkResultVec_11_3_1 = checkVec_checkResultVec_dataGroup_27[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_27 = checkVec_checkResultVec_dataGroup_27[3:1];
  wire [2:0]        checkVec_checkResultVec_11_4_1 = checkVec_checkResultVec_accessRegGrowth_27;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_27 = {checkVec_checkResultVec_11_3_1, checkVec_checkResultVec_11_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_27 = checkVec_checkResultVec_decimalProportion_27[4:2];
  wire              checkVec_checkResultVec_overlap_27 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_27 >= checkVec_checkResultVec_intLMULInput_27[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_27} >= checkVec_checkResultVec_intLMULInput_27,
      source_11[31:10]};
  wire              checkVec_checkResultVec_11_5_1 = checkVec_checkResultVec_overlap_27 | ~checkVec_checkResultVec_11_6_1;
  wire              checkVec_checkResultVec_12_6_1 = checkVec_validVec_1[12];
  wire [9:0]        checkVec_checkResultVec_dataPosition_28 = {source_12[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_227 = 2'h1 << checkVec_checkResultVec_dataPosition_28[1];
  wire [3:0]        checkVec_checkResultVec_12_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_227[1]}}, {2{_checkVec_checkResultVec_accessMask_T_227[0]}}};
  wire [1:0]        checkVec_checkResultVec_12_1_1 = {checkVec_checkResultVec_dataPosition_28[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_12_2_1 = checkVec_checkResultVec_dataPosition_28[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_28 = checkVec_checkResultVec_dataPosition_28[9:6];
  wire              checkVec_checkResultVec_12_3_1 = checkVec_checkResultVec_dataGroup_28[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_28 = checkVec_checkResultVec_dataGroup_28[3:1];
  wire [2:0]        checkVec_checkResultVec_12_4_1 = checkVec_checkResultVec_accessRegGrowth_28;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_28 = {checkVec_checkResultVec_12_3_1, checkVec_checkResultVec_12_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_28 = checkVec_checkResultVec_decimalProportion_28[4:2];
  wire              checkVec_checkResultVec_overlap_28 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_28 >= checkVec_checkResultVec_intLMULInput_28[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_28} >= checkVec_checkResultVec_intLMULInput_28,
      source_12[31:10]};
  wire              checkVec_checkResultVec_12_5_1 = checkVec_checkResultVec_overlap_28 | ~checkVec_checkResultVec_12_6_1;
  wire              checkVec_checkResultVec_13_6_1 = checkVec_validVec_1[13];
  wire [9:0]        checkVec_checkResultVec_dataPosition_29 = {source_13[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_235 = 2'h1 << checkVec_checkResultVec_dataPosition_29[1];
  wire [3:0]        checkVec_checkResultVec_13_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_235[1]}}, {2{_checkVec_checkResultVec_accessMask_T_235[0]}}};
  wire [1:0]        checkVec_checkResultVec_13_1_1 = {checkVec_checkResultVec_dataPosition_29[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_13_2_1 = checkVec_checkResultVec_dataPosition_29[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_29 = checkVec_checkResultVec_dataPosition_29[9:6];
  wire              checkVec_checkResultVec_13_3_1 = checkVec_checkResultVec_dataGroup_29[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_29 = checkVec_checkResultVec_dataGroup_29[3:1];
  wire [2:0]        checkVec_checkResultVec_13_4_1 = checkVec_checkResultVec_accessRegGrowth_29;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_29 = {checkVec_checkResultVec_13_3_1, checkVec_checkResultVec_13_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_29 = checkVec_checkResultVec_decimalProportion_29[4:2];
  wire              checkVec_checkResultVec_overlap_29 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_29 >= checkVec_checkResultVec_intLMULInput_29[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_29} >= checkVec_checkResultVec_intLMULInput_29,
      source_13[31:10]};
  wire              checkVec_checkResultVec_13_5_1 = checkVec_checkResultVec_overlap_29 | ~checkVec_checkResultVec_13_6_1;
  wire              checkVec_checkResultVec_14_6_1 = checkVec_validVec_1[14];
  wire [9:0]        checkVec_checkResultVec_dataPosition_30 = {source_14[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_243 = 2'h1 << checkVec_checkResultVec_dataPosition_30[1];
  wire [3:0]        checkVec_checkResultVec_14_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_243[1]}}, {2{_checkVec_checkResultVec_accessMask_T_243[0]}}};
  wire [1:0]        checkVec_checkResultVec_14_1_1 = {checkVec_checkResultVec_dataPosition_30[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_14_2_1 = checkVec_checkResultVec_dataPosition_30[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_30 = checkVec_checkResultVec_dataPosition_30[9:6];
  wire              checkVec_checkResultVec_14_3_1 = checkVec_checkResultVec_dataGroup_30[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_30 = checkVec_checkResultVec_dataGroup_30[3:1];
  wire [2:0]        checkVec_checkResultVec_14_4_1 = checkVec_checkResultVec_accessRegGrowth_30;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_30 = {checkVec_checkResultVec_14_3_1, checkVec_checkResultVec_14_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_30 = checkVec_checkResultVec_decimalProportion_30[4:2];
  wire              checkVec_checkResultVec_overlap_30 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_30 >= checkVec_checkResultVec_intLMULInput_30[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_30} >= checkVec_checkResultVec_intLMULInput_30,
      source_14[31:10]};
  wire              checkVec_checkResultVec_14_5_1 = checkVec_checkResultVec_overlap_30 | ~checkVec_checkResultVec_14_6_1;
  wire              checkVec_checkResultVec_15_6_1 = checkVec_validVec_1[15];
  wire [9:0]        checkVec_checkResultVec_dataPosition_31 = {source_15[8:0], 1'h0};
  wire [1:0]        _checkVec_checkResultVec_accessMask_T_251 = 2'h1 << checkVec_checkResultVec_dataPosition_31[1];
  wire [3:0]        checkVec_checkResultVec_15_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_251[1]}}, {2{_checkVec_checkResultVec_accessMask_T_251[0]}}};
  wire [1:0]        checkVec_checkResultVec_15_1_1 = {checkVec_checkResultVec_dataPosition_31[1], 1'h0};
  wire [3:0]        checkVec_checkResultVec_15_2_1 = checkVec_checkResultVec_dataPosition_31[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_31 = checkVec_checkResultVec_dataPosition_31[9:6];
  wire              checkVec_checkResultVec_15_3_1 = checkVec_checkResultVec_dataGroup_31[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_31 = checkVec_checkResultVec_dataGroup_31[3:1];
  wire [2:0]        checkVec_checkResultVec_15_4_1 = checkVec_checkResultVec_accessRegGrowth_31;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_31 = {checkVec_checkResultVec_15_3_1, checkVec_checkResultVec_15_2_1};
  wire [2:0]        checkVec_checkResultVec_decimal_31 = checkVec_checkResultVec_decimalProportion_31[4:2];
  wire              checkVec_checkResultVec_overlap_31 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_31 >= checkVec_checkResultVec_intLMULInput_31[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_31} >= checkVec_checkResultVec_intLMULInput_31,
      source_15[31:10]};
  wire              checkVec_checkResultVec_15_5_1 = checkVec_checkResultVec_overlap_31 | ~checkVec_checkResultVec_15_6_1;
  wire [7:0]        checkVec_checkResult_lo_lo_lo_7 = {checkVec_checkResultVec_1_0_1, checkVec_checkResultVec_0_0_1};
  wire [7:0]        checkVec_checkResult_lo_lo_hi_7 = {checkVec_checkResultVec_3_0_1, checkVec_checkResultVec_2_0_1};
  wire [15:0]       checkVec_checkResult_lo_lo_7 = {checkVec_checkResult_lo_lo_hi_7, checkVec_checkResult_lo_lo_lo_7};
  wire [7:0]        checkVec_checkResult_lo_hi_lo_7 = {checkVec_checkResultVec_5_0_1, checkVec_checkResultVec_4_0_1};
  wire [7:0]        checkVec_checkResult_lo_hi_hi_7 = {checkVec_checkResultVec_7_0_1, checkVec_checkResultVec_6_0_1};
  wire [15:0]       checkVec_checkResult_lo_hi_7 = {checkVec_checkResult_lo_hi_hi_7, checkVec_checkResult_lo_hi_lo_7};
  wire [31:0]       checkVec_checkResult_lo_7 = {checkVec_checkResult_lo_hi_7, checkVec_checkResult_lo_lo_7};
  wire [7:0]        checkVec_checkResult_hi_lo_lo_7 = {checkVec_checkResultVec_9_0_1, checkVec_checkResultVec_8_0_1};
  wire [7:0]        checkVec_checkResult_hi_lo_hi_7 = {checkVec_checkResultVec_11_0_1, checkVec_checkResultVec_10_0_1};
  wire [15:0]       checkVec_checkResult_hi_lo_7 = {checkVec_checkResult_hi_lo_hi_7, checkVec_checkResult_hi_lo_lo_7};
  wire [7:0]        checkVec_checkResult_hi_hi_lo_7 = {checkVec_checkResultVec_13_0_1, checkVec_checkResultVec_12_0_1};
  wire [7:0]        checkVec_checkResult_hi_hi_hi_7 = {checkVec_checkResultVec_15_0_1, checkVec_checkResultVec_14_0_1};
  wire [15:0]       checkVec_checkResult_hi_hi_7 = {checkVec_checkResult_hi_hi_hi_7, checkVec_checkResult_hi_hi_lo_7};
  wire [31:0]       checkVec_checkResult_hi_7 = {checkVec_checkResult_hi_hi_7, checkVec_checkResult_hi_lo_7};
  wire [63:0]       checkVec_1_0 = {checkVec_checkResult_hi_7, checkVec_checkResult_lo_7};
  wire [3:0]        checkVec_checkResult_lo_lo_lo_8 = {checkVec_checkResultVec_1_1_1, checkVec_checkResultVec_0_1_1};
  wire [3:0]        checkVec_checkResult_lo_lo_hi_8 = {checkVec_checkResultVec_3_1_1, checkVec_checkResultVec_2_1_1};
  wire [7:0]        checkVec_checkResult_lo_lo_8 = {checkVec_checkResult_lo_lo_hi_8, checkVec_checkResult_lo_lo_lo_8};
  wire [3:0]        checkVec_checkResult_lo_hi_lo_8 = {checkVec_checkResultVec_5_1_1, checkVec_checkResultVec_4_1_1};
  wire [3:0]        checkVec_checkResult_lo_hi_hi_8 = {checkVec_checkResultVec_7_1_1, checkVec_checkResultVec_6_1_1};
  wire [7:0]        checkVec_checkResult_lo_hi_8 = {checkVec_checkResult_lo_hi_hi_8, checkVec_checkResult_lo_hi_lo_8};
  wire [15:0]       checkVec_checkResult_lo_8 = {checkVec_checkResult_lo_hi_8, checkVec_checkResult_lo_lo_8};
  wire [3:0]        checkVec_checkResult_hi_lo_lo_8 = {checkVec_checkResultVec_9_1_1, checkVec_checkResultVec_8_1_1};
  wire [3:0]        checkVec_checkResult_hi_lo_hi_8 = {checkVec_checkResultVec_11_1_1, checkVec_checkResultVec_10_1_1};
  wire [7:0]        checkVec_checkResult_hi_lo_8 = {checkVec_checkResult_hi_lo_hi_8, checkVec_checkResult_hi_lo_lo_8};
  wire [3:0]        checkVec_checkResult_hi_hi_lo_8 = {checkVec_checkResultVec_13_1_1, checkVec_checkResultVec_12_1_1};
  wire [3:0]        checkVec_checkResult_hi_hi_hi_8 = {checkVec_checkResultVec_15_1_1, checkVec_checkResultVec_14_1_1};
  wire [7:0]        checkVec_checkResult_hi_hi_8 = {checkVec_checkResult_hi_hi_hi_8, checkVec_checkResult_hi_hi_lo_8};
  wire [15:0]       checkVec_checkResult_hi_8 = {checkVec_checkResult_hi_hi_8, checkVec_checkResult_hi_lo_8};
  wire [31:0]       checkVec_1_1 = {checkVec_checkResult_hi_8, checkVec_checkResult_lo_8};
  wire [7:0]        checkVec_checkResult_lo_lo_lo_9 = {checkVec_checkResultVec_1_2_1, checkVec_checkResultVec_0_2_1};
  wire [7:0]        checkVec_checkResult_lo_lo_hi_9 = {checkVec_checkResultVec_3_2_1, checkVec_checkResultVec_2_2_1};
  wire [15:0]       checkVec_checkResult_lo_lo_9 = {checkVec_checkResult_lo_lo_hi_9, checkVec_checkResult_lo_lo_lo_9};
  wire [7:0]        checkVec_checkResult_lo_hi_lo_9 = {checkVec_checkResultVec_5_2_1, checkVec_checkResultVec_4_2_1};
  wire [7:0]        checkVec_checkResult_lo_hi_hi_9 = {checkVec_checkResultVec_7_2_1, checkVec_checkResultVec_6_2_1};
  wire [15:0]       checkVec_checkResult_lo_hi_9 = {checkVec_checkResult_lo_hi_hi_9, checkVec_checkResult_lo_hi_lo_9};
  wire [31:0]       checkVec_checkResult_lo_9 = {checkVec_checkResult_lo_hi_9, checkVec_checkResult_lo_lo_9};
  wire [7:0]        checkVec_checkResult_hi_lo_lo_9 = {checkVec_checkResultVec_9_2_1, checkVec_checkResultVec_8_2_1};
  wire [7:0]        checkVec_checkResult_hi_lo_hi_9 = {checkVec_checkResultVec_11_2_1, checkVec_checkResultVec_10_2_1};
  wire [15:0]       checkVec_checkResult_hi_lo_9 = {checkVec_checkResult_hi_lo_hi_9, checkVec_checkResult_hi_lo_lo_9};
  wire [7:0]        checkVec_checkResult_hi_hi_lo_9 = {checkVec_checkResultVec_13_2_1, checkVec_checkResultVec_12_2_1};
  wire [7:0]        checkVec_checkResult_hi_hi_hi_9 = {checkVec_checkResultVec_15_2_1, checkVec_checkResultVec_14_2_1};
  wire [15:0]       checkVec_checkResult_hi_hi_9 = {checkVec_checkResult_hi_hi_hi_9, checkVec_checkResult_hi_hi_lo_9};
  wire [31:0]       checkVec_checkResult_hi_9 = {checkVec_checkResult_hi_hi_9, checkVec_checkResult_hi_lo_9};
  wire [63:0]       checkVec_1_2 = {checkVec_checkResult_hi_9, checkVec_checkResult_lo_9};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_10 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_0_3_1};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_10 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_2_3_1};
  wire [3:0]        checkVec_checkResult_lo_lo_10 = {checkVec_checkResult_lo_lo_hi_10, checkVec_checkResult_lo_lo_lo_10};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_10 = {checkVec_checkResultVec_5_3_1, checkVec_checkResultVec_4_3_1};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_10 = {checkVec_checkResultVec_7_3_1, checkVec_checkResultVec_6_3_1};
  wire [3:0]        checkVec_checkResult_lo_hi_10 = {checkVec_checkResult_lo_hi_hi_10, checkVec_checkResult_lo_hi_lo_10};
  wire [7:0]        checkVec_checkResult_lo_10 = {checkVec_checkResult_lo_hi_10, checkVec_checkResult_lo_lo_10};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_10 = {checkVec_checkResultVec_9_3_1, checkVec_checkResultVec_8_3_1};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_10 = {checkVec_checkResultVec_11_3_1, checkVec_checkResultVec_10_3_1};
  wire [3:0]        checkVec_checkResult_hi_lo_10 = {checkVec_checkResult_hi_lo_hi_10, checkVec_checkResult_hi_lo_lo_10};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_10 = {checkVec_checkResultVec_13_3_1, checkVec_checkResultVec_12_3_1};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_10 = {checkVec_checkResultVec_15_3_1, checkVec_checkResultVec_14_3_1};
  wire [3:0]        checkVec_checkResult_hi_hi_10 = {checkVec_checkResult_hi_hi_hi_10, checkVec_checkResult_hi_hi_lo_10};
  wire [7:0]        checkVec_checkResult_hi_10 = {checkVec_checkResult_hi_hi_10, checkVec_checkResult_hi_lo_10};
  wire [15:0]       checkVec_1_3 = {checkVec_checkResult_hi_10, checkVec_checkResult_lo_10};
  wire [5:0]        checkVec_checkResult_lo_lo_lo_11 = {checkVec_checkResultVec_1_4_1, checkVec_checkResultVec_0_4_1};
  wire [5:0]        checkVec_checkResult_lo_lo_hi_11 = {checkVec_checkResultVec_3_4_1, checkVec_checkResultVec_2_4_1};
  wire [11:0]       checkVec_checkResult_lo_lo_11 = {checkVec_checkResult_lo_lo_hi_11, checkVec_checkResult_lo_lo_lo_11};
  wire [5:0]        checkVec_checkResult_lo_hi_lo_11 = {checkVec_checkResultVec_5_4_1, checkVec_checkResultVec_4_4_1};
  wire [5:0]        checkVec_checkResult_lo_hi_hi_11 = {checkVec_checkResultVec_7_4_1, checkVec_checkResultVec_6_4_1};
  wire [11:0]       checkVec_checkResult_lo_hi_11 = {checkVec_checkResult_lo_hi_hi_11, checkVec_checkResult_lo_hi_lo_11};
  wire [23:0]       checkVec_checkResult_lo_11 = {checkVec_checkResult_lo_hi_11, checkVec_checkResult_lo_lo_11};
  wire [5:0]        checkVec_checkResult_hi_lo_lo_11 = {checkVec_checkResultVec_9_4_1, checkVec_checkResultVec_8_4_1};
  wire [5:0]        checkVec_checkResult_hi_lo_hi_11 = {checkVec_checkResultVec_11_4_1, checkVec_checkResultVec_10_4_1};
  wire [11:0]       checkVec_checkResult_hi_lo_11 = {checkVec_checkResult_hi_lo_hi_11, checkVec_checkResult_hi_lo_lo_11};
  wire [5:0]        checkVec_checkResult_hi_hi_lo_11 = {checkVec_checkResultVec_13_4_1, checkVec_checkResultVec_12_4_1};
  wire [5:0]        checkVec_checkResult_hi_hi_hi_11 = {checkVec_checkResultVec_15_4_1, checkVec_checkResultVec_14_4_1};
  wire [11:0]       checkVec_checkResult_hi_hi_11 = {checkVec_checkResult_hi_hi_hi_11, checkVec_checkResult_hi_hi_lo_11};
  wire [23:0]       checkVec_checkResult_hi_11 = {checkVec_checkResult_hi_hi_11, checkVec_checkResult_hi_lo_11};
  wire [47:0]       checkVec_1_4 = {checkVec_checkResult_hi_11, checkVec_checkResult_lo_11};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_12 = {checkVec_checkResultVec_1_5_1, checkVec_checkResultVec_0_5_1};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_12 = {checkVec_checkResultVec_3_5_1, checkVec_checkResultVec_2_5_1};
  wire [3:0]        checkVec_checkResult_lo_lo_12 = {checkVec_checkResult_lo_lo_hi_12, checkVec_checkResult_lo_lo_lo_12};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_12 = {checkVec_checkResultVec_5_5_1, checkVec_checkResultVec_4_5_1};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_12 = {checkVec_checkResultVec_7_5_1, checkVec_checkResultVec_6_5_1};
  wire [3:0]        checkVec_checkResult_lo_hi_12 = {checkVec_checkResult_lo_hi_hi_12, checkVec_checkResult_lo_hi_lo_12};
  wire [7:0]        checkVec_checkResult_lo_12 = {checkVec_checkResult_lo_hi_12, checkVec_checkResult_lo_lo_12};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_12 = {checkVec_checkResultVec_9_5_1, checkVec_checkResultVec_8_5_1};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_12 = {checkVec_checkResultVec_11_5_1, checkVec_checkResultVec_10_5_1};
  wire [3:0]        checkVec_checkResult_hi_lo_12 = {checkVec_checkResult_hi_lo_hi_12, checkVec_checkResult_hi_lo_lo_12};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_12 = {checkVec_checkResultVec_13_5_1, checkVec_checkResultVec_12_5_1};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_12 = {checkVec_checkResultVec_15_5_1, checkVec_checkResultVec_14_5_1};
  wire [3:0]        checkVec_checkResult_hi_hi_12 = {checkVec_checkResult_hi_hi_hi_12, checkVec_checkResult_hi_hi_lo_12};
  wire [7:0]        checkVec_checkResult_hi_12 = {checkVec_checkResult_hi_hi_12, checkVec_checkResult_hi_lo_12};
  wire [15:0]       checkVec_1_5 = {checkVec_checkResult_hi_12, checkVec_checkResult_lo_12};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_13 = {checkVec_checkResultVec_1_6_1, checkVec_checkResultVec_0_6_1};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_13 = {checkVec_checkResultVec_3_6_1, checkVec_checkResultVec_2_6_1};
  wire [3:0]        checkVec_checkResult_lo_lo_13 = {checkVec_checkResult_lo_lo_hi_13, checkVec_checkResult_lo_lo_lo_13};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_13 = {checkVec_checkResultVec_5_6_1, checkVec_checkResultVec_4_6_1};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_13 = {checkVec_checkResultVec_7_6_1, checkVec_checkResultVec_6_6_1};
  wire [3:0]        checkVec_checkResult_lo_hi_13 = {checkVec_checkResult_lo_hi_hi_13, checkVec_checkResult_lo_hi_lo_13};
  wire [7:0]        checkVec_checkResult_lo_13 = {checkVec_checkResult_lo_hi_13, checkVec_checkResult_lo_lo_13};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_13 = {checkVec_checkResultVec_9_6_1, checkVec_checkResultVec_8_6_1};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_13 = {checkVec_checkResultVec_11_6_1, checkVec_checkResultVec_10_6_1};
  wire [3:0]        checkVec_checkResult_hi_lo_13 = {checkVec_checkResult_hi_lo_hi_13, checkVec_checkResult_hi_lo_lo_13};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_13 = {checkVec_checkResultVec_13_6_1, checkVec_checkResultVec_12_6_1};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_13 = {checkVec_checkResultVec_15_6_1, checkVec_checkResultVec_14_6_1};
  wire [3:0]        checkVec_checkResult_hi_hi_13 = {checkVec_checkResult_hi_hi_hi_13, checkVec_checkResult_hi_hi_lo_13};
  wire [7:0]        checkVec_checkResult_hi_13 = {checkVec_checkResult_hi_hi_13, checkVec_checkResult_hi_lo_13};
  wire [15:0]       checkVec_1_6 = {checkVec_checkResult_hi_13, checkVec_checkResult_lo_13};
  wire              checkVec_checkResultVec_0_6_2 = checkVec_validVec_2[0];
  wire [9:0]        checkVec_checkResultVec_dataPosition_32 = {source_0[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_0_2_2 = checkVec_checkResultVec_dataPosition_32[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_32 = checkVec_checkResultVec_dataPosition_32[9:6];
  wire              checkVec_checkResultVec_0_3_2 = checkVec_checkResultVec_dataGroup_32[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_32 = checkVec_checkResultVec_dataGroup_32[3:1];
  wire [2:0]        checkVec_checkResultVec_0_4_2 = checkVec_checkResultVec_accessRegGrowth_32;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_32 = {checkVec_checkResultVec_0_3_2, checkVec_checkResultVec_0_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_32 = checkVec_checkResultVec_decimalProportion_32[4:2];
  wire              checkVec_checkResultVec_overlap_32 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_32 >= checkVec_checkResultVec_intLMULInput_32[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_32} >= checkVec_checkResultVec_intLMULInput_32,
      source_0[31:10]};
  wire              checkVec_checkResultVec_0_5_2 = checkVec_checkResultVec_overlap_32 | ~checkVec_checkResultVec_0_6_2;
  wire              checkVec_checkResultVec_1_6_2 = checkVec_validVec_2[1];
  wire [9:0]        checkVec_checkResultVec_dataPosition_33 = {source_1[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_1_2_2 = checkVec_checkResultVec_dataPosition_33[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_33 = checkVec_checkResultVec_dataPosition_33[9:6];
  wire              checkVec_checkResultVec_1_3_2 = checkVec_checkResultVec_dataGroup_33[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_33 = checkVec_checkResultVec_dataGroup_33[3:1];
  wire [2:0]        checkVec_checkResultVec_1_4_2 = checkVec_checkResultVec_accessRegGrowth_33;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_33 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_1_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_33 = checkVec_checkResultVec_decimalProportion_33[4:2];
  wire              checkVec_checkResultVec_overlap_33 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_33 >= checkVec_checkResultVec_intLMULInput_33[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_33} >= checkVec_checkResultVec_intLMULInput_33,
      source_1[31:10]};
  wire              checkVec_checkResultVec_1_5_2 = checkVec_checkResultVec_overlap_33 | ~checkVec_checkResultVec_1_6_2;
  wire              checkVec_checkResultVec_2_6_2 = checkVec_validVec_2[2];
  wire [9:0]        checkVec_checkResultVec_dataPosition_34 = {source_2[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_2_2_2 = checkVec_checkResultVec_dataPosition_34[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_34 = checkVec_checkResultVec_dataPosition_34[9:6];
  wire              checkVec_checkResultVec_2_3_2 = checkVec_checkResultVec_dataGroup_34[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_34 = checkVec_checkResultVec_dataGroup_34[3:1];
  wire [2:0]        checkVec_checkResultVec_2_4_2 = checkVec_checkResultVec_accessRegGrowth_34;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_34 = {checkVec_checkResultVec_2_3_2, checkVec_checkResultVec_2_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_34 = checkVec_checkResultVec_decimalProportion_34[4:2];
  wire              checkVec_checkResultVec_overlap_34 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_34 >= checkVec_checkResultVec_intLMULInput_34[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_34} >= checkVec_checkResultVec_intLMULInput_34,
      source_2[31:10]};
  wire              checkVec_checkResultVec_2_5_2 = checkVec_checkResultVec_overlap_34 | ~checkVec_checkResultVec_2_6_2;
  wire              checkVec_checkResultVec_3_6_2 = checkVec_validVec_2[3];
  wire [9:0]        checkVec_checkResultVec_dataPosition_35 = {source_3[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_3_2_2 = checkVec_checkResultVec_dataPosition_35[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_35 = checkVec_checkResultVec_dataPosition_35[9:6];
  wire              checkVec_checkResultVec_3_3_2 = checkVec_checkResultVec_dataGroup_35[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_35 = checkVec_checkResultVec_dataGroup_35[3:1];
  wire [2:0]        checkVec_checkResultVec_3_4_2 = checkVec_checkResultVec_accessRegGrowth_35;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_35 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_3_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_35 = checkVec_checkResultVec_decimalProportion_35[4:2];
  wire              checkVec_checkResultVec_overlap_35 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_35 >= checkVec_checkResultVec_intLMULInput_35[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_35} >= checkVec_checkResultVec_intLMULInput_35,
      source_3[31:10]};
  wire              checkVec_checkResultVec_3_5_2 = checkVec_checkResultVec_overlap_35 | ~checkVec_checkResultVec_3_6_2;
  wire              checkVec_checkResultVec_4_6_2 = checkVec_validVec_2[4];
  wire [9:0]        checkVec_checkResultVec_dataPosition_36 = {source_4[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_4_2_2 = checkVec_checkResultVec_dataPosition_36[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_36 = checkVec_checkResultVec_dataPosition_36[9:6];
  wire              checkVec_checkResultVec_4_3_2 = checkVec_checkResultVec_dataGroup_36[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_36 = checkVec_checkResultVec_dataGroup_36[3:1];
  wire [2:0]        checkVec_checkResultVec_4_4_2 = checkVec_checkResultVec_accessRegGrowth_36;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_36 = {checkVec_checkResultVec_4_3_2, checkVec_checkResultVec_4_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_36 = checkVec_checkResultVec_decimalProportion_36[4:2];
  wire              checkVec_checkResultVec_overlap_36 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_36 >= checkVec_checkResultVec_intLMULInput_36[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_36} >= checkVec_checkResultVec_intLMULInput_36,
      source_4[31:10]};
  wire              checkVec_checkResultVec_4_5_2 = checkVec_checkResultVec_overlap_36 | ~checkVec_checkResultVec_4_6_2;
  wire              checkVec_checkResultVec_5_6_2 = checkVec_validVec_2[5];
  wire [9:0]        checkVec_checkResultVec_dataPosition_37 = {source_5[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_5_2_2 = checkVec_checkResultVec_dataPosition_37[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_37 = checkVec_checkResultVec_dataPosition_37[9:6];
  wire              checkVec_checkResultVec_5_3_2 = checkVec_checkResultVec_dataGroup_37[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_37 = checkVec_checkResultVec_dataGroup_37[3:1];
  wire [2:0]        checkVec_checkResultVec_5_4_2 = checkVec_checkResultVec_accessRegGrowth_37;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_37 = {checkVec_checkResultVec_5_3_2, checkVec_checkResultVec_5_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_37 = checkVec_checkResultVec_decimalProportion_37[4:2];
  wire              checkVec_checkResultVec_overlap_37 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_37 >= checkVec_checkResultVec_intLMULInput_37[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_37} >= checkVec_checkResultVec_intLMULInput_37,
      source_5[31:10]};
  wire              checkVec_checkResultVec_5_5_2 = checkVec_checkResultVec_overlap_37 | ~checkVec_checkResultVec_5_6_2;
  wire              checkVec_checkResultVec_6_6_2 = checkVec_validVec_2[6];
  wire [9:0]        checkVec_checkResultVec_dataPosition_38 = {source_6[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_6_2_2 = checkVec_checkResultVec_dataPosition_38[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_38 = checkVec_checkResultVec_dataPosition_38[9:6];
  wire              checkVec_checkResultVec_6_3_2 = checkVec_checkResultVec_dataGroup_38[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_38 = checkVec_checkResultVec_dataGroup_38[3:1];
  wire [2:0]        checkVec_checkResultVec_6_4_2 = checkVec_checkResultVec_accessRegGrowth_38;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_38 = {checkVec_checkResultVec_6_3_2, checkVec_checkResultVec_6_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_38 = checkVec_checkResultVec_decimalProportion_38[4:2];
  wire              checkVec_checkResultVec_overlap_38 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_38 >= checkVec_checkResultVec_intLMULInput_38[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_38} >= checkVec_checkResultVec_intLMULInput_38,
      source_6[31:10]};
  wire              checkVec_checkResultVec_6_5_2 = checkVec_checkResultVec_overlap_38 | ~checkVec_checkResultVec_6_6_2;
  wire              checkVec_checkResultVec_7_6_2 = checkVec_validVec_2[7];
  wire [9:0]        checkVec_checkResultVec_dataPosition_39 = {source_7[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_7_2_2 = checkVec_checkResultVec_dataPosition_39[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_39 = checkVec_checkResultVec_dataPosition_39[9:6];
  wire              checkVec_checkResultVec_7_3_2 = checkVec_checkResultVec_dataGroup_39[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_39 = checkVec_checkResultVec_dataGroup_39[3:1];
  wire [2:0]        checkVec_checkResultVec_7_4_2 = checkVec_checkResultVec_accessRegGrowth_39;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_39 = {checkVec_checkResultVec_7_3_2, checkVec_checkResultVec_7_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_39 = checkVec_checkResultVec_decimalProportion_39[4:2];
  wire              checkVec_checkResultVec_overlap_39 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_39 >= checkVec_checkResultVec_intLMULInput_39[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_39} >= checkVec_checkResultVec_intLMULInput_39,
      source_7[31:10]};
  wire              checkVec_checkResultVec_7_5_2 = checkVec_checkResultVec_overlap_39 | ~checkVec_checkResultVec_7_6_2;
  wire              checkVec_checkResultVec_8_6_2 = checkVec_validVec_2[8];
  wire [9:0]        checkVec_checkResultVec_dataPosition_40 = {source_8[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_8_2_2 = checkVec_checkResultVec_dataPosition_40[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_40 = checkVec_checkResultVec_dataPosition_40[9:6];
  wire              checkVec_checkResultVec_8_3_2 = checkVec_checkResultVec_dataGroup_40[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_40 = checkVec_checkResultVec_dataGroup_40[3:1];
  wire [2:0]        checkVec_checkResultVec_8_4_2 = checkVec_checkResultVec_accessRegGrowth_40;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_40 = {checkVec_checkResultVec_8_3_2, checkVec_checkResultVec_8_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_40 = checkVec_checkResultVec_decimalProportion_40[4:2];
  wire              checkVec_checkResultVec_overlap_40 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_40 >= checkVec_checkResultVec_intLMULInput_40[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_40} >= checkVec_checkResultVec_intLMULInput_40,
      source_8[31:10]};
  wire              checkVec_checkResultVec_8_5_2 = checkVec_checkResultVec_overlap_40 | ~checkVec_checkResultVec_8_6_2;
  wire              checkVec_checkResultVec_9_6_2 = checkVec_validVec_2[9];
  wire [9:0]        checkVec_checkResultVec_dataPosition_41 = {source_9[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_9_2_2 = checkVec_checkResultVec_dataPosition_41[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_41 = checkVec_checkResultVec_dataPosition_41[9:6];
  wire              checkVec_checkResultVec_9_3_2 = checkVec_checkResultVec_dataGroup_41[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_41 = checkVec_checkResultVec_dataGroup_41[3:1];
  wire [2:0]        checkVec_checkResultVec_9_4_2 = checkVec_checkResultVec_accessRegGrowth_41;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_41 = {checkVec_checkResultVec_9_3_2, checkVec_checkResultVec_9_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_41 = checkVec_checkResultVec_decimalProportion_41[4:2];
  wire              checkVec_checkResultVec_overlap_41 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_41 >= checkVec_checkResultVec_intLMULInput_41[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_41} >= checkVec_checkResultVec_intLMULInput_41,
      source_9[31:10]};
  wire              checkVec_checkResultVec_9_5_2 = checkVec_checkResultVec_overlap_41 | ~checkVec_checkResultVec_9_6_2;
  wire              checkVec_checkResultVec_10_6_2 = checkVec_validVec_2[10];
  wire [9:0]        checkVec_checkResultVec_dataPosition_42 = {source_10[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_10_2_2 = checkVec_checkResultVec_dataPosition_42[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_42 = checkVec_checkResultVec_dataPosition_42[9:6];
  wire              checkVec_checkResultVec_10_3_2 = checkVec_checkResultVec_dataGroup_42[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_42 = checkVec_checkResultVec_dataGroup_42[3:1];
  wire [2:0]        checkVec_checkResultVec_10_4_2 = checkVec_checkResultVec_accessRegGrowth_42;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_42 = {checkVec_checkResultVec_10_3_2, checkVec_checkResultVec_10_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_42 = checkVec_checkResultVec_decimalProportion_42[4:2];
  wire              checkVec_checkResultVec_overlap_42 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_42 >= checkVec_checkResultVec_intLMULInput_42[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_42} >= checkVec_checkResultVec_intLMULInput_42,
      source_10[31:10]};
  wire              checkVec_checkResultVec_10_5_2 = checkVec_checkResultVec_overlap_42 | ~checkVec_checkResultVec_10_6_2;
  wire              checkVec_checkResultVec_11_6_2 = checkVec_validVec_2[11];
  wire [9:0]        checkVec_checkResultVec_dataPosition_43 = {source_11[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_11_2_2 = checkVec_checkResultVec_dataPosition_43[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_43 = checkVec_checkResultVec_dataPosition_43[9:6];
  wire              checkVec_checkResultVec_11_3_2 = checkVec_checkResultVec_dataGroup_43[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_43 = checkVec_checkResultVec_dataGroup_43[3:1];
  wire [2:0]        checkVec_checkResultVec_11_4_2 = checkVec_checkResultVec_accessRegGrowth_43;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_43 = {checkVec_checkResultVec_11_3_2, checkVec_checkResultVec_11_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_43 = checkVec_checkResultVec_decimalProportion_43[4:2];
  wire              checkVec_checkResultVec_overlap_43 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_43 >= checkVec_checkResultVec_intLMULInput_43[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_43} >= checkVec_checkResultVec_intLMULInput_43,
      source_11[31:10]};
  wire              checkVec_checkResultVec_11_5_2 = checkVec_checkResultVec_overlap_43 | ~checkVec_checkResultVec_11_6_2;
  wire              checkVec_checkResultVec_12_6_2 = checkVec_validVec_2[12];
  wire [9:0]        checkVec_checkResultVec_dataPosition_44 = {source_12[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_12_2_2 = checkVec_checkResultVec_dataPosition_44[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_44 = checkVec_checkResultVec_dataPosition_44[9:6];
  wire              checkVec_checkResultVec_12_3_2 = checkVec_checkResultVec_dataGroup_44[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_44 = checkVec_checkResultVec_dataGroup_44[3:1];
  wire [2:0]        checkVec_checkResultVec_12_4_2 = checkVec_checkResultVec_accessRegGrowth_44;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_44 = {checkVec_checkResultVec_12_3_2, checkVec_checkResultVec_12_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_44 = checkVec_checkResultVec_decimalProportion_44[4:2];
  wire              checkVec_checkResultVec_overlap_44 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_44 >= checkVec_checkResultVec_intLMULInput_44[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_44} >= checkVec_checkResultVec_intLMULInput_44,
      source_12[31:10]};
  wire              checkVec_checkResultVec_12_5_2 = checkVec_checkResultVec_overlap_44 | ~checkVec_checkResultVec_12_6_2;
  wire              checkVec_checkResultVec_13_6_2 = checkVec_validVec_2[13];
  wire [9:0]        checkVec_checkResultVec_dataPosition_45 = {source_13[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_13_2_2 = checkVec_checkResultVec_dataPosition_45[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_45 = checkVec_checkResultVec_dataPosition_45[9:6];
  wire              checkVec_checkResultVec_13_3_2 = checkVec_checkResultVec_dataGroup_45[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_45 = checkVec_checkResultVec_dataGroup_45[3:1];
  wire [2:0]        checkVec_checkResultVec_13_4_2 = checkVec_checkResultVec_accessRegGrowth_45;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_45 = {checkVec_checkResultVec_13_3_2, checkVec_checkResultVec_13_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_45 = checkVec_checkResultVec_decimalProportion_45[4:2];
  wire              checkVec_checkResultVec_overlap_45 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_45 >= checkVec_checkResultVec_intLMULInput_45[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_45} >= checkVec_checkResultVec_intLMULInput_45,
      source_13[31:10]};
  wire              checkVec_checkResultVec_13_5_2 = checkVec_checkResultVec_overlap_45 | ~checkVec_checkResultVec_13_6_2;
  wire              checkVec_checkResultVec_14_6_2 = checkVec_validVec_2[14];
  wire [9:0]        checkVec_checkResultVec_dataPosition_46 = {source_14[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_14_2_2 = checkVec_checkResultVec_dataPosition_46[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_46 = checkVec_checkResultVec_dataPosition_46[9:6];
  wire              checkVec_checkResultVec_14_3_2 = checkVec_checkResultVec_dataGroup_46[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_46 = checkVec_checkResultVec_dataGroup_46[3:1];
  wire [2:0]        checkVec_checkResultVec_14_4_2 = checkVec_checkResultVec_accessRegGrowth_46;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_46 = {checkVec_checkResultVec_14_3_2, checkVec_checkResultVec_14_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_46 = checkVec_checkResultVec_decimalProportion_46[4:2];
  wire              checkVec_checkResultVec_overlap_46 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_46 >= checkVec_checkResultVec_intLMULInput_46[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_46} >= checkVec_checkResultVec_intLMULInput_46,
      source_14[31:10]};
  wire              checkVec_checkResultVec_14_5_2 = checkVec_checkResultVec_overlap_46 | ~checkVec_checkResultVec_14_6_2;
  wire              checkVec_checkResultVec_15_6_2 = checkVec_validVec_2[15];
  wire [9:0]        checkVec_checkResultVec_dataPosition_47 = {source_15[7:0], 2'h0};
  wire [3:0]        checkVec_checkResultVec_15_2_2 = checkVec_checkResultVec_dataPosition_47[5:2];
  wire [3:0]        checkVec_checkResultVec_dataGroup_47 = checkVec_checkResultVec_dataPosition_47[9:6];
  wire              checkVec_checkResultVec_15_3_2 = checkVec_checkResultVec_dataGroup_47[0];
  wire [2:0]        checkVec_checkResultVec_accessRegGrowth_47 = checkVec_checkResultVec_dataGroup_47[3:1];
  wire [2:0]        checkVec_checkResultVec_15_4_2 = checkVec_checkResultVec_accessRegGrowth_47;
  wire [4:0]        checkVec_checkResultVec_decimalProportion_47 = {checkVec_checkResultVec_15_3_2, checkVec_checkResultVec_15_2_2};
  wire [2:0]        checkVec_checkResultVec_decimal_47 = checkVec_checkResultVec_decimalProportion_47[4:2];
  wire              checkVec_checkResultVec_overlap_47 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_47 >= checkVec_checkResultVec_intLMULInput_47[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_47} >= checkVec_checkResultVec_intLMULInput_47,
      source_15[31:10]};
  wire              checkVec_checkResultVec_15_5_2 = checkVec_checkResultVec_overlap_47 | ~checkVec_checkResultVec_15_6_2;
  wire [7:0]        checkVec_checkResult_lo_lo_lo_16 = {checkVec_checkResultVec_1_2_2, checkVec_checkResultVec_0_2_2};
  wire [7:0]        checkVec_checkResult_lo_lo_hi_16 = {checkVec_checkResultVec_3_2_2, checkVec_checkResultVec_2_2_2};
  wire [15:0]       checkVec_checkResult_lo_lo_16 = {checkVec_checkResult_lo_lo_hi_16, checkVec_checkResult_lo_lo_lo_16};
  wire [7:0]        checkVec_checkResult_lo_hi_lo_16 = {checkVec_checkResultVec_5_2_2, checkVec_checkResultVec_4_2_2};
  wire [7:0]        checkVec_checkResult_lo_hi_hi_16 = {checkVec_checkResultVec_7_2_2, checkVec_checkResultVec_6_2_2};
  wire [15:0]       checkVec_checkResult_lo_hi_16 = {checkVec_checkResult_lo_hi_hi_16, checkVec_checkResult_lo_hi_lo_16};
  wire [31:0]       checkVec_checkResult_lo_16 = {checkVec_checkResult_lo_hi_16, checkVec_checkResult_lo_lo_16};
  wire [7:0]        checkVec_checkResult_hi_lo_lo_16 = {checkVec_checkResultVec_9_2_2, checkVec_checkResultVec_8_2_2};
  wire [7:0]        checkVec_checkResult_hi_lo_hi_16 = {checkVec_checkResultVec_11_2_2, checkVec_checkResultVec_10_2_2};
  wire [15:0]       checkVec_checkResult_hi_lo_16 = {checkVec_checkResult_hi_lo_hi_16, checkVec_checkResult_hi_lo_lo_16};
  wire [7:0]        checkVec_checkResult_hi_hi_lo_16 = {checkVec_checkResultVec_13_2_2, checkVec_checkResultVec_12_2_2};
  wire [7:0]        checkVec_checkResult_hi_hi_hi_16 = {checkVec_checkResultVec_15_2_2, checkVec_checkResultVec_14_2_2};
  wire [15:0]       checkVec_checkResult_hi_hi_16 = {checkVec_checkResult_hi_hi_hi_16, checkVec_checkResult_hi_hi_lo_16};
  wire [31:0]       checkVec_checkResult_hi_16 = {checkVec_checkResult_hi_hi_16, checkVec_checkResult_hi_lo_16};
  wire [63:0]       checkVec_2_2 = {checkVec_checkResult_hi_16, checkVec_checkResult_lo_16};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_17 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_0_3_2};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_17 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_2_3_2};
  wire [3:0]        checkVec_checkResult_lo_lo_17 = {checkVec_checkResult_lo_lo_hi_17, checkVec_checkResult_lo_lo_lo_17};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_17 = {checkVec_checkResultVec_5_3_2, checkVec_checkResultVec_4_3_2};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_17 = {checkVec_checkResultVec_7_3_2, checkVec_checkResultVec_6_3_2};
  wire [3:0]        checkVec_checkResult_lo_hi_17 = {checkVec_checkResult_lo_hi_hi_17, checkVec_checkResult_lo_hi_lo_17};
  wire [7:0]        checkVec_checkResult_lo_17 = {checkVec_checkResult_lo_hi_17, checkVec_checkResult_lo_lo_17};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_17 = {checkVec_checkResultVec_9_3_2, checkVec_checkResultVec_8_3_2};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_17 = {checkVec_checkResultVec_11_3_2, checkVec_checkResultVec_10_3_2};
  wire [3:0]        checkVec_checkResult_hi_lo_17 = {checkVec_checkResult_hi_lo_hi_17, checkVec_checkResult_hi_lo_lo_17};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_17 = {checkVec_checkResultVec_13_3_2, checkVec_checkResultVec_12_3_2};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_17 = {checkVec_checkResultVec_15_3_2, checkVec_checkResultVec_14_3_2};
  wire [3:0]        checkVec_checkResult_hi_hi_17 = {checkVec_checkResult_hi_hi_hi_17, checkVec_checkResult_hi_hi_lo_17};
  wire [7:0]        checkVec_checkResult_hi_17 = {checkVec_checkResult_hi_hi_17, checkVec_checkResult_hi_lo_17};
  wire [15:0]       checkVec_2_3 = {checkVec_checkResult_hi_17, checkVec_checkResult_lo_17};
  wire [5:0]        checkVec_checkResult_lo_lo_lo_18 = {checkVec_checkResultVec_1_4_2, checkVec_checkResultVec_0_4_2};
  wire [5:0]        checkVec_checkResult_lo_lo_hi_18 = {checkVec_checkResultVec_3_4_2, checkVec_checkResultVec_2_4_2};
  wire [11:0]       checkVec_checkResult_lo_lo_18 = {checkVec_checkResult_lo_lo_hi_18, checkVec_checkResult_lo_lo_lo_18};
  wire [5:0]        checkVec_checkResult_lo_hi_lo_18 = {checkVec_checkResultVec_5_4_2, checkVec_checkResultVec_4_4_2};
  wire [5:0]        checkVec_checkResult_lo_hi_hi_18 = {checkVec_checkResultVec_7_4_2, checkVec_checkResultVec_6_4_2};
  wire [11:0]       checkVec_checkResult_lo_hi_18 = {checkVec_checkResult_lo_hi_hi_18, checkVec_checkResult_lo_hi_lo_18};
  wire [23:0]       checkVec_checkResult_lo_18 = {checkVec_checkResult_lo_hi_18, checkVec_checkResult_lo_lo_18};
  wire [5:0]        checkVec_checkResult_hi_lo_lo_18 = {checkVec_checkResultVec_9_4_2, checkVec_checkResultVec_8_4_2};
  wire [5:0]        checkVec_checkResult_hi_lo_hi_18 = {checkVec_checkResultVec_11_4_2, checkVec_checkResultVec_10_4_2};
  wire [11:0]       checkVec_checkResult_hi_lo_18 = {checkVec_checkResult_hi_lo_hi_18, checkVec_checkResult_hi_lo_lo_18};
  wire [5:0]        checkVec_checkResult_hi_hi_lo_18 = {checkVec_checkResultVec_13_4_2, checkVec_checkResultVec_12_4_2};
  wire [5:0]        checkVec_checkResult_hi_hi_hi_18 = {checkVec_checkResultVec_15_4_2, checkVec_checkResultVec_14_4_2};
  wire [11:0]       checkVec_checkResult_hi_hi_18 = {checkVec_checkResult_hi_hi_hi_18, checkVec_checkResult_hi_hi_lo_18};
  wire [23:0]       checkVec_checkResult_hi_18 = {checkVec_checkResult_hi_hi_18, checkVec_checkResult_hi_lo_18};
  wire [47:0]       checkVec_2_4 = {checkVec_checkResult_hi_18, checkVec_checkResult_lo_18};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_19 = {checkVec_checkResultVec_1_5_2, checkVec_checkResultVec_0_5_2};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_19 = {checkVec_checkResultVec_3_5_2, checkVec_checkResultVec_2_5_2};
  wire [3:0]        checkVec_checkResult_lo_lo_19 = {checkVec_checkResult_lo_lo_hi_19, checkVec_checkResult_lo_lo_lo_19};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_19 = {checkVec_checkResultVec_5_5_2, checkVec_checkResultVec_4_5_2};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_19 = {checkVec_checkResultVec_7_5_2, checkVec_checkResultVec_6_5_2};
  wire [3:0]        checkVec_checkResult_lo_hi_19 = {checkVec_checkResult_lo_hi_hi_19, checkVec_checkResult_lo_hi_lo_19};
  wire [7:0]        checkVec_checkResult_lo_19 = {checkVec_checkResult_lo_hi_19, checkVec_checkResult_lo_lo_19};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_19 = {checkVec_checkResultVec_9_5_2, checkVec_checkResultVec_8_5_2};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_19 = {checkVec_checkResultVec_11_5_2, checkVec_checkResultVec_10_5_2};
  wire [3:0]        checkVec_checkResult_hi_lo_19 = {checkVec_checkResult_hi_lo_hi_19, checkVec_checkResult_hi_lo_lo_19};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_19 = {checkVec_checkResultVec_13_5_2, checkVec_checkResultVec_12_5_2};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_19 = {checkVec_checkResultVec_15_5_2, checkVec_checkResultVec_14_5_2};
  wire [3:0]        checkVec_checkResult_hi_hi_19 = {checkVec_checkResult_hi_hi_hi_19, checkVec_checkResult_hi_hi_lo_19};
  wire [7:0]        checkVec_checkResult_hi_19 = {checkVec_checkResult_hi_hi_19, checkVec_checkResult_hi_lo_19};
  wire [15:0]       checkVec_2_5 = {checkVec_checkResult_hi_19, checkVec_checkResult_lo_19};
  wire [1:0]        checkVec_checkResult_lo_lo_lo_20 = {checkVec_checkResultVec_1_6_2, checkVec_checkResultVec_0_6_2};
  wire [1:0]        checkVec_checkResult_lo_lo_hi_20 = {checkVec_checkResultVec_3_6_2, checkVec_checkResultVec_2_6_2};
  wire [3:0]        checkVec_checkResult_lo_lo_20 = {checkVec_checkResult_lo_lo_hi_20, checkVec_checkResult_lo_lo_lo_20};
  wire [1:0]        checkVec_checkResult_lo_hi_lo_20 = {checkVec_checkResultVec_5_6_2, checkVec_checkResultVec_4_6_2};
  wire [1:0]        checkVec_checkResult_lo_hi_hi_20 = {checkVec_checkResultVec_7_6_2, checkVec_checkResultVec_6_6_2};
  wire [3:0]        checkVec_checkResult_lo_hi_20 = {checkVec_checkResult_lo_hi_hi_20, checkVec_checkResult_lo_hi_lo_20};
  wire [7:0]        checkVec_checkResult_lo_20 = {checkVec_checkResult_lo_hi_20, checkVec_checkResult_lo_lo_20};
  wire [1:0]        checkVec_checkResult_hi_lo_lo_20 = {checkVec_checkResultVec_9_6_2, checkVec_checkResultVec_8_6_2};
  wire [1:0]        checkVec_checkResult_hi_lo_hi_20 = {checkVec_checkResultVec_11_6_2, checkVec_checkResultVec_10_6_2};
  wire [3:0]        checkVec_checkResult_hi_lo_20 = {checkVec_checkResult_hi_lo_hi_20, checkVec_checkResult_hi_lo_lo_20};
  wire [1:0]        checkVec_checkResult_hi_hi_lo_20 = {checkVec_checkResultVec_13_6_2, checkVec_checkResultVec_12_6_2};
  wire [1:0]        checkVec_checkResult_hi_hi_hi_20 = {checkVec_checkResultVec_15_6_2, checkVec_checkResultVec_14_6_2};
  wire [3:0]        checkVec_checkResult_hi_hi_20 = {checkVec_checkResult_hi_hi_hi_20, checkVec_checkResult_hi_hi_lo_20};
  wire [7:0]        checkVec_checkResult_hi_20 = {checkVec_checkResult_hi_hi_20, checkVec_checkResult_hi_lo_20};
  wire [15:0]       checkVec_2_6 = {checkVec_checkResult_hi_20, checkVec_checkResult_lo_20};
  wire [31:0]       dataOffsetSelect = (sew1H[0] ? checkVec_0_1 : 32'h0) | (sew1H[1] ? checkVec_1_1 : 32'h0);
  wire [63:0]       accessLaneSelect = (sew1H[0] ? checkVec_0_2 : 64'h0) | (sew1H[1] ? checkVec_1_2 : 64'h0) | (sew1H[2] ? checkVec_2_2 : 64'h0);
  wire [15:0]       offsetSelect = (sew1H[0] ? checkVec_0_3 : 16'h0) | (sew1H[1] ? checkVec_1_3 : 16'h0) | (sew1H[2] ? checkVec_2_3 : 16'h0);
  wire [47:0]       growthSelect = (sew1H[0] ? checkVec_0_4 : 48'h0) | (sew1H[1] ? checkVec_1_4 : 48'h0) | (sew1H[2] ? checkVec_2_4 : 48'h0);
  wire [15:0]       notReadSelect = (sew1H[0] ? checkVec_0_5 : 16'h0) | (sew1H[1] ? checkVec_1_5 : 16'h0) | (sew1H[2] ? checkVec_2_5 : 16'h0);
  wire [15:0]       elementValidSelect = (sew1H[0] ? checkVec_0_6 : 16'h0) | (sew1H[1] ? checkVec_1_6 : 16'h0) | (sew1H[2] ? checkVec_2_6 : 16'h0);
  wire              readTypeRequestDeq;
  wire              waiteStageEnqReady;
  wire              readWaitQueue_deq_valid;
  assign readWaitQueue_deq_valid = ~_readWaitQueue_fifo_empty;
  wire [6:0]        readWaitQueue_dataOut_executeGroup;
  wire [15:0]       readWaitQueue_dataOut_sourceValid;
  wire [15:0]       readWaitQueue_dataOut_replaceVs1;
  wire [15:0]       readWaitQueue_dataOut_needRead;
  wire              readWaitQueue_dataOut_last;
  wire [16:0]       readWaitQueue_dataIn_lo = {readWaitQueue_enq_bits_needRead, readWaitQueue_enq_bits_last};
  wire [22:0]       readWaitQueue_dataIn_hi_hi = {readWaitQueue_enq_bits_executeGroup, readWaitQueue_enq_bits_sourceValid};
  wire [38:0]       readWaitQueue_dataIn_hi = {readWaitQueue_dataIn_hi_hi, readWaitQueue_enq_bits_replaceVs1};
  wire [55:0]       readWaitQueue_dataIn = {readWaitQueue_dataIn_hi, readWaitQueue_dataIn_lo};
  assign readWaitQueue_dataOut_last = _readWaitQueue_fifo_data_out[0];
  assign readWaitQueue_dataOut_needRead = _readWaitQueue_fifo_data_out[16:1];
  assign readWaitQueue_dataOut_replaceVs1 = _readWaitQueue_fifo_data_out[32:17];
  assign readWaitQueue_dataOut_sourceValid = _readWaitQueue_fifo_data_out[48:33];
  assign readWaitQueue_dataOut_executeGroup = _readWaitQueue_fifo_data_out[55:49];
  wire [6:0]        readWaitQueue_deq_bits_executeGroup = readWaitQueue_dataOut_executeGroup;
  wire [15:0]       readWaitQueue_deq_bits_sourceValid = readWaitQueue_dataOut_sourceValid;
  wire [15:0]       readWaitQueue_deq_bits_replaceVs1 = readWaitQueue_dataOut_replaceVs1;
  wire [15:0]       readWaitQueue_deq_bits_needRead = readWaitQueue_dataOut_needRead;
  wire              readWaitQueue_deq_bits_last = readWaitQueue_dataOut_last;
  wire              readWaitQueue_enq_ready = ~_readWaitQueue_fifo_full;
  wire              readWaitQueue_enq_valid;
  wire              readWaitQueue_deq_ready;
  wire              _GEN_78 = lastExecuteGroupDeq | viota;
  assign exeRequestQueue_0_deq_ready = ~exeReqReg_0_valid | _GEN_78;
  assign exeRequestQueue_1_deq_ready = ~exeReqReg_1_valid | _GEN_78;
  assign exeRequestQueue_2_deq_ready = ~exeReqReg_2_valid | _GEN_78;
  assign exeRequestQueue_3_deq_ready = ~exeReqReg_3_valid | _GEN_78;
  assign exeRequestQueue_4_deq_ready = ~exeReqReg_4_valid | _GEN_78;
  assign exeRequestQueue_5_deq_ready = ~exeReqReg_5_valid | _GEN_78;
  assign exeRequestQueue_6_deq_ready = ~exeReqReg_6_valid | _GEN_78;
  assign exeRequestQueue_7_deq_ready = ~exeReqReg_7_valid | _GEN_78;
  assign exeRequestQueue_8_deq_ready = ~exeReqReg_8_valid | _GEN_78;
  assign exeRequestQueue_9_deq_ready = ~exeReqReg_9_valid | _GEN_78;
  assign exeRequestQueue_10_deq_ready = ~exeReqReg_10_valid | _GEN_78;
  assign exeRequestQueue_11_deq_ready = ~exeReqReg_11_valid | _GEN_78;
  assign exeRequestQueue_12_deq_ready = ~exeReqReg_12_valid | _GEN_78;
  assign exeRequestQueue_13_deq_ready = ~exeReqReg_13_valid | _GEN_78;
  assign exeRequestQueue_14_deq_ready = ~exeReqReg_14_valid | _GEN_78;
  assign exeRequestQueue_15_deq_ready = ~exeReqReg_15_valid | _GEN_78;
  wire              isLastExecuteGroup = executeIndex == lastExecuteIndex;
  wire              allDataValid =
    (exeReqReg_0_valid | ~(groupDataNeed[0])) & (exeReqReg_1_valid | ~(groupDataNeed[1])) & (exeReqReg_2_valid | ~(groupDataNeed[2])) & (exeReqReg_3_valid | ~(groupDataNeed[3])) & (exeReqReg_4_valid | ~(groupDataNeed[4]))
    & (exeReqReg_5_valid | ~(groupDataNeed[5])) & (exeReqReg_6_valid | ~(groupDataNeed[6])) & (exeReqReg_7_valid | ~(groupDataNeed[7])) & (exeReqReg_8_valid | ~(groupDataNeed[8])) & (exeReqReg_9_valid | ~(groupDataNeed[9]))
    & (exeReqReg_10_valid | ~(groupDataNeed[10])) & (exeReqReg_11_valid | ~(groupDataNeed[11])) & (exeReqReg_12_valid | ~(groupDataNeed[12])) & (exeReqReg_13_valid | ~(groupDataNeed[13])) & (exeReqReg_14_valid | ~(groupDataNeed[14]))
    & (exeReqReg_15_valid | ~(groupDataNeed[15]));
  wire              anyDataValid =
    exeReqReg_0_valid | exeReqReg_1_valid | exeReqReg_2_valid | exeReqReg_3_valid | exeReqReg_4_valid | exeReqReg_5_valid | exeReqReg_6_valid | exeReqReg_7_valid | exeReqReg_8_valid | exeReqReg_9_valid | exeReqReg_10_valid
    | exeReqReg_11_valid | exeReqReg_12_valid | exeReqReg_13_valid | exeReqReg_14_valid | exeReqReg_15_valid;
  wire              _GEN_79 = compress | mvRd;
  wire              readVs1Valid = (unitType[2] | _GEN_79) & ~readVS1Reg_requestSend | gatherSRead;
  wire              _GEN_80 = compress | ~gatherSRead;
  wire [4:0]        readVS1Req_vs = _GEN_80 ? instReg_vs1 : instReg_vs1 + {2'h0, gatherGrowth};
  wire              readVS1Req_offset = ~compress & gatherSRead & gatherOffset;
  wire [3:0]        readVS1Req_readLane = compress ? readVS1Reg_readIndex : gatherSRead ? gatherLane : 4'h0;
  wire [1:0]        readVS1Req_dataOffset = _GEN_80 ? 2'h0 : gatherDatOffset;
  wire              selectExecuteReq_1_bits_offset = readIssueStageState_readOffset[1];
  wire              selectExecuteReq_2_bits_offset = readIssueStageState_readOffset[2];
  wire              selectExecuteReq_3_bits_offset = readIssueStageState_readOffset[3];
  wire              selectExecuteReq_4_bits_offset = readIssueStageState_readOffset[4];
  wire              selectExecuteReq_5_bits_offset = readIssueStageState_readOffset[5];
  wire              selectExecuteReq_6_bits_offset = readIssueStageState_readOffset[6];
  wire              selectExecuteReq_7_bits_offset = readIssueStageState_readOffset[7];
  wire              selectExecuteReq_8_bits_offset = readIssueStageState_readOffset[8];
  wire              selectExecuteReq_9_bits_offset = readIssueStageState_readOffset[9];
  wire              selectExecuteReq_10_bits_offset = readIssueStageState_readOffset[10];
  wire              selectExecuteReq_11_bits_offset = readIssueStageState_readOffset[11];
  wire              selectExecuteReq_12_bits_offset = readIssueStageState_readOffset[12];
  wire              selectExecuteReq_13_bits_offset = readIssueStageState_readOffset[13];
  wire              selectExecuteReq_14_bits_offset = readIssueStageState_readOffset[14];
  wire              selectExecuteReq_15_bits_offset = readIssueStageState_readOffset[15];
  wire [1:0]        selectExecuteReq_1_bits_dataOffset = readIssueStageState_readDataOffset[3:2];
  wire [1:0]        selectExecuteReq_2_bits_dataOffset = readIssueStageState_readDataOffset[5:4];
  wire [1:0]        selectExecuteReq_3_bits_dataOffset = readIssueStageState_readDataOffset[7:6];
  wire [1:0]        selectExecuteReq_4_bits_dataOffset = readIssueStageState_readDataOffset[9:8];
  wire [1:0]        selectExecuteReq_5_bits_dataOffset = readIssueStageState_readDataOffset[11:10];
  wire [1:0]        selectExecuteReq_6_bits_dataOffset = readIssueStageState_readDataOffset[13:12];
  wire [1:0]        selectExecuteReq_7_bits_dataOffset = readIssueStageState_readDataOffset[15:14];
  wire [1:0]        selectExecuteReq_8_bits_dataOffset = readIssueStageState_readDataOffset[17:16];
  wire [1:0]        selectExecuteReq_9_bits_dataOffset = readIssueStageState_readDataOffset[19:18];
  wire [1:0]        selectExecuteReq_10_bits_dataOffset = readIssueStageState_readDataOffset[21:20];
  wire [1:0]        selectExecuteReq_11_bits_dataOffset = readIssueStageState_readDataOffset[23:22];
  wire [1:0]        selectExecuteReq_12_bits_dataOffset = readIssueStageState_readDataOffset[25:24];
  wire [1:0]        selectExecuteReq_13_bits_dataOffset = readIssueStageState_readDataOffset[27:26];
  wire [1:0]        selectExecuteReq_14_bits_dataOffset = readIssueStageState_readDataOffset[29:28];
  wire [1:0]        selectExecuteReq_15_bits_dataOffset = readIssueStageState_readDataOffset[31:30];
  wire              selectExecuteReq_0_valid = readVs1Valid | readIssueStageValid & ~(readIssueStageState_groupReadState[0]) & readIssueStageState_needRead[0] & readType;
  wire [4:0]        selectExecuteReq_0_bits_vs = readVs1Valid ? readVS1Req_vs : instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_0};
  wire              selectExecuteReq_0_bits_offset = readVs1Valid ? readVS1Req_offset : readIssueStageState_readOffset[0];
  wire [3:0]        selectExecuteReq_0_bits_readLane = readVs1Valid ? readVS1Req_readLane : readIssueStageState_accessLane_0;
  wire [1:0]        selectExecuteReq_0_bits_dataOffset = readVs1Valid ? readVS1Req_dataOffset : readIssueStageState_readDataOffset[1:0];
  wire              _tokenCheck_T = _readCrossBar_input_0_ready & readCrossBar_input_0_valid;
  wire              pipeReadFire_0 = ~readVs1Valid & _tokenCheck_T;
  wire [4:0]        selectExecuteReq_1_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_1};
  wire              selectExecuteReq_1_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[1]) & readIssueStageState_needRead[1] & readType;
  wire              pipeReadFire_1 = _readCrossBar_input_1_ready & readCrossBar_input_1_valid;
  wire [4:0]        selectExecuteReq_2_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_2};
  wire              selectExecuteReq_2_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[2]) & readIssueStageState_needRead[2] & readType;
  wire              pipeReadFire_2 = _readCrossBar_input_2_ready & readCrossBar_input_2_valid;
  wire [4:0]        selectExecuteReq_3_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_3};
  wire              selectExecuteReq_3_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[3]) & readIssueStageState_needRead[3] & readType;
  wire              pipeReadFire_3 = _readCrossBar_input_3_ready & readCrossBar_input_3_valid;
  wire [4:0]        selectExecuteReq_4_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_4};
  wire              selectExecuteReq_4_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[4]) & readIssueStageState_needRead[4] & readType;
  wire              pipeReadFire_4 = _readCrossBar_input_4_ready & readCrossBar_input_4_valid;
  wire [4:0]        selectExecuteReq_5_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_5};
  wire              selectExecuteReq_5_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[5]) & readIssueStageState_needRead[5] & readType;
  wire              pipeReadFire_5 = _readCrossBar_input_5_ready & readCrossBar_input_5_valid;
  wire [4:0]        selectExecuteReq_6_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_6};
  wire              selectExecuteReq_6_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[6]) & readIssueStageState_needRead[6] & readType;
  wire              pipeReadFire_6 = _readCrossBar_input_6_ready & readCrossBar_input_6_valid;
  wire [4:0]        selectExecuteReq_7_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_7};
  wire              selectExecuteReq_7_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[7]) & readIssueStageState_needRead[7] & readType;
  wire              pipeReadFire_7 = _readCrossBar_input_7_ready & readCrossBar_input_7_valid;
  wire [4:0]        selectExecuteReq_8_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_8};
  wire              selectExecuteReq_8_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[8]) & readIssueStageState_needRead[8] & readType;
  wire              pipeReadFire_8 = _readCrossBar_input_8_ready & readCrossBar_input_8_valid;
  wire [4:0]        selectExecuteReq_9_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_9};
  wire              selectExecuteReq_9_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[9]) & readIssueStageState_needRead[9] & readType;
  wire              pipeReadFire_9 = _readCrossBar_input_9_ready & readCrossBar_input_9_valid;
  wire [4:0]        selectExecuteReq_10_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_10};
  wire              selectExecuteReq_10_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[10]) & readIssueStageState_needRead[10] & readType;
  wire              pipeReadFire_10 = _readCrossBar_input_10_ready & readCrossBar_input_10_valid;
  wire [4:0]        selectExecuteReq_11_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_11};
  wire              selectExecuteReq_11_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[11]) & readIssueStageState_needRead[11] & readType;
  wire              pipeReadFire_11 = _readCrossBar_input_11_ready & readCrossBar_input_11_valid;
  wire [4:0]        selectExecuteReq_12_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_12};
  wire              selectExecuteReq_12_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[12]) & readIssueStageState_needRead[12] & readType;
  wire              pipeReadFire_12 = _readCrossBar_input_12_ready & readCrossBar_input_12_valid;
  wire [4:0]        selectExecuteReq_13_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_13};
  wire              selectExecuteReq_13_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[13]) & readIssueStageState_needRead[13] & readType;
  wire              pipeReadFire_13 = _readCrossBar_input_13_ready & readCrossBar_input_13_valid;
  wire [4:0]        selectExecuteReq_14_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_14};
  wire              selectExecuteReq_14_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[14]) & readIssueStageState_needRead[14] & readType;
  wire              pipeReadFire_14 = _readCrossBar_input_14_ready & readCrossBar_input_14_valid;
  wire [4:0]        selectExecuteReq_15_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_15};
  wire              selectExecuteReq_15_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[15]) & readIssueStageState_needRead[15] & readType;
  wire              pipeReadFire_15 = _readCrossBar_input_15_ready & readCrossBar_input_15_valid;
  reg  [3:0]        tokenCheck_counter;
  wire [3:0]        tokenCheck_counterChange = _tokenCheck_T ? 4'h1 : 4'hF;
  wire              tokenCheck = ~(tokenCheck_counter[3]);
  assign readCrossBar_input_0_valid = selectExecuteReq_0_valid & tokenCheck;
  reg  [3:0]        tokenCheck_counter_1;
  wire [3:0]        tokenCheck_counterChange_1 = pipeReadFire_1 ? 4'h1 : 4'hF;
  wire              tokenCheck_1 = ~(tokenCheck_counter_1[3]);
  assign readCrossBar_input_1_valid = selectExecuteReq_1_valid & tokenCheck_1;
  reg  [3:0]        tokenCheck_counter_2;
  wire [3:0]        tokenCheck_counterChange_2 = pipeReadFire_2 ? 4'h1 : 4'hF;
  wire              tokenCheck_2 = ~(tokenCheck_counter_2[3]);
  assign readCrossBar_input_2_valid = selectExecuteReq_2_valid & tokenCheck_2;
  reg  [3:0]        tokenCheck_counter_3;
  wire [3:0]        tokenCheck_counterChange_3 = pipeReadFire_3 ? 4'h1 : 4'hF;
  wire              tokenCheck_3 = ~(tokenCheck_counter_3[3]);
  assign readCrossBar_input_3_valid = selectExecuteReq_3_valid & tokenCheck_3;
  reg  [3:0]        tokenCheck_counter_4;
  wire [3:0]        tokenCheck_counterChange_4 = pipeReadFire_4 ? 4'h1 : 4'hF;
  wire              tokenCheck_4 = ~(tokenCheck_counter_4[3]);
  assign readCrossBar_input_4_valid = selectExecuteReq_4_valid & tokenCheck_4;
  reg  [3:0]        tokenCheck_counter_5;
  wire [3:0]        tokenCheck_counterChange_5 = pipeReadFire_5 ? 4'h1 : 4'hF;
  wire              tokenCheck_5 = ~(tokenCheck_counter_5[3]);
  assign readCrossBar_input_5_valid = selectExecuteReq_5_valid & tokenCheck_5;
  reg  [3:0]        tokenCheck_counter_6;
  wire [3:0]        tokenCheck_counterChange_6 = pipeReadFire_6 ? 4'h1 : 4'hF;
  wire              tokenCheck_6 = ~(tokenCheck_counter_6[3]);
  assign readCrossBar_input_6_valid = selectExecuteReq_6_valid & tokenCheck_6;
  reg  [3:0]        tokenCheck_counter_7;
  wire [3:0]        tokenCheck_counterChange_7 = pipeReadFire_7 ? 4'h1 : 4'hF;
  wire              tokenCheck_7 = ~(tokenCheck_counter_7[3]);
  assign readCrossBar_input_7_valid = selectExecuteReq_7_valid & tokenCheck_7;
  reg  [3:0]        tokenCheck_counter_8;
  wire [3:0]        tokenCheck_counterChange_8 = pipeReadFire_8 ? 4'h1 : 4'hF;
  wire              tokenCheck_8 = ~(tokenCheck_counter_8[3]);
  assign readCrossBar_input_8_valid = selectExecuteReq_8_valid & tokenCheck_8;
  reg  [3:0]        tokenCheck_counter_9;
  wire [3:0]        tokenCheck_counterChange_9 = pipeReadFire_9 ? 4'h1 : 4'hF;
  wire              tokenCheck_9 = ~(tokenCheck_counter_9[3]);
  assign readCrossBar_input_9_valid = selectExecuteReq_9_valid & tokenCheck_9;
  reg  [3:0]        tokenCheck_counter_10;
  wire [3:0]        tokenCheck_counterChange_10 = pipeReadFire_10 ? 4'h1 : 4'hF;
  wire              tokenCheck_10 = ~(tokenCheck_counter_10[3]);
  assign readCrossBar_input_10_valid = selectExecuteReq_10_valid & tokenCheck_10;
  reg  [3:0]        tokenCheck_counter_11;
  wire [3:0]        tokenCheck_counterChange_11 = pipeReadFire_11 ? 4'h1 : 4'hF;
  wire              tokenCheck_11 = ~(tokenCheck_counter_11[3]);
  assign readCrossBar_input_11_valid = selectExecuteReq_11_valid & tokenCheck_11;
  reg  [3:0]        tokenCheck_counter_12;
  wire [3:0]        tokenCheck_counterChange_12 = pipeReadFire_12 ? 4'h1 : 4'hF;
  wire              tokenCheck_12 = ~(tokenCheck_counter_12[3]);
  assign readCrossBar_input_12_valid = selectExecuteReq_12_valid & tokenCheck_12;
  reg  [3:0]        tokenCheck_counter_13;
  wire [3:0]        tokenCheck_counterChange_13 = pipeReadFire_13 ? 4'h1 : 4'hF;
  wire              tokenCheck_13 = ~(tokenCheck_counter_13[3]);
  assign readCrossBar_input_13_valid = selectExecuteReq_13_valid & tokenCheck_13;
  reg  [3:0]        tokenCheck_counter_14;
  wire [3:0]        tokenCheck_counterChange_14 = pipeReadFire_14 ? 4'h1 : 4'hF;
  wire              tokenCheck_14 = ~(tokenCheck_counter_14[3]);
  assign readCrossBar_input_14_valid = selectExecuteReq_14_valid & tokenCheck_14;
  reg  [3:0]        tokenCheck_counter_15;
  wire [3:0]        tokenCheck_counterChange_15 = pipeReadFire_15 ? 4'h1 : 4'hF;
  wire              tokenCheck_15 = ~(tokenCheck_counter_15[3]);
  assign readCrossBar_input_15_valid = selectExecuteReq_15_valid & tokenCheck_15;
  wire [1:0]        readFire_lo_lo_lo = {pipeReadFire_1, pipeReadFire_0};
  wire [1:0]        readFire_lo_lo_hi = {pipeReadFire_3, pipeReadFire_2};
  wire [3:0]        readFire_lo_lo = {readFire_lo_lo_hi, readFire_lo_lo_lo};
  wire [1:0]        readFire_lo_hi_lo = {pipeReadFire_5, pipeReadFire_4};
  wire [1:0]        readFire_lo_hi_hi = {pipeReadFire_7, pipeReadFire_6};
  wire [3:0]        readFire_lo_hi = {readFire_lo_hi_hi, readFire_lo_hi_lo};
  wire [7:0]        readFire_lo = {readFire_lo_hi, readFire_lo_lo};
  wire [1:0]        readFire_hi_lo_lo = {pipeReadFire_9, pipeReadFire_8};
  wire [1:0]        readFire_hi_lo_hi = {pipeReadFire_11, pipeReadFire_10};
  wire [3:0]        readFire_hi_lo = {readFire_hi_lo_hi, readFire_hi_lo_lo};
  wire [1:0]        readFire_hi_hi_lo = {pipeReadFire_13, pipeReadFire_12};
  wire [1:0]        readFire_hi_hi_hi = {pipeReadFire_15, pipeReadFire_14};
  wire [3:0]        readFire_hi_hi = {readFire_hi_hi_hi, readFire_hi_hi_lo};
  wire [7:0]        readFire_hi = {readFire_hi_hi, readFire_hi_lo};
  wire [15:0]       readFire = {readFire_hi, readFire_lo};
  wire              anyReadFire = |readFire;
  wire [15:0]       readStateUpdate = readFire | readIssueStageState_groupReadState;
  wire              groupReadFinish = readStateUpdate == readIssueStageState_needRead;
  assign readTypeRequestDeq = anyReadFire & groupReadFinish | readIssueStageValid & readIssueStageState_needRead == 16'h0;
  assign readWaitQueue_enq_valid = readTypeRequestDeq;
  wire [15:0]       compressUnitResultQueue_enq_bits_ffoOutput;
  wire              compressUnitResultQueue_enq_bits_compressValid;
  wire [16:0]       compressUnitResultQueue_dataIn_lo = {compressUnitResultQueue_enq_bits_ffoOutput, compressUnitResultQueue_enq_bits_compressValid};
  wire [511:0]      compressUnitResultQueue_enq_bits_data;
  wire [63:0]       compressUnitResultQueue_enq_bits_mask;
  wire [575:0]      compressUnitResultQueue_dataIn_hi_hi = {compressUnitResultQueue_enq_bits_data, compressUnitResultQueue_enq_bits_mask};
  wire [4:0]        compressUnitResultQueue_enq_bits_groupCounter;
  wire [580:0]      compressUnitResultQueue_dataIn_hi = {compressUnitResultQueue_dataIn_hi_hi, compressUnitResultQueue_enq_bits_groupCounter};
  wire [597:0]      compressUnitResultQueue_dataIn = {compressUnitResultQueue_dataIn_hi, compressUnitResultQueue_dataIn_lo};
  wire              compressUnitResultQueue_dataOut_compressValid = _compressUnitResultQueue_fifo_data_out[0];
  wire [15:0]       compressUnitResultQueue_dataOut_ffoOutput = _compressUnitResultQueue_fifo_data_out[16:1];
  wire [4:0]        compressUnitResultQueue_dataOut_groupCounter = _compressUnitResultQueue_fifo_data_out[21:17];
  wire [63:0]       compressUnitResultQueue_dataOut_mask = _compressUnitResultQueue_fifo_data_out[85:22];
  wire [511:0]      compressUnitResultQueue_dataOut_data = _compressUnitResultQueue_fifo_data_out[597:86];
  wire              compressUnitResultQueue_enq_ready = ~_compressUnitResultQueue_fifo_full;
  wire              compressUnitResultQueue_deq_ready;
  wire              compressUnitResultQueue_enq_valid;
  wire              compressUnitResultQueue_deq_valid = ~_compressUnitResultQueue_fifo_empty | compressUnitResultQueue_enq_valid;
  wire [511:0]      compressUnitResultQueue_deq_bits_data = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_data : compressUnitResultQueue_dataOut_data;
  wire [63:0]       compressUnitResultQueue_deq_bits_mask = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_mask : compressUnitResultQueue_dataOut_mask;
  wire [4:0]        compressUnitResultQueue_deq_bits_groupCounter = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_groupCounter : compressUnitResultQueue_dataOut_groupCounter;
  wire [15:0]       compressUnitResultQueue_deq_bits_ffoOutput = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_ffoOutput : compressUnitResultQueue_dataOut_ffoOutput;
  wire              compressUnitResultQueue_deq_bits_compressValid = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_compressValid : compressUnitResultQueue_dataOut_compressValid;
  wire              noSourceValid = noSource & counterValid & ((|instReg_vl) | mvRd & ~readVS1Reg_sendToExecution);
  wire              vs1DataValid = readVS1Reg_dataValid | ~(unitType[2] | _GEN_79);
  wire [1:0]        _GEN_81 = {_maskedWrite_in_1_ready, _maskedWrite_in_0_ready};
  wire [1:0]        executeDeqReady_lo_lo_lo;
  assign executeDeqReady_lo_lo_lo = _GEN_81;
  wire [1:0]        compressUnitResultQueue_deq_ready_lo_lo_lo;
  assign compressUnitResultQueue_deq_ready_lo_lo_lo = _GEN_81;
  wire [1:0]        _GEN_82 = {_maskedWrite_in_3_ready, _maskedWrite_in_2_ready};
  wire [1:0]        executeDeqReady_lo_lo_hi;
  assign executeDeqReady_lo_lo_hi = _GEN_82;
  wire [1:0]        compressUnitResultQueue_deq_ready_lo_lo_hi;
  assign compressUnitResultQueue_deq_ready_lo_lo_hi = _GEN_82;
  wire [3:0]        executeDeqReady_lo_lo = {executeDeqReady_lo_lo_hi, executeDeqReady_lo_lo_lo};
  wire [1:0]        _GEN_83 = {_maskedWrite_in_5_ready, _maskedWrite_in_4_ready};
  wire [1:0]        executeDeqReady_lo_hi_lo;
  assign executeDeqReady_lo_hi_lo = _GEN_83;
  wire [1:0]        compressUnitResultQueue_deq_ready_lo_hi_lo;
  assign compressUnitResultQueue_deq_ready_lo_hi_lo = _GEN_83;
  wire [1:0]        _GEN_84 = {_maskedWrite_in_7_ready, _maskedWrite_in_6_ready};
  wire [1:0]        executeDeqReady_lo_hi_hi;
  assign executeDeqReady_lo_hi_hi = _GEN_84;
  wire [1:0]        compressUnitResultQueue_deq_ready_lo_hi_hi;
  assign compressUnitResultQueue_deq_ready_lo_hi_hi = _GEN_84;
  wire [3:0]        executeDeqReady_lo_hi = {executeDeqReady_lo_hi_hi, executeDeqReady_lo_hi_lo};
  wire [7:0]        executeDeqReady_lo = {executeDeqReady_lo_hi, executeDeqReady_lo_lo};
  wire [1:0]        _GEN_85 = {_maskedWrite_in_9_ready, _maskedWrite_in_8_ready};
  wire [1:0]        executeDeqReady_hi_lo_lo;
  assign executeDeqReady_hi_lo_lo = _GEN_85;
  wire [1:0]        compressUnitResultQueue_deq_ready_hi_lo_lo;
  assign compressUnitResultQueue_deq_ready_hi_lo_lo = _GEN_85;
  wire [1:0]        _GEN_86 = {_maskedWrite_in_11_ready, _maskedWrite_in_10_ready};
  wire [1:0]        executeDeqReady_hi_lo_hi;
  assign executeDeqReady_hi_lo_hi = _GEN_86;
  wire [1:0]        compressUnitResultQueue_deq_ready_hi_lo_hi;
  assign compressUnitResultQueue_deq_ready_hi_lo_hi = _GEN_86;
  wire [3:0]        executeDeqReady_hi_lo = {executeDeqReady_hi_lo_hi, executeDeqReady_hi_lo_lo};
  wire [1:0]        _GEN_87 = {_maskedWrite_in_13_ready, _maskedWrite_in_12_ready};
  wire [1:0]        executeDeqReady_hi_hi_lo;
  assign executeDeqReady_hi_hi_lo = _GEN_87;
  wire [1:0]        compressUnitResultQueue_deq_ready_hi_hi_lo;
  assign compressUnitResultQueue_deq_ready_hi_hi_lo = _GEN_87;
  wire [1:0]        _GEN_88 = {_maskedWrite_in_15_ready, _maskedWrite_in_14_ready};
  wire [1:0]        executeDeqReady_hi_hi_hi;
  assign executeDeqReady_hi_hi_hi = _GEN_88;
  wire [1:0]        compressUnitResultQueue_deq_ready_hi_hi_hi;
  assign compressUnitResultQueue_deq_ready_hi_hi_hi = _GEN_88;
  wire [3:0]        executeDeqReady_hi_hi = {executeDeqReady_hi_hi_hi, executeDeqReady_hi_hi_lo};
  wire [7:0]        executeDeqReady_hi = {executeDeqReady_hi_hi, executeDeqReady_hi_lo};
  wire              compressUnitResultQueue_empty;
  wire              executeDeqReady = (&{executeDeqReady_hi, executeDeqReady_lo}) & compressUnitResultQueue_empty;
  wire              otherTypeRequestDeq = (noSource ? noSourceValid : allDataValid) & vs1DataValid & instVlValid & executeDeqReady;
  wire              reorderQueueAllocate;
  wire              _GEN_89 = accessCountQueue_enq_ready & reorderQueueAllocate;
  assign readIssueStageEnq = (allDataValid | _slideAddressGen_indexDeq_valid) & (readTypeRequestDeq | ~readIssueStageValid) & instVlValid & readType & _GEN_89;
  assign accessCountQueue_enq_valid = readIssueStageEnq;
  wire              executeReady;
  wire              requestStageDeq = readType ? readIssueStageEnq : otherTypeRequestDeq & executeReady;
  wire              slideAddressGen_indexDeq_ready = (readTypeRequestDeq | ~readIssueStageValid) & _GEN_89;
  wire              _GEN_90 = slideAddressGen_indexDeq_ready & _slideAddressGen_indexDeq_valid;
  wire              _GEN_91 = readIssueStageEnq & _GEN_90;
  assign accessCountEnq_0 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h0 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h0 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h0 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h0 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h0 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h0 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h0 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h0 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h0 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h0 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h0 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h0 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h0 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h0 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h0 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h0 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h0 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_1 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h1 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h1 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h1 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h1 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h1 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h1 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h1 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h1 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h1 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h1 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h1 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h1 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h1 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h1 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h1 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h1 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h1 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_2 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h2 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h2 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h2 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h2 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h2 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h2 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h2 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h2 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h2 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h2 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h2 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h2 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h2 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h2 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h2 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h2 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h2 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_3 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h3 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h3 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h3 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h3 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h3 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h3 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h3 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h3 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h3 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h3 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h3 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h3 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h3 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h3 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h3 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h3 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h3 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_4 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h4 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h4 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h4 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h4 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h4 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h4 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h4 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h4 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h4 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h4 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h4 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h4 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h4 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h4 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h4 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h4 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h4 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_5 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h5 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h5 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h5 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h5 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h5 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h5 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h5 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h5 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h5 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h5 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h5 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h5 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h5 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h5 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h5 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h5 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h5 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_6 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h6 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h6 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h6 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h6 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h6 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h6 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h6 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h6 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h6 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h6 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h6 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h6 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h6 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h6 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h6 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h6 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h6 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_7 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h7 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h7 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h7 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h7 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h7 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h7 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h7 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h7 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h7 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h7 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h7 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h7 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h7 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h7 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h7 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h7 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h7 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_8 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h8 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h8 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h8 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h8 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h8 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h8 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h8 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h8 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h8 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h8 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h8 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h8 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h8 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h8 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h8 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h8 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h8 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_9 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'h9 & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'h9 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'h9 & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'h9 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'h9 & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'h9 & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'h9 & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'h9 & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'h9 & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'h9 & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'h9 & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'h9 & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'h9 & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'h9 & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'h9 & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'h9 & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'h9 & ~(notReadSelect[15])}}}};
  assign accessCountEnq_10 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'hA & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'hA & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'hA & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'hA & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'hA & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'hA & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'hA & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'hA & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'hA & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'hA & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'hA & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'hA & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'hA & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'hA & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'hA & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'hA & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'hA & ~(notReadSelect[15])}}}};
  assign accessCountEnq_11 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'hB & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'hB & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'hB & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'hB & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'hB & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'hB & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'hB & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'hB & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'hB & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'hB & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'hB & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'hB & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'hB & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'hB & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'hB & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'hB & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'hB & ~(notReadSelect[15])}}}};
  assign accessCountEnq_12 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'hC & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'hC & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'hC & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'hC & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'hC & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'hC & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'hC & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'hC & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'hC & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'hC & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'hC & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'hC & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'hC & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'hC & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'hC & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'hC & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'hC & ~(notReadSelect[15])}}}};
  assign accessCountEnq_13 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'hD & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'hD & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'hD & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'hD & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'hD & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'hD & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'hD & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'hD & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'hD & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'hD & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'hD & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'hD & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'hD & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'hD & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'hD & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'hD & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'hD & ~(notReadSelect[15])}}}};
  assign accessCountEnq_14 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_4 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_5 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_6 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_7 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_8 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_9 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_10 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_11 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_12 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_13 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0,
                     {1'h0, _slideAddressGen_indexDeq_bits_accessLane_14 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_15 == 4'hE & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, accessLaneSelect[3:0] == 4'hE & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[7:4] == 4'hE & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, accessLaneSelect[11:8] == 4'hE & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[15:12] == 4'hE & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, accessLaneSelect[19:16] == 4'hE & ~(notReadSelect[4])} + {1'h0, accessLaneSelect[23:20] == 4'hE & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, accessLaneSelect[27:24] == 4'hE & ~(notReadSelect[6])} + {1'h0, accessLaneSelect[31:28] == 4'hE & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, accessLaneSelect[35:32] == 4'hE & ~(notReadSelect[8])} + {1'h0, accessLaneSelect[39:36] == 4'hE & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, accessLaneSelect[43:40] == 4'hE & ~(notReadSelect[10])} + {1'h0, accessLaneSelect[47:44] == 4'hE & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, accessLaneSelect[51:48] == 4'hE & ~(notReadSelect[12])} + {1'h0, accessLaneSelect[55:52] == 4'hE & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, accessLaneSelect[59:56] == 4'hE & ~(notReadSelect[14])} + {1'h0, accessLaneSelect[63:60] == 4'hE & ~(notReadSelect[15])}}}};
  assign accessCountEnq_15 =
    _GEN_91
      ? {1'h0,
         {1'h0,
          {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_0) & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_1) & _slideAddressGen_indexDeq_bits_needRead[1]}}
            + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_2) & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_3) & _slideAddressGen_indexDeq_bits_needRead[3]}}}
           + {1'h0,
              {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_4) & _slideAddressGen_indexDeq_bits_needRead[4]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_5) & _slideAddressGen_indexDeq_bits_needRead[5]}}
                + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_6) & _slideAddressGen_indexDeq_bits_needRead[6]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_7) & _slideAddressGen_indexDeq_bits_needRead[7]}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_8) & _slideAddressGen_indexDeq_bits_needRead[8]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_9) & _slideAddressGen_indexDeq_bits_needRead[9]}}
              + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_10) & _slideAddressGen_indexDeq_bits_needRead[10]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_11) & _slideAddressGen_indexDeq_bits_needRead[11]}}}
             + {1'h0,
                {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_12) & _slideAddressGen_indexDeq_bits_needRead[12]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_13) & _slideAddressGen_indexDeq_bits_needRead[13]}}
                  + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_14) & _slideAddressGen_indexDeq_bits_needRead[14]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_15) & _slideAddressGen_indexDeq_bits_needRead[15]}}}}
      : {1'h0,
         {1'h0,
          {1'h0, {1'h0, (&(accessLaneSelect[3:0])) & ~(notReadSelect[0])} + {1'h0, (&(accessLaneSelect[7:4])) & ~(notReadSelect[1])}}
            + {1'h0, {1'h0, (&(accessLaneSelect[11:8])) & ~(notReadSelect[2])} + {1'h0, (&(accessLaneSelect[15:12])) & ~(notReadSelect[3])}}}
           + {1'h0,
              {1'h0, {1'h0, (&(accessLaneSelect[19:16])) & ~(notReadSelect[4])} + {1'h0, (&(accessLaneSelect[23:20])) & ~(notReadSelect[5])}}
                + {1'h0, {1'h0, (&(accessLaneSelect[27:24])) & ~(notReadSelect[6])} + {1'h0, (&(accessLaneSelect[31:28])) & ~(notReadSelect[7])}}}}
        + {1'h0,
           {1'h0,
            {1'h0, {1'h0, (&(accessLaneSelect[35:32])) & ~(notReadSelect[8])} + {1'h0, (&(accessLaneSelect[39:36])) & ~(notReadSelect[9])}}
              + {1'h0, {1'h0, (&(accessLaneSelect[43:40])) & ~(notReadSelect[10])} + {1'h0, (&(accessLaneSelect[47:44])) & ~(notReadSelect[11])}}}
             + {1'h0,
                {1'h0, {1'h0, (&(accessLaneSelect[51:48])) & ~(notReadSelect[12])} + {1'h0, (&(accessLaneSelect[55:52])) & ~(notReadSelect[13])}}
                  + {1'h0, {1'h0, (&(accessLaneSelect[59:56])) & ~(notReadSelect[14])} + {1'h0, (&(accessLaneSelect[63:60])) & ~(notReadSelect[15])}}}};
  assign lastExecuteGroupDeq = requestStageDeq & isLastExecuteGroup;
  wire [15:0]       readMessageQueue_deq_bits_readSource;
  wire              deqAllocate;
  wire              reorderQueueVec_0_deq_valid;
  assign reorderQueueVec_0_deq_valid = ~_reorderQueueVec_fifo_empty;
  wire [31:0]       reorderQueueVec_dataOut_data;
  wire [15:0]       reorderQueueVec_dataOut_write1H;
  wire [31:0]       dataAfterReorderCheck_0 = reorderQueueVec_0_deq_bits_data;
  wire [31:0]       reorderQueueVec_0_enq_bits_data;
  wire [15:0]       reorderQueueVec_0_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn = {reorderQueueVec_0_enq_bits_data, reorderQueueVec_0_enq_bits_write1H};
  assign reorderQueueVec_dataOut_write1H = _reorderQueueVec_fifo_data_out[15:0];
  assign reorderQueueVec_dataOut_data = _reorderQueueVec_fifo_data_out[47:16];
  assign reorderQueueVec_0_deq_bits_data = reorderQueueVec_dataOut_data;
  wire [15:0]       reorderQueueVec_0_deq_bits_write1H = reorderQueueVec_dataOut_write1H;
  wire              reorderQueueVec_0_enq_ready = ~_reorderQueueVec_fifo_full;
  wire              reorderQueueVec_0_deq_ready;
  wire [15:0]       readMessageQueue_1_deq_bits_readSource;
  wire              deqAllocate_1;
  wire              reorderQueueVec_1_deq_valid;
  assign reorderQueueVec_1_deq_valid = ~_reorderQueueVec_fifo_1_empty;
  wire [31:0]       reorderQueueVec_dataOut_1_data;
  wire [15:0]       reorderQueueVec_dataOut_1_write1H;
  wire [31:0]       dataAfterReorderCheck_1 = reorderQueueVec_1_deq_bits_data;
  wire [31:0]       reorderQueueVec_1_enq_bits_data;
  wire [15:0]       reorderQueueVec_1_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_1 = {reorderQueueVec_1_enq_bits_data, reorderQueueVec_1_enq_bits_write1H};
  assign reorderQueueVec_dataOut_1_write1H = _reorderQueueVec_fifo_1_data_out[15:0];
  assign reorderQueueVec_dataOut_1_data = _reorderQueueVec_fifo_1_data_out[47:16];
  assign reorderQueueVec_1_deq_bits_data = reorderQueueVec_dataOut_1_data;
  wire [15:0]       reorderQueueVec_1_deq_bits_write1H = reorderQueueVec_dataOut_1_write1H;
  wire              reorderQueueVec_1_enq_ready = ~_reorderQueueVec_fifo_1_full;
  wire              reorderQueueVec_1_deq_ready;
  wire [15:0]       readMessageQueue_2_deq_bits_readSource;
  wire              deqAllocate_2;
  wire              reorderQueueVec_2_deq_valid;
  assign reorderQueueVec_2_deq_valid = ~_reorderQueueVec_fifo_2_empty;
  wire [31:0]       reorderQueueVec_dataOut_2_data;
  wire [15:0]       reorderQueueVec_dataOut_2_write1H;
  wire [31:0]       dataAfterReorderCheck_2 = reorderQueueVec_2_deq_bits_data;
  wire [31:0]       reorderQueueVec_2_enq_bits_data;
  wire [15:0]       reorderQueueVec_2_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_2 = {reorderQueueVec_2_enq_bits_data, reorderQueueVec_2_enq_bits_write1H};
  assign reorderQueueVec_dataOut_2_write1H = _reorderQueueVec_fifo_2_data_out[15:0];
  assign reorderQueueVec_dataOut_2_data = _reorderQueueVec_fifo_2_data_out[47:16];
  assign reorderQueueVec_2_deq_bits_data = reorderQueueVec_dataOut_2_data;
  wire [15:0]       reorderQueueVec_2_deq_bits_write1H = reorderQueueVec_dataOut_2_write1H;
  wire              reorderQueueVec_2_enq_ready = ~_reorderQueueVec_fifo_2_full;
  wire              reorderQueueVec_2_deq_ready;
  wire [15:0]       readMessageQueue_3_deq_bits_readSource;
  wire              deqAllocate_3;
  wire              reorderQueueVec_3_deq_valid;
  assign reorderQueueVec_3_deq_valid = ~_reorderQueueVec_fifo_3_empty;
  wire [31:0]       reorderQueueVec_dataOut_3_data;
  wire [15:0]       reorderQueueVec_dataOut_3_write1H;
  wire [31:0]       dataAfterReorderCheck_3 = reorderQueueVec_3_deq_bits_data;
  wire [31:0]       reorderQueueVec_3_enq_bits_data;
  wire [15:0]       reorderQueueVec_3_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_3 = {reorderQueueVec_3_enq_bits_data, reorderQueueVec_3_enq_bits_write1H};
  assign reorderQueueVec_dataOut_3_write1H = _reorderQueueVec_fifo_3_data_out[15:0];
  assign reorderQueueVec_dataOut_3_data = _reorderQueueVec_fifo_3_data_out[47:16];
  assign reorderQueueVec_3_deq_bits_data = reorderQueueVec_dataOut_3_data;
  wire [15:0]       reorderQueueVec_3_deq_bits_write1H = reorderQueueVec_dataOut_3_write1H;
  wire              reorderQueueVec_3_enq_ready = ~_reorderQueueVec_fifo_3_full;
  wire              reorderQueueVec_3_deq_ready;
  wire [15:0]       readMessageQueue_4_deq_bits_readSource;
  wire              deqAllocate_4;
  wire              reorderQueueVec_4_deq_valid;
  assign reorderQueueVec_4_deq_valid = ~_reorderQueueVec_fifo_4_empty;
  wire [31:0]       reorderQueueVec_dataOut_4_data;
  wire [15:0]       reorderQueueVec_dataOut_4_write1H;
  wire [31:0]       dataAfterReorderCheck_4 = reorderQueueVec_4_deq_bits_data;
  wire [31:0]       reorderQueueVec_4_enq_bits_data;
  wire [15:0]       reorderQueueVec_4_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_4 = {reorderQueueVec_4_enq_bits_data, reorderQueueVec_4_enq_bits_write1H};
  assign reorderQueueVec_dataOut_4_write1H = _reorderQueueVec_fifo_4_data_out[15:0];
  assign reorderQueueVec_dataOut_4_data = _reorderQueueVec_fifo_4_data_out[47:16];
  assign reorderQueueVec_4_deq_bits_data = reorderQueueVec_dataOut_4_data;
  wire [15:0]       reorderQueueVec_4_deq_bits_write1H = reorderQueueVec_dataOut_4_write1H;
  wire              reorderQueueVec_4_enq_ready = ~_reorderQueueVec_fifo_4_full;
  wire              reorderQueueVec_4_deq_ready;
  wire [15:0]       readMessageQueue_5_deq_bits_readSource;
  wire              deqAllocate_5;
  wire              reorderQueueVec_5_deq_valid;
  assign reorderQueueVec_5_deq_valid = ~_reorderQueueVec_fifo_5_empty;
  wire [31:0]       reorderQueueVec_dataOut_5_data;
  wire [15:0]       reorderQueueVec_dataOut_5_write1H;
  wire [31:0]       dataAfterReorderCheck_5 = reorderQueueVec_5_deq_bits_data;
  wire [31:0]       reorderQueueVec_5_enq_bits_data;
  wire [15:0]       reorderQueueVec_5_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_5 = {reorderQueueVec_5_enq_bits_data, reorderQueueVec_5_enq_bits_write1H};
  assign reorderQueueVec_dataOut_5_write1H = _reorderQueueVec_fifo_5_data_out[15:0];
  assign reorderQueueVec_dataOut_5_data = _reorderQueueVec_fifo_5_data_out[47:16];
  assign reorderQueueVec_5_deq_bits_data = reorderQueueVec_dataOut_5_data;
  wire [15:0]       reorderQueueVec_5_deq_bits_write1H = reorderQueueVec_dataOut_5_write1H;
  wire              reorderQueueVec_5_enq_ready = ~_reorderQueueVec_fifo_5_full;
  wire              reorderQueueVec_5_deq_ready;
  wire [15:0]       readMessageQueue_6_deq_bits_readSource;
  wire              deqAllocate_6;
  wire              reorderQueueVec_6_deq_valid;
  assign reorderQueueVec_6_deq_valid = ~_reorderQueueVec_fifo_6_empty;
  wire [31:0]       reorderQueueVec_dataOut_6_data;
  wire [15:0]       reorderQueueVec_dataOut_6_write1H;
  wire [31:0]       dataAfterReorderCheck_6 = reorderQueueVec_6_deq_bits_data;
  wire [31:0]       reorderQueueVec_6_enq_bits_data;
  wire [15:0]       reorderQueueVec_6_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_6 = {reorderQueueVec_6_enq_bits_data, reorderQueueVec_6_enq_bits_write1H};
  assign reorderQueueVec_dataOut_6_write1H = _reorderQueueVec_fifo_6_data_out[15:0];
  assign reorderQueueVec_dataOut_6_data = _reorderQueueVec_fifo_6_data_out[47:16];
  assign reorderQueueVec_6_deq_bits_data = reorderQueueVec_dataOut_6_data;
  wire [15:0]       reorderQueueVec_6_deq_bits_write1H = reorderQueueVec_dataOut_6_write1H;
  wire              reorderQueueVec_6_enq_ready = ~_reorderQueueVec_fifo_6_full;
  wire              reorderQueueVec_6_deq_ready;
  wire [15:0]       readMessageQueue_7_deq_bits_readSource;
  wire              deqAllocate_7;
  wire              reorderQueueVec_7_deq_valid;
  assign reorderQueueVec_7_deq_valid = ~_reorderQueueVec_fifo_7_empty;
  wire [31:0]       reorderQueueVec_dataOut_7_data;
  wire [15:0]       reorderQueueVec_dataOut_7_write1H;
  wire [31:0]       dataAfterReorderCheck_7 = reorderQueueVec_7_deq_bits_data;
  wire [31:0]       reorderQueueVec_7_enq_bits_data;
  wire [15:0]       reorderQueueVec_7_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_7 = {reorderQueueVec_7_enq_bits_data, reorderQueueVec_7_enq_bits_write1H};
  assign reorderQueueVec_dataOut_7_write1H = _reorderQueueVec_fifo_7_data_out[15:0];
  assign reorderQueueVec_dataOut_7_data = _reorderQueueVec_fifo_7_data_out[47:16];
  assign reorderQueueVec_7_deq_bits_data = reorderQueueVec_dataOut_7_data;
  wire [15:0]       reorderQueueVec_7_deq_bits_write1H = reorderQueueVec_dataOut_7_write1H;
  wire              reorderQueueVec_7_enq_ready = ~_reorderQueueVec_fifo_7_full;
  wire              reorderQueueVec_7_deq_ready;
  wire [15:0]       readMessageQueue_8_deq_bits_readSource;
  wire              deqAllocate_8;
  wire              reorderQueueVec_8_deq_valid;
  assign reorderQueueVec_8_deq_valid = ~_reorderQueueVec_fifo_8_empty;
  wire [31:0]       reorderQueueVec_dataOut_8_data;
  wire [15:0]       reorderQueueVec_dataOut_8_write1H;
  wire [31:0]       dataAfterReorderCheck_8 = reorderQueueVec_8_deq_bits_data;
  wire [31:0]       reorderQueueVec_8_enq_bits_data;
  wire [15:0]       reorderQueueVec_8_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_8 = {reorderQueueVec_8_enq_bits_data, reorderQueueVec_8_enq_bits_write1H};
  assign reorderQueueVec_dataOut_8_write1H = _reorderQueueVec_fifo_8_data_out[15:0];
  assign reorderQueueVec_dataOut_8_data = _reorderQueueVec_fifo_8_data_out[47:16];
  assign reorderQueueVec_8_deq_bits_data = reorderQueueVec_dataOut_8_data;
  wire [15:0]       reorderQueueVec_8_deq_bits_write1H = reorderQueueVec_dataOut_8_write1H;
  wire              reorderQueueVec_8_enq_ready = ~_reorderQueueVec_fifo_8_full;
  wire              reorderQueueVec_8_deq_ready;
  wire [15:0]       readMessageQueue_9_deq_bits_readSource;
  wire              deqAllocate_9;
  wire              reorderQueueVec_9_deq_valid;
  assign reorderQueueVec_9_deq_valid = ~_reorderQueueVec_fifo_9_empty;
  wire [31:0]       reorderQueueVec_dataOut_9_data;
  wire [15:0]       reorderQueueVec_dataOut_9_write1H;
  wire [31:0]       dataAfterReorderCheck_9 = reorderQueueVec_9_deq_bits_data;
  wire [31:0]       reorderQueueVec_9_enq_bits_data;
  wire [15:0]       reorderQueueVec_9_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_9 = {reorderQueueVec_9_enq_bits_data, reorderQueueVec_9_enq_bits_write1H};
  assign reorderQueueVec_dataOut_9_write1H = _reorderQueueVec_fifo_9_data_out[15:0];
  assign reorderQueueVec_dataOut_9_data = _reorderQueueVec_fifo_9_data_out[47:16];
  assign reorderQueueVec_9_deq_bits_data = reorderQueueVec_dataOut_9_data;
  wire [15:0]       reorderQueueVec_9_deq_bits_write1H = reorderQueueVec_dataOut_9_write1H;
  wire              reorderQueueVec_9_enq_ready = ~_reorderQueueVec_fifo_9_full;
  wire              reorderQueueVec_9_deq_ready;
  wire [15:0]       readMessageQueue_10_deq_bits_readSource;
  wire              deqAllocate_10;
  wire              reorderQueueVec_10_deq_valid;
  assign reorderQueueVec_10_deq_valid = ~_reorderQueueVec_fifo_10_empty;
  wire [31:0]       reorderQueueVec_dataOut_10_data;
  wire [15:0]       reorderQueueVec_dataOut_10_write1H;
  wire [31:0]       dataAfterReorderCheck_10 = reorderQueueVec_10_deq_bits_data;
  wire [31:0]       reorderQueueVec_10_enq_bits_data;
  wire [15:0]       reorderQueueVec_10_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_10 = {reorderQueueVec_10_enq_bits_data, reorderQueueVec_10_enq_bits_write1H};
  assign reorderQueueVec_dataOut_10_write1H = _reorderQueueVec_fifo_10_data_out[15:0];
  assign reorderQueueVec_dataOut_10_data = _reorderQueueVec_fifo_10_data_out[47:16];
  assign reorderQueueVec_10_deq_bits_data = reorderQueueVec_dataOut_10_data;
  wire [15:0]       reorderQueueVec_10_deq_bits_write1H = reorderQueueVec_dataOut_10_write1H;
  wire              reorderQueueVec_10_enq_ready = ~_reorderQueueVec_fifo_10_full;
  wire              reorderQueueVec_10_deq_ready;
  wire [15:0]       readMessageQueue_11_deq_bits_readSource;
  wire              deqAllocate_11;
  wire              reorderQueueVec_11_deq_valid;
  assign reorderQueueVec_11_deq_valid = ~_reorderQueueVec_fifo_11_empty;
  wire [31:0]       reorderQueueVec_dataOut_11_data;
  wire [15:0]       reorderQueueVec_dataOut_11_write1H;
  wire [31:0]       dataAfterReorderCheck_11 = reorderQueueVec_11_deq_bits_data;
  wire [31:0]       reorderQueueVec_11_enq_bits_data;
  wire [15:0]       reorderQueueVec_11_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_11 = {reorderQueueVec_11_enq_bits_data, reorderQueueVec_11_enq_bits_write1H};
  assign reorderQueueVec_dataOut_11_write1H = _reorderQueueVec_fifo_11_data_out[15:0];
  assign reorderQueueVec_dataOut_11_data = _reorderQueueVec_fifo_11_data_out[47:16];
  assign reorderQueueVec_11_deq_bits_data = reorderQueueVec_dataOut_11_data;
  wire [15:0]       reorderQueueVec_11_deq_bits_write1H = reorderQueueVec_dataOut_11_write1H;
  wire              reorderQueueVec_11_enq_ready = ~_reorderQueueVec_fifo_11_full;
  wire              reorderQueueVec_11_deq_ready;
  wire [15:0]       readMessageQueue_12_deq_bits_readSource;
  wire              deqAllocate_12;
  wire              reorderQueueVec_12_deq_valid;
  assign reorderQueueVec_12_deq_valid = ~_reorderQueueVec_fifo_12_empty;
  wire [31:0]       reorderQueueVec_dataOut_12_data;
  wire [15:0]       reorderQueueVec_dataOut_12_write1H;
  wire [31:0]       dataAfterReorderCheck_12 = reorderQueueVec_12_deq_bits_data;
  wire [31:0]       reorderQueueVec_12_enq_bits_data;
  wire [15:0]       reorderQueueVec_12_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_12 = {reorderQueueVec_12_enq_bits_data, reorderQueueVec_12_enq_bits_write1H};
  assign reorderQueueVec_dataOut_12_write1H = _reorderQueueVec_fifo_12_data_out[15:0];
  assign reorderQueueVec_dataOut_12_data = _reorderQueueVec_fifo_12_data_out[47:16];
  assign reorderQueueVec_12_deq_bits_data = reorderQueueVec_dataOut_12_data;
  wire [15:0]       reorderQueueVec_12_deq_bits_write1H = reorderQueueVec_dataOut_12_write1H;
  wire              reorderQueueVec_12_enq_ready = ~_reorderQueueVec_fifo_12_full;
  wire              reorderQueueVec_12_deq_ready;
  wire [15:0]       readMessageQueue_13_deq_bits_readSource;
  wire              deqAllocate_13;
  wire              reorderQueueVec_13_deq_valid;
  assign reorderQueueVec_13_deq_valid = ~_reorderQueueVec_fifo_13_empty;
  wire [31:0]       reorderQueueVec_dataOut_13_data;
  wire [15:0]       reorderQueueVec_dataOut_13_write1H;
  wire [31:0]       dataAfterReorderCheck_13 = reorderQueueVec_13_deq_bits_data;
  wire [31:0]       reorderQueueVec_13_enq_bits_data;
  wire [15:0]       reorderQueueVec_13_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_13 = {reorderQueueVec_13_enq_bits_data, reorderQueueVec_13_enq_bits_write1H};
  assign reorderQueueVec_dataOut_13_write1H = _reorderQueueVec_fifo_13_data_out[15:0];
  assign reorderQueueVec_dataOut_13_data = _reorderQueueVec_fifo_13_data_out[47:16];
  assign reorderQueueVec_13_deq_bits_data = reorderQueueVec_dataOut_13_data;
  wire [15:0]       reorderQueueVec_13_deq_bits_write1H = reorderQueueVec_dataOut_13_write1H;
  wire              reorderQueueVec_13_enq_ready = ~_reorderQueueVec_fifo_13_full;
  wire              reorderQueueVec_13_deq_ready;
  wire [15:0]       readMessageQueue_14_deq_bits_readSource;
  wire              deqAllocate_14;
  wire              reorderQueueVec_14_deq_valid;
  assign reorderQueueVec_14_deq_valid = ~_reorderQueueVec_fifo_14_empty;
  wire [31:0]       reorderQueueVec_dataOut_14_data;
  wire [15:0]       reorderQueueVec_dataOut_14_write1H;
  wire [31:0]       dataAfterReorderCheck_14 = reorderQueueVec_14_deq_bits_data;
  wire [31:0]       reorderQueueVec_14_enq_bits_data;
  wire [15:0]       reorderQueueVec_14_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_14 = {reorderQueueVec_14_enq_bits_data, reorderQueueVec_14_enq_bits_write1H};
  assign reorderQueueVec_dataOut_14_write1H = _reorderQueueVec_fifo_14_data_out[15:0];
  assign reorderQueueVec_dataOut_14_data = _reorderQueueVec_fifo_14_data_out[47:16];
  assign reorderQueueVec_14_deq_bits_data = reorderQueueVec_dataOut_14_data;
  wire [15:0]       reorderQueueVec_14_deq_bits_write1H = reorderQueueVec_dataOut_14_write1H;
  wire              reorderQueueVec_14_enq_ready = ~_reorderQueueVec_fifo_14_full;
  wire              reorderQueueVec_14_deq_ready;
  wire [15:0]       readMessageQueue_15_deq_bits_readSource;
  wire              deqAllocate_15;
  wire              reorderQueueVec_15_deq_valid;
  assign reorderQueueVec_15_deq_valid = ~_reorderQueueVec_fifo_15_empty;
  wire [31:0]       reorderQueueVec_dataOut_15_data;
  wire [15:0]       reorderQueueVec_dataOut_15_write1H;
  wire [31:0]       dataAfterReorderCheck_15 = reorderQueueVec_15_deq_bits_data;
  wire [31:0]       reorderQueueVec_15_enq_bits_data;
  wire [15:0]       reorderQueueVec_15_enq_bits_write1H;
  wire [47:0]       reorderQueueVec_dataIn_15 = {reorderQueueVec_15_enq_bits_data, reorderQueueVec_15_enq_bits_write1H};
  assign reorderQueueVec_dataOut_15_write1H = _reorderQueueVec_fifo_15_data_out[15:0];
  assign reorderQueueVec_dataOut_15_data = _reorderQueueVec_fifo_15_data_out[47:16];
  assign reorderQueueVec_15_deq_bits_data = reorderQueueVec_dataOut_15_data;
  wire [15:0]       reorderQueueVec_15_deq_bits_write1H = reorderQueueVec_dataOut_15_write1H;
  wire              reorderQueueVec_15_enq_ready = ~_reorderQueueVec_fifo_15_full;
  wire              reorderQueueVec_15_deq_ready;
  reg  [5:0]        reorderQueueAllocate_counter;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate;
  wire              _write1HPipe_0_T = reorderQueueVec_0_deq_ready & reorderQueueVec_0_deq_valid;
  wire              reorderQueueAllocate_release = _write1HPipe_0_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate = readIssueStageEnq ? accessCountEnq_0 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate = reorderQueueAllocate_counter + {1'h0, reorderQueueAllocate_allocate} - {5'h0, reorderQueueAllocate_release};
  reg  [5:0]        reorderQueueAllocate_counter_1;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_1;
  wire              _write1HPipe_1_T = reorderQueueVec_1_deq_ready & reorderQueueVec_1_deq_valid;
  wire              reorderQueueAllocate_release_1 = _write1HPipe_1_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_1 = readIssueStageEnq ? accessCountEnq_1 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_1 = reorderQueueAllocate_counter_1 + {1'h0, reorderQueueAllocate_allocate_1} - {5'h0, reorderQueueAllocate_release_1};
  reg  [5:0]        reorderQueueAllocate_counter_2;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_2;
  wire              _write1HPipe_2_T = reorderQueueVec_2_deq_ready & reorderQueueVec_2_deq_valid;
  wire              reorderQueueAllocate_release_2 = _write1HPipe_2_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_2 = readIssueStageEnq ? accessCountEnq_2 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_2 = reorderQueueAllocate_counter_2 + {1'h0, reorderQueueAllocate_allocate_2} - {5'h0, reorderQueueAllocate_release_2};
  reg  [5:0]        reorderQueueAllocate_counter_3;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_3;
  wire              _write1HPipe_3_T = reorderQueueVec_3_deq_ready & reorderQueueVec_3_deq_valid;
  wire              reorderQueueAllocate_release_3 = _write1HPipe_3_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_3 = readIssueStageEnq ? accessCountEnq_3 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_3 = reorderQueueAllocate_counter_3 + {1'h0, reorderQueueAllocate_allocate_3} - {5'h0, reorderQueueAllocate_release_3};
  reg  [5:0]        reorderQueueAllocate_counter_4;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_4;
  wire              _write1HPipe_4_T = reorderQueueVec_4_deq_ready & reorderQueueVec_4_deq_valid;
  wire              reorderQueueAllocate_release_4 = _write1HPipe_4_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_4 = readIssueStageEnq ? accessCountEnq_4 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_4 = reorderQueueAllocate_counter_4 + {1'h0, reorderQueueAllocate_allocate_4} - {5'h0, reorderQueueAllocate_release_4};
  reg  [5:0]        reorderQueueAllocate_counter_5;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_5;
  wire              _write1HPipe_5_T = reorderQueueVec_5_deq_ready & reorderQueueVec_5_deq_valid;
  wire              reorderQueueAllocate_release_5 = _write1HPipe_5_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_5 = readIssueStageEnq ? accessCountEnq_5 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_5 = reorderQueueAllocate_counter_5 + {1'h0, reorderQueueAllocate_allocate_5} - {5'h0, reorderQueueAllocate_release_5};
  reg  [5:0]        reorderQueueAllocate_counter_6;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_6;
  wire              _write1HPipe_6_T = reorderQueueVec_6_deq_ready & reorderQueueVec_6_deq_valid;
  wire              reorderQueueAllocate_release_6 = _write1HPipe_6_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_6 = readIssueStageEnq ? accessCountEnq_6 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_6 = reorderQueueAllocate_counter_6 + {1'h0, reorderQueueAllocate_allocate_6} - {5'h0, reorderQueueAllocate_release_6};
  reg  [5:0]        reorderQueueAllocate_counter_7;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_7;
  wire              _write1HPipe_7_T = reorderQueueVec_7_deq_ready & reorderQueueVec_7_deq_valid;
  wire              reorderQueueAllocate_release_7 = _write1HPipe_7_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_7 = readIssueStageEnq ? accessCountEnq_7 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_7 = reorderQueueAllocate_counter_7 + {1'h0, reorderQueueAllocate_allocate_7} - {5'h0, reorderQueueAllocate_release_7};
  reg  [5:0]        reorderQueueAllocate_counter_8;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_8;
  wire              _write1HPipe_8_T = reorderQueueVec_8_deq_ready & reorderQueueVec_8_deq_valid;
  wire              reorderQueueAllocate_release_8 = _write1HPipe_8_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_8 = readIssueStageEnq ? accessCountEnq_8 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_8 = reorderQueueAllocate_counter_8 + {1'h0, reorderQueueAllocate_allocate_8} - {5'h0, reorderQueueAllocate_release_8};
  reg  [5:0]        reorderQueueAllocate_counter_9;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_9;
  wire              _write1HPipe_9_T = reorderQueueVec_9_deq_ready & reorderQueueVec_9_deq_valid;
  wire              reorderQueueAllocate_release_9 = _write1HPipe_9_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_9 = readIssueStageEnq ? accessCountEnq_9 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_9 = reorderQueueAllocate_counter_9 + {1'h0, reorderQueueAllocate_allocate_9} - {5'h0, reorderQueueAllocate_release_9};
  reg  [5:0]        reorderQueueAllocate_counter_10;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_10;
  wire              _write1HPipe_10_T = reorderQueueVec_10_deq_ready & reorderQueueVec_10_deq_valid;
  wire              reorderQueueAllocate_release_10 = _write1HPipe_10_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_10 = readIssueStageEnq ? accessCountEnq_10 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_10 = reorderQueueAllocate_counter_10 + {1'h0, reorderQueueAllocate_allocate_10} - {5'h0, reorderQueueAllocate_release_10};
  reg  [5:0]        reorderQueueAllocate_counter_11;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_11;
  wire              _write1HPipe_11_T = reorderQueueVec_11_deq_ready & reorderQueueVec_11_deq_valid;
  wire              reorderQueueAllocate_release_11 = _write1HPipe_11_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_11 = readIssueStageEnq ? accessCountEnq_11 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_11 = reorderQueueAllocate_counter_11 + {1'h0, reorderQueueAllocate_allocate_11} - {5'h0, reorderQueueAllocate_release_11};
  reg  [5:0]        reorderQueueAllocate_counter_12;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_12;
  wire              _write1HPipe_12_T = reorderQueueVec_12_deq_ready & reorderQueueVec_12_deq_valid;
  wire              reorderQueueAllocate_release_12 = _write1HPipe_12_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_12 = readIssueStageEnq ? accessCountEnq_12 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_12 = reorderQueueAllocate_counter_12 + {1'h0, reorderQueueAllocate_allocate_12} - {5'h0, reorderQueueAllocate_release_12};
  reg  [5:0]        reorderQueueAllocate_counter_13;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_13;
  wire              _write1HPipe_13_T = reorderQueueVec_13_deq_ready & reorderQueueVec_13_deq_valid;
  wire              reorderQueueAllocate_release_13 = _write1HPipe_13_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_13 = readIssueStageEnq ? accessCountEnq_13 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_13 = reorderQueueAllocate_counter_13 + {1'h0, reorderQueueAllocate_allocate_13} - {5'h0, reorderQueueAllocate_release_13};
  reg  [5:0]        reorderQueueAllocate_counter_14;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_14;
  wire              _write1HPipe_14_T = reorderQueueVec_14_deq_ready & reorderQueueVec_14_deq_valid;
  wire              reorderQueueAllocate_release_14 = _write1HPipe_14_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_14 = readIssueStageEnq ? accessCountEnq_14 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_14 = reorderQueueAllocate_counter_14 + {1'h0, reorderQueueAllocate_allocate_14} - {5'h0, reorderQueueAllocate_release_14};
  reg  [5:0]        reorderQueueAllocate_counter_15;
  reg  [5:0]        reorderQueueAllocate_counterWillUpdate_15;
  wire              _write1HPipe_15_T = reorderQueueVec_15_deq_ready & reorderQueueVec_15_deq_valid;
  wire              reorderQueueAllocate_release_15 = _write1HPipe_15_T & readValid;
  wire [4:0]        reorderQueueAllocate_allocate_15 = readIssueStageEnq ? accessCountEnq_15 : 5'h0;
  wire [5:0]        reorderQueueAllocate_counterUpdate_15 = reorderQueueAllocate_counter_15 + {1'h0, reorderQueueAllocate_allocate_15} - {5'h0, reorderQueueAllocate_release_15};
  assign reorderQueueAllocate =
    ~(reorderQueueAllocate_counterWillUpdate[5]) & ~(reorderQueueAllocate_counterWillUpdate_1[5]) & ~(reorderQueueAllocate_counterWillUpdate_2[5]) & ~(reorderQueueAllocate_counterWillUpdate_3[5])
    & ~(reorderQueueAllocate_counterWillUpdate_4[5]) & ~(reorderQueueAllocate_counterWillUpdate_5[5]) & ~(reorderQueueAllocate_counterWillUpdate_6[5]) & ~(reorderQueueAllocate_counterWillUpdate_7[5])
    & ~(reorderQueueAllocate_counterWillUpdate_8[5]) & ~(reorderQueueAllocate_counterWillUpdate_9[5]) & ~(reorderQueueAllocate_counterWillUpdate_10[5]) & ~(reorderQueueAllocate_counterWillUpdate_11[5])
    & ~(reorderQueueAllocate_counterWillUpdate_12[5]) & ~(reorderQueueAllocate_counterWillUpdate_13[5]) & ~(reorderQueueAllocate_counterWillUpdate_14[5]) & ~(reorderQueueAllocate_counterWillUpdate_15[5]);
  reg               reorderStageValid;
  reg  [4:0]        reorderStageState_0;
  reg  [4:0]        reorderStageState_1;
  reg  [4:0]        reorderStageState_2;
  reg  [4:0]        reorderStageState_3;
  reg  [4:0]        reorderStageState_4;
  reg  [4:0]        reorderStageState_5;
  reg  [4:0]        reorderStageState_6;
  reg  [4:0]        reorderStageState_7;
  reg  [4:0]        reorderStageState_8;
  reg  [4:0]        reorderStageState_9;
  reg  [4:0]        reorderStageState_10;
  reg  [4:0]        reorderStageState_11;
  reg  [4:0]        reorderStageState_12;
  reg  [4:0]        reorderStageState_13;
  reg  [4:0]        reorderStageState_14;
  reg  [4:0]        reorderStageState_15;
  reg  [4:0]        reorderStageNeed_0;
  reg  [4:0]        reorderStageNeed_1;
  reg  [4:0]        reorderStageNeed_2;
  reg  [4:0]        reorderStageNeed_3;
  reg  [4:0]        reorderStageNeed_4;
  reg  [4:0]        reorderStageNeed_5;
  reg  [4:0]        reorderStageNeed_6;
  reg  [4:0]        reorderStageNeed_7;
  reg  [4:0]        reorderStageNeed_8;
  reg  [4:0]        reorderStageNeed_9;
  reg  [4:0]        reorderStageNeed_10;
  reg  [4:0]        reorderStageNeed_11;
  reg  [4:0]        reorderStageNeed_12;
  reg  [4:0]        reorderStageNeed_13;
  reg  [4:0]        reorderStageNeed_14;
  reg  [4:0]        reorderStageNeed_15;
  wire              stateCheck =
    reorderStageState_0 == reorderStageNeed_0 & reorderStageState_1 == reorderStageNeed_1 & reorderStageState_2 == reorderStageNeed_2 & reorderStageState_3 == reorderStageNeed_3 & reorderStageState_4 == reorderStageNeed_4
    & reorderStageState_5 == reorderStageNeed_5 & reorderStageState_6 == reorderStageNeed_6 & reorderStageState_7 == reorderStageNeed_7 & reorderStageState_8 == reorderStageNeed_8 & reorderStageState_9 == reorderStageNeed_9
    & reorderStageState_10 == reorderStageNeed_10 & reorderStageState_11 == reorderStageNeed_11 & reorderStageState_12 == reorderStageNeed_12 & reorderStageState_13 == reorderStageNeed_13 & reorderStageState_14 == reorderStageNeed_14
    & reorderStageState_15 == reorderStageNeed_15;
  assign accessCountQueue_deq_ready = ~reorderStageValid | stateCheck;
  wire              reorderStageEnqFire = accessCountQueue_deq_ready & accessCountQueue_deq_valid;
  wire              reorderStageDeqFire = stateCheck & reorderStageValid;
  wire [15:0]       sourceLane;
  wire              readMessageQueue_deq_valid;
  assign readMessageQueue_deq_valid = ~_readMessageQueue_fifo_empty;
  wire [15:0]       readMessageQueue_dataOut_readSource;
  assign reorderQueueVec_0_enq_bits_write1H = readMessageQueue_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_dataOffset;
  wire [15:0]       readMessageQueue_enq_bits_readSource;
  wire [1:0]        readMessageQueue_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn = {readMessageQueue_enq_bits_readSource, readMessageQueue_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_dataOffset = _readMessageQueue_fifo_data_out[1:0];
  assign readMessageQueue_dataOut_readSource = _readMessageQueue_fifo_data_out[17:2];
  assign readMessageQueue_deq_bits_readSource = readMessageQueue_dataOut_readSource;
  wire [1:0]        readMessageQueue_deq_bits_dataOffset = readMessageQueue_dataOut_dataOffset;
  wire              readMessageQueue_enq_ready = ~_readMessageQueue_fifo_full;
  wire              readMessageQueue_enq_valid;
  assign deqAllocate = ~readValid | reorderStageValid & reorderStageState_0 != reorderStageNeed_0;
  assign reorderQueueVec_0_deq_ready = deqAllocate;
  assign sourceLane = 16'h1 << _readCrossBar_output_0_bits_writeIndex;
  assign readMessageQueue_enq_bits_readSource = sourceLane;
  wire              readChannel_0_valid_0 = maskDestinationType ? _maskedWrite_readChannel_0_valid : _readCrossBar_output_0_valid & readMessageQueue_enq_ready;
  wire [4:0]        readChannel_0_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_vs : _readCrossBar_output_0_bits_vs;
  wire              readChannel_0_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_offset : _readCrossBar_output_0_bits_offset;
  assign readMessageQueue_enq_valid = readChannel_0_ready_0 & readChannel_0_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_0_enq_bits_data = readResult_0_bits >> {27'h0, readMessageQueue_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_0 = _write1HPipe_0_T & ~maskDestinationType ? reorderQueueVec_0_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_1;
  wire              readMessageQueue_1_deq_valid;
  assign readMessageQueue_1_deq_valid = ~_readMessageQueue_fifo_1_empty;
  wire [15:0]       readMessageQueue_dataOut_1_readSource;
  assign reorderQueueVec_1_enq_bits_write1H = readMessageQueue_1_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_1_dataOffset;
  wire [15:0]       readMessageQueue_1_enq_bits_readSource;
  wire [1:0]        readMessageQueue_1_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_1 = {readMessageQueue_1_enq_bits_readSource, readMessageQueue_1_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_1_dataOffset = _readMessageQueue_fifo_1_data_out[1:0];
  assign readMessageQueue_dataOut_1_readSource = _readMessageQueue_fifo_1_data_out[17:2];
  assign readMessageQueue_1_deq_bits_readSource = readMessageQueue_dataOut_1_readSource;
  wire [1:0]        readMessageQueue_1_deq_bits_dataOffset = readMessageQueue_dataOut_1_dataOffset;
  wire              readMessageQueue_1_enq_ready = ~_readMessageQueue_fifo_1_full;
  wire              readMessageQueue_1_enq_valid;
  assign deqAllocate_1 = ~readValid | reorderStageValid & reorderStageState_1 != reorderStageNeed_1;
  assign reorderQueueVec_1_deq_ready = deqAllocate_1;
  assign sourceLane_1 = 16'h1 << _readCrossBar_output_1_bits_writeIndex;
  assign readMessageQueue_1_enq_bits_readSource = sourceLane_1;
  wire              readChannel_1_valid_0 = maskDestinationType ? _maskedWrite_readChannel_1_valid : _readCrossBar_output_1_valid & readMessageQueue_1_enq_ready;
  wire [4:0]        readChannel_1_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_vs : _readCrossBar_output_1_bits_vs;
  wire              readChannel_1_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_offset : _readCrossBar_output_1_bits_offset;
  assign readMessageQueue_1_enq_valid = readChannel_1_ready_0 & readChannel_1_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_1_enq_bits_data = readResult_1_bits >> {27'h0, readMessageQueue_1_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_1 = _write1HPipe_1_T & ~maskDestinationType ? reorderQueueVec_1_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_2;
  wire              readMessageQueue_2_deq_valid;
  assign readMessageQueue_2_deq_valid = ~_readMessageQueue_fifo_2_empty;
  wire [15:0]       readMessageQueue_dataOut_2_readSource;
  assign reorderQueueVec_2_enq_bits_write1H = readMessageQueue_2_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_2_dataOffset;
  wire [15:0]       readMessageQueue_2_enq_bits_readSource;
  wire [1:0]        readMessageQueue_2_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_2 = {readMessageQueue_2_enq_bits_readSource, readMessageQueue_2_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_2_dataOffset = _readMessageQueue_fifo_2_data_out[1:0];
  assign readMessageQueue_dataOut_2_readSource = _readMessageQueue_fifo_2_data_out[17:2];
  assign readMessageQueue_2_deq_bits_readSource = readMessageQueue_dataOut_2_readSource;
  wire [1:0]        readMessageQueue_2_deq_bits_dataOffset = readMessageQueue_dataOut_2_dataOffset;
  wire              readMessageQueue_2_enq_ready = ~_readMessageQueue_fifo_2_full;
  wire              readMessageQueue_2_enq_valid;
  assign deqAllocate_2 = ~readValid | reorderStageValid & reorderStageState_2 != reorderStageNeed_2;
  assign reorderQueueVec_2_deq_ready = deqAllocate_2;
  assign sourceLane_2 = 16'h1 << _readCrossBar_output_2_bits_writeIndex;
  assign readMessageQueue_2_enq_bits_readSource = sourceLane_2;
  wire              readChannel_2_valid_0 = maskDestinationType ? _maskedWrite_readChannel_2_valid : _readCrossBar_output_2_valid & readMessageQueue_2_enq_ready;
  wire [4:0]        readChannel_2_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_vs : _readCrossBar_output_2_bits_vs;
  wire              readChannel_2_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_offset : _readCrossBar_output_2_bits_offset;
  assign readMessageQueue_2_enq_valid = readChannel_2_ready_0 & readChannel_2_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_2_enq_bits_data = readResult_2_bits >> {27'h0, readMessageQueue_2_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_2 = _write1HPipe_2_T & ~maskDestinationType ? reorderQueueVec_2_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_3;
  wire              readMessageQueue_3_deq_valid;
  assign readMessageQueue_3_deq_valid = ~_readMessageQueue_fifo_3_empty;
  wire [15:0]       readMessageQueue_dataOut_3_readSource;
  assign reorderQueueVec_3_enq_bits_write1H = readMessageQueue_3_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_3_dataOffset;
  wire [15:0]       readMessageQueue_3_enq_bits_readSource;
  wire [1:0]        readMessageQueue_3_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_3 = {readMessageQueue_3_enq_bits_readSource, readMessageQueue_3_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_3_dataOffset = _readMessageQueue_fifo_3_data_out[1:0];
  assign readMessageQueue_dataOut_3_readSource = _readMessageQueue_fifo_3_data_out[17:2];
  assign readMessageQueue_3_deq_bits_readSource = readMessageQueue_dataOut_3_readSource;
  wire [1:0]        readMessageQueue_3_deq_bits_dataOffset = readMessageQueue_dataOut_3_dataOffset;
  wire              readMessageQueue_3_enq_ready = ~_readMessageQueue_fifo_3_full;
  wire              readMessageQueue_3_enq_valid;
  assign deqAllocate_3 = ~readValid | reorderStageValid & reorderStageState_3 != reorderStageNeed_3;
  assign reorderQueueVec_3_deq_ready = deqAllocate_3;
  assign sourceLane_3 = 16'h1 << _readCrossBar_output_3_bits_writeIndex;
  assign readMessageQueue_3_enq_bits_readSource = sourceLane_3;
  wire              readChannel_3_valid_0 = maskDestinationType ? _maskedWrite_readChannel_3_valid : _readCrossBar_output_3_valid & readMessageQueue_3_enq_ready;
  wire [4:0]        readChannel_3_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_vs : _readCrossBar_output_3_bits_vs;
  wire              readChannel_3_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_offset : _readCrossBar_output_3_bits_offset;
  assign readMessageQueue_3_enq_valid = readChannel_3_ready_0 & readChannel_3_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_3_enq_bits_data = readResult_3_bits >> {27'h0, readMessageQueue_3_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_3 = _write1HPipe_3_T & ~maskDestinationType ? reorderQueueVec_3_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_4;
  wire              readMessageQueue_4_deq_valid;
  assign readMessageQueue_4_deq_valid = ~_readMessageQueue_fifo_4_empty;
  wire [15:0]       readMessageQueue_dataOut_4_readSource;
  assign reorderQueueVec_4_enq_bits_write1H = readMessageQueue_4_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_4_dataOffset;
  wire [15:0]       readMessageQueue_4_enq_bits_readSource;
  wire [1:0]        readMessageQueue_4_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_4 = {readMessageQueue_4_enq_bits_readSource, readMessageQueue_4_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_4_dataOffset = _readMessageQueue_fifo_4_data_out[1:0];
  assign readMessageQueue_dataOut_4_readSource = _readMessageQueue_fifo_4_data_out[17:2];
  assign readMessageQueue_4_deq_bits_readSource = readMessageQueue_dataOut_4_readSource;
  wire [1:0]        readMessageQueue_4_deq_bits_dataOffset = readMessageQueue_dataOut_4_dataOffset;
  wire              readMessageQueue_4_enq_ready = ~_readMessageQueue_fifo_4_full;
  wire              readMessageQueue_4_enq_valid;
  assign deqAllocate_4 = ~readValid | reorderStageValid & reorderStageState_4 != reorderStageNeed_4;
  assign reorderQueueVec_4_deq_ready = deqAllocate_4;
  assign sourceLane_4 = 16'h1 << _readCrossBar_output_4_bits_writeIndex;
  assign readMessageQueue_4_enq_bits_readSource = sourceLane_4;
  wire              readChannel_4_valid_0 = maskDestinationType ? _maskedWrite_readChannel_4_valid : _readCrossBar_output_4_valid & readMessageQueue_4_enq_ready;
  wire [4:0]        readChannel_4_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_4_bits_vs : _readCrossBar_output_4_bits_vs;
  wire              readChannel_4_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_4_bits_offset : _readCrossBar_output_4_bits_offset;
  assign readMessageQueue_4_enq_valid = readChannel_4_ready_0 & readChannel_4_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_4_enq_bits_data = readResult_4_bits >> {27'h0, readMessageQueue_4_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_4 = _write1HPipe_4_T & ~maskDestinationType ? reorderQueueVec_4_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_5;
  wire              readMessageQueue_5_deq_valid;
  assign readMessageQueue_5_deq_valid = ~_readMessageQueue_fifo_5_empty;
  wire [15:0]       readMessageQueue_dataOut_5_readSource;
  assign reorderQueueVec_5_enq_bits_write1H = readMessageQueue_5_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_5_dataOffset;
  wire [15:0]       readMessageQueue_5_enq_bits_readSource;
  wire [1:0]        readMessageQueue_5_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_5 = {readMessageQueue_5_enq_bits_readSource, readMessageQueue_5_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_5_dataOffset = _readMessageQueue_fifo_5_data_out[1:0];
  assign readMessageQueue_dataOut_5_readSource = _readMessageQueue_fifo_5_data_out[17:2];
  assign readMessageQueue_5_deq_bits_readSource = readMessageQueue_dataOut_5_readSource;
  wire [1:0]        readMessageQueue_5_deq_bits_dataOffset = readMessageQueue_dataOut_5_dataOffset;
  wire              readMessageQueue_5_enq_ready = ~_readMessageQueue_fifo_5_full;
  wire              readMessageQueue_5_enq_valid;
  assign deqAllocate_5 = ~readValid | reorderStageValid & reorderStageState_5 != reorderStageNeed_5;
  assign reorderQueueVec_5_deq_ready = deqAllocate_5;
  assign sourceLane_5 = 16'h1 << _readCrossBar_output_5_bits_writeIndex;
  assign readMessageQueue_5_enq_bits_readSource = sourceLane_5;
  wire              readChannel_5_valid_0 = maskDestinationType ? _maskedWrite_readChannel_5_valid : _readCrossBar_output_5_valid & readMessageQueue_5_enq_ready;
  wire [4:0]        readChannel_5_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_5_bits_vs : _readCrossBar_output_5_bits_vs;
  wire              readChannel_5_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_5_bits_offset : _readCrossBar_output_5_bits_offset;
  assign readMessageQueue_5_enq_valid = readChannel_5_ready_0 & readChannel_5_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_5_enq_bits_data = readResult_5_bits >> {27'h0, readMessageQueue_5_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_5 = _write1HPipe_5_T & ~maskDestinationType ? reorderQueueVec_5_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_6;
  wire              readMessageQueue_6_deq_valid;
  assign readMessageQueue_6_deq_valid = ~_readMessageQueue_fifo_6_empty;
  wire [15:0]       readMessageQueue_dataOut_6_readSource;
  assign reorderQueueVec_6_enq_bits_write1H = readMessageQueue_6_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_6_dataOffset;
  wire [15:0]       readMessageQueue_6_enq_bits_readSource;
  wire [1:0]        readMessageQueue_6_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_6 = {readMessageQueue_6_enq_bits_readSource, readMessageQueue_6_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_6_dataOffset = _readMessageQueue_fifo_6_data_out[1:0];
  assign readMessageQueue_dataOut_6_readSource = _readMessageQueue_fifo_6_data_out[17:2];
  assign readMessageQueue_6_deq_bits_readSource = readMessageQueue_dataOut_6_readSource;
  wire [1:0]        readMessageQueue_6_deq_bits_dataOffset = readMessageQueue_dataOut_6_dataOffset;
  wire              readMessageQueue_6_enq_ready = ~_readMessageQueue_fifo_6_full;
  wire              readMessageQueue_6_enq_valid;
  assign deqAllocate_6 = ~readValid | reorderStageValid & reorderStageState_6 != reorderStageNeed_6;
  assign reorderQueueVec_6_deq_ready = deqAllocate_6;
  assign sourceLane_6 = 16'h1 << _readCrossBar_output_6_bits_writeIndex;
  assign readMessageQueue_6_enq_bits_readSource = sourceLane_6;
  wire              readChannel_6_valid_0 = maskDestinationType ? _maskedWrite_readChannel_6_valid : _readCrossBar_output_6_valid & readMessageQueue_6_enq_ready;
  wire [4:0]        readChannel_6_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_6_bits_vs : _readCrossBar_output_6_bits_vs;
  wire              readChannel_6_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_6_bits_offset : _readCrossBar_output_6_bits_offset;
  assign readMessageQueue_6_enq_valid = readChannel_6_ready_0 & readChannel_6_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_6_enq_bits_data = readResult_6_bits >> {27'h0, readMessageQueue_6_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_6 = _write1HPipe_6_T & ~maskDestinationType ? reorderQueueVec_6_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_7;
  wire              readMessageQueue_7_deq_valid;
  assign readMessageQueue_7_deq_valid = ~_readMessageQueue_fifo_7_empty;
  wire [15:0]       readMessageQueue_dataOut_7_readSource;
  assign reorderQueueVec_7_enq_bits_write1H = readMessageQueue_7_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_7_dataOffset;
  wire [15:0]       readMessageQueue_7_enq_bits_readSource;
  wire [1:0]        readMessageQueue_7_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_7 = {readMessageQueue_7_enq_bits_readSource, readMessageQueue_7_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_7_dataOffset = _readMessageQueue_fifo_7_data_out[1:0];
  assign readMessageQueue_dataOut_7_readSource = _readMessageQueue_fifo_7_data_out[17:2];
  assign readMessageQueue_7_deq_bits_readSource = readMessageQueue_dataOut_7_readSource;
  wire [1:0]        readMessageQueue_7_deq_bits_dataOffset = readMessageQueue_dataOut_7_dataOffset;
  wire              readMessageQueue_7_enq_ready = ~_readMessageQueue_fifo_7_full;
  wire              readMessageQueue_7_enq_valid;
  assign deqAllocate_7 = ~readValid | reorderStageValid & reorderStageState_7 != reorderStageNeed_7;
  assign reorderQueueVec_7_deq_ready = deqAllocate_7;
  assign sourceLane_7 = 16'h1 << _readCrossBar_output_7_bits_writeIndex;
  assign readMessageQueue_7_enq_bits_readSource = sourceLane_7;
  wire              readChannel_7_valid_0 = maskDestinationType ? _maskedWrite_readChannel_7_valid : _readCrossBar_output_7_valid & readMessageQueue_7_enq_ready;
  wire [4:0]        readChannel_7_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_7_bits_vs : _readCrossBar_output_7_bits_vs;
  wire              readChannel_7_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_7_bits_offset : _readCrossBar_output_7_bits_offset;
  assign readMessageQueue_7_enq_valid = readChannel_7_ready_0 & readChannel_7_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_7_enq_bits_data = readResult_7_bits >> {27'h0, readMessageQueue_7_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_7 = _write1HPipe_7_T & ~maskDestinationType ? reorderQueueVec_7_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_8;
  wire              readMessageQueue_8_deq_valid;
  assign readMessageQueue_8_deq_valid = ~_readMessageQueue_fifo_8_empty;
  wire [15:0]       readMessageQueue_dataOut_8_readSource;
  assign reorderQueueVec_8_enq_bits_write1H = readMessageQueue_8_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_8_dataOffset;
  wire [15:0]       readMessageQueue_8_enq_bits_readSource;
  wire [1:0]        readMessageQueue_8_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_8 = {readMessageQueue_8_enq_bits_readSource, readMessageQueue_8_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_8_dataOffset = _readMessageQueue_fifo_8_data_out[1:0];
  assign readMessageQueue_dataOut_8_readSource = _readMessageQueue_fifo_8_data_out[17:2];
  assign readMessageQueue_8_deq_bits_readSource = readMessageQueue_dataOut_8_readSource;
  wire [1:0]        readMessageQueue_8_deq_bits_dataOffset = readMessageQueue_dataOut_8_dataOffset;
  wire              readMessageQueue_8_enq_ready = ~_readMessageQueue_fifo_8_full;
  wire              readMessageQueue_8_enq_valid;
  assign deqAllocate_8 = ~readValid | reorderStageValid & reorderStageState_8 != reorderStageNeed_8;
  assign reorderQueueVec_8_deq_ready = deqAllocate_8;
  assign sourceLane_8 = 16'h1 << _readCrossBar_output_8_bits_writeIndex;
  assign readMessageQueue_8_enq_bits_readSource = sourceLane_8;
  wire              readChannel_8_valid_0 = maskDestinationType ? _maskedWrite_readChannel_8_valid : _readCrossBar_output_8_valid & readMessageQueue_8_enq_ready;
  wire [4:0]        readChannel_8_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_8_bits_vs : _readCrossBar_output_8_bits_vs;
  wire              readChannel_8_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_8_bits_offset : _readCrossBar_output_8_bits_offset;
  assign readMessageQueue_8_enq_valid = readChannel_8_ready_0 & readChannel_8_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_8_enq_bits_data = readResult_8_bits >> {27'h0, readMessageQueue_8_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_8 = _write1HPipe_8_T & ~maskDestinationType ? reorderQueueVec_8_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_9;
  wire              readMessageQueue_9_deq_valid;
  assign readMessageQueue_9_deq_valid = ~_readMessageQueue_fifo_9_empty;
  wire [15:0]       readMessageQueue_dataOut_9_readSource;
  assign reorderQueueVec_9_enq_bits_write1H = readMessageQueue_9_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_9_dataOffset;
  wire [15:0]       readMessageQueue_9_enq_bits_readSource;
  wire [1:0]        readMessageQueue_9_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_9 = {readMessageQueue_9_enq_bits_readSource, readMessageQueue_9_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_9_dataOffset = _readMessageQueue_fifo_9_data_out[1:0];
  assign readMessageQueue_dataOut_9_readSource = _readMessageQueue_fifo_9_data_out[17:2];
  assign readMessageQueue_9_deq_bits_readSource = readMessageQueue_dataOut_9_readSource;
  wire [1:0]        readMessageQueue_9_deq_bits_dataOffset = readMessageQueue_dataOut_9_dataOffset;
  wire              readMessageQueue_9_enq_ready = ~_readMessageQueue_fifo_9_full;
  wire              readMessageQueue_9_enq_valid;
  assign deqAllocate_9 = ~readValid | reorderStageValid & reorderStageState_9 != reorderStageNeed_9;
  assign reorderQueueVec_9_deq_ready = deqAllocate_9;
  assign sourceLane_9 = 16'h1 << _readCrossBar_output_9_bits_writeIndex;
  assign readMessageQueue_9_enq_bits_readSource = sourceLane_9;
  wire              readChannel_9_valid_0 = maskDestinationType ? _maskedWrite_readChannel_9_valid : _readCrossBar_output_9_valid & readMessageQueue_9_enq_ready;
  wire [4:0]        readChannel_9_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_9_bits_vs : _readCrossBar_output_9_bits_vs;
  wire              readChannel_9_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_9_bits_offset : _readCrossBar_output_9_bits_offset;
  assign readMessageQueue_9_enq_valid = readChannel_9_ready_0 & readChannel_9_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_9_enq_bits_data = readResult_9_bits >> {27'h0, readMessageQueue_9_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_9 = _write1HPipe_9_T & ~maskDestinationType ? reorderQueueVec_9_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_10;
  wire              readMessageQueue_10_deq_valid;
  assign readMessageQueue_10_deq_valid = ~_readMessageQueue_fifo_10_empty;
  wire [15:0]       readMessageQueue_dataOut_10_readSource;
  assign reorderQueueVec_10_enq_bits_write1H = readMessageQueue_10_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_10_dataOffset;
  wire [15:0]       readMessageQueue_10_enq_bits_readSource;
  wire [1:0]        readMessageQueue_10_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_10 = {readMessageQueue_10_enq_bits_readSource, readMessageQueue_10_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_10_dataOffset = _readMessageQueue_fifo_10_data_out[1:0];
  assign readMessageQueue_dataOut_10_readSource = _readMessageQueue_fifo_10_data_out[17:2];
  assign readMessageQueue_10_deq_bits_readSource = readMessageQueue_dataOut_10_readSource;
  wire [1:0]        readMessageQueue_10_deq_bits_dataOffset = readMessageQueue_dataOut_10_dataOffset;
  wire              readMessageQueue_10_enq_ready = ~_readMessageQueue_fifo_10_full;
  wire              readMessageQueue_10_enq_valid;
  assign deqAllocate_10 = ~readValid | reorderStageValid & reorderStageState_10 != reorderStageNeed_10;
  assign reorderQueueVec_10_deq_ready = deqAllocate_10;
  assign sourceLane_10 = 16'h1 << _readCrossBar_output_10_bits_writeIndex;
  assign readMessageQueue_10_enq_bits_readSource = sourceLane_10;
  wire              readChannel_10_valid_0 = maskDestinationType ? _maskedWrite_readChannel_10_valid : _readCrossBar_output_10_valid & readMessageQueue_10_enq_ready;
  wire [4:0]        readChannel_10_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_10_bits_vs : _readCrossBar_output_10_bits_vs;
  wire              readChannel_10_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_10_bits_offset : _readCrossBar_output_10_bits_offset;
  assign readMessageQueue_10_enq_valid = readChannel_10_ready_0 & readChannel_10_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_10_enq_bits_data = readResult_10_bits >> {27'h0, readMessageQueue_10_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_10 = _write1HPipe_10_T & ~maskDestinationType ? reorderQueueVec_10_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_11;
  wire              readMessageQueue_11_deq_valid;
  assign readMessageQueue_11_deq_valid = ~_readMessageQueue_fifo_11_empty;
  wire [15:0]       readMessageQueue_dataOut_11_readSource;
  assign reorderQueueVec_11_enq_bits_write1H = readMessageQueue_11_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_11_dataOffset;
  wire [15:0]       readMessageQueue_11_enq_bits_readSource;
  wire [1:0]        readMessageQueue_11_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_11 = {readMessageQueue_11_enq_bits_readSource, readMessageQueue_11_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_11_dataOffset = _readMessageQueue_fifo_11_data_out[1:0];
  assign readMessageQueue_dataOut_11_readSource = _readMessageQueue_fifo_11_data_out[17:2];
  assign readMessageQueue_11_deq_bits_readSource = readMessageQueue_dataOut_11_readSource;
  wire [1:0]        readMessageQueue_11_deq_bits_dataOffset = readMessageQueue_dataOut_11_dataOffset;
  wire              readMessageQueue_11_enq_ready = ~_readMessageQueue_fifo_11_full;
  wire              readMessageQueue_11_enq_valid;
  assign deqAllocate_11 = ~readValid | reorderStageValid & reorderStageState_11 != reorderStageNeed_11;
  assign reorderQueueVec_11_deq_ready = deqAllocate_11;
  assign sourceLane_11 = 16'h1 << _readCrossBar_output_11_bits_writeIndex;
  assign readMessageQueue_11_enq_bits_readSource = sourceLane_11;
  wire              readChannel_11_valid_0 = maskDestinationType ? _maskedWrite_readChannel_11_valid : _readCrossBar_output_11_valid & readMessageQueue_11_enq_ready;
  wire [4:0]        readChannel_11_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_11_bits_vs : _readCrossBar_output_11_bits_vs;
  wire              readChannel_11_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_11_bits_offset : _readCrossBar_output_11_bits_offset;
  assign readMessageQueue_11_enq_valid = readChannel_11_ready_0 & readChannel_11_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_11_enq_bits_data = readResult_11_bits >> {27'h0, readMessageQueue_11_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_11 = _write1HPipe_11_T & ~maskDestinationType ? reorderQueueVec_11_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_12;
  wire              readMessageQueue_12_deq_valid;
  assign readMessageQueue_12_deq_valid = ~_readMessageQueue_fifo_12_empty;
  wire [15:0]       readMessageQueue_dataOut_12_readSource;
  assign reorderQueueVec_12_enq_bits_write1H = readMessageQueue_12_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_12_dataOffset;
  wire [15:0]       readMessageQueue_12_enq_bits_readSource;
  wire [1:0]        readMessageQueue_12_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_12 = {readMessageQueue_12_enq_bits_readSource, readMessageQueue_12_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_12_dataOffset = _readMessageQueue_fifo_12_data_out[1:0];
  assign readMessageQueue_dataOut_12_readSource = _readMessageQueue_fifo_12_data_out[17:2];
  assign readMessageQueue_12_deq_bits_readSource = readMessageQueue_dataOut_12_readSource;
  wire [1:0]        readMessageQueue_12_deq_bits_dataOffset = readMessageQueue_dataOut_12_dataOffset;
  wire              readMessageQueue_12_enq_ready = ~_readMessageQueue_fifo_12_full;
  wire              readMessageQueue_12_enq_valid;
  assign deqAllocate_12 = ~readValid | reorderStageValid & reorderStageState_12 != reorderStageNeed_12;
  assign reorderQueueVec_12_deq_ready = deqAllocate_12;
  assign sourceLane_12 = 16'h1 << _readCrossBar_output_12_bits_writeIndex;
  assign readMessageQueue_12_enq_bits_readSource = sourceLane_12;
  wire              readChannel_12_valid_0 = maskDestinationType ? _maskedWrite_readChannel_12_valid : _readCrossBar_output_12_valid & readMessageQueue_12_enq_ready;
  wire [4:0]        readChannel_12_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_12_bits_vs : _readCrossBar_output_12_bits_vs;
  wire              readChannel_12_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_12_bits_offset : _readCrossBar_output_12_bits_offset;
  assign readMessageQueue_12_enq_valid = readChannel_12_ready_0 & readChannel_12_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_12_enq_bits_data = readResult_12_bits >> {27'h0, readMessageQueue_12_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_12 = _write1HPipe_12_T & ~maskDestinationType ? reorderQueueVec_12_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_13;
  wire              readMessageQueue_13_deq_valid;
  assign readMessageQueue_13_deq_valid = ~_readMessageQueue_fifo_13_empty;
  wire [15:0]       readMessageQueue_dataOut_13_readSource;
  assign reorderQueueVec_13_enq_bits_write1H = readMessageQueue_13_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_13_dataOffset;
  wire [15:0]       readMessageQueue_13_enq_bits_readSource;
  wire [1:0]        readMessageQueue_13_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_13 = {readMessageQueue_13_enq_bits_readSource, readMessageQueue_13_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_13_dataOffset = _readMessageQueue_fifo_13_data_out[1:0];
  assign readMessageQueue_dataOut_13_readSource = _readMessageQueue_fifo_13_data_out[17:2];
  assign readMessageQueue_13_deq_bits_readSource = readMessageQueue_dataOut_13_readSource;
  wire [1:0]        readMessageQueue_13_deq_bits_dataOffset = readMessageQueue_dataOut_13_dataOffset;
  wire              readMessageQueue_13_enq_ready = ~_readMessageQueue_fifo_13_full;
  wire              readMessageQueue_13_enq_valid;
  assign deqAllocate_13 = ~readValid | reorderStageValid & reorderStageState_13 != reorderStageNeed_13;
  assign reorderQueueVec_13_deq_ready = deqAllocate_13;
  assign sourceLane_13 = 16'h1 << _readCrossBar_output_13_bits_writeIndex;
  assign readMessageQueue_13_enq_bits_readSource = sourceLane_13;
  wire              readChannel_13_valid_0 = maskDestinationType ? _maskedWrite_readChannel_13_valid : _readCrossBar_output_13_valid & readMessageQueue_13_enq_ready;
  wire [4:0]        readChannel_13_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_13_bits_vs : _readCrossBar_output_13_bits_vs;
  wire              readChannel_13_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_13_bits_offset : _readCrossBar_output_13_bits_offset;
  assign readMessageQueue_13_enq_valid = readChannel_13_ready_0 & readChannel_13_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_13_enq_bits_data = readResult_13_bits >> {27'h0, readMessageQueue_13_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_13 = _write1HPipe_13_T & ~maskDestinationType ? reorderQueueVec_13_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_14;
  wire              readMessageQueue_14_deq_valid;
  assign readMessageQueue_14_deq_valid = ~_readMessageQueue_fifo_14_empty;
  wire [15:0]       readMessageQueue_dataOut_14_readSource;
  assign reorderQueueVec_14_enq_bits_write1H = readMessageQueue_14_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_14_dataOffset;
  wire [15:0]       readMessageQueue_14_enq_bits_readSource;
  wire [1:0]        readMessageQueue_14_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_14 = {readMessageQueue_14_enq_bits_readSource, readMessageQueue_14_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_14_dataOffset = _readMessageQueue_fifo_14_data_out[1:0];
  assign readMessageQueue_dataOut_14_readSource = _readMessageQueue_fifo_14_data_out[17:2];
  assign readMessageQueue_14_deq_bits_readSource = readMessageQueue_dataOut_14_readSource;
  wire [1:0]        readMessageQueue_14_deq_bits_dataOffset = readMessageQueue_dataOut_14_dataOffset;
  wire              readMessageQueue_14_enq_ready = ~_readMessageQueue_fifo_14_full;
  wire              readMessageQueue_14_enq_valid;
  assign deqAllocate_14 = ~readValid | reorderStageValid & reorderStageState_14 != reorderStageNeed_14;
  assign reorderQueueVec_14_deq_ready = deqAllocate_14;
  assign sourceLane_14 = 16'h1 << _readCrossBar_output_14_bits_writeIndex;
  assign readMessageQueue_14_enq_bits_readSource = sourceLane_14;
  wire              readChannel_14_valid_0 = maskDestinationType ? _maskedWrite_readChannel_14_valid : _readCrossBar_output_14_valid & readMessageQueue_14_enq_ready;
  wire [4:0]        readChannel_14_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_14_bits_vs : _readCrossBar_output_14_bits_vs;
  wire              readChannel_14_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_14_bits_offset : _readCrossBar_output_14_bits_offset;
  assign readMessageQueue_14_enq_valid = readChannel_14_ready_0 & readChannel_14_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_14_enq_bits_data = readResult_14_bits >> {27'h0, readMessageQueue_14_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_14 = _write1HPipe_14_T & ~maskDestinationType ? reorderQueueVec_14_deq_bits_write1H : 16'h0;
  wire [15:0]       sourceLane_15;
  wire              readMessageQueue_15_deq_valid;
  assign readMessageQueue_15_deq_valid = ~_readMessageQueue_fifo_15_empty;
  wire [15:0]       readMessageQueue_dataOut_15_readSource;
  assign reorderQueueVec_15_enq_bits_write1H = readMessageQueue_15_deq_bits_readSource;
  wire [1:0]        readMessageQueue_dataOut_15_dataOffset;
  wire [15:0]       readMessageQueue_15_enq_bits_readSource;
  wire [1:0]        readMessageQueue_15_enq_bits_dataOffset;
  wire [17:0]       readMessageQueue_dataIn_15 = {readMessageQueue_15_enq_bits_readSource, readMessageQueue_15_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_15_dataOffset = _readMessageQueue_fifo_15_data_out[1:0];
  assign readMessageQueue_dataOut_15_readSource = _readMessageQueue_fifo_15_data_out[17:2];
  assign readMessageQueue_15_deq_bits_readSource = readMessageQueue_dataOut_15_readSource;
  wire [1:0]        readMessageQueue_15_deq_bits_dataOffset = readMessageQueue_dataOut_15_dataOffset;
  wire              readMessageQueue_15_enq_ready = ~_readMessageQueue_fifo_15_full;
  wire              readMessageQueue_15_enq_valid;
  assign deqAllocate_15 = ~readValid | reorderStageValid & reorderStageState_15 != reorderStageNeed_15;
  assign reorderQueueVec_15_deq_ready = deqAllocate_15;
  assign sourceLane_15 = 16'h1 << _readCrossBar_output_15_bits_writeIndex;
  assign readMessageQueue_15_enq_bits_readSource = sourceLane_15;
  wire              readChannel_15_valid_0 = maskDestinationType ? _maskedWrite_readChannel_15_valid : _readCrossBar_output_15_valid & readMessageQueue_15_enq_ready;
  wire [4:0]        readChannel_15_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_15_bits_vs : _readCrossBar_output_15_bits_vs;
  wire              readChannel_15_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_15_bits_offset : _readCrossBar_output_15_bits_offset;
  assign readMessageQueue_15_enq_valid = readChannel_15_ready_0 & readChannel_15_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_15_enq_bits_data = readResult_15_bits >> {27'h0, readMessageQueue_15_deq_bits_dataOffset, 3'h0};
  wire [15:0]       write1HPipe_15 = _write1HPipe_15_T & ~maskDestinationType ? reorderQueueVec_15_deq_bits_write1H : 16'h0;
  wire [31:0]       readData_data;
  wire              readData_readDataQueue_enq_ready = ~_readData_readDataQueue_fifo_full;
  wire              readData_readDataQueue_deq_ready;
  wire              readData_readDataQueue_enq_valid;
  wire              readData_readDataQueue_deq_valid = ~_readData_readDataQueue_fifo_empty | readData_readDataQueue_enq_valid;
  wire [31:0]       readData_readDataQueue_enq_bits;
  wire [31:0]       readData_readDataQueue_deq_bits = _readData_readDataQueue_fifo_empty ? readData_readDataQueue_enq_bits : _readData_readDataQueue_fifo_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo = {write1HPipe_1[0], write1HPipe_0[0]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi = {write1HPipe_3[0], write1HPipe_2[0]};
  wire [3:0]        readData_readResultSelect_lo_lo = {readData_readResultSelect_lo_lo_hi, readData_readResultSelect_lo_lo_lo};
  wire [1:0]        readData_readResultSelect_lo_hi_lo = {write1HPipe_5[0], write1HPipe_4[0]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi = {write1HPipe_7[0], write1HPipe_6[0]};
  wire [3:0]        readData_readResultSelect_lo_hi = {readData_readResultSelect_lo_hi_hi, readData_readResultSelect_lo_hi_lo};
  wire [7:0]        readData_readResultSelect_lo = {readData_readResultSelect_lo_hi, readData_readResultSelect_lo_lo};
  wire [1:0]        readData_readResultSelect_hi_lo_lo = {write1HPipe_9[0], write1HPipe_8[0]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi = {write1HPipe_11[0], write1HPipe_10[0]};
  wire [3:0]        readData_readResultSelect_hi_lo = {readData_readResultSelect_hi_lo_hi, readData_readResultSelect_hi_lo_lo};
  wire [1:0]        readData_readResultSelect_hi_hi_lo = {write1HPipe_13[0], write1HPipe_12[0]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi = {write1HPipe_15[0], write1HPipe_14[0]};
  wire [3:0]        readData_readResultSelect_hi_hi = {readData_readResultSelect_hi_hi_hi, readData_readResultSelect_hi_hi_lo};
  wire [7:0]        readData_readResultSelect_hi = {readData_readResultSelect_hi_hi, readData_readResultSelect_hi_lo};
  wire [15:0]       readData_readResultSelect = {readData_readResultSelect_hi, readData_readResultSelect_lo};
  assign readData_data =
    (readData_readResultSelect[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_enq_bits = readData_data;
  wire              readTokenRelease_0 = readData_readDataQueue_deq_ready & readData_readDataQueue_deq_valid;
  assign readData_readDataQueue_enq_valid = |readData_readResultSelect;
  wire [31:0]       readData_data_1;
  wire              isWaiteForThisData_1;
  wire              readData_readDataQueue_1_enq_ready = ~_readData_readDataQueue_fifo_1_full;
  wire              readData_readDataQueue_1_deq_ready;
  wire              readData_readDataQueue_1_enq_valid;
  wire              readData_readDataQueue_1_deq_valid = ~_readData_readDataQueue_fifo_1_empty | readData_readDataQueue_1_enq_valid;
  wire [31:0]       readData_readDataQueue_1_enq_bits;
  wire [31:0]       readData_readDataQueue_1_deq_bits = _readData_readDataQueue_fifo_1_empty ? readData_readDataQueue_1_enq_bits : _readData_readDataQueue_fifo_1_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_1 = {write1HPipe_1[1], write1HPipe_0[1]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_1 = {write1HPipe_3[1], write1HPipe_2[1]};
  wire [3:0]        readData_readResultSelect_lo_lo_1 = {readData_readResultSelect_lo_lo_hi_1, readData_readResultSelect_lo_lo_lo_1};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_1 = {write1HPipe_5[1], write1HPipe_4[1]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_1 = {write1HPipe_7[1], write1HPipe_6[1]};
  wire [3:0]        readData_readResultSelect_lo_hi_1 = {readData_readResultSelect_lo_hi_hi_1, readData_readResultSelect_lo_hi_lo_1};
  wire [7:0]        readData_readResultSelect_lo_1 = {readData_readResultSelect_lo_hi_1, readData_readResultSelect_lo_lo_1};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_1 = {write1HPipe_9[1], write1HPipe_8[1]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_1 = {write1HPipe_11[1], write1HPipe_10[1]};
  wire [3:0]        readData_readResultSelect_hi_lo_1 = {readData_readResultSelect_hi_lo_hi_1, readData_readResultSelect_hi_lo_lo_1};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_1 = {write1HPipe_13[1], write1HPipe_12[1]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_1 = {write1HPipe_15[1], write1HPipe_14[1]};
  wire [3:0]        readData_readResultSelect_hi_hi_1 = {readData_readResultSelect_hi_hi_hi_1, readData_readResultSelect_hi_hi_lo_1};
  wire [7:0]        readData_readResultSelect_hi_1 = {readData_readResultSelect_hi_hi_1, readData_readResultSelect_hi_lo_1};
  wire [15:0]       readData_readResultSelect_1 = {readData_readResultSelect_hi_1, readData_readResultSelect_lo_1};
  assign readData_data_1 =
    (readData_readResultSelect_1[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_1[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_1[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_1[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_1[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_1[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_1[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_1[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_1[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_1[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_1[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_1[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_1[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_1[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_1[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_1[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_1_enq_bits = readData_data_1;
  wire              readTokenRelease_1 = readData_readDataQueue_1_deq_ready & readData_readDataQueue_1_deq_valid;
  assign readData_readDataQueue_1_enq_valid = |readData_readResultSelect_1;
  wire [31:0]       readData_data_2;
  wire              isWaiteForThisData_2;
  wire              readData_readDataQueue_2_enq_ready = ~_readData_readDataQueue_fifo_2_full;
  wire              readData_readDataQueue_2_deq_ready;
  wire              readData_readDataQueue_2_enq_valid;
  wire              readData_readDataQueue_2_deq_valid = ~_readData_readDataQueue_fifo_2_empty | readData_readDataQueue_2_enq_valid;
  wire [31:0]       readData_readDataQueue_2_enq_bits;
  wire [31:0]       readData_readDataQueue_2_deq_bits = _readData_readDataQueue_fifo_2_empty ? readData_readDataQueue_2_enq_bits : _readData_readDataQueue_fifo_2_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_2 = {write1HPipe_1[2], write1HPipe_0[2]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_2 = {write1HPipe_3[2], write1HPipe_2[2]};
  wire [3:0]        readData_readResultSelect_lo_lo_2 = {readData_readResultSelect_lo_lo_hi_2, readData_readResultSelect_lo_lo_lo_2};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_2 = {write1HPipe_5[2], write1HPipe_4[2]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_2 = {write1HPipe_7[2], write1HPipe_6[2]};
  wire [3:0]        readData_readResultSelect_lo_hi_2 = {readData_readResultSelect_lo_hi_hi_2, readData_readResultSelect_lo_hi_lo_2};
  wire [7:0]        readData_readResultSelect_lo_2 = {readData_readResultSelect_lo_hi_2, readData_readResultSelect_lo_lo_2};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_2 = {write1HPipe_9[2], write1HPipe_8[2]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_2 = {write1HPipe_11[2], write1HPipe_10[2]};
  wire [3:0]        readData_readResultSelect_hi_lo_2 = {readData_readResultSelect_hi_lo_hi_2, readData_readResultSelect_hi_lo_lo_2};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_2 = {write1HPipe_13[2], write1HPipe_12[2]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_2 = {write1HPipe_15[2], write1HPipe_14[2]};
  wire [3:0]        readData_readResultSelect_hi_hi_2 = {readData_readResultSelect_hi_hi_hi_2, readData_readResultSelect_hi_hi_lo_2};
  wire [7:0]        readData_readResultSelect_hi_2 = {readData_readResultSelect_hi_hi_2, readData_readResultSelect_hi_lo_2};
  wire [15:0]       readData_readResultSelect_2 = {readData_readResultSelect_hi_2, readData_readResultSelect_lo_2};
  assign readData_data_2 =
    (readData_readResultSelect_2[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_2[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_2[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_2[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_2[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_2[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_2[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_2[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_2[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_2[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_2[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_2[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_2[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_2[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_2[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_2[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_2_enq_bits = readData_data_2;
  wire              readTokenRelease_2 = readData_readDataQueue_2_deq_ready & readData_readDataQueue_2_deq_valid;
  assign readData_readDataQueue_2_enq_valid = |readData_readResultSelect_2;
  wire [31:0]       readData_data_3;
  wire              isWaiteForThisData_3;
  wire              readData_readDataQueue_3_enq_ready = ~_readData_readDataQueue_fifo_3_full;
  wire              readData_readDataQueue_3_deq_ready;
  wire              readData_readDataQueue_3_enq_valid;
  wire              readData_readDataQueue_3_deq_valid = ~_readData_readDataQueue_fifo_3_empty | readData_readDataQueue_3_enq_valid;
  wire [31:0]       readData_readDataQueue_3_enq_bits;
  wire [31:0]       readData_readDataQueue_3_deq_bits = _readData_readDataQueue_fifo_3_empty ? readData_readDataQueue_3_enq_bits : _readData_readDataQueue_fifo_3_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_3 = {write1HPipe_1[3], write1HPipe_0[3]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_3 = {write1HPipe_3[3], write1HPipe_2[3]};
  wire [3:0]        readData_readResultSelect_lo_lo_3 = {readData_readResultSelect_lo_lo_hi_3, readData_readResultSelect_lo_lo_lo_3};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_3 = {write1HPipe_5[3], write1HPipe_4[3]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_3 = {write1HPipe_7[3], write1HPipe_6[3]};
  wire [3:0]        readData_readResultSelect_lo_hi_3 = {readData_readResultSelect_lo_hi_hi_3, readData_readResultSelect_lo_hi_lo_3};
  wire [7:0]        readData_readResultSelect_lo_3 = {readData_readResultSelect_lo_hi_3, readData_readResultSelect_lo_lo_3};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_3 = {write1HPipe_9[3], write1HPipe_8[3]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_3 = {write1HPipe_11[3], write1HPipe_10[3]};
  wire [3:0]        readData_readResultSelect_hi_lo_3 = {readData_readResultSelect_hi_lo_hi_3, readData_readResultSelect_hi_lo_lo_3};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_3 = {write1HPipe_13[3], write1HPipe_12[3]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_3 = {write1HPipe_15[3], write1HPipe_14[3]};
  wire [3:0]        readData_readResultSelect_hi_hi_3 = {readData_readResultSelect_hi_hi_hi_3, readData_readResultSelect_hi_hi_lo_3};
  wire [7:0]        readData_readResultSelect_hi_3 = {readData_readResultSelect_hi_hi_3, readData_readResultSelect_hi_lo_3};
  wire [15:0]       readData_readResultSelect_3 = {readData_readResultSelect_hi_3, readData_readResultSelect_lo_3};
  assign readData_data_3 =
    (readData_readResultSelect_3[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_3[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_3[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_3[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_3[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_3[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_3[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_3[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_3[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_3[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_3[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_3[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_3[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_3[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_3[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_3[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_3_enq_bits = readData_data_3;
  wire              readTokenRelease_3 = readData_readDataQueue_3_deq_ready & readData_readDataQueue_3_deq_valid;
  assign readData_readDataQueue_3_enq_valid = |readData_readResultSelect_3;
  wire [31:0]       readData_data_4;
  wire              isWaiteForThisData_4;
  wire              readData_readDataQueue_4_enq_ready = ~_readData_readDataQueue_fifo_4_full;
  wire              readData_readDataQueue_4_deq_ready;
  wire              readData_readDataQueue_4_enq_valid;
  wire              readData_readDataQueue_4_deq_valid = ~_readData_readDataQueue_fifo_4_empty | readData_readDataQueue_4_enq_valid;
  wire [31:0]       readData_readDataQueue_4_enq_bits;
  wire [31:0]       readData_readDataQueue_4_deq_bits = _readData_readDataQueue_fifo_4_empty ? readData_readDataQueue_4_enq_bits : _readData_readDataQueue_fifo_4_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_4 = {write1HPipe_1[4], write1HPipe_0[4]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_4 = {write1HPipe_3[4], write1HPipe_2[4]};
  wire [3:0]        readData_readResultSelect_lo_lo_4 = {readData_readResultSelect_lo_lo_hi_4, readData_readResultSelect_lo_lo_lo_4};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_4 = {write1HPipe_5[4], write1HPipe_4[4]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_4 = {write1HPipe_7[4], write1HPipe_6[4]};
  wire [3:0]        readData_readResultSelect_lo_hi_4 = {readData_readResultSelect_lo_hi_hi_4, readData_readResultSelect_lo_hi_lo_4};
  wire [7:0]        readData_readResultSelect_lo_4 = {readData_readResultSelect_lo_hi_4, readData_readResultSelect_lo_lo_4};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_4 = {write1HPipe_9[4], write1HPipe_8[4]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_4 = {write1HPipe_11[4], write1HPipe_10[4]};
  wire [3:0]        readData_readResultSelect_hi_lo_4 = {readData_readResultSelect_hi_lo_hi_4, readData_readResultSelect_hi_lo_lo_4};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_4 = {write1HPipe_13[4], write1HPipe_12[4]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_4 = {write1HPipe_15[4], write1HPipe_14[4]};
  wire [3:0]        readData_readResultSelect_hi_hi_4 = {readData_readResultSelect_hi_hi_hi_4, readData_readResultSelect_hi_hi_lo_4};
  wire [7:0]        readData_readResultSelect_hi_4 = {readData_readResultSelect_hi_hi_4, readData_readResultSelect_hi_lo_4};
  wire [15:0]       readData_readResultSelect_4 = {readData_readResultSelect_hi_4, readData_readResultSelect_lo_4};
  assign readData_data_4 =
    (readData_readResultSelect_4[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_4[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_4[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_4[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_4[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_4[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_4[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_4[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_4[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_4[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_4[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_4[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_4[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_4[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_4[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_4[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_4_enq_bits = readData_data_4;
  wire              readTokenRelease_4 = readData_readDataQueue_4_deq_ready & readData_readDataQueue_4_deq_valid;
  assign readData_readDataQueue_4_enq_valid = |readData_readResultSelect_4;
  wire [31:0]       readData_data_5;
  wire              isWaiteForThisData_5;
  wire              readData_readDataQueue_5_enq_ready = ~_readData_readDataQueue_fifo_5_full;
  wire              readData_readDataQueue_5_deq_ready;
  wire              readData_readDataQueue_5_enq_valid;
  wire              readData_readDataQueue_5_deq_valid = ~_readData_readDataQueue_fifo_5_empty | readData_readDataQueue_5_enq_valid;
  wire [31:0]       readData_readDataQueue_5_enq_bits;
  wire [31:0]       readData_readDataQueue_5_deq_bits = _readData_readDataQueue_fifo_5_empty ? readData_readDataQueue_5_enq_bits : _readData_readDataQueue_fifo_5_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_5 = {write1HPipe_1[5], write1HPipe_0[5]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_5 = {write1HPipe_3[5], write1HPipe_2[5]};
  wire [3:0]        readData_readResultSelect_lo_lo_5 = {readData_readResultSelect_lo_lo_hi_5, readData_readResultSelect_lo_lo_lo_5};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_5 = {write1HPipe_5[5], write1HPipe_4[5]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_5 = {write1HPipe_7[5], write1HPipe_6[5]};
  wire [3:0]        readData_readResultSelect_lo_hi_5 = {readData_readResultSelect_lo_hi_hi_5, readData_readResultSelect_lo_hi_lo_5};
  wire [7:0]        readData_readResultSelect_lo_5 = {readData_readResultSelect_lo_hi_5, readData_readResultSelect_lo_lo_5};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_5 = {write1HPipe_9[5], write1HPipe_8[5]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_5 = {write1HPipe_11[5], write1HPipe_10[5]};
  wire [3:0]        readData_readResultSelect_hi_lo_5 = {readData_readResultSelect_hi_lo_hi_5, readData_readResultSelect_hi_lo_lo_5};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_5 = {write1HPipe_13[5], write1HPipe_12[5]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_5 = {write1HPipe_15[5], write1HPipe_14[5]};
  wire [3:0]        readData_readResultSelect_hi_hi_5 = {readData_readResultSelect_hi_hi_hi_5, readData_readResultSelect_hi_hi_lo_5};
  wire [7:0]        readData_readResultSelect_hi_5 = {readData_readResultSelect_hi_hi_5, readData_readResultSelect_hi_lo_5};
  wire [15:0]       readData_readResultSelect_5 = {readData_readResultSelect_hi_5, readData_readResultSelect_lo_5};
  assign readData_data_5 =
    (readData_readResultSelect_5[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_5[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_5[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_5[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_5[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_5[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_5[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_5[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_5[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_5[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_5[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_5[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_5[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_5[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_5[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_5[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_5_enq_bits = readData_data_5;
  wire              readTokenRelease_5 = readData_readDataQueue_5_deq_ready & readData_readDataQueue_5_deq_valid;
  assign readData_readDataQueue_5_enq_valid = |readData_readResultSelect_5;
  wire [31:0]       readData_data_6;
  wire              isWaiteForThisData_6;
  wire              readData_readDataQueue_6_enq_ready = ~_readData_readDataQueue_fifo_6_full;
  wire              readData_readDataQueue_6_deq_ready;
  wire              readData_readDataQueue_6_enq_valid;
  wire              readData_readDataQueue_6_deq_valid = ~_readData_readDataQueue_fifo_6_empty | readData_readDataQueue_6_enq_valid;
  wire [31:0]       readData_readDataQueue_6_enq_bits;
  wire [31:0]       readData_readDataQueue_6_deq_bits = _readData_readDataQueue_fifo_6_empty ? readData_readDataQueue_6_enq_bits : _readData_readDataQueue_fifo_6_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_6 = {write1HPipe_1[6], write1HPipe_0[6]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_6 = {write1HPipe_3[6], write1HPipe_2[6]};
  wire [3:0]        readData_readResultSelect_lo_lo_6 = {readData_readResultSelect_lo_lo_hi_6, readData_readResultSelect_lo_lo_lo_6};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_6 = {write1HPipe_5[6], write1HPipe_4[6]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_6 = {write1HPipe_7[6], write1HPipe_6[6]};
  wire [3:0]        readData_readResultSelect_lo_hi_6 = {readData_readResultSelect_lo_hi_hi_6, readData_readResultSelect_lo_hi_lo_6};
  wire [7:0]        readData_readResultSelect_lo_6 = {readData_readResultSelect_lo_hi_6, readData_readResultSelect_lo_lo_6};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_6 = {write1HPipe_9[6], write1HPipe_8[6]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_6 = {write1HPipe_11[6], write1HPipe_10[6]};
  wire [3:0]        readData_readResultSelect_hi_lo_6 = {readData_readResultSelect_hi_lo_hi_6, readData_readResultSelect_hi_lo_lo_6};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_6 = {write1HPipe_13[6], write1HPipe_12[6]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_6 = {write1HPipe_15[6], write1HPipe_14[6]};
  wire [3:0]        readData_readResultSelect_hi_hi_6 = {readData_readResultSelect_hi_hi_hi_6, readData_readResultSelect_hi_hi_lo_6};
  wire [7:0]        readData_readResultSelect_hi_6 = {readData_readResultSelect_hi_hi_6, readData_readResultSelect_hi_lo_6};
  wire [15:0]       readData_readResultSelect_6 = {readData_readResultSelect_hi_6, readData_readResultSelect_lo_6};
  assign readData_data_6 =
    (readData_readResultSelect_6[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_6[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_6[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_6[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_6[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_6[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_6[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_6[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_6[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_6[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_6[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_6[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_6[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_6[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_6[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_6[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_6_enq_bits = readData_data_6;
  wire              readTokenRelease_6 = readData_readDataQueue_6_deq_ready & readData_readDataQueue_6_deq_valid;
  assign readData_readDataQueue_6_enq_valid = |readData_readResultSelect_6;
  wire [31:0]       readData_data_7;
  wire              isWaiteForThisData_7;
  wire              readData_readDataQueue_7_enq_ready = ~_readData_readDataQueue_fifo_7_full;
  wire              readData_readDataQueue_7_deq_ready;
  wire              readData_readDataQueue_7_enq_valid;
  wire              readData_readDataQueue_7_deq_valid = ~_readData_readDataQueue_fifo_7_empty | readData_readDataQueue_7_enq_valid;
  wire [31:0]       readData_readDataQueue_7_enq_bits;
  wire [31:0]       readData_readDataQueue_7_deq_bits = _readData_readDataQueue_fifo_7_empty ? readData_readDataQueue_7_enq_bits : _readData_readDataQueue_fifo_7_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_7 = {write1HPipe_1[7], write1HPipe_0[7]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_7 = {write1HPipe_3[7], write1HPipe_2[7]};
  wire [3:0]        readData_readResultSelect_lo_lo_7 = {readData_readResultSelect_lo_lo_hi_7, readData_readResultSelect_lo_lo_lo_7};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_7 = {write1HPipe_5[7], write1HPipe_4[7]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_7 = {write1HPipe_7[7], write1HPipe_6[7]};
  wire [3:0]        readData_readResultSelect_lo_hi_7 = {readData_readResultSelect_lo_hi_hi_7, readData_readResultSelect_lo_hi_lo_7};
  wire [7:0]        readData_readResultSelect_lo_7 = {readData_readResultSelect_lo_hi_7, readData_readResultSelect_lo_lo_7};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_7 = {write1HPipe_9[7], write1HPipe_8[7]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_7 = {write1HPipe_11[7], write1HPipe_10[7]};
  wire [3:0]        readData_readResultSelect_hi_lo_7 = {readData_readResultSelect_hi_lo_hi_7, readData_readResultSelect_hi_lo_lo_7};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_7 = {write1HPipe_13[7], write1HPipe_12[7]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_7 = {write1HPipe_15[7], write1HPipe_14[7]};
  wire [3:0]        readData_readResultSelect_hi_hi_7 = {readData_readResultSelect_hi_hi_hi_7, readData_readResultSelect_hi_hi_lo_7};
  wire [7:0]        readData_readResultSelect_hi_7 = {readData_readResultSelect_hi_hi_7, readData_readResultSelect_hi_lo_7};
  wire [15:0]       readData_readResultSelect_7 = {readData_readResultSelect_hi_7, readData_readResultSelect_lo_7};
  assign readData_data_7 =
    (readData_readResultSelect_7[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_7[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_7[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_7[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_7[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_7[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_7[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_7[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_7[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_7[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_7[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_7[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_7[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_7[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_7[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_7[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_7_enq_bits = readData_data_7;
  wire              readTokenRelease_7 = readData_readDataQueue_7_deq_ready & readData_readDataQueue_7_deq_valid;
  assign readData_readDataQueue_7_enq_valid = |readData_readResultSelect_7;
  wire [31:0]       readData_data_8;
  wire              isWaiteForThisData_8;
  wire              readData_readDataQueue_8_enq_ready = ~_readData_readDataQueue_fifo_8_full;
  wire              readData_readDataQueue_8_deq_ready;
  wire              readData_readDataQueue_8_enq_valid;
  wire              readData_readDataQueue_8_deq_valid = ~_readData_readDataQueue_fifo_8_empty | readData_readDataQueue_8_enq_valid;
  wire [31:0]       readData_readDataQueue_8_enq_bits;
  wire [31:0]       readData_readDataQueue_8_deq_bits = _readData_readDataQueue_fifo_8_empty ? readData_readDataQueue_8_enq_bits : _readData_readDataQueue_fifo_8_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_8 = {write1HPipe_1[8], write1HPipe_0[8]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_8 = {write1HPipe_3[8], write1HPipe_2[8]};
  wire [3:0]        readData_readResultSelect_lo_lo_8 = {readData_readResultSelect_lo_lo_hi_8, readData_readResultSelect_lo_lo_lo_8};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_8 = {write1HPipe_5[8], write1HPipe_4[8]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_8 = {write1HPipe_7[8], write1HPipe_6[8]};
  wire [3:0]        readData_readResultSelect_lo_hi_8 = {readData_readResultSelect_lo_hi_hi_8, readData_readResultSelect_lo_hi_lo_8};
  wire [7:0]        readData_readResultSelect_lo_8 = {readData_readResultSelect_lo_hi_8, readData_readResultSelect_lo_lo_8};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_8 = {write1HPipe_9[8], write1HPipe_8[8]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_8 = {write1HPipe_11[8], write1HPipe_10[8]};
  wire [3:0]        readData_readResultSelect_hi_lo_8 = {readData_readResultSelect_hi_lo_hi_8, readData_readResultSelect_hi_lo_lo_8};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_8 = {write1HPipe_13[8], write1HPipe_12[8]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_8 = {write1HPipe_15[8], write1HPipe_14[8]};
  wire [3:0]        readData_readResultSelect_hi_hi_8 = {readData_readResultSelect_hi_hi_hi_8, readData_readResultSelect_hi_hi_lo_8};
  wire [7:0]        readData_readResultSelect_hi_8 = {readData_readResultSelect_hi_hi_8, readData_readResultSelect_hi_lo_8};
  wire [15:0]       readData_readResultSelect_8 = {readData_readResultSelect_hi_8, readData_readResultSelect_lo_8};
  assign readData_data_8 =
    (readData_readResultSelect_8[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_8[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_8[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_8[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_8[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_8[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_8[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_8[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_8[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_8[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_8[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_8[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_8[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_8[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_8[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_8[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_8_enq_bits = readData_data_8;
  wire              readTokenRelease_8 = readData_readDataQueue_8_deq_ready & readData_readDataQueue_8_deq_valid;
  assign readData_readDataQueue_8_enq_valid = |readData_readResultSelect_8;
  wire [31:0]       readData_data_9;
  wire              isWaiteForThisData_9;
  wire              readData_readDataQueue_9_enq_ready = ~_readData_readDataQueue_fifo_9_full;
  wire              readData_readDataQueue_9_deq_ready;
  wire              readData_readDataQueue_9_enq_valid;
  wire              readData_readDataQueue_9_deq_valid = ~_readData_readDataQueue_fifo_9_empty | readData_readDataQueue_9_enq_valid;
  wire [31:0]       readData_readDataQueue_9_enq_bits;
  wire [31:0]       readData_readDataQueue_9_deq_bits = _readData_readDataQueue_fifo_9_empty ? readData_readDataQueue_9_enq_bits : _readData_readDataQueue_fifo_9_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_9 = {write1HPipe_1[9], write1HPipe_0[9]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_9 = {write1HPipe_3[9], write1HPipe_2[9]};
  wire [3:0]        readData_readResultSelect_lo_lo_9 = {readData_readResultSelect_lo_lo_hi_9, readData_readResultSelect_lo_lo_lo_9};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_9 = {write1HPipe_5[9], write1HPipe_4[9]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_9 = {write1HPipe_7[9], write1HPipe_6[9]};
  wire [3:0]        readData_readResultSelect_lo_hi_9 = {readData_readResultSelect_lo_hi_hi_9, readData_readResultSelect_lo_hi_lo_9};
  wire [7:0]        readData_readResultSelect_lo_9 = {readData_readResultSelect_lo_hi_9, readData_readResultSelect_lo_lo_9};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_9 = {write1HPipe_9[9], write1HPipe_8[9]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_9 = {write1HPipe_11[9], write1HPipe_10[9]};
  wire [3:0]        readData_readResultSelect_hi_lo_9 = {readData_readResultSelect_hi_lo_hi_9, readData_readResultSelect_hi_lo_lo_9};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_9 = {write1HPipe_13[9], write1HPipe_12[9]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_9 = {write1HPipe_15[9], write1HPipe_14[9]};
  wire [3:0]        readData_readResultSelect_hi_hi_9 = {readData_readResultSelect_hi_hi_hi_9, readData_readResultSelect_hi_hi_lo_9};
  wire [7:0]        readData_readResultSelect_hi_9 = {readData_readResultSelect_hi_hi_9, readData_readResultSelect_hi_lo_9};
  wire [15:0]       readData_readResultSelect_9 = {readData_readResultSelect_hi_9, readData_readResultSelect_lo_9};
  assign readData_data_9 =
    (readData_readResultSelect_9[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_9[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_9[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_9[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_9[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_9[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_9[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_9[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_9[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_9[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_9[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_9[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_9[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_9[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_9[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_9[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_9_enq_bits = readData_data_9;
  wire              readTokenRelease_9 = readData_readDataQueue_9_deq_ready & readData_readDataQueue_9_deq_valid;
  assign readData_readDataQueue_9_enq_valid = |readData_readResultSelect_9;
  wire [31:0]       readData_data_10;
  wire              isWaiteForThisData_10;
  wire              readData_readDataQueue_10_enq_ready = ~_readData_readDataQueue_fifo_10_full;
  wire              readData_readDataQueue_10_deq_ready;
  wire              readData_readDataQueue_10_enq_valid;
  wire              readData_readDataQueue_10_deq_valid = ~_readData_readDataQueue_fifo_10_empty | readData_readDataQueue_10_enq_valid;
  wire [31:0]       readData_readDataQueue_10_enq_bits;
  wire [31:0]       readData_readDataQueue_10_deq_bits = _readData_readDataQueue_fifo_10_empty ? readData_readDataQueue_10_enq_bits : _readData_readDataQueue_fifo_10_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_10 = {write1HPipe_1[10], write1HPipe_0[10]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_10 = {write1HPipe_3[10], write1HPipe_2[10]};
  wire [3:0]        readData_readResultSelect_lo_lo_10 = {readData_readResultSelect_lo_lo_hi_10, readData_readResultSelect_lo_lo_lo_10};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_10 = {write1HPipe_5[10], write1HPipe_4[10]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_10 = {write1HPipe_7[10], write1HPipe_6[10]};
  wire [3:0]        readData_readResultSelect_lo_hi_10 = {readData_readResultSelect_lo_hi_hi_10, readData_readResultSelect_lo_hi_lo_10};
  wire [7:0]        readData_readResultSelect_lo_10 = {readData_readResultSelect_lo_hi_10, readData_readResultSelect_lo_lo_10};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_10 = {write1HPipe_9[10], write1HPipe_8[10]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_10 = {write1HPipe_11[10], write1HPipe_10[10]};
  wire [3:0]        readData_readResultSelect_hi_lo_10 = {readData_readResultSelect_hi_lo_hi_10, readData_readResultSelect_hi_lo_lo_10};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_10 = {write1HPipe_13[10], write1HPipe_12[10]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_10 = {write1HPipe_15[10], write1HPipe_14[10]};
  wire [3:0]        readData_readResultSelect_hi_hi_10 = {readData_readResultSelect_hi_hi_hi_10, readData_readResultSelect_hi_hi_lo_10};
  wire [7:0]        readData_readResultSelect_hi_10 = {readData_readResultSelect_hi_hi_10, readData_readResultSelect_hi_lo_10};
  wire [15:0]       readData_readResultSelect_10 = {readData_readResultSelect_hi_10, readData_readResultSelect_lo_10};
  assign readData_data_10 =
    (readData_readResultSelect_10[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_10[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_10[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_10[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_10[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_10[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_10[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_10[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_10[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_10[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_10[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_10[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_10[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_10[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_10[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_10[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_10_enq_bits = readData_data_10;
  wire              readTokenRelease_10 = readData_readDataQueue_10_deq_ready & readData_readDataQueue_10_deq_valid;
  assign readData_readDataQueue_10_enq_valid = |readData_readResultSelect_10;
  wire [31:0]       readData_data_11;
  wire              isWaiteForThisData_11;
  wire              readData_readDataQueue_11_enq_ready = ~_readData_readDataQueue_fifo_11_full;
  wire              readData_readDataQueue_11_deq_ready;
  wire              readData_readDataQueue_11_enq_valid;
  wire              readData_readDataQueue_11_deq_valid = ~_readData_readDataQueue_fifo_11_empty | readData_readDataQueue_11_enq_valid;
  wire [31:0]       readData_readDataQueue_11_enq_bits;
  wire [31:0]       readData_readDataQueue_11_deq_bits = _readData_readDataQueue_fifo_11_empty ? readData_readDataQueue_11_enq_bits : _readData_readDataQueue_fifo_11_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_11 = {write1HPipe_1[11], write1HPipe_0[11]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_11 = {write1HPipe_3[11], write1HPipe_2[11]};
  wire [3:0]        readData_readResultSelect_lo_lo_11 = {readData_readResultSelect_lo_lo_hi_11, readData_readResultSelect_lo_lo_lo_11};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_11 = {write1HPipe_5[11], write1HPipe_4[11]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_11 = {write1HPipe_7[11], write1HPipe_6[11]};
  wire [3:0]        readData_readResultSelect_lo_hi_11 = {readData_readResultSelect_lo_hi_hi_11, readData_readResultSelect_lo_hi_lo_11};
  wire [7:0]        readData_readResultSelect_lo_11 = {readData_readResultSelect_lo_hi_11, readData_readResultSelect_lo_lo_11};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_11 = {write1HPipe_9[11], write1HPipe_8[11]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_11 = {write1HPipe_11[11], write1HPipe_10[11]};
  wire [3:0]        readData_readResultSelect_hi_lo_11 = {readData_readResultSelect_hi_lo_hi_11, readData_readResultSelect_hi_lo_lo_11};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_11 = {write1HPipe_13[11], write1HPipe_12[11]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_11 = {write1HPipe_15[11], write1HPipe_14[11]};
  wire [3:0]        readData_readResultSelect_hi_hi_11 = {readData_readResultSelect_hi_hi_hi_11, readData_readResultSelect_hi_hi_lo_11};
  wire [7:0]        readData_readResultSelect_hi_11 = {readData_readResultSelect_hi_hi_11, readData_readResultSelect_hi_lo_11};
  wire [15:0]       readData_readResultSelect_11 = {readData_readResultSelect_hi_11, readData_readResultSelect_lo_11};
  assign readData_data_11 =
    (readData_readResultSelect_11[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_11[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_11[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_11[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_11[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_11[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_11[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_11[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_11[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_11[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_11[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_11[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_11[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_11[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_11[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_11[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_11_enq_bits = readData_data_11;
  wire              readTokenRelease_11 = readData_readDataQueue_11_deq_ready & readData_readDataQueue_11_deq_valid;
  assign readData_readDataQueue_11_enq_valid = |readData_readResultSelect_11;
  wire [31:0]       readData_data_12;
  wire              isWaiteForThisData_12;
  wire              readData_readDataQueue_12_enq_ready = ~_readData_readDataQueue_fifo_12_full;
  wire              readData_readDataQueue_12_deq_ready;
  wire              readData_readDataQueue_12_enq_valid;
  wire              readData_readDataQueue_12_deq_valid = ~_readData_readDataQueue_fifo_12_empty | readData_readDataQueue_12_enq_valid;
  wire [31:0]       readData_readDataQueue_12_enq_bits;
  wire [31:0]       readData_readDataQueue_12_deq_bits = _readData_readDataQueue_fifo_12_empty ? readData_readDataQueue_12_enq_bits : _readData_readDataQueue_fifo_12_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_12 = {write1HPipe_1[12], write1HPipe_0[12]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_12 = {write1HPipe_3[12], write1HPipe_2[12]};
  wire [3:0]        readData_readResultSelect_lo_lo_12 = {readData_readResultSelect_lo_lo_hi_12, readData_readResultSelect_lo_lo_lo_12};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_12 = {write1HPipe_5[12], write1HPipe_4[12]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_12 = {write1HPipe_7[12], write1HPipe_6[12]};
  wire [3:0]        readData_readResultSelect_lo_hi_12 = {readData_readResultSelect_lo_hi_hi_12, readData_readResultSelect_lo_hi_lo_12};
  wire [7:0]        readData_readResultSelect_lo_12 = {readData_readResultSelect_lo_hi_12, readData_readResultSelect_lo_lo_12};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_12 = {write1HPipe_9[12], write1HPipe_8[12]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_12 = {write1HPipe_11[12], write1HPipe_10[12]};
  wire [3:0]        readData_readResultSelect_hi_lo_12 = {readData_readResultSelect_hi_lo_hi_12, readData_readResultSelect_hi_lo_lo_12};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_12 = {write1HPipe_13[12], write1HPipe_12[12]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_12 = {write1HPipe_15[12], write1HPipe_14[12]};
  wire [3:0]        readData_readResultSelect_hi_hi_12 = {readData_readResultSelect_hi_hi_hi_12, readData_readResultSelect_hi_hi_lo_12};
  wire [7:0]        readData_readResultSelect_hi_12 = {readData_readResultSelect_hi_hi_12, readData_readResultSelect_hi_lo_12};
  wire [15:0]       readData_readResultSelect_12 = {readData_readResultSelect_hi_12, readData_readResultSelect_lo_12};
  assign readData_data_12 =
    (readData_readResultSelect_12[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_12[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_12[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_12[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_12[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_12[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_12[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_12[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_12[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_12[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_12[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_12[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_12[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_12[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_12[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_12[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_12_enq_bits = readData_data_12;
  wire              readTokenRelease_12 = readData_readDataQueue_12_deq_ready & readData_readDataQueue_12_deq_valid;
  assign readData_readDataQueue_12_enq_valid = |readData_readResultSelect_12;
  wire [31:0]       readData_data_13;
  wire              isWaiteForThisData_13;
  wire              readData_readDataQueue_13_enq_ready = ~_readData_readDataQueue_fifo_13_full;
  wire              readData_readDataQueue_13_deq_ready;
  wire              readData_readDataQueue_13_enq_valid;
  wire              readData_readDataQueue_13_deq_valid = ~_readData_readDataQueue_fifo_13_empty | readData_readDataQueue_13_enq_valid;
  wire [31:0]       readData_readDataQueue_13_enq_bits;
  wire [31:0]       readData_readDataQueue_13_deq_bits = _readData_readDataQueue_fifo_13_empty ? readData_readDataQueue_13_enq_bits : _readData_readDataQueue_fifo_13_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_13 = {write1HPipe_1[13], write1HPipe_0[13]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_13 = {write1HPipe_3[13], write1HPipe_2[13]};
  wire [3:0]        readData_readResultSelect_lo_lo_13 = {readData_readResultSelect_lo_lo_hi_13, readData_readResultSelect_lo_lo_lo_13};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_13 = {write1HPipe_5[13], write1HPipe_4[13]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_13 = {write1HPipe_7[13], write1HPipe_6[13]};
  wire [3:0]        readData_readResultSelect_lo_hi_13 = {readData_readResultSelect_lo_hi_hi_13, readData_readResultSelect_lo_hi_lo_13};
  wire [7:0]        readData_readResultSelect_lo_13 = {readData_readResultSelect_lo_hi_13, readData_readResultSelect_lo_lo_13};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_13 = {write1HPipe_9[13], write1HPipe_8[13]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_13 = {write1HPipe_11[13], write1HPipe_10[13]};
  wire [3:0]        readData_readResultSelect_hi_lo_13 = {readData_readResultSelect_hi_lo_hi_13, readData_readResultSelect_hi_lo_lo_13};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_13 = {write1HPipe_13[13], write1HPipe_12[13]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_13 = {write1HPipe_15[13], write1HPipe_14[13]};
  wire [3:0]        readData_readResultSelect_hi_hi_13 = {readData_readResultSelect_hi_hi_hi_13, readData_readResultSelect_hi_hi_lo_13};
  wire [7:0]        readData_readResultSelect_hi_13 = {readData_readResultSelect_hi_hi_13, readData_readResultSelect_hi_lo_13};
  wire [15:0]       readData_readResultSelect_13 = {readData_readResultSelect_hi_13, readData_readResultSelect_lo_13};
  assign readData_data_13 =
    (readData_readResultSelect_13[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_13[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_13[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_13[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_13[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_13[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_13[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_13[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_13[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_13[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_13[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_13[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_13[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_13[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_13[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_13[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_13_enq_bits = readData_data_13;
  wire              readTokenRelease_13 = readData_readDataQueue_13_deq_ready & readData_readDataQueue_13_deq_valid;
  assign readData_readDataQueue_13_enq_valid = |readData_readResultSelect_13;
  wire [31:0]       readData_data_14;
  wire              isWaiteForThisData_14;
  wire              readData_readDataQueue_14_enq_ready = ~_readData_readDataQueue_fifo_14_full;
  wire              readData_readDataQueue_14_deq_ready;
  wire              readData_readDataQueue_14_enq_valid;
  wire              readData_readDataQueue_14_deq_valid = ~_readData_readDataQueue_fifo_14_empty | readData_readDataQueue_14_enq_valid;
  wire [31:0]       readData_readDataQueue_14_enq_bits;
  wire [31:0]       readData_readDataQueue_14_deq_bits = _readData_readDataQueue_fifo_14_empty ? readData_readDataQueue_14_enq_bits : _readData_readDataQueue_fifo_14_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_14 = {write1HPipe_1[14], write1HPipe_0[14]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_14 = {write1HPipe_3[14], write1HPipe_2[14]};
  wire [3:0]        readData_readResultSelect_lo_lo_14 = {readData_readResultSelect_lo_lo_hi_14, readData_readResultSelect_lo_lo_lo_14};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_14 = {write1HPipe_5[14], write1HPipe_4[14]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_14 = {write1HPipe_7[14], write1HPipe_6[14]};
  wire [3:0]        readData_readResultSelect_lo_hi_14 = {readData_readResultSelect_lo_hi_hi_14, readData_readResultSelect_lo_hi_lo_14};
  wire [7:0]        readData_readResultSelect_lo_14 = {readData_readResultSelect_lo_hi_14, readData_readResultSelect_lo_lo_14};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_14 = {write1HPipe_9[14], write1HPipe_8[14]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_14 = {write1HPipe_11[14], write1HPipe_10[14]};
  wire [3:0]        readData_readResultSelect_hi_lo_14 = {readData_readResultSelect_hi_lo_hi_14, readData_readResultSelect_hi_lo_lo_14};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_14 = {write1HPipe_13[14], write1HPipe_12[14]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_14 = {write1HPipe_15[14], write1HPipe_14[14]};
  wire [3:0]        readData_readResultSelect_hi_hi_14 = {readData_readResultSelect_hi_hi_hi_14, readData_readResultSelect_hi_hi_lo_14};
  wire [7:0]        readData_readResultSelect_hi_14 = {readData_readResultSelect_hi_hi_14, readData_readResultSelect_hi_lo_14};
  wire [15:0]       readData_readResultSelect_14 = {readData_readResultSelect_hi_14, readData_readResultSelect_lo_14};
  assign readData_data_14 =
    (readData_readResultSelect_14[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_14[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_14[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_14[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_14[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_14[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_14[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_14[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_14[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_14[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_14[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_14[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_14[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_14[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_14[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_14[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_14_enq_bits = readData_data_14;
  wire              readTokenRelease_14 = readData_readDataQueue_14_deq_ready & readData_readDataQueue_14_deq_valid;
  assign readData_readDataQueue_14_enq_valid = |readData_readResultSelect_14;
  wire [31:0]       readData_data_15;
  wire              isWaiteForThisData_15;
  wire              readData_readDataQueue_15_enq_ready = ~_readData_readDataQueue_fifo_15_full;
  wire              readData_readDataQueue_15_deq_ready;
  wire              readData_readDataQueue_15_enq_valid;
  wire              readData_readDataQueue_15_deq_valid = ~_readData_readDataQueue_fifo_15_empty | readData_readDataQueue_15_enq_valid;
  wire [31:0]       readData_readDataQueue_15_enq_bits;
  wire [31:0]       readData_readDataQueue_15_deq_bits = _readData_readDataQueue_fifo_15_empty ? readData_readDataQueue_15_enq_bits : _readData_readDataQueue_fifo_15_data_out;
  wire [1:0]        readData_readResultSelect_lo_lo_lo_15 = {write1HPipe_1[15], write1HPipe_0[15]};
  wire [1:0]        readData_readResultSelect_lo_lo_hi_15 = {write1HPipe_3[15], write1HPipe_2[15]};
  wire [3:0]        readData_readResultSelect_lo_lo_15 = {readData_readResultSelect_lo_lo_hi_15, readData_readResultSelect_lo_lo_lo_15};
  wire [1:0]        readData_readResultSelect_lo_hi_lo_15 = {write1HPipe_5[15], write1HPipe_4[15]};
  wire [1:0]        readData_readResultSelect_lo_hi_hi_15 = {write1HPipe_7[15], write1HPipe_6[15]};
  wire [3:0]        readData_readResultSelect_lo_hi_15 = {readData_readResultSelect_lo_hi_hi_15, readData_readResultSelect_lo_hi_lo_15};
  wire [7:0]        readData_readResultSelect_lo_15 = {readData_readResultSelect_lo_hi_15, readData_readResultSelect_lo_lo_15};
  wire [1:0]        readData_readResultSelect_hi_lo_lo_15 = {write1HPipe_9[15], write1HPipe_8[15]};
  wire [1:0]        readData_readResultSelect_hi_lo_hi_15 = {write1HPipe_11[15], write1HPipe_10[15]};
  wire [3:0]        readData_readResultSelect_hi_lo_15 = {readData_readResultSelect_hi_lo_hi_15, readData_readResultSelect_hi_lo_lo_15};
  wire [1:0]        readData_readResultSelect_hi_hi_lo_15 = {write1HPipe_13[15], write1HPipe_12[15]};
  wire [1:0]        readData_readResultSelect_hi_hi_hi_15 = {write1HPipe_15[15], write1HPipe_14[15]};
  wire [3:0]        readData_readResultSelect_hi_hi_15 = {readData_readResultSelect_hi_hi_hi_15, readData_readResultSelect_hi_hi_lo_15};
  wire [7:0]        readData_readResultSelect_hi_15 = {readData_readResultSelect_hi_hi_15, readData_readResultSelect_hi_lo_15};
  wire [15:0]       readData_readResultSelect_15 = {readData_readResultSelect_hi_15, readData_readResultSelect_lo_15};
  assign readData_data_15 =
    (readData_readResultSelect_15[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_15[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_15[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_15[3] ? dataAfterReorderCheck_3 : 32'h0) | (readData_readResultSelect_15[4] ? dataAfterReorderCheck_4 : 32'h0) | (readData_readResultSelect_15[5] ? dataAfterReorderCheck_5 : 32'h0)
    | (readData_readResultSelect_15[6] ? dataAfterReorderCheck_6 : 32'h0) | (readData_readResultSelect_15[7] ? dataAfterReorderCheck_7 : 32'h0) | (readData_readResultSelect_15[8] ? dataAfterReorderCheck_8 : 32'h0)
    | (readData_readResultSelect_15[9] ? dataAfterReorderCheck_9 : 32'h0) | (readData_readResultSelect_15[10] ? dataAfterReorderCheck_10 : 32'h0) | (readData_readResultSelect_15[11] ? dataAfterReorderCheck_11 : 32'h0)
    | (readData_readResultSelect_15[12] ? dataAfterReorderCheck_12 : 32'h0) | (readData_readResultSelect_15[13] ? dataAfterReorderCheck_13 : 32'h0) | (readData_readResultSelect_15[14] ? dataAfterReorderCheck_14 : 32'h0)
    | (readData_readResultSelect_15[15] ? dataAfterReorderCheck_15 : 32'h0);
  assign readData_readDataQueue_15_enq_bits = readData_data_15;
  wire              readTokenRelease_15 = readData_readDataQueue_15_deq_ready & readData_readDataQueue_15_deq_valid;
  assign readData_readDataQueue_15_enq_valid = |readData_readResultSelect_15;
  reg  [6:0]        waiteReadDataPipeReg_executeGroup;
  reg  [15:0]       waiteReadDataPipeReg_sourceValid;
  reg  [15:0]       waiteReadDataPipeReg_replaceVs1;
  reg  [15:0]       waiteReadDataPipeReg_needRead;
  reg               waiteReadDataPipeReg_last;
  reg  [31:0]       waiteReadData_0;
  reg  [31:0]       waiteReadData_1;
  reg  [31:0]       waiteReadData_2;
  reg  [31:0]       waiteReadData_3;
  reg  [31:0]       waiteReadData_4;
  reg  [31:0]       waiteReadData_5;
  reg  [31:0]       waiteReadData_6;
  reg  [31:0]       waiteReadData_7;
  reg  [31:0]       waiteReadData_8;
  reg  [31:0]       waiteReadData_9;
  reg  [31:0]       waiteReadData_10;
  reg  [31:0]       waiteReadData_11;
  reg  [31:0]       waiteReadData_12;
  reg  [31:0]       waiteReadData_13;
  reg  [31:0]       waiteReadData_14;
  reg  [31:0]       waiteReadData_15;
  reg  [15:0]       waiteReadSate;
  reg               waiteReadStageValid;
  wire [1:0]        executeIndexVec_0 = waiteReadDataPipeReg_executeGroup[1:0];
  wire [1:0]        executeIndexVec_1 = {waiteReadDataPipeReg_executeGroup[0], 1'h0};
  wire              writeDataVec_data_dataIsRead = waiteReadDataPipeReg_needRead[0];
  wire              writeDataVec_data_dataIsRead_16 = waiteReadDataPipeReg_needRead[0];
  wire              writeDataVec_data_dataIsRead_32 = waiteReadDataPipeReg_needRead[0];
  wire [31:0]       _GEN_92 = waiteReadDataPipeReg_replaceVs1[0] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData;
  assign writeDataVec_data_unreadData = _GEN_92;
  wire [31:0]       writeDataVec_data_unreadData_16;
  assign writeDataVec_data_unreadData_16 = _GEN_92;
  wire [31:0]       writeDataVec_data_unreadData_32;
  assign writeDataVec_data_unreadData_32 = _GEN_92;
  wire [7:0]        writeDataVec_data_dataElement = writeDataVec_data_dataIsRead ? waiteReadData_0[7:0] : writeDataVec_data_unreadData[7:0];
  wire              writeDataVec_data_dataIsRead_1 = waiteReadDataPipeReg_needRead[1];
  wire              writeDataVec_data_dataIsRead_17 = waiteReadDataPipeReg_needRead[1];
  wire              writeDataVec_data_dataIsRead_33 = waiteReadDataPipeReg_needRead[1];
  wire [31:0]       _GEN_93 = waiteReadDataPipeReg_replaceVs1[1] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_1;
  assign writeDataVec_data_unreadData_1 = _GEN_93;
  wire [31:0]       writeDataVec_data_unreadData_17;
  assign writeDataVec_data_unreadData_17 = _GEN_93;
  wire [31:0]       writeDataVec_data_unreadData_33;
  assign writeDataVec_data_unreadData_33 = _GEN_93;
  wire [7:0]        writeDataVec_data_dataElement_1 = writeDataVec_data_dataIsRead_1 ? waiteReadData_1[7:0] : writeDataVec_data_unreadData_1[7:0];
  wire              writeDataVec_data_dataIsRead_2 = waiteReadDataPipeReg_needRead[2];
  wire              writeDataVec_data_dataIsRead_18 = waiteReadDataPipeReg_needRead[2];
  wire              writeDataVec_data_dataIsRead_34 = waiteReadDataPipeReg_needRead[2];
  wire [31:0]       _GEN_94 = waiteReadDataPipeReg_replaceVs1[2] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_2;
  assign writeDataVec_data_unreadData_2 = _GEN_94;
  wire [31:0]       writeDataVec_data_unreadData_18;
  assign writeDataVec_data_unreadData_18 = _GEN_94;
  wire [31:0]       writeDataVec_data_unreadData_34;
  assign writeDataVec_data_unreadData_34 = _GEN_94;
  wire [7:0]        writeDataVec_data_dataElement_2 = writeDataVec_data_dataIsRead_2 ? waiteReadData_2[7:0] : writeDataVec_data_unreadData_2[7:0];
  wire              writeDataVec_data_dataIsRead_3 = waiteReadDataPipeReg_needRead[3];
  wire              writeDataVec_data_dataIsRead_19 = waiteReadDataPipeReg_needRead[3];
  wire              writeDataVec_data_dataIsRead_35 = waiteReadDataPipeReg_needRead[3];
  wire [31:0]       _GEN_95 = waiteReadDataPipeReg_replaceVs1[3] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_3;
  assign writeDataVec_data_unreadData_3 = _GEN_95;
  wire [31:0]       writeDataVec_data_unreadData_19;
  assign writeDataVec_data_unreadData_19 = _GEN_95;
  wire [31:0]       writeDataVec_data_unreadData_35;
  assign writeDataVec_data_unreadData_35 = _GEN_95;
  wire [7:0]        writeDataVec_data_dataElement_3 = writeDataVec_data_dataIsRead_3 ? waiteReadData_3[7:0] : writeDataVec_data_unreadData_3[7:0];
  wire              writeDataVec_data_dataIsRead_4 = waiteReadDataPipeReg_needRead[4];
  wire              writeDataVec_data_dataIsRead_20 = waiteReadDataPipeReg_needRead[4];
  wire              writeDataVec_data_dataIsRead_36 = waiteReadDataPipeReg_needRead[4];
  wire [31:0]       _GEN_96 = waiteReadDataPipeReg_replaceVs1[4] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_4;
  assign writeDataVec_data_unreadData_4 = _GEN_96;
  wire [31:0]       writeDataVec_data_unreadData_20;
  assign writeDataVec_data_unreadData_20 = _GEN_96;
  wire [31:0]       writeDataVec_data_unreadData_36;
  assign writeDataVec_data_unreadData_36 = _GEN_96;
  wire [7:0]        writeDataVec_data_dataElement_4 = writeDataVec_data_dataIsRead_4 ? waiteReadData_4[7:0] : writeDataVec_data_unreadData_4[7:0];
  wire              writeDataVec_data_dataIsRead_5 = waiteReadDataPipeReg_needRead[5];
  wire              writeDataVec_data_dataIsRead_21 = waiteReadDataPipeReg_needRead[5];
  wire              writeDataVec_data_dataIsRead_37 = waiteReadDataPipeReg_needRead[5];
  wire [31:0]       _GEN_97 = waiteReadDataPipeReg_replaceVs1[5] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_5;
  assign writeDataVec_data_unreadData_5 = _GEN_97;
  wire [31:0]       writeDataVec_data_unreadData_21;
  assign writeDataVec_data_unreadData_21 = _GEN_97;
  wire [31:0]       writeDataVec_data_unreadData_37;
  assign writeDataVec_data_unreadData_37 = _GEN_97;
  wire [7:0]        writeDataVec_data_dataElement_5 = writeDataVec_data_dataIsRead_5 ? waiteReadData_5[7:0] : writeDataVec_data_unreadData_5[7:0];
  wire              writeDataVec_data_dataIsRead_6 = waiteReadDataPipeReg_needRead[6];
  wire              writeDataVec_data_dataIsRead_22 = waiteReadDataPipeReg_needRead[6];
  wire              writeDataVec_data_dataIsRead_38 = waiteReadDataPipeReg_needRead[6];
  wire [31:0]       _GEN_98 = waiteReadDataPipeReg_replaceVs1[6] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_6;
  assign writeDataVec_data_unreadData_6 = _GEN_98;
  wire [31:0]       writeDataVec_data_unreadData_22;
  assign writeDataVec_data_unreadData_22 = _GEN_98;
  wire [31:0]       writeDataVec_data_unreadData_38;
  assign writeDataVec_data_unreadData_38 = _GEN_98;
  wire [7:0]        writeDataVec_data_dataElement_6 = writeDataVec_data_dataIsRead_6 ? waiteReadData_6[7:0] : writeDataVec_data_unreadData_6[7:0];
  wire              writeDataVec_data_dataIsRead_7 = waiteReadDataPipeReg_needRead[7];
  wire              writeDataVec_data_dataIsRead_23 = waiteReadDataPipeReg_needRead[7];
  wire              writeDataVec_data_dataIsRead_39 = waiteReadDataPipeReg_needRead[7];
  wire [31:0]       _GEN_99 = waiteReadDataPipeReg_replaceVs1[7] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_7;
  assign writeDataVec_data_unreadData_7 = _GEN_99;
  wire [31:0]       writeDataVec_data_unreadData_23;
  assign writeDataVec_data_unreadData_23 = _GEN_99;
  wire [31:0]       writeDataVec_data_unreadData_39;
  assign writeDataVec_data_unreadData_39 = _GEN_99;
  wire [7:0]        writeDataVec_data_dataElement_7 = writeDataVec_data_dataIsRead_7 ? waiteReadData_7[7:0] : writeDataVec_data_unreadData_7[7:0];
  wire              writeDataVec_data_dataIsRead_8 = waiteReadDataPipeReg_needRead[8];
  wire              writeDataVec_data_dataIsRead_24 = waiteReadDataPipeReg_needRead[8];
  wire              writeDataVec_data_dataIsRead_40 = waiteReadDataPipeReg_needRead[8];
  wire [31:0]       _GEN_100 = waiteReadDataPipeReg_replaceVs1[8] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_8;
  assign writeDataVec_data_unreadData_8 = _GEN_100;
  wire [31:0]       writeDataVec_data_unreadData_24;
  assign writeDataVec_data_unreadData_24 = _GEN_100;
  wire [31:0]       writeDataVec_data_unreadData_40;
  assign writeDataVec_data_unreadData_40 = _GEN_100;
  wire [7:0]        writeDataVec_data_dataElement_8 = writeDataVec_data_dataIsRead_8 ? waiteReadData_8[7:0] : writeDataVec_data_unreadData_8[7:0];
  wire              writeDataVec_data_dataIsRead_9 = waiteReadDataPipeReg_needRead[9];
  wire              writeDataVec_data_dataIsRead_25 = waiteReadDataPipeReg_needRead[9];
  wire              writeDataVec_data_dataIsRead_41 = waiteReadDataPipeReg_needRead[9];
  wire [31:0]       _GEN_101 = waiteReadDataPipeReg_replaceVs1[9] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_9;
  assign writeDataVec_data_unreadData_9 = _GEN_101;
  wire [31:0]       writeDataVec_data_unreadData_25;
  assign writeDataVec_data_unreadData_25 = _GEN_101;
  wire [31:0]       writeDataVec_data_unreadData_41;
  assign writeDataVec_data_unreadData_41 = _GEN_101;
  wire [7:0]        writeDataVec_data_dataElement_9 = writeDataVec_data_dataIsRead_9 ? waiteReadData_9[7:0] : writeDataVec_data_unreadData_9[7:0];
  wire              writeDataVec_data_dataIsRead_10 = waiteReadDataPipeReg_needRead[10];
  wire              writeDataVec_data_dataIsRead_26 = waiteReadDataPipeReg_needRead[10];
  wire              writeDataVec_data_dataIsRead_42 = waiteReadDataPipeReg_needRead[10];
  wire [31:0]       _GEN_102 = waiteReadDataPipeReg_replaceVs1[10] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_10;
  assign writeDataVec_data_unreadData_10 = _GEN_102;
  wire [31:0]       writeDataVec_data_unreadData_26;
  assign writeDataVec_data_unreadData_26 = _GEN_102;
  wire [31:0]       writeDataVec_data_unreadData_42;
  assign writeDataVec_data_unreadData_42 = _GEN_102;
  wire [7:0]        writeDataVec_data_dataElement_10 = writeDataVec_data_dataIsRead_10 ? waiteReadData_10[7:0] : writeDataVec_data_unreadData_10[7:0];
  wire              writeDataVec_data_dataIsRead_11 = waiteReadDataPipeReg_needRead[11];
  wire              writeDataVec_data_dataIsRead_27 = waiteReadDataPipeReg_needRead[11];
  wire              writeDataVec_data_dataIsRead_43 = waiteReadDataPipeReg_needRead[11];
  wire [31:0]       _GEN_103 = waiteReadDataPipeReg_replaceVs1[11] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_11;
  assign writeDataVec_data_unreadData_11 = _GEN_103;
  wire [31:0]       writeDataVec_data_unreadData_27;
  assign writeDataVec_data_unreadData_27 = _GEN_103;
  wire [31:0]       writeDataVec_data_unreadData_43;
  assign writeDataVec_data_unreadData_43 = _GEN_103;
  wire [7:0]        writeDataVec_data_dataElement_11 = writeDataVec_data_dataIsRead_11 ? waiteReadData_11[7:0] : writeDataVec_data_unreadData_11[7:0];
  wire              writeDataVec_data_dataIsRead_12 = waiteReadDataPipeReg_needRead[12];
  wire              writeDataVec_data_dataIsRead_28 = waiteReadDataPipeReg_needRead[12];
  wire              writeDataVec_data_dataIsRead_44 = waiteReadDataPipeReg_needRead[12];
  wire [31:0]       _GEN_104 = waiteReadDataPipeReg_replaceVs1[12] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_12;
  assign writeDataVec_data_unreadData_12 = _GEN_104;
  wire [31:0]       writeDataVec_data_unreadData_28;
  assign writeDataVec_data_unreadData_28 = _GEN_104;
  wire [31:0]       writeDataVec_data_unreadData_44;
  assign writeDataVec_data_unreadData_44 = _GEN_104;
  wire [7:0]        writeDataVec_data_dataElement_12 = writeDataVec_data_dataIsRead_12 ? waiteReadData_12[7:0] : writeDataVec_data_unreadData_12[7:0];
  wire              writeDataVec_data_dataIsRead_13 = waiteReadDataPipeReg_needRead[13];
  wire              writeDataVec_data_dataIsRead_29 = waiteReadDataPipeReg_needRead[13];
  wire              writeDataVec_data_dataIsRead_45 = waiteReadDataPipeReg_needRead[13];
  wire [31:0]       _GEN_105 = waiteReadDataPipeReg_replaceVs1[13] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_13;
  assign writeDataVec_data_unreadData_13 = _GEN_105;
  wire [31:0]       writeDataVec_data_unreadData_29;
  assign writeDataVec_data_unreadData_29 = _GEN_105;
  wire [31:0]       writeDataVec_data_unreadData_45;
  assign writeDataVec_data_unreadData_45 = _GEN_105;
  wire [7:0]        writeDataVec_data_dataElement_13 = writeDataVec_data_dataIsRead_13 ? waiteReadData_13[7:0] : writeDataVec_data_unreadData_13[7:0];
  wire              writeDataVec_data_dataIsRead_14 = waiteReadDataPipeReg_needRead[14];
  wire              writeDataVec_data_dataIsRead_30 = waiteReadDataPipeReg_needRead[14];
  wire              writeDataVec_data_dataIsRead_46 = waiteReadDataPipeReg_needRead[14];
  wire [31:0]       _GEN_109 = waiteReadDataPipeReg_replaceVs1[14] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_14;
  assign writeDataVec_data_unreadData_14 = _GEN_109;
  wire [31:0]       writeDataVec_data_unreadData_30;
  assign writeDataVec_data_unreadData_30 = _GEN_109;
  wire [31:0]       writeDataVec_data_unreadData_46;
  assign writeDataVec_data_unreadData_46 = _GEN_109;
  wire [7:0]        writeDataVec_data_dataElement_14 = writeDataVec_data_dataIsRead_14 ? waiteReadData_14[7:0] : writeDataVec_data_unreadData_14[7:0];
  wire              writeDataVec_data_dataIsRead_15 = waiteReadDataPipeReg_needRead[15];
  wire              writeDataVec_data_dataIsRead_31 = waiteReadDataPipeReg_needRead[15];
  wire              writeDataVec_data_dataIsRead_47 = waiteReadDataPipeReg_needRead[15];
  wire [31:0]       _GEN_110 = waiteReadDataPipeReg_replaceVs1[15] ? instReg_readFromScala : 32'h0;
  wire [31:0]       writeDataVec_data_unreadData_15;
  assign writeDataVec_data_unreadData_15 = _GEN_110;
  wire [31:0]       writeDataVec_data_unreadData_31;
  assign writeDataVec_data_unreadData_31 = _GEN_110;
  wire [31:0]       writeDataVec_data_unreadData_47;
  assign writeDataVec_data_unreadData_47 = _GEN_110;
  wire [7:0]        writeDataVec_data_dataElement_15 = writeDataVec_data_dataIsRead_15 ? waiteReadData_15[7:0] : writeDataVec_data_unreadData_15[7:0];
  wire [15:0]       writeDataVec_data_lo_lo_lo = {writeDataVec_data_dataElement_1, writeDataVec_data_dataElement};
  wire [15:0]       writeDataVec_data_lo_lo_hi = {writeDataVec_data_dataElement_3, writeDataVec_data_dataElement_2};
  wire [31:0]       writeDataVec_data_lo_lo = {writeDataVec_data_lo_lo_hi, writeDataVec_data_lo_lo_lo};
  wire [15:0]       writeDataVec_data_lo_hi_lo = {writeDataVec_data_dataElement_5, writeDataVec_data_dataElement_4};
  wire [15:0]       writeDataVec_data_lo_hi_hi = {writeDataVec_data_dataElement_7, writeDataVec_data_dataElement_6};
  wire [31:0]       writeDataVec_data_lo_hi = {writeDataVec_data_lo_hi_hi, writeDataVec_data_lo_hi_lo};
  wire [63:0]       writeDataVec_data_lo = {writeDataVec_data_lo_hi, writeDataVec_data_lo_lo};
  wire [15:0]       writeDataVec_data_hi_lo_lo = {writeDataVec_data_dataElement_9, writeDataVec_data_dataElement_8};
  wire [15:0]       writeDataVec_data_hi_lo_hi = {writeDataVec_data_dataElement_11, writeDataVec_data_dataElement_10};
  wire [31:0]       writeDataVec_data_hi_lo = {writeDataVec_data_hi_lo_hi, writeDataVec_data_hi_lo_lo};
  wire [15:0]       writeDataVec_data_hi_hi_lo = {writeDataVec_data_dataElement_13, writeDataVec_data_dataElement_12};
  wire [15:0]       writeDataVec_data_hi_hi_hi = {writeDataVec_data_dataElement_15, writeDataVec_data_dataElement_14};
  wire [31:0]       writeDataVec_data_hi_hi = {writeDataVec_data_hi_hi_hi, writeDataVec_data_hi_hi_lo};
  wire [63:0]       writeDataVec_data_hi = {writeDataVec_data_hi_hi, writeDataVec_data_hi_lo};
  wire [127:0]      writeDataVec_data = {writeDataVec_data_hi, writeDataVec_data_lo};
  wire [638:0]      writeDataVec_shifterData = {511'h0, writeDataVec_data} << {630'h0, executeIndexVec_0, 7'h0};
  wire [511:0]      writeDataVec_0 = writeDataVec_shifterData[511:0];
  wire [15:0]       writeDataVec_data_dataElement_16 = writeDataVec_data_dataIsRead_16 ? waiteReadData_0[15:0] : writeDataVec_data_unreadData_16[15:0];
  wire [15:0]       writeDataVec_data_dataElement_17 = writeDataVec_data_dataIsRead_17 ? waiteReadData_1[15:0] : writeDataVec_data_unreadData_17[15:0];
  wire [15:0]       writeDataVec_data_dataElement_18 = writeDataVec_data_dataIsRead_18 ? waiteReadData_2[15:0] : writeDataVec_data_unreadData_18[15:0];
  wire [15:0]       writeDataVec_data_dataElement_19 = writeDataVec_data_dataIsRead_19 ? waiteReadData_3[15:0] : writeDataVec_data_unreadData_19[15:0];
  wire [15:0]       writeDataVec_data_dataElement_20 = writeDataVec_data_dataIsRead_20 ? waiteReadData_4[15:0] : writeDataVec_data_unreadData_20[15:0];
  wire [15:0]       writeDataVec_data_dataElement_21 = writeDataVec_data_dataIsRead_21 ? waiteReadData_5[15:0] : writeDataVec_data_unreadData_21[15:0];
  wire [15:0]       writeDataVec_data_dataElement_22 = writeDataVec_data_dataIsRead_22 ? waiteReadData_6[15:0] : writeDataVec_data_unreadData_22[15:0];
  wire [15:0]       writeDataVec_data_dataElement_23 = writeDataVec_data_dataIsRead_23 ? waiteReadData_7[15:0] : writeDataVec_data_unreadData_23[15:0];
  wire [15:0]       writeDataVec_data_dataElement_24 = writeDataVec_data_dataIsRead_24 ? waiteReadData_8[15:0] : writeDataVec_data_unreadData_24[15:0];
  wire [15:0]       writeDataVec_data_dataElement_25 = writeDataVec_data_dataIsRead_25 ? waiteReadData_9[15:0] : writeDataVec_data_unreadData_25[15:0];
  wire [15:0]       writeDataVec_data_dataElement_26 = writeDataVec_data_dataIsRead_26 ? waiteReadData_10[15:0] : writeDataVec_data_unreadData_26[15:0];
  wire [15:0]       writeDataVec_data_dataElement_27 = writeDataVec_data_dataIsRead_27 ? waiteReadData_11[15:0] : writeDataVec_data_unreadData_27[15:0];
  wire [15:0]       writeDataVec_data_dataElement_28 = writeDataVec_data_dataIsRead_28 ? waiteReadData_12[15:0] : writeDataVec_data_unreadData_28[15:0];
  wire [15:0]       writeDataVec_data_dataElement_29 = writeDataVec_data_dataIsRead_29 ? waiteReadData_13[15:0] : writeDataVec_data_unreadData_29[15:0];
  wire [15:0]       writeDataVec_data_dataElement_30 = writeDataVec_data_dataIsRead_30 ? waiteReadData_14[15:0] : writeDataVec_data_unreadData_30[15:0];
  wire [15:0]       writeDataVec_data_dataElement_31 = writeDataVec_data_dataIsRead_31 ? waiteReadData_15[15:0] : writeDataVec_data_unreadData_31[15:0];
  wire [31:0]       writeDataVec_data_lo_lo_lo_1 = {writeDataVec_data_dataElement_17, writeDataVec_data_dataElement_16};
  wire [31:0]       writeDataVec_data_lo_lo_hi_1 = {writeDataVec_data_dataElement_19, writeDataVec_data_dataElement_18};
  wire [63:0]       writeDataVec_data_lo_lo_1 = {writeDataVec_data_lo_lo_hi_1, writeDataVec_data_lo_lo_lo_1};
  wire [31:0]       writeDataVec_data_lo_hi_lo_1 = {writeDataVec_data_dataElement_21, writeDataVec_data_dataElement_20};
  wire [31:0]       writeDataVec_data_lo_hi_hi_1 = {writeDataVec_data_dataElement_23, writeDataVec_data_dataElement_22};
  wire [63:0]       writeDataVec_data_lo_hi_1 = {writeDataVec_data_lo_hi_hi_1, writeDataVec_data_lo_hi_lo_1};
  wire [127:0]      writeDataVec_data_lo_1 = {writeDataVec_data_lo_hi_1, writeDataVec_data_lo_lo_1};
  wire [31:0]       writeDataVec_data_hi_lo_lo_1 = {writeDataVec_data_dataElement_25, writeDataVec_data_dataElement_24};
  wire [31:0]       writeDataVec_data_hi_lo_hi_1 = {writeDataVec_data_dataElement_27, writeDataVec_data_dataElement_26};
  wire [63:0]       writeDataVec_data_hi_lo_1 = {writeDataVec_data_hi_lo_hi_1, writeDataVec_data_hi_lo_lo_1};
  wire [31:0]       writeDataVec_data_hi_hi_lo_1 = {writeDataVec_data_dataElement_29, writeDataVec_data_dataElement_28};
  wire [31:0]       writeDataVec_data_hi_hi_hi_1 = {writeDataVec_data_dataElement_31, writeDataVec_data_dataElement_30};
  wire [63:0]       writeDataVec_data_hi_hi_1 = {writeDataVec_data_hi_hi_hi_1, writeDataVec_data_hi_hi_lo_1};
  wire [127:0]      writeDataVec_data_hi_1 = {writeDataVec_data_hi_hi_1, writeDataVec_data_hi_lo_1};
  wire [255:0]      writeDataVec_data_1 = {writeDataVec_data_hi_1, writeDataVec_data_lo_1};
  wire [766:0]      writeDataVec_shifterData_1 = {511'h0, writeDataVec_data_1} << {758'h0, executeIndexVec_1, 7'h0};
  wire [511:0]      writeDataVec_1 = writeDataVec_shifterData_1[511:0];
  wire [31:0]       writeDataVec_data_dataElement_32 = writeDataVec_data_dataIsRead_32 ? waiteReadData_0 : writeDataVec_data_unreadData_32;
  wire [31:0]       writeDataVec_data_dataElement_33 = writeDataVec_data_dataIsRead_33 ? waiteReadData_1 : writeDataVec_data_unreadData_33;
  wire [31:0]       writeDataVec_data_dataElement_34 = writeDataVec_data_dataIsRead_34 ? waiteReadData_2 : writeDataVec_data_unreadData_34;
  wire [31:0]       writeDataVec_data_dataElement_35 = writeDataVec_data_dataIsRead_35 ? waiteReadData_3 : writeDataVec_data_unreadData_35;
  wire [31:0]       writeDataVec_data_dataElement_36 = writeDataVec_data_dataIsRead_36 ? waiteReadData_4 : writeDataVec_data_unreadData_36;
  wire [31:0]       writeDataVec_data_dataElement_37 = writeDataVec_data_dataIsRead_37 ? waiteReadData_5 : writeDataVec_data_unreadData_37;
  wire [31:0]       writeDataVec_data_dataElement_38 = writeDataVec_data_dataIsRead_38 ? waiteReadData_6 : writeDataVec_data_unreadData_38;
  wire [31:0]       writeDataVec_data_dataElement_39 = writeDataVec_data_dataIsRead_39 ? waiteReadData_7 : writeDataVec_data_unreadData_39;
  wire [31:0]       writeDataVec_data_dataElement_40 = writeDataVec_data_dataIsRead_40 ? waiteReadData_8 : writeDataVec_data_unreadData_40;
  wire [31:0]       writeDataVec_data_dataElement_41 = writeDataVec_data_dataIsRead_41 ? waiteReadData_9 : writeDataVec_data_unreadData_41;
  wire [31:0]       writeDataVec_data_dataElement_42 = writeDataVec_data_dataIsRead_42 ? waiteReadData_10 : writeDataVec_data_unreadData_42;
  wire [31:0]       writeDataVec_data_dataElement_43 = writeDataVec_data_dataIsRead_43 ? waiteReadData_11 : writeDataVec_data_unreadData_43;
  wire [31:0]       writeDataVec_data_dataElement_44 = writeDataVec_data_dataIsRead_44 ? waiteReadData_12 : writeDataVec_data_unreadData_44;
  wire [31:0]       writeDataVec_data_dataElement_45 = writeDataVec_data_dataIsRead_45 ? waiteReadData_13 : writeDataVec_data_unreadData_45;
  wire [31:0]       writeDataVec_data_dataElement_46 = writeDataVec_data_dataIsRead_46 ? waiteReadData_14 : writeDataVec_data_unreadData_46;
  wire [31:0]       writeDataVec_data_dataElement_47 = writeDataVec_data_dataIsRead_47 ? waiteReadData_15 : writeDataVec_data_unreadData_47;
  wire [63:0]       writeDataVec_data_lo_lo_lo_2 = {writeDataVec_data_dataElement_33, writeDataVec_data_dataElement_32};
  wire [63:0]       writeDataVec_data_lo_lo_hi_2 = {writeDataVec_data_dataElement_35, writeDataVec_data_dataElement_34};
  wire [127:0]      writeDataVec_data_lo_lo_2 = {writeDataVec_data_lo_lo_hi_2, writeDataVec_data_lo_lo_lo_2};
  wire [63:0]       writeDataVec_data_lo_hi_lo_2 = {writeDataVec_data_dataElement_37, writeDataVec_data_dataElement_36};
  wire [63:0]       writeDataVec_data_lo_hi_hi_2 = {writeDataVec_data_dataElement_39, writeDataVec_data_dataElement_38};
  wire [127:0]      writeDataVec_data_lo_hi_2 = {writeDataVec_data_lo_hi_hi_2, writeDataVec_data_lo_hi_lo_2};
  wire [255:0]      writeDataVec_data_lo_2 = {writeDataVec_data_lo_hi_2, writeDataVec_data_lo_lo_2};
  wire [63:0]       writeDataVec_data_hi_lo_lo_2 = {writeDataVec_data_dataElement_41, writeDataVec_data_dataElement_40};
  wire [63:0]       writeDataVec_data_hi_lo_hi_2 = {writeDataVec_data_dataElement_43, writeDataVec_data_dataElement_42};
  wire [127:0]      writeDataVec_data_hi_lo_2 = {writeDataVec_data_hi_lo_hi_2, writeDataVec_data_hi_lo_lo_2};
  wire [63:0]       writeDataVec_data_hi_hi_lo_2 = {writeDataVec_data_dataElement_45, writeDataVec_data_dataElement_44};
  wire [63:0]       writeDataVec_data_hi_hi_hi_2 = {writeDataVec_data_dataElement_47, writeDataVec_data_dataElement_46};
  wire [127:0]      writeDataVec_data_hi_hi_2 = {writeDataVec_data_hi_hi_hi_2, writeDataVec_data_hi_hi_lo_2};
  wire [255:0]      writeDataVec_data_hi_2 = {writeDataVec_data_hi_hi_2, writeDataVec_data_hi_lo_2};
  wire [511:0]      writeDataVec_data_2 = {writeDataVec_data_hi_2, writeDataVec_data_lo_2};
  wire [766:0]      writeDataVec_shifterData_2 = {255'h0, writeDataVec_data_2};
  wire [511:0]      writeDataVec_2 = writeDataVec_shifterData_2[511:0];
  wire [511:0]      writeData = (sew1H[0] ? writeDataVec_0 : 512'h0) | (sew1H[1] ? writeDataVec_1 : 512'h0) | (sew1H[2] ? writeDataVec_2 : 512'h0);
  wire [1:0]        writeMaskVec_mask_lo_lo_lo = waiteReadDataPipeReg_sourceValid[1:0];
  wire [1:0]        writeMaskVec_mask_lo_lo_hi = waiteReadDataPipeReg_sourceValid[3:2];
  wire [3:0]        writeMaskVec_mask_lo_lo = {writeMaskVec_mask_lo_lo_hi, writeMaskVec_mask_lo_lo_lo};
  wire [1:0]        writeMaskVec_mask_lo_hi_lo = waiteReadDataPipeReg_sourceValid[5:4];
  wire [1:0]        writeMaskVec_mask_lo_hi_hi = waiteReadDataPipeReg_sourceValid[7:6];
  wire [3:0]        writeMaskVec_mask_lo_hi = {writeMaskVec_mask_lo_hi_hi, writeMaskVec_mask_lo_hi_lo};
  wire [7:0]        writeMaskVec_mask_lo = {writeMaskVec_mask_lo_hi, writeMaskVec_mask_lo_lo};
  wire [1:0]        writeMaskVec_mask_hi_lo_lo = waiteReadDataPipeReg_sourceValid[9:8];
  wire [1:0]        writeMaskVec_mask_hi_lo_hi = waiteReadDataPipeReg_sourceValid[11:10];
  wire [3:0]        writeMaskVec_mask_hi_lo = {writeMaskVec_mask_hi_lo_hi, writeMaskVec_mask_hi_lo_lo};
  wire [1:0]        writeMaskVec_mask_hi_hi_lo = waiteReadDataPipeReg_sourceValid[13:12];
  wire [1:0]        writeMaskVec_mask_hi_hi_hi = waiteReadDataPipeReg_sourceValid[15:14];
  wire [3:0]        writeMaskVec_mask_hi_hi = {writeMaskVec_mask_hi_hi_hi, writeMaskVec_mask_hi_hi_lo};
  wire [7:0]        writeMaskVec_mask_hi = {writeMaskVec_mask_hi_hi, writeMaskVec_mask_hi_lo};
  wire [15:0]       writeMaskVec_mask = {writeMaskVec_mask_hi, writeMaskVec_mask_lo};
  wire [78:0]       writeMaskVec_shifterMask = {63'h0, writeMaskVec_mask} << {73'h0, executeIndexVec_0, 4'h0};
  wire [63:0]       writeMaskVec_0 = writeMaskVec_shifterMask[63:0];
  wire [3:0]        writeMaskVec_mask_lo_lo_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[1]}}, {2{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [3:0]        writeMaskVec_mask_lo_lo_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[3]}}, {2{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [7:0]        writeMaskVec_mask_lo_lo_1 = {writeMaskVec_mask_lo_lo_hi_1, writeMaskVec_mask_lo_lo_lo_1};
  wire [3:0]        writeMaskVec_mask_lo_hi_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[5]}}, {2{waiteReadDataPipeReg_sourceValid[4]}}};
  wire [3:0]        writeMaskVec_mask_lo_hi_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[7]}}, {2{waiteReadDataPipeReg_sourceValid[6]}}};
  wire [7:0]        writeMaskVec_mask_lo_hi_1 = {writeMaskVec_mask_lo_hi_hi_1, writeMaskVec_mask_lo_hi_lo_1};
  wire [15:0]       writeMaskVec_mask_lo_1 = {writeMaskVec_mask_lo_hi_1, writeMaskVec_mask_lo_lo_1};
  wire [3:0]        writeMaskVec_mask_hi_lo_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[9]}}, {2{waiteReadDataPipeReg_sourceValid[8]}}};
  wire [3:0]        writeMaskVec_mask_hi_lo_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[11]}}, {2{waiteReadDataPipeReg_sourceValid[10]}}};
  wire [7:0]        writeMaskVec_mask_hi_lo_1 = {writeMaskVec_mask_hi_lo_hi_1, writeMaskVec_mask_hi_lo_lo_1};
  wire [3:0]        writeMaskVec_mask_hi_hi_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[13]}}, {2{waiteReadDataPipeReg_sourceValid[12]}}};
  wire [3:0]        writeMaskVec_mask_hi_hi_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[15]}}, {2{waiteReadDataPipeReg_sourceValid[14]}}};
  wire [7:0]        writeMaskVec_mask_hi_hi_1 = {writeMaskVec_mask_hi_hi_hi_1, writeMaskVec_mask_hi_hi_lo_1};
  wire [15:0]       writeMaskVec_mask_hi_1 = {writeMaskVec_mask_hi_hi_1, writeMaskVec_mask_hi_lo_1};
  wire [31:0]       writeMaskVec_mask_1 = {writeMaskVec_mask_hi_1, writeMaskVec_mask_lo_1};
  wire [94:0]       writeMaskVec_shifterMask_1 = {63'h0, writeMaskVec_mask_1} << {89'h0, executeIndexVec_1, 4'h0};
  wire [63:0]       writeMaskVec_1 = writeMaskVec_shifterMask_1[63:0];
  wire [7:0]        writeMaskVec_mask_lo_lo_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[1]}}, {4{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [7:0]        writeMaskVec_mask_lo_lo_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[3]}}, {4{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [15:0]       writeMaskVec_mask_lo_lo_2 = {writeMaskVec_mask_lo_lo_hi_2, writeMaskVec_mask_lo_lo_lo_2};
  wire [7:0]        writeMaskVec_mask_lo_hi_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[5]}}, {4{waiteReadDataPipeReg_sourceValid[4]}}};
  wire [7:0]        writeMaskVec_mask_lo_hi_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[7]}}, {4{waiteReadDataPipeReg_sourceValid[6]}}};
  wire [15:0]       writeMaskVec_mask_lo_hi_2 = {writeMaskVec_mask_lo_hi_hi_2, writeMaskVec_mask_lo_hi_lo_2};
  wire [31:0]       writeMaskVec_mask_lo_2 = {writeMaskVec_mask_lo_hi_2, writeMaskVec_mask_lo_lo_2};
  wire [7:0]        writeMaskVec_mask_hi_lo_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[9]}}, {4{waiteReadDataPipeReg_sourceValid[8]}}};
  wire [7:0]        writeMaskVec_mask_hi_lo_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[11]}}, {4{waiteReadDataPipeReg_sourceValid[10]}}};
  wire [15:0]       writeMaskVec_mask_hi_lo_2 = {writeMaskVec_mask_hi_lo_hi_2, writeMaskVec_mask_hi_lo_lo_2};
  wire [7:0]        writeMaskVec_mask_hi_hi_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[13]}}, {4{waiteReadDataPipeReg_sourceValid[12]}}};
  wire [7:0]        writeMaskVec_mask_hi_hi_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[15]}}, {4{waiteReadDataPipeReg_sourceValid[14]}}};
  wire [15:0]       writeMaskVec_mask_hi_hi_2 = {writeMaskVec_mask_hi_hi_hi_2, writeMaskVec_mask_hi_hi_lo_2};
  wire [31:0]       writeMaskVec_mask_hi_2 = {writeMaskVec_mask_hi_hi_2, writeMaskVec_mask_hi_lo_2};
  wire [63:0]       writeMaskVec_mask_2 = {writeMaskVec_mask_hi_2, writeMaskVec_mask_lo_2};
  wire [94:0]       writeMaskVec_shifterMask_2 = {31'h0, writeMaskVec_mask_2};
  wire [63:0]       writeMaskVec_2 = writeMaskVec_shifterMask_2[63:0];
  wire [63:0]       writeMask = (sew1H[0] ? writeMaskVec_0 : 64'h0) | (sew1H[1] ? writeMaskVec_1 : 64'h0) | (sew1H[2] ? writeMaskVec_2 : 64'h0);
  wire [9:0]        _writeRequest_res_writeData_groupCounter_T_30 = {3'h0, waiteReadDataPipeReg_executeGroup} << instReg_sew;
  wire [4:0]        writeRequest_0_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_1_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_2_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_3_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_4_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_5_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_6_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_7_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_8_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_9_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_10_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_11_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_12_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_13_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_14_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [4:0]        writeRequest_15_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_30[6:2];
  wire [31:0]       writeRequest_0_writeData_data = writeData[31:0];
  wire [31:0]       writeRequest_1_writeData_data = writeData[63:32];
  wire [31:0]       writeRequest_2_writeData_data = writeData[95:64];
  wire [31:0]       writeRequest_3_writeData_data = writeData[127:96];
  wire [31:0]       writeRequest_4_writeData_data = writeData[159:128];
  wire [31:0]       writeRequest_5_writeData_data = writeData[191:160];
  wire [31:0]       writeRequest_6_writeData_data = writeData[223:192];
  wire [31:0]       writeRequest_7_writeData_data = writeData[255:224];
  wire [31:0]       writeRequest_8_writeData_data = writeData[287:256];
  wire [31:0]       writeRequest_9_writeData_data = writeData[319:288];
  wire [31:0]       writeRequest_10_writeData_data = writeData[351:320];
  wire [31:0]       writeRequest_11_writeData_data = writeData[383:352];
  wire [31:0]       writeRequest_12_writeData_data = writeData[415:384];
  wire [31:0]       writeRequest_13_writeData_data = writeData[447:416];
  wire [31:0]       writeRequest_14_writeData_data = writeData[479:448];
  wire [31:0]       writeRequest_15_writeData_data = writeData[511:480];
  wire [3:0]        writeRequest_0_writeData_mask = writeMask[3:0];
  wire [3:0]        writeRequest_1_writeData_mask = writeMask[7:4];
  wire [3:0]        writeRequest_2_writeData_mask = writeMask[11:8];
  wire [3:0]        writeRequest_3_writeData_mask = writeMask[15:12];
  wire [3:0]        writeRequest_4_writeData_mask = writeMask[19:16];
  wire [3:0]        writeRequest_5_writeData_mask = writeMask[23:20];
  wire [3:0]        writeRequest_6_writeData_mask = writeMask[27:24];
  wire [3:0]        writeRequest_7_writeData_mask = writeMask[31:28];
  wire [3:0]        writeRequest_8_writeData_mask = writeMask[35:32];
  wire [3:0]        writeRequest_9_writeData_mask = writeMask[39:36];
  wire [3:0]        writeRequest_10_writeData_mask = writeMask[43:40];
  wire [3:0]        writeRequest_11_writeData_mask = writeMask[47:44];
  wire [3:0]        writeRequest_12_writeData_mask = writeMask[51:48];
  wire [3:0]        writeRequest_13_writeData_mask = writeMask[55:52];
  wire [3:0]        writeRequest_14_writeData_mask = writeMask[59:56];
  wire [3:0]        writeRequest_15_writeData_mask = writeMask[63:60];
  wire [1:0]        WillWriteLane_lo_lo_lo = {|writeRequest_1_writeData_mask, |writeRequest_0_writeData_mask};
  wire [1:0]        WillWriteLane_lo_lo_hi = {|writeRequest_3_writeData_mask, |writeRequest_2_writeData_mask};
  wire [3:0]        WillWriteLane_lo_lo = {WillWriteLane_lo_lo_hi, WillWriteLane_lo_lo_lo};
  wire [1:0]        WillWriteLane_lo_hi_lo = {|writeRequest_5_writeData_mask, |writeRequest_4_writeData_mask};
  wire [1:0]        WillWriteLane_lo_hi_hi = {|writeRequest_7_writeData_mask, |writeRequest_6_writeData_mask};
  wire [3:0]        WillWriteLane_lo_hi = {WillWriteLane_lo_hi_hi, WillWriteLane_lo_hi_lo};
  wire [7:0]        WillWriteLane_lo = {WillWriteLane_lo_hi, WillWriteLane_lo_lo};
  wire [1:0]        WillWriteLane_hi_lo_lo = {|writeRequest_9_writeData_mask, |writeRequest_8_writeData_mask};
  wire [1:0]        WillWriteLane_hi_lo_hi = {|writeRequest_11_writeData_mask, |writeRequest_10_writeData_mask};
  wire [3:0]        WillWriteLane_hi_lo = {WillWriteLane_hi_lo_hi, WillWriteLane_hi_lo_lo};
  wire [1:0]        WillWriteLane_hi_hi_lo = {|writeRequest_13_writeData_mask, |writeRequest_12_writeData_mask};
  wire [1:0]        WillWriteLane_hi_hi_hi = {|writeRequest_15_writeData_mask, |writeRequest_14_writeData_mask};
  wire [3:0]        WillWriteLane_hi_hi = {WillWriteLane_hi_hi_hi, WillWriteLane_hi_hi_lo};
  wire [7:0]        WillWriteLane_hi = {WillWriteLane_hi_hi, WillWriteLane_hi_lo};
  wire [15:0]       WillWriteLane = {WillWriteLane_hi, WillWriteLane_lo};
  wire              waiteStageDeqValid = waiteReadStageValid & (waiteReadSate == waiteReadDataPipeReg_needRead | waiteReadDataPipeReg_needRead == 16'h0);
  wire              waiteStageDeqReady;
  wire              waiteStageDeqFire = waiteStageDeqValid & waiteStageDeqReady;
  assign waiteStageEnqReady = ~waiteReadStageValid | waiteStageDeqFire;
  assign readWaitQueue_deq_ready = waiteStageEnqReady;
  wire              waiteStageEnqFire = readWaitQueue_deq_valid & waiteStageEnqReady;
  wire              isWaiteForThisData = waiteReadDataPipeReg_needRead[0] & ~(waiteReadSate[0]) & waiteReadStageValid;
  assign readData_readDataQueue_deq_ready = isWaiteForThisData | unitType[2] | compress | gatherWaiteRead | mvRd;
  assign isWaiteForThisData_1 = waiteReadDataPipeReg_needRead[1] & ~(waiteReadSate[1]) & waiteReadStageValid;
  assign readData_readDataQueue_1_deq_ready = isWaiteForThisData_1;
  assign isWaiteForThisData_2 = waiteReadDataPipeReg_needRead[2] & ~(waiteReadSate[2]) & waiteReadStageValid;
  assign readData_readDataQueue_2_deq_ready = isWaiteForThisData_2;
  assign isWaiteForThisData_3 = waiteReadDataPipeReg_needRead[3] & ~(waiteReadSate[3]) & waiteReadStageValid;
  assign readData_readDataQueue_3_deq_ready = isWaiteForThisData_3;
  assign isWaiteForThisData_4 = waiteReadDataPipeReg_needRead[4] & ~(waiteReadSate[4]) & waiteReadStageValid;
  assign readData_readDataQueue_4_deq_ready = isWaiteForThisData_4;
  assign isWaiteForThisData_5 = waiteReadDataPipeReg_needRead[5] & ~(waiteReadSate[5]) & waiteReadStageValid;
  assign readData_readDataQueue_5_deq_ready = isWaiteForThisData_5;
  assign isWaiteForThisData_6 = waiteReadDataPipeReg_needRead[6] & ~(waiteReadSate[6]) & waiteReadStageValid;
  assign readData_readDataQueue_6_deq_ready = isWaiteForThisData_6;
  assign isWaiteForThisData_7 = waiteReadDataPipeReg_needRead[7] & ~(waiteReadSate[7]) & waiteReadStageValid;
  assign readData_readDataQueue_7_deq_ready = isWaiteForThisData_7;
  assign isWaiteForThisData_8 = waiteReadDataPipeReg_needRead[8] & ~(waiteReadSate[8]) & waiteReadStageValid;
  assign readData_readDataQueue_8_deq_ready = isWaiteForThisData_8;
  assign isWaiteForThisData_9 = waiteReadDataPipeReg_needRead[9] & ~(waiteReadSate[9]) & waiteReadStageValid;
  assign readData_readDataQueue_9_deq_ready = isWaiteForThisData_9;
  assign isWaiteForThisData_10 = waiteReadDataPipeReg_needRead[10] & ~(waiteReadSate[10]) & waiteReadStageValid;
  assign readData_readDataQueue_10_deq_ready = isWaiteForThisData_10;
  assign isWaiteForThisData_11 = waiteReadDataPipeReg_needRead[11] & ~(waiteReadSate[11]) & waiteReadStageValid;
  assign readData_readDataQueue_11_deq_ready = isWaiteForThisData_11;
  assign isWaiteForThisData_12 = waiteReadDataPipeReg_needRead[12] & ~(waiteReadSate[12]) & waiteReadStageValid;
  assign readData_readDataQueue_12_deq_ready = isWaiteForThisData_12;
  assign isWaiteForThisData_13 = waiteReadDataPipeReg_needRead[13] & ~(waiteReadSate[13]) & waiteReadStageValid;
  assign readData_readDataQueue_13_deq_ready = isWaiteForThisData_13;
  assign isWaiteForThisData_14 = waiteReadDataPipeReg_needRead[14] & ~(waiteReadSate[14]) & waiteReadStageValid;
  assign readData_readDataQueue_14_deq_ready = isWaiteForThisData_14;
  assign isWaiteForThisData_15 = waiteReadDataPipeReg_needRead[15] & ~(waiteReadSate[15]) & waiteReadStageValid;
  assign readData_readDataQueue_15_deq_ready = isWaiteForThisData_15;
  wire [1:0]        readResultValid_lo_lo_lo = {readTokenRelease_1, readTokenRelease_0};
  wire [1:0]        readResultValid_lo_lo_hi = {readTokenRelease_3, readTokenRelease_2};
  wire [3:0]        readResultValid_lo_lo = {readResultValid_lo_lo_hi, readResultValid_lo_lo_lo};
  wire [1:0]        readResultValid_lo_hi_lo = {readTokenRelease_5, readTokenRelease_4};
  wire [1:0]        readResultValid_lo_hi_hi = {readTokenRelease_7, readTokenRelease_6};
  wire [3:0]        readResultValid_lo_hi = {readResultValid_lo_hi_hi, readResultValid_lo_hi_lo};
  wire [7:0]        readResultValid_lo = {readResultValid_lo_hi, readResultValid_lo_lo};
  wire [1:0]        readResultValid_hi_lo_lo = {readTokenRelease_9, readTokenRelease_8};
  wire [1:0]        readResultValid_hi_lo_hi = {readTokenRelease_11, readTokenRelease_10};
  wire [3:0]        readResultValid_hi_lo = {readResultValid_hi_lo_hi, readResultValid_hi_lo_lo};
  wire [1:0]        readResultValid_hi_hi_lo = {readTokenRelease_13, readTokenRelease_12};
  wire [1:0]        readResultValid_hi_hi_hi = {readTokenRelease_15, readTokenRelease_14};
  wire [3:0]        readResultValid_hi_hi = {readResultValid_hi_hi_hi, readResultValid_hi_hi_lo};
  wire [7:0]        readResultValid_hi = {readResultValid_hi_hi, readResultValid_hi_lo};
  wire [15:0]       readResultValid = {readResultValid_hi, readResultValid_lo};
  wire              executeEnqValid = otherTypeRequestDeq & ~readType;
  wire [63:0]       source2_lo_lo_lo = {exeReqReg_1_bits_source2, exeReqReg_0_bits_source2};
  wire [63:0]       source2_lo_lo_hi = {exeReqReg_3_bits_source2, exeReqReg_2_bits_source2};
  wire [127:0]      source2_lo_lo = {source2_lo_lo_hi, source2_lo_lo_lo};
  wire [63:0]       source2_lo_hi_lo = {exeReqReg_5_bits_source2, exeReqReg_4_bits_source2};
  wire [63:0]       source2_lo_hi_hi = {exeReqReg_7_bits_source2, exeReqReg_6_bits_source2};
  wire [127:0]      source2_lo_hi = {source2_lo_hi_hi, source2_lo_hi_lo};
  wire [255:0]      source2_lo = {source2_lo_hi, source2_lo_lo};
  wire [63:0]       source2_hi_lo_lo = {exeReqReg_9_bits_source2, exeReqReg_8_bits_source2};
  wire [63:0]       source2_hi_lo_hi = {exeReqReg_11_bits_source2, exeReqReg_10_bits_source2};
  wire [127:0]      source2_hi_lo = {source2_hi_lo_hi, source2_hi_lo_lo};
  wire [63:0]       source2_hi_hi_lo = {exeReqReg_13_bits_source2, exeReqReg_12_bits_source2};
  wire [63:0]       source2_hi_hi_hi = {exeReqReg_15_bits_source2, exeReqReg_14_bits_source2};
  wire [127:0]      source2_hi_hi = {source2_hi_hi_hi, source2_hi_hi_lo};
  wire [255:0]      source2_hi = {source2_hi_hi, source2_hi_lo};
  wire [511:0]      source2 = {source2_hi, source2_lo};
  wire [127:0]      source1_lo_lo = {source1_lo_lo_hi, source1_lo_lo_lo};
  wire [127:0]      source1_lo_hi = {source1_lo_hi_hi, source1_lo_hi_lo};
  wire [255:0]      source1_lo = {source1_lo_hi, source1_lo_lo};
  wire [127:0]      source1_hi_lo = {source1_hi_lo_hi, source1_hi_lo_lo};
  wire [127:0]      source1_hi_hi = {source1_hi_hi_hi, source1_hi_hi_lo};
  wire [255:0]      source1_hi = {source1_hi_hi, source1_hi_lo};
  wire [511:0]      source1 = {source1_hi, source1_lo};
  wire              vs1Split_2_2 = vs1Split_vs1SetIndex;
  wire [31:0]       _compressSource1_T_6 = sew1H[0] | sew1H[1] ? readVS1Reg_data : 32'h0;
  wire [31:0]       compressSource1 = {_compressSource1_T_6[31:16], _compressSource1_T_6[15:0] | (sew1H[2] ? (vs1Split_vs1SetIndex ? readVS1Reg_data[31:16] : readVS1Reg_data[15:0]) : 16'h0)};
  wire [31:0]       source1Select = mv ? readVS1Reg_data : compressSource1;
  wire              source1Change = sew1H[0] | sew1H[1] | sew1H[2] & vs1Split_2_2;
  assign viotaCounterAdd = executeEnqValid & unitType[1];
  wire [1:0]        view__in_bits_ffoInput_lo_lo_lo = {exeReqReg_1_bits_ffo, exeReqReg_0_bits_ffo};
  wire [1:0]        view__in_bits_ffoInput_lo_lo_hi = {exeReqReg_3_bits_ffo, exeReqReg_2_bits_ffo};
  wire [3:0]        view__in_bits_ffoInput_lo_lo = {view__in_bits_ffoInput_lo_lo_hi, view__in_bits_ffoInput_lo_lo_lo};
  wire [1:0]        view__in_bits_ffoInput_lo_hi_lo = {exeReqReg_5_bits_ffo, exeReqReg_4_bits_ffo};
  wire [1:0]        view__in_bits_ffoInput_lo_hi_hi = {exeReqReg_7_bits_ffo, exeReqReg_6_bits_ffo};
  wire [3:0]        view__in_bits_ffoInput_lo_hi = {view__in_bits_ffoInput_lo_hi_hi, view__in_bits_ffoInput_lo_hi_lo};
  wire [7:0]        view__in_bits_ffoInput_lo = {view__in_bits_ffoInput_lo_hi, view__in_bits_ffoInput_lo_lo};
  wire [1:0]        view__in_bits_ffoInput_hi_lo_lo = {exeReqReg_9_bits_ffo, exeReqReg_8_bits_ffo};
  wire [1:0]        view__in_bits_ffoInput_hi_lo_hi = {exeReqReg_11_bits_ffo, exeReqReg_10_bits_ffo};
  wire [3:0]        view__in_bits_ffoInput_hi_lo = {view__in_bits_ffoInput_hi_lo_hi, view__in_bits_ffoInput_hi_lo_lo};
  wire [1:0]        view__in_bits_ffoInput_hi_hi_lo = {exeReqReg_13_bits_ffo, exeReqReg_12_bits_ffo};
  wire [1:0]        view__in_bits_ffoInput_hi_hi_hi = {exeReqReg_15_bits_ffo, exeReqReg_14_bits_ffo};
  wire [3:0]        view__in_bits_ffoInput_hi_hi = {view__in_bits_ffoInput_hi_hi_hi, view__in_bits_ffoInput_hi_hi_lo};
  wire [7:0]        view__in_bits_ffoInput_hi = {view__in_bits_ffoInput_hi_hi, view__in_bits_ffoInput_hi_lo};
  wire [3:0]        view__in_bits_validInput_lo_lo = {view__in_bits_validInput_lo_lo_hi, view__in_bits_validInput_lo_lo_lo};
  wire [3:0]        view__in_bits_validInput_lo_hi = {view__in_bits_validInput_lo_hi_hi, view__in_bits_validInput_lo_hi_lo};
  wire [7:0]        view__in_bits_validInput_lo = {view__in_bits_validInput_lo_hi, view__in_bits_validInput_lo_lo};
  wire [3:0]        view__in_bits_validInput_hi_lo = {view__in_bits_validInput_hi_lo_hi, view__in_bits_validInput_hi_lo_lo};
  wire [3:0]        view__in_bits_validInput_hi_hi = {view__in_bits_validInput_hi_hi_hi, view__in_bits_validInput_hi_hi_lo};
  wire [7:0]        view__in_bits_validInput_hi = {view__in_bits_validInput_hi_hi, view__in_bits_validInput_hi_lo};
  wire              reduceUnit_in_valid = executeEnqValid & unitType[2];
  wire [3:0]        view__in_bits_sourceValid_lo_lo = {view__in_bits_sourceValid_lo_lo_hi, view__in_bits_sourceValid_lo_lo_lo};
  wire [3:0]        view__in_bits_sourceValid_lo_hi = {view__in_bits_sourceValid_lo_hi_hi, view__in_bits_sourceValid_lo_hi_lo};
  wire [7:0]        view__in_bits_sourceValid_lo = {view__in_bits_sourceValid_lo_hi, view__in_bits_sourceValid_lo_lo};
  wire [3:0]        view__in_bits_sourceValid_hi_lo = {view__in_bits_sourceValid_hi_lo_hi, view__in_bits_sourceValid_hi_lo_lo};
  wire [3:0]        view__in_bits_sourceValid_hi_hi = {view__in_bits_sourceValid_hi_hi_hi, view__in_bits_sourceValid_hi_hi_lo};
  wire [7:0]        view__in_bits_sourceValid_hi = {view__in_bits_sourceValid_hi_hi, view__in_bits_sourceValid_hi_lo};
  wire              _view__firstGroup_T_1 = _reduceUnit_in_ready & reduceUnit_in_valid;
  wire [1:0]        view__in_bits_fpSourceValid_lo_lo_lo = {exeReqReg_1_bits_fpReduceValid, exeReqReg_0_bits_fpReduceValid};
  wire [1:0]        view__in_bits_fpSourceValid_lo_lo_hi = {exeReqReg_3_bits_fpReduceValid, exeReqReg_2_bits_fpReduceValid};
  wire [3:0]        view__in_bits_fpSourceValid_lo_lo = {view__in_bits_fpSourceValid_lo_lo_hi, view__in_bits_fpSourceValid_lo_lo_lo};
  wire [1:0]        view__in_bits_fpSourceValid_lo_hi_lo = {exeReqReg_5_bits_fpReduceValid, exeReqReg_4_bits_fpReduceValid};
  wire [1:0]        view__in_bits_fpSourceValid_lo_hi_hi = {exeReqReg_7_bits_fpReduceValid, exeReqReg_6_bits_fpReduceValid};
  wire [3:0]        view__in_bits_fpSourceValid_lo_hi = {view__in_bits_fpSourceValid_lo_hi_hi, view__in_bits_fpSourceValid_lo_hi_lo};
  wire [7:0]        view__in_bits_fpSourceValid_lo = {view__in_bits_fpSourceValid_lo_hi, view__in_bits_fpSourceValid_lo_lo};
  wire [1:0]        view__in_bits_fpSourceValid_hi_lo_lo = {exeReqReg_9_bits_fpReduceValid, exeReqReg_8_bits_fpReduceValid};
  wire [1:0]        view__in_bits_fpSourceValid_hi_lo_hi = {exeReqReg_11_bits_fpReduceValid, exeReqReg_10_bits_fpReduceValid};
  wire [3:0]        view__in_bits_fpSourceValid_hi_lo = {view__in_bits_fpSourceValid_hi_lo_hi, view__in_bits_fpSourceValid_hi_lo_lo};
  wire [1:0]        view__in_bits_fpSourceValid_hi_hi_lo = {exeReqReg_13_bits_fpReduceValid, exeReqReg_12_bits_fpReduceValid};
  wire [1:0]        view__in_bits_fpSourceValid_hi_hi_hi = {exeReqReg_15_bits_fpReduceValid, exeReqReg_14_bits_fpReduceValid};
  wire [3:0]        view__in_bits_fpSourceValid_hi_hi = {view__in_bits_fpSourceValid_hi_hi_hi, view__in_bits_fpSourceValid_hi_hi_lo};
  wire [7:0]        view__in_bits_fpSourceValid_hi = {view__in_bits_fpSourceValid_hi_hi, view__in_bits_fpSourceValid_hi_lo};
  wire [6:0]        extendGroupCount = extendType ? (subType[2] ? _extendGroupCount_T_1 : {1'h0, requestCounter, executeIndex[1]}) : {2'h0, requestCounter};
  wire [511:0]      _executeResult_T_4 = unitType[1] ? compressUnitResultQueue_deq_bits_data : 512'h0;
  wire [511:0]      executeResult = {_executeResult_T_4[511:32], _executeResult_T_4[31:0] | (unitType[2] ? _reduceUnit_out_bits_data : 32'h0)} | (unitType[3] ? _extendUnit_out : 512'h0);
  assign executeReady = readType | unitType[1] | unitType[2] & _reduceUnit_in_ready & readVS1Reg_dataValid | unitType[3] & executeEnqValid;
  wire [3:0]        compressUnitResultQueue_deq_ready_lo_lo = {compressUnitResultQueue_deq_ready_lo_lo_hi, compressUnitResultQueue_deq_ready_lo_lo_lo};
  wire [3:0]        compressUnitResultQueue_deq_ready_lo_hi = {compressUnitResultQueue_deq_ready_lo_hi_hi, compressUnitResultQueue_deq_ready_lo_hi_lo};
  wire [7:0]        compressUnitResultQueue_deq_ready_lo = {compressUnitResultQueue_deq_ready_lo_hi, compressUnitResultQueue_deq_ready_lo_lo};
  wire [3:0]        compressUnitResultQueue_deq_ready_hi_lo = {compressUnitResultQueue_deq_ready_hi_lo_hi, compressUnitResultQueue_deq_ready_hi_lo_lo};
  wire [3:0]        compressUnitResultQueue_deq_ready_hi_hi = {compressUnitResultQueue_deq_ready_hi_hi_hi, compressUnitResultQueue_deq_ready_hi_hi_lo};
  wire [7:0]        compressUnitResultQueue_deq_ready_hi = {compressUnitResultQueue_deq_ready_hi_hi, compressUnitResultQueue_deq_ready_hi_lo};
  assign compressUnitResultQueue_deq_ready = &{compressUnitResultQueue_deq_ready_hi, compressUnitResultQueue_deq_ready_lo};
  wire              compressDeq = compressUnitResultQueue_deq_ready & compressUnitResultQueue_deq_valid;
  wire              executeValid = unitType[1] & compressDeq | unitType[3] & executeEnqValid;
  assign executeGroupCounter = (unitType[1] | unitType[2] ? requestCounter : 5'h0) | (unitType[3] ? extendGroupCount[4:0] : 5'h0);
  wire [6:0]        executeDeqGroupCounter = {2'h0, (unitType[1] ? compressUnitResultQueue_deq_bits_groupCounter : 5'h0) | (unitType[2] ? requestCounter : 5'h0)} | (unitType[3] ? extendGroupCount : 7'h0);
  wire [63:0]       executeWriteByteMask = compress | ffo | mvVd ? compressUnitResultQueue_deq_bits_mask : executeByteMask;
  wire              maskFilter = |{~maskDestinationType, currentMaskGroupForDestination[31:0]};
  wire              maskFilter_1 = |{~maskDestinationType, currentMaskGroupForDestination[63:32]};
  wire              maskFilter_2 = |{~maskDestinationType, currentMaskGroupForDestination[95:64]};
  wire              maskFilter_3 = |{~maskDestinationType, currentMaskGroupForDestination[127:96]};
  wire              maskFilter_4 = |{~maskDestinationType, currentMaskGroupForDestination[159:128]};
  wire              maskFilter_5 = |{~maskDestinationType, currentMaskGroupForDestination[191:160]};
  wire              maskFilter_6 = |{~maskDestinationType, currentMaskGroupForDestination[223:192]};
  wire              maskFilter_7 = |{~maskDestinationType, currentMaskGroupForDestination[255:224]};
  wire              maskFilter_8 = |{~maskDestinationType, currentMaskGroupForDestination[287:256]};
  wire              maskFilter_9 = |{~maskDestinationType, currentMaskGroupForDestination[319:288]};
  wire              maskFilter_10 = |{~maskDestinationType, currentMaskGroupForDestination[351:320]};
  wire              maskFilter_11 = |{~maskDestinationType, currentMaskGroupForDestination[383:352]};
  wire              maskFilter_12 = |{~maskDestinationType, currentMaskGroupForDestination[415:384]};
  wire              maskFilter_13 = |{~maskDestinationType, currentMaskGroupForDestination[447:416]};
  wire              maskFilter_14 = |{~maskDestinationType, currentMaskGroupForDestination[479:448]};
  wire              maskFilter_15 = |{~maskDestinationType, currentMaskGroupForDestination[511:480]};
  assign writeQueue_0_deq_valid = ~_writeQueue_fifo_empty;
  wire              exeResp_0_valid_0 = writeQueue_0_deq_valid;
  wire              writeQueue_dataOut_ffoByOther;
  wire [31:0]       writeQueue_dataOut_writeData_data;
  wire [31:0]       exeResp_0_bits_data_0 = writeQueue_0_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_writeData_mask;
  wire [3:0]        exeResp_0_bits_mask_0 = writeQueue_0_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_writeData_vd;
  wire [2:0]        writeQueue_dataOut_index;
  wire [4:0]        writeQueue_0_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_0_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo = {writeQueue_0_enq_bits_writeData_groupCounter, writeQueue_0_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_0_enq_bits_writeData_data;
  wire [3:0]        writeQueue_0_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi = {writeQueue_0_enq_bits_writeData_data, writeQueue_0_enq_bits_writeData_mask};
  wire              writeQueue_0_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_1 = {writeQueue_0_enq_bits_ffoByOther, writeQueue_dataIn_hi, writeQueue_dataIn_lo};
  wire [49:0]       writeQueue_dataIn = {writeQueue_dataIn_hi_1, writeQueue_0_enq_bits_index};
  assign writeQueue_dataOut_index = _writeQueue_fifo_data_out[2:0];
  assign writeQueue_dataOut_writeData_vd = _writeQueue_fifo_data_out[7:3];
  assign writeQueue_dataOut_writeData_groupCounter = _writeQueue_fifo_data_out[12:8];
  assign writeQueue_dataOut_writeData_mask = _writeQueue_fifo_data_out[16:13];
  assign writeQueue_dataOut_writeData_data = _writeQueue_fifo_data_out[48:17];
  assign writeQueue_dataOut_ffoByOther = _writeQueue_fifo_data_out[49];
  wire              writeQueue_0_deq_bits_ffoByOther = writeQueue_dataOut_ffoByOther;
  assign writeQueue_0_deq_bits_writeData_data = writeQueue_dataOut_writeData_data;
  assign writeQueue_0_deq_bits_writeData_mask = writeQueue_dataOut_writeData_mask;
  wire [4:0]        writeQueue_0_deq_bits_writeData_groupCounter = writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]        writeQueue_0_deq_bits_writeData_vd = writeQueue_dataOut_writeData_vd;
  wire [2:0]        writeQueue_0_deq_bits_index = writeQueue_dataOut_index;
  wire              writeQueue_0_enq_ready = ~_writeQueue_fifo_full;
  wire              writeQueue_0_enq_valid;
  assign writeQueue_1_deq_valid = ~_writeQueue_fifo_1_empty;
  wire              exeResp_1_valid_0 = writeQueue_1_deq_valid;
  wire              writeQueue_dataOut_1_ffoByOther;
  wire [31:0]       writeQueue_dataOut_1_writeData_data;
  wire [31:0]       exeResp_1_bits_data_0 = writeQueue_1_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_1_writeData_mask;
  wire [3:0]        exeResp_1_bits_mask_0 = writeQueue_1_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_1_writeData_vd;
  wire [2:0]        writeQueue_dataOut_1_index;
  wire [4:0]        writeQueue_1_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_1_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_1 = {writeQueue_1_enq_bits_writeData_groupCounter, writeQueue_1_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_1_enq_bits_writeData_data;
  wire [3:0]        writeQueue_1_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_2 = {writeQueue_1_enq_bits_writeData_data, writeQueue_1_enq_bits_writeData_mask};
  wire              writeQueue_1_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_3 = {writeQueue_1_enq_bits_ffoByOther, writeQueue_dataIn_hi_2, writeQueue_dataIn_lo_1};
  wire [49:0]       writeQueue_dataIn_1 = {writeQueue_dataIn_hi_3, writeQueue_1_enq_bits_index};
  assign writeQueue_dataOut_1_index = _writeQueue_fifo_1_data_out[2:0];
  assign writeQueue_dataOut_1_writeData_vd = _writeQueue_fifo_1_data_out[7:3];
  assign writeQueue_dataOut_1_writeData_groupCounter = _writeQueue_fifo_1_data_out[12:8];
  assign writeQueue_dataOut_1_writeData_mask = _writeQueue_fifo_1_data_out[16:13];
  assign writeQueue_dataOut_1_writeData_data = _writeQueue_fifo_1_data_out[48:17];
  assign writeQueue_dataOut_1_ffoByOther = _writeQueue_fifo_1_data_out[49];
  wire              writeQueue_1_deq_bits_ffoByOther = writeQueue_dataOut_1_ffoByOther;
  assign writeQueue_1_deq_bits_writeData_data = writeQueue_dataOut_1_writeData_data;
  assign writeQueue_1_deq_bits_writeData_mask = writeQueue_dataOut_1_writeData_mask;
  wire [4:0]        writeQueue_1_deq_bits_writeData_groupCounter = writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]        writeQueue_1_deq_bits_writeData_vd = writeQueue_dataOut_1_writeData_vd;
  wire [2:0]        writeQueue_1_deq_bits_index = writeQueue_dataOut_1_index;
  wire              writeQueue_1_enq_ready = ~_writeQueue_fifo_1_full;
  wire              writeQueue_1_enq_valid;
  assign writeQueue_2_deq_valid = ~_writeQueue_fifo_2_empty;
  wire              exeResp_2_valid_0 = writeQueue_2_deq_valid;
  wire              writeQueue_dataOut_2_ffoByOther;
  wire [31:0]       writeQueue_dataOut_2_writeData_data;
  wire [31:0]       exeResp_2_bits_data_0 = writeQueue_2_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_2_writeData_mask;
  wire [3:0]        exeResp_2_bits_mask_0 = writeQueue_2_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_2_writeData_vd;
  wire [2:0]        writeQueue_dataOut_2_index;
  wire [4:0]        writeQueue_2_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_2_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_2 = {writeQueue_2_enq_bits_writeData_groupCounter, writeQueue_2_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_2_enq_bits_writeData_data;
  wire [3:0]        writeQueue_2_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_4 = {writeQueue_2_enq_bits_writeData_data, writeQueue_2_enq_bits_writeData_mask};
  wire              writeQueue_2_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_5 = {writeQueue_2_enq_bits_ffoByOther, writeQueue_dataIn_hi_4, writeQueue_dataIn_lo_2};
  wire [49:0]       writeQueue_dataIn_2 = {writeQueue_dataIn_hi_5, writeQueue_2_enq_bits_index};
  assign writeQueue_dataOut_2_index = _writeQueue_fifo_2_data_out[2:0];
  assign writeQueue_dataOut_2_writeData_vd = _writeQueue_fifo_2_data_out[7:3];
  assign writeQueue_dataOut_2_writeData_groupCounter = _writeQueue_fifo_2_data_out[12:8];
  assign writeQueue_dataOut_2_writeData_mask = _writeQueue_fifo_2_data_out[16:13];
  assign writeQueue_dataOut_2_writeData_data = _writeQueue_fifo_2_data_out[48:17];
  assign writeQueue_dataOut_2_ffoByOther = _writeQueue_fifo_2_data_out[49];
  wire              writeQueue_2_deq_bits_ffoByOther = writeQueue_dataOut_2_ffoByOther;
  assign writeQueue_2_deq_bits_writeData_data = writeQueue_dataOut_2_writeData_data;
  assign writeQueue_2_deq_bits_writeData_mask = writeQueue_dataOut_2_writeData_mask;
  wire [4:0]        writeQueue_2_deq_bits_writeData_groupCounter = writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]        writeQueue_2_deq_bits_writeData_vd = writeQueue_dataOut_2_writeData_vd;
  wire [2:0]        writeQueue_2_deq_bits_index = writeQueue_dataOut_2_index;
  wire              writeQueue_2_enq_ready = ~_writeQueue_fifo_2_full;
  wire              writeQueue_2_enq_valid;
  assign writeQueue_3_deq_valid = ~_writeQueue_fifo_3_empty;
  wire              exeResp_3_valid_0 = writeQueue_3_deq_valid;
  wire              writeQueue_dataOut_3_ffoByOther;
  wire [31:0]       writeQueue_dataOut_3_writeData_data;
  wire [31:0]       exeResp_3_bits_data_0 = writeQueue_3_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_3_writeData_mask;
  wire [3:0]        exeResp_3_bits_mask_0 = writeQueue_3_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_3_writeData_vd;
  wire [2:0]        writeQueue_dataOut_3_index;
  wire [4:0]        writeQueue_3_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_3_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_3 = {writeQueue_3_enq_bits_writeData_groupCounter, writeQueue_3_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_3_enq_bits_writeData_data;
  wire [3:0]        writeQueue_3_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_6 = {writeQueue_3_enq_bits_writeData_data, writeQueue_3_enq_bits_writeData_mask};
  wire              writeQueue_3_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_7 = {writeQueue_3_enq_bits_ffoByOther, writeQueue_dataIn_hi_6, writeQueue_dataIn_lo_3};
  wire [49:0]       writeQueue_dataIn_3 = {writeQueue_dataIn_hi_7, writeQueue_3_enq_bits_index};
  assign writeQueue_dataOut_3_index = _writeQueue_fifo_3_data_out[2:0];
  assign writeQueue_dataOut_3_writeData_vd = _writeQueue_fifo_3_data_out[7:3];
  assign writeQueue_dataOut_3_writeData_groupCounter = _writeQueue_fifo_3_data_out[12:8];
  assign writeQueue_dataOut_3_writeData_mask = _writeQueue_fifo_3_data_out[16:13];
  assign writeQueue_dataOut_3_writeData_data = _writeQueue_fifo_3_data_out[48:17];
  assign writeQueue_dataOut_3_ffoByOther = _writeQueue_fifo_3_data_out[49];
  wire              writeQueue_3_deq_bits_ffoByOther = writeQueue_dataOut_3_ffoByOther;
  assign writeQueue_3_deq_bits_writeData_data = writeQueue_dataOut_3_writeData_data;
  assign writeQueue_3_deq_bits_writeData_mask = writeQueue_dataOut_3_writeData_mask;
  wire [4:0]        writeQueue_3_deq_bits_writeData_groupCounter = writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]        writeQueue_3_deq_bits_writeData_vd = writeQueue_dataOut_3_writeData_vd;
  wire [2:0]        writeQueue_3_deq_bits_index = writeQueue_dataOut_3_index;
  wire              writeQueue_3_enq_ready = ~_writeQueue_fifo_3_full;
  wire              writeQueue_3_enq_valid;
  assign writeQueue_4_deq_valid = ~_writeQueue_fifo_4_empty;
  wire              exeResp_4_valid_0 = writeQueue_4_deq_valid;
  wire              writeQueue_dataOut_4_ffoByOther;
  wire [31:0]       writeQueue_dataOut_4_writeData_data;
  wire [31:0]       exeResp_4_bits_data_0 = writeQueue_4_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_4_writeData_mask;
  wire [3:0]        exeResp_4_bits_mask_0 = writeQueue_4_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_4_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_4_writeData_vd;
  wire [2:0]        writeQueue_dataOut_4_index;
  wire [4:0]        writeQueue_4_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_4_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_4 = {writeQueue_4_enq_bits_writeData_groupCounter, writeQueue_4_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_4_enq_bits_writeData_data;
  wire [3:0]        writeQueue_4_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_8 = {writeQueue_4_enq_bits_writeData_data, writeQueue_4_enq_bits_writeData_mask};
  wire              writeQueue_4_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_9 = {writeQueue_4_enq_bits_ffoByOther, writeQueue_dataIn_hi_8, writeQueue_dataIn_lo_4};
  wire [49:0]       writeQueue_dataIn_4 = {writeQueue_dataIn_hi_9, writeQueue_4_enq_bits_index};
  assign writeQueue_dataOut_4_index = _writeQueue_fifo_4_data_out[2:0];
  assign writeQueue_dataOut_4_writeData_vd = _writeQueue_fifo_4_data_out[7:3];
  assign writeQueue_dataOut_4_writeData_groupCounter = _writeQueue_fifo_4_data_out[12:8];
  assign writeQueue_dataOut_4_writeData_mask = _writeQueue_fifo_4_data_out[16:13];
  assign writeQueue_dataOut_4_writeData_data = _writeQueue_fifo_4_data_out[48:17];
  assign writeQueue_dataOut_4_ffoByOther = _writeQueue_fifo_4_data_out[49];
  wire              writeQueue_4_deq_bits_ffoByOther = writeQueue_dataOut_4_ffoByOther;
  assign writeQueue_4_deq_bits_writeData_data = writeQueue_dataOut_4_writeData_data;
  assign writeQueue_4_deq_bits_writeData_mask = writeQueue_dataOut_4_writeData_mask;
  wire [4:0]        writeQueue_4_deq_bits_writeData_groupCounter = writeQueue_dataOut_4_writeData_groupCounter;
  wire [4:0]        writeQueue_4_deq_bits_writeData_vd = writeQueue_dataOut_4_writeData_vd;
  wire [2:0]        writeQueue_4_deq_bits_index = writeQueue_dataOut_4_index;
  wire              writeQueue_4_enq_ready = ~_writeQueue_fifo_4_full;
  wire              writeQueue_4_enq_valid;
  assign writeQueue_5_deq_valid = ~_writeQueue_fifo_5_empty;
  wire              exeResp_5_valid_0 = writeQueue_5_deq_valid;
  wire              writeQueue_dataOut_5_ffoByOther;
  wire [31:0]       writeQueue_dataOut_5_writeData_data;
  wire [31:0]       exeResp_5_bits_data_0 = writeQueue_5_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_5_writeData_mask;
  wire [3:0]        exeResp_5_bits_mask_0 = writeQueue_5_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_5_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_5_writeData_vd;
  wire [2:0]        writeQueue_dataOut_5_index;
  wire [4:0]        writeQueue_5_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_5_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_5 = {writeQueue_5_enq_bits_writeData_groupCounter, writeQueue_5_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_5_enq_bits_writeData_data;
  wire [3:0]        writeQueue_5_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_10 = {writeQueue_5_enq_bits_writeData_data, writeQueue_5_enq_bits_writeData_mask};
  wire              writeQueue_5_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_11 = {writeQueue_5_enq_bits_ffoByOther, writeQueue_dataIn_hi_10, writeQueue_dataIn_lo_5};
  wire [49:0]       writeQueue_dataIn_5 = {writeQueue_dataIn_hi_11, writeQueue_5_enq_bits_index};
  assign writeQueue_dataOut_5_index = _writeQueue_fifo_5_data_out[2:0];
  assign writeQueue_dataOut_5_writeData_vd = _writeQueue_fifo_5_data_out[7:3];
  assign writeQueue_dataOut_5_writeData_groupCounter = _writeQueue_fifo_5_data_out[12:8];
  assign writeQueue_dataOut_5_writeData_mask = _writeQueue_fifo_5_data_out[16:13];
  assign writeQueue_dataOut_5_writeData_data = _writeQueue_fifo_5_data_out[48:17];
  assign writeQueue_dataOut_5_ffoByOther = _writeQueue_fifo_5_data_out[49];
  wire              writeQueue_5_deq_bits_ffoByOther = writeQueue_dataOut_5_ffoByOther;
  assign writeQueue_5_deq_bits_writeData_data = writeQueue_dataOut_5_writeData_data;
  assign writeQueue_5_deq_bits_writeData_mask = writeQueue_dataOut_5_writeData_mask;
  wire [4:0]        writeQueue_5_deq_bits_writeData_groupCounter = writeQueue_dataOut_5_writeData_groupCounter;
  wire [4:0]        writeQueue_5_deq_bits_writeData_vd = writeQueue_dataOut_5_writeData_vd;
  wire [2:0]        writeQueue_5_deq_bits_index = writeQueue_dataOut_5_index;
  wire              writeQueue_5_enq_ready = ~_writeQueue_fifo_5_full;
  wire              writeQueue_5_enq_valid;
  assign writeQueue_6_deq_valid = ~_writeQueue_fifo_6_empty;
  wire              exeResp_6_valid_0 = writeQueue_6_deq_valid;
  wire              writeQueue_dataOut_6_ffoByOther;
  wire [31:0]       writeQueue_dataOut_6_writeData_data;
  wire [31:0]       exeResp_6_bits_data_0 = writeQueue_6_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_6_writeData_mask;
  wire [3:0]        exeResp_6_bits_mask_0 = writeQueue_6_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_6_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_6_writeData_vd;
  wire [2:0]        writeQueue_dataOut_6_index;
  wire [4:0]        writeQueue_6_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_6_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_6 = {writeQueue_6_enq_bits_writeData_groupCounter, writeQueue_6_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_6_enq_bits_writeData_data;
  wire [3:0]        writeQueue_6_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_12 = {writeQueue_6_enq_bits_writeData_data, writeQueue_6_enq_bits_writeData_mask};
  wire              writeQueue_6_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_13 = {writeQueue_6_enq_bits_ffoByOther, writeQueue_dataIn_hi_12, writeQueue_dataIn_lo_6};
  wire [49:0]       writeQueue_dataIn_6 = {writeQueue_dataIn_hi_13, writeQueue_6_enq_bits_index};
  assign writeQueue_dataOut_6_index = _writeQueue_fifo_6_data_out[2:0];
  assign writeQueue_dataOut_6_writeData_vd = _writeQueue_fifo_6_data_out[7:3];
  assign writeQueue_dataOut_6_writeData_groupCounter = _writeQueue_fifo_6_data_out[12:8];
  assign writeQueue_dataOut_6_writeData_mask = _writeQueue_fifo_6_data_out[16:13];
  assign writeQueue_dataOut_6_writeData_data = _writeQueue_fifo_6_data_out[48:17];
  assign writeQueue_dataOut_6_ffoByOther = _writeQueue_fifo_6_data_out[49];
  wire              writeQueue_6_deq_bits_ffoByOther = writeQueue_dataOut_6_ffoByOther;
  assign writeQueue_6_deq_bits_writeData_data = writeQueue_dataOut_6_writeData_data;
  assign writeQueue_6_deq_bits_writeData_mask = writeQueue_dataOut_6_writeData_mask;
  wire [4:0]        writeQueue_6_deq_bits_writeData_groupCounter = writeQueue_dataOut_6_writeData_groupCounter;
  wire [4:0]        writeQueue_6_deq_bits_writeData_vd = writeQueue_dataOut_6_writeData_vd;
  wire [2:0]        writeQueue_6_deq_bits_index = writeQueue_dataOut_6_index;
  wire              writeQueue_6_enq_ready = ~_writeQueue_fifo_6_full;
  wire              writeQueue_6_enq_valid;
  assign writeQueue_7_deq_valid = ~_writeQueue_fifo_7_empty;
  wire              exeResp_7_valid_0 = writeQueue_7_deq_valid;
  wire              writeQueue_dataOut_7_ffoByOther;
  wire [31:0]       writeQueue_dataOut_7_writeData_data;
  wire [31:0]       exeResp_7_bits_data_0 = writeQueue_7_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_7_writeData_mask;
  wire [3:0]        exeResp_7_bits_mask_0 = writeQueue_7_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_7_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_7_writeData_vd;
  wire [2:0]        writeQueue_dataOut_7_index;
  wire [4:0]        writeQueue_7_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_7_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_7 = {writeQueue_7_enq_bits_writeData_groupCounter, writeQueue_7_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_7_enq_bits_writeData_data;
  wire [3:0]        writeQueue_7_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_14 = {writeQueue_7_enq_bits_writeData_data, writeQueue_7_enq_bits_writeData_mask};
  wire              writeQueue_7_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_15 = {writeQueue_7_enq_bits_ffoByOther, writeQueue_dataIn_hi_14, writeQueue_dataIn_lo_7};
  wire [49:0]       writeQueue_dataIn_7 = {writeQueue_dataIn_hi_15, writeQueue_7_enq_bits_index};
  assign writeQueue_dataOut_7_index = _writeQueue_fifo_7_data_out[2:0];
  assign writeQueue_dataOut_7_writeData_vd = _writeQueue_fifo_7_data_out[7:3];
  assign writeQueue_dataOut_7_writeData_groupCounter = _writeQueue_fifo_7_data_out[12:8];
  assign writeQueue_dataOut_7_writeData_mask = _writeQueue_fifo_7_data_out[16:13];
  assign writeQueue_dataOut_7_writeData_data = _writeQueue_fifo_7_data_out[48:17];
  assign writeQueue_dataOut_7_ffoByOther = _writeQueue_fifo_7_data_out[49];
  wire              writeQueue_7_deq_bits_ffoByOther = writeQueue_dataOut_7_ffoByOther;
  assign writeQueue_7_deq_bits_writeData_data = writeQueue_dataOut_7_writeData_data;
  assign writeQueue_7_deq_bits_writeData_mask = writeQueue_dataOut_7_writeData_mask;
  wire [4:0]        writeQueue_7_deq_bits_writeData_groupCounter = writeQueue_dataOut_7_writeData_groupCounter;
  wire [4:0]        writeQueue_7_deq_bits_writeData_vd = writeQueue_dataOut_7_writeData_vd;
  wire [2:0]        writeQueue_7_deq_bits_index = writeQueue_dataOut_7_index;
  wire              writeQueue_7_enq_ready = ~_writeQueue_fifo_7_full;
  wire              writeQueue_7_enq_valid;
  assign writeQueue_8_deq_valid = ~_writeQueue_fifo_8_empty;
  wire              exeResp_8_valid_0 = writeQueue_8_deq_valid;
  wire              writeQueue_dataOut_8_ffoByOther;
  wire [31:0]       writeQueue_dataOut_8_writeData_data;
  wire [31:0]       exeResp_8_bits_data_0 = writeQueue_8_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_8_writeData_mask;
  wire [3:0]        exeResp_8_bits_mask_0 = writeQueue_8_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_8_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_8_writeData_vd;
  wire [2:0]        writeQueue_dataOut_8_index;
  wire [4:0]        writeQueue_8_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_8_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_8 = {writeQueue_8_enq_bits_writeData_groupCounter, writeQueue_8_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_8_enq_bits_writeData_data;
  wire [3:0]        writeQueue_8_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_16 = {writeQueue_8_enq_bits_writeData_data, writeQueue_8_enq_bits_writeData_mask};
  wire              writeQueue_8_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_17 = {writeQueue_8_enq_bits_ffoByOther, writeQueue_dataIn_hi_16, writeQueue_dataIn_lo_8};
  wire [49:0]       writeQueue_dataIn_8 = {writeQueue_dataIn_hi_17, writeQueue_8_enq_bits_index};
  assign writeQueue_dataOut_8_index = _writeQueue_fifo_8_data_out[2:0];
  assign writeQueue_dataOut_8_writeData_vd = _writeQueue_fifo_8_data_out[7:3];
  assign writeQueue_dataOut_8_writeData_groupCounter = _writeQueue_fifo_8_data_out[12:8];
  assign writeQueue_dataOut_8_writeData_mask = _writeQueue_fifo_8_data_out[16:13];
  assign writeQueue_dataOut_8_writeData_data = _writeQueue_fifo_8_data_out[48:17];
  assign writeQueue_dataOut_8_ffoByOther = _writeQueue_fifo_8_data_out[49];
  wire              writeQueue_8_deq_bits_ffoByOther = writeQueue_dataOut_8_ffoByOther;
  assign writeQueue_8_deq_bits_writeData_data = writeQueue_dataOut_8_writeData_data;
  assign writeQueue_8_deq_bits_writeData_mask = writeQueue_dataOut_8_writeData_mask;
  wire [4:0]        writeQueue_8_deq_bits_writeData_groupCounter = writeQueue_dataOut_8_writeData_groupCounter;
  wire [4:0]        writeQueue_8_deq_bits_writeData_vd = writeQueue_dataOut_8_writeData_vd;
  wire [2:0]        writeQueue_8_deq_bits_index = writeQueue_dataOut_8_index;
  wire              writeQueue_8_enq_ready = ~_writeQueue_fifo_8_full;
  wire              writeQueue_8_enq_valid;
  assign writeQueue_9_deq_valid = ~_writeQueue_fifo_9_empty;
  wire              exeResp_9_valid_0 = writeQueue_9_deq_valid;
  wire              writeQueue_dataOut_9_ffoByOther;
  wire [31:0]       writeQueue_dataOut_9_writeData_data;
  wire [31:0]       exeResp_9_bits_data_0 = writeQueue_9_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_9_writeData_mask;
  wire [3:0]        exeResp_9_bits_mask_0 = writeQueue_9_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_9_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_9_writeData_vd;
  wire [2:0]        writeQueue_dataOut_9_index;
  wire [4:0]        writeQueue_9_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_9_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_9 = {writeQueue_9_enq_bits_writeData_groupCounter, writeQueue_9_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_9_enq_bits_writeData_data;
  wire [3:0]        writeQueue_9_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_18 = {writeQueue_9_enq_bits_writeData_data, writeQueue_9_enq_bits_writeData_mask};
  wire              writeQueue_9_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_19 = {writeQueue_9_enq_bits_ffoByOther, writeQueue_dataIn_hi_18, writeQueue_dataIn_lo_9};
  wire [49:0]       writeQueue_dataIn_9 = {writeQueue_dataIn_hi_19, writeQueue_9_enq_bits_index};
  assign writeQueue_dataOut_9_index = _writeQueue_fifo_9_data_out[2:0];
  assign writeQueue_dataOut_9_writeData_vd = _writeQueue_fifo_9_data_out[7:3];
  assign writeQueue_dataOut_9_writeData_groupCounter = _writeQueue_fifo_9_data_out[12:8];
  assign writeQueue_dataOut_9_writeData_mask = _writeQueue_fifo_9_data_out[16:13];
  assign writeQueue_dataOut_9_writeData_data = _writeQueue_fifo_9_data_out[48:17];
  assign writeQueue_dataOut_9_ffoByOther = _writeQueue_fifo_9_data_out[49];
  wire              writeQueue_9_deq_bits_ffoByOther = writeQueue_dataOut_9_ffoByOther;
  assign writeQueue_9_deq_bits_writeData_data = writeQueue_dataOut_9_writeData_data;
  assign writeQueue_9_deq_bits_writeData_mask = writeQueue_dataOut_9_writeData_mask;
  wire [4:0]        writeQueue_9_deq_bits_writeData_groupCounter = writeQueue_dataOut_9_writeData_groupCounter;
  wire [4:0]        writeQueue_9_deq_bits_writeData_vd = writeQueue_dataOut_9_writeData_vd;
  wire [2:0]        writeQueue_9_deq_bits_index = writeQueue_dataOut_9_index;
  wire              writeQueue_9_enq_ready = ~_writeQueue_fifo_9_full;
  wire              writeQueue_9_enq_valid;
  assign writeQueue_10_deq_valid = ~_writeQueue_fifo_10_empty;
  wire              exeResp_10_valid_0 = writeQueue_10_deq_valid;
  wire              writeQueue_dataOut_10_ffoByOther;
  wire [31:0]       writeQueue_dataOut_10_writeData_data;
  wire [31:0]       exeResp_10_bits_data_0 = writeQueue_10_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_10_writeData_mask;
  wire [3:0]        exeResp_10_bits_mask_0 = writeQueue_10_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_10_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_10_writeData_vd;
  wire [2:0]        writeQueue_dataOut_10_index;
  wire [4:0]        writeQueue_10_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_10_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_10 = {writeQueue_10_enq_bits_writeData_groupCounter, writeQueue_10_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_10_enq_bits_writeData_data;
  wire [3:0]        writeQueue_10_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_20 = {writeQueue_10_enq_bits_writeData_data, writeQueue_10_enq_bits_writeData_mask};
  wire              writeQueue_10_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_21 = {writeQueue_10_enq_bits_ffoByOther, writeQueue_dataIn_hi_20, writeQueue_dataIn_lo_10};
  wire [49:0]       writeQueue_dataIn_10 = {writeQueue_dataIn_hi_21, writeQueue_10_enq_bits_index};
  assign writeQueue_dataOut_10_index = _writeQueue_fifo_10_data_out[2:0];
  assign writeQueue_dataOut_10_writeData_vd = _writeQueue_fifo_10_data_out[7:3];
  assign writeQueue_dataOut_10_writeData_groupCounter = _writeQueue_fifo_10_data_out[12:8];
  assign writeQueue_dataOut_10_writeData_mask = _writeQueue_fifo_10_data_out[16:13];
  assign writeQueue_dataOut_10_writeData_data = _writeQueue_fifo_10_data_out[48:17];
  assign writeQueue_dataOut_10_ffoByOther = _writeQueue_fifo_10_data_out[49];
  wire              writeQueue_10_deq_bits_ffoByOther = writeQueue_dataOut_10_ffoByOther;
  assign writeQueue_10_deq_bits_writeData_data = writeQueue_dataOut_10_writeData_data;
  assign writeQueue_10_deq_bits_writeData_mask = writeQueue_dataOut_10_writeData_mask;
  wire [4:0]        writeQueue_10_deq_bits_writeData_groupCounter = writeQueue_dataOut_10_writeData_groupCounter;
  wire [4:0]        writeQueue_10_deq_bits_writeData_vd = writeQueue_dataOut_10_writeData_vd;
  wire [2:0]        writeQueue_10_deq_bits_index = writeQueue_dataOut_10_index;
  wire              writeQueue_10_enq_ready = ~_writeQueue_fifo_10_full;
  wire              writeQueue_10_enq_valid;
  assign writeQueue_11_deq_valid = ~_writeQueue_fifo_11_empty;
  wire              exeResp_11_valid_0 = writeQueue_11_deq_valid;
  wire              writeQueue_dataOut_11_ffoByOther;
  wire [31:0]       writeQueue_dataOut_11_writeData_data;
  wire [31:0]       exeResp_11_bits_data_0 = writeQueue_11_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_11_writeData_mask;
  wire [3:0]        exeResp_11_bits_mask_0 = writeQueue_11_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_11_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_11_writeData_vd;
  wire [2:0]        writeQueue_dataOut_11_index;
  wire [4:0]        writeQueue_11_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_11_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_11 = {writeQueue_11_enq_bits_writeData_groupCounter, writeQueue_11_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_11_enq_bits_writeData_data;
  wire [3:0]        writeQueue_11_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_22 = {writeQueue_11_enq_bits_writeData_data, writeQueue_11_enq_bits_writeData_mask};
  wire              writeQueue_11_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_23 = {writeQueue_11_enq_bits_ffoByOther, writeQueue_dataIn_hi_22, writeQueue_dataIn_lo_11};
  wire [49:0]       writeQueue_dataIn_11 = {writeQueue_dataIn_hi_23, writeQueue_11_enq_bits_index};
  assign writeQueue_dataOut_11_index = _writeQueue_fifo_11_data_out[2:0];
  assign writeQueue_dataOut_11_writeData_vd = _writeQueue_fifo_11_data_out[7:3];
  assign writeQueue_dataOut_11_writeData_groupCounter = _writeQueue_fifo_11_data_out[12:8];
  assign writeQueue_dataOut_11_writeData_mask = _writeQueue_fifo_11_data_out[16:13];
  assign writeQueue_dataOut_11_writeData_data = _writeQueue_fifo_11_data_out[48:17];
  assign writeQueue_dataOut_11_ffoByOther = _writeQueue_fifo_11_data_out[49];
  wire              writeQueue_11_deq_bits_ffoByOther = writeQueue_dataOut_11_ffoByOther;
  assign writeQueue_11_deq_bits_writeData_data = writeQueue_dataOut_11_writeData_data;
  assign writeQueue_11_deq_bits_writeData_mask = writeQueue_dataOut_11_writeData_mask;
  wire [4:0]        writeQueue_11_deq_bits_writeData_groupCounter = writeQueue_dataOut_11_writeData_groupCounter;
  wire [4:0]        writeQueue_11_deq_bits_writeData_vd = writeQueue_dataOut_11_writeData_vd;
  wire [2:0]        writeQueue_11_deq_bits_index = writeQueue_dataOut_11_index;
  wire              writeQueue_11_enq_ready = ~_writeQueue_fifo_11_full;
  wire              writeQueue_11_enq_valid;
  assign writeQueue_12_deq_valid = ~_writeQueue_fifo_12_empty;
  wire              exeResp_12_valid_0 = writeQueue_12_deq_valid;
  wire              writeQueue_dataOut_12_ffoByOther;
  wire [31:0]       writeQueue_dataOut_12_writeData_data;
  wire [31:0]       exeResp_12_bits_data_0 = writeQueue_12_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_12_writeData_mask;
  wire [3:0]        exeResp_12_bits_mask_0 = writeQueue_12_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_12_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_12_writeData_vd;
  wire [2:0]        writeQueue_dataOut_12_index;
  wire [4:0]        writeQueue_12_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_12_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_12 = {writeQueue_12_enq_bits_writeData_groupCounter, writeQueue_12_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_12_enq_bits_writeData_data;
  wire [3:0]        writeQueue_12_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_24 = {writeQueue_12_enq_bits_writeData_data, writeQueue_12_enq_bits_writeData_mask};
  wire              writeQueue_12_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_25 = {writeQueue_12_enq_bits_ffoByOther, writeQueue_dataIn_hi_24, writeQueue_dataIn_lo_12};
  wire [49:0]       writeQueue_dataIn_12 = {writeQueue_dataIn_hi_25, writeQueue_12_enq_bits_index};
  assign writeQueue_dataOut_12_index = _writeQueue_fifo_12_data_out[2:0];
  assign writeQueue_dataOut_12_writeData_vd = _writeQueue_fifo_12_data_out[7:3];
  assign writeQueue_dataOut_12_writeData_groupCounter = _writeQueue_fifo_12_data_out[12:8];
  assign writeQueue_dataOut_12_writeData_mask = _writeQueue_fifo_12_data_out[16:13];
  assign writeQueue_dataOut_12_writeData_data = _writeQueue_fifo_12_data_out[48:17];
  assign writeQueue_dataOut_12_ffoByOther = _writeQueue_fifo_12_data_out[49];
  wire              writeQueue_12_deq_bits_ffoByOther = writeQueue_dataOut_12_ffoByOther;
  assign writeQueue_12_deq_bits_writeData_data = writeQueue_dataOut_12_writeData_data;
  assign writeQueue_12_deq_bits_writeData_mask = writeQueue_dataOut_12_writeData_mask;
  wire [4:0]        writeQueue_12_deq_bits_writeData_groupCounter = writeQueue_dataOut_12_writeData_groupCounter;
  wire [4:0]        writeQueue_12_deq_bits_writeData_vd = writeQueue_dataOut_12_writeData_vd;
  wire [2:0]        writeQueue_12_deq_bits_index = writeQueue_dataOut_12_index;
  wire              writeQueue_12_enq_ready = ~_writeQueue_fifo_12_full;
  wire              writeQueue_12_enq_valid;
  assign writeQueue_13_deq_valid = ~_writeQueue_fifo_13_empty;
  wire              exeResp_13_valid_0 = writeQueue_13_deq_valid;
  wire              writeQueue_dataOut_13_ffoByOther;
  wire [31:0]       writeQueue_dataOut_13_writeData_data;
  wire [31:0]       exeResp_13_bits_data_0 = writeQueue_13_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_13_writeData_mask;
  wire [3:0]        exeResp_13_bits_mask_0 = writeQueue_13_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_13_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_13_writeData_vd;
  wire [2:0]        writeQueue_dataOut_13_index;
  wire [4:0]        writeQueue_13_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_13_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_13 = {writeQueue_13_enq_bits_writeData_groupCounter, writeQueue_13_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_13_enq_bits_writeData_data;
  wire [3:0]        writeQueue_13_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_26 = {writeQueue_13_enq_bits_writeData_data, writeQueue_13_enq_bits_writeData_mask};
  wire              writeQueue_13_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_27 = {writeQueue_13_enq_bits_ffoByOther, writeQueue_dataIn_hi_26, writeQueue_dataIn_lo_13};
  wire [49:0]       writeQueue_dataIn_13 = {writeQueue_dataIn_hi_27, writeQueue_13_enq_bits_index};
  assign writeQueue_dataOut_13_index = _writeQueue_fifo_13_data_out[2:0];
  assign writeQueue_dataOut_13_writeData_vd = _writeQueue_fifo_13_data_out[7:3];
  assign writeQueue_dataOut_13_writeData_groupCounter = _writeQueue_fifo_13_data_out[12:8];
  assign writeQueue_dataOut_13_writeData_mask = _writeQueue_fifo_13_data_out[16:13];
  assign writeQueue_dataOut_13_writeData_data = _writeQueue_fifo_13_data_out[48:17];
  assign writeQueue_dataOut_13_ffoByOther = _writeQueue_fifo_13_data_out[49];
  wire              writeQueue_13_deq_bits_ffoByOther = writeQueue_dataOut_13_ffoByOther;
  assign writeQueue_13_deq_bits_writeData_data = writeQueue_dataOut_13_writeData_data;
  assign writeQueue_13_deq_bits_writeData_mask = writeQueue_dataOut_13_writeData_mask;
  wire [4:0]        writeQueue_13_deq_bits_writeData_groupCounter = writeQueue_dataOut_13_writeData_groupCounter;
  wire [4:0]        writeQueue_13_deq_bits_writeData_vd = writeQueue_dataOut_13_writeData_vd;
  wire [2:0]        writeQueue_13_deq_bits_index = writeQueue_dataOut_13_index;
  wire              writeQueue_13_enq_ready = ~_writeQueue_fifo_13_full;
  wire              writeQueue_13_enq_valid;
  assign writeQueue_14_deq_valid = ~_writeQueue_fifo_14_empty;
  wire              exeResp_14_valid_0 = writeQueue_14_deq_valid;
  wire              writeQueue_dataOut_14_ffoByOther;
  wire [31:0]       writeQueue_dataOut_14_writeData_data;
  wire [31:0]       exeResp_14_bits_data_0 = writeQueue_14_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_14_writeData_mask;
  wire [3:0]        exeResp_14_bits_mask_0 = writeQueue_14_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_14_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_14_writeData_vd;
  wire [2:0]        writeQueue_dataOut_14_index;
  wire [4:0]        writeQueue_14_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_14_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_14 = {writeQueue_14_enq_bits_writeData_groupCounter, writeQueue_14_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_14_enq_bits_writeData_data;
  wire [3:0]        writeQueue_14_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_28 = {writeQueue_14_enq_bits_writeData_data, writeQueue_14_enq_bits_writeData_mask};
  wire              writeQueue_14_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_29 = {writeQueue_14_enq_bits_ffoByOther, writeQueue_dataIn_hi_28, writeQueue_dataIn_lo_14};
  wire [49:0]       writeQueue_dataIn_14 = {writeQueue_dataIn_hi_29, writeQueue_14_enq_bits_index};
  assign writeQueue_dataOut_14_index = _writeQueue_fifo_14_data_out[2:0];
  assign writeQueue_dataOut_14_writeData_vd = _writeQueue_fifo_14_data_out[7:3];
  assign writeQueue_dataOut_14_writeData_groupCounter = _writeQueue_fifo_14_data_out[12:8];
  assign writeQueue_dataOut_14_writeData_mask = _writeQueue_fifo_14_data_out[16:13];
  assign writeQueue_dataOut_14_writeData_data = _writeQueue_fifo_14_data_out[48:17];
  assign writeQueue_dataOut_14_ffoByOther = _writeQueue_fifo_14_data_out[49];
  wire              writeQueue_14_deq_bits_ffoByOther = writeQueue_dataOut_14_ffoByOther;
  assign writeQueue_14_deq_bits_writeData_data = writeQueue_dataOut_14_writeData_data;
  assign writeQueue_14_deq_bits_writeData_mask = writeQueue_dataOut_14_writeData_mask;
  wire [4:0]        writeQueue_14_deq_bits_writeData_groupCounter = writeQueue_dataOut_14_writeData_groupCounter;
  wire [4:0]        writeQueue_14_deq_bits_writeData_vd = writeQueue_dataOut_14_writeData_vd;
  wire [2:0]        writeQueue_14_deq_bits_index = writeQueue_dataOut_14_index;
  wire              writeQueue_14_enq_ready = ~_writeQueue_fifo_14_full;
  wire              writeQueue_14_enq_valid;
  assign writeQueue_15_deq_valid = ~_writeQueue_fifo_15_empty;
  wire              exeResp_15_valid_0 = writeQueue_15_deq_valid;
  wire              writeQueue_dataOut_15_ffoByOther;
  wire [31:0]       writeQueue_dataOut_15_writeData_data;
  wire [31:0]       exeResp_15_bits_data_0 = writeQueue_15_deq_bits_writeData_data;
  wire [3:0]        writeQueue_dataOut_15_writeData_mask;
  wire [3:0]        exeResp_15_bits_mask_0 = writeQueue_15_deq_bits_writeData_mask;
  wire [4:0]        writeQueue_dataOut_15_writeData_groupCounter;
  wire [4:0]        writeQueue_dataOut_15_writeData_vd;
  wire [2:0]        writeQueue_dataOut_15_index;
  wire [4:0]        writeQueue_15_enq_bits_writeData_groupCounter;
  wire [4:0]        writeQueue_15_enq_bits_writeData_vd;
  wire [9:0]        writeQueue_dataIn_lo_15 = {writeQueue_15_enq_bits_writeData_groupCounter, writeQueue_15_enq_bits_writeData_vd};
  wire [31:0]       writeQueue_15_enq_bits_writeData_data;
  wire [3:0]        writeQueue_15_enq_bits_writeData_mask;
  wire [35:0]       writeQueue_dataIn_hi_30 = {writeQueue_15_enq_bits_writeData_data, writeQueue_15_enq_bits_writeData_mask};
  wire              writeQueue_15_enq_bits_ffoByOther;
  wire [46:0]       writeQueue_dataIn_hi_31 = {writeQueue_15_enq_bits_ffoByOther, writeQueue_dataIn_hi_30, writeQueue_dataIn_lo_15};
  wire [49:0]       writeQueue_dataIn_15 = {writeQueue_dataIn_hi_31, writeQueue_15_enq_bits_index};
  assign writeQueue_dataOut_15_index = _writeQueue_fifo_15_data_out[2:0];
  assign writeQueue_dataOut_15_writeData_vd = _writeQueue_fifo_15_data_out[7:3];
  assign writeQueue_dataOut_15_writeData_groupCounter = _writeQueue_fifo_15_data_out[12:8];
  assign writeQueue_dataOut_15_writeData_mask = _writeQueue_fifo_15_data_out[16:13];
  assign writeQueue_dataOut_15_writeData_data = _writeQueue_fifo_15_data_out[48:17];
  assign writeQueue_dataOut_15_ffoByOther = _writeQueue_fifo_15_data_out[49];
  wire              writeQueue_15_deq_bits_ffoByOther = writeQueue_dataOut_15_ffoByOther;
  assign writeQueue_15_deq_bits_writeData_data = writeQueue_dataOut_15_writeData_data;
  assign writeQueue_15_deq_bits_writeData_mask = writeQueue_dataOut_15_writeData_mask;
  wire [4:0]        writeQueue_15_deq_bits_writeData_groupCounter = writeQueue_dataOut_15_writeData_groupCounter;
  wire [4:0]        writeQueue_15_deq_bits_writeData_vd = writeQueue_dataOut_15_writeData_vd;
  wire [2:0]        writeQueue_15_deq_bits_index = writeQueue_dataOut_15_index;
  wire              writeQueue_15_enq_ready = ~_writeQueue_fifo_15_full;
  wire              writeQueue_15_enq_valid;
  wire              dataNotInShifter_readTypeWriteVrf = waiteStageDeqFire & WillWriteLane[0];
  assign writeQueue_0_enq_valid = _maskedWrite_out_0_valid | dataNotInShifter_readTypeWriteVrf;
  assign writeQueue_0_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_vd : 5'h0;
  assign writeQueue_0_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_groupCounter : _maskedWrite_out_0_bits_writeData_groupCounter;
  assign writeQueue_0_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_mask : _maskedWrite_out_0_bits_writeData_mask;
  assign writeQueue_0_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_data : _maskedWrite_out_0_bits_writeData_data;
  assign writeQueue_0_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf & _maskedWrite_out_0_bits_ffoByOther;
  wire [4:0]        exeResp_0_bits_vd_0 = instReg_vd + {1'h0, writeQueue_0_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_0_bits_offset_0 = writeQueue_0_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter;
  wire              _dataNotInShifter_T = exeResp_0_ready_0 & exeResp_0_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange = _dataNotInShifter_T ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_1 = waiteStageDeqFire & WillWriteLane[1];
  assign writeQueue_1_enq_valid = _maskedWrite_out_1_valid | dataNotInShifter_readTypeWriteVrf_1;
  assign writeQueue_1_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_vd : 5'h0;
  assign writeQueue_1_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_groupCounter : _maskedWrite_out_1_bits_writeData_groupCounter;
  assign writeQueue_1_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_mask : _maskedWrite_out_1_bits_writeData_mask;
  assign writeQueue_1_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_data : _maskedWrite_out_1_bits_writeData_data;
  assign writeQueue_1_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_1 & _maskedWrite_out_1_bits_ffoByOther;
  wire [4:0]        exeResp_1_bits_vd_0 = instReg_vd + {1'h0, writeQueue_1_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_1_bits_offset_0 = writeQueue_1_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_1;
  wire              _dataNotInShifter_T_3 = exeResp_1_ready_0 & exeResp_1_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_1 = _dataNotInShifter_T_3 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_2 = waiteStageDeqFire & WillWriteLane[2];
  assign writeQueue_2_enq_valid = _maskedWrite_out_2_valid | dataNotInShifter_readTypeWriteVrf_2;
  assign writeQueue_2_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_vd : 5'h0;
  assign writeQueue_2_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_groupCounter : _maskedWrite_out_2_bits_writeData_groupCounter;
  assign writeQueue_2_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_mask : _maskedWrite_out_2_bits_writeData_mask;
  assign writeQueue_2_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_data : _maskedWrite_out_2_bits_writeData_data;
  assign writeQueue_2_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_2 & _maskedWrite_out_2_bits_ffoByOther;
  wire [4:0]        exeResp_2_bits_vd_0 = instReg_vd + {1'h0, writeQueue_2_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_2_bits_offset_0 = writeQueue_2_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_2;
  wire              _dataNotInShifter_T_6 = exeResp_2_ready_0 & exeResp_2_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_2 = _dataNotInShifter_T_6 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_3 = waiteStageDeqFire & WillWriteLane[3];
  assign writeQueue_3_enq_valid = _maskedWrite_out_3_valid | dataNotInShifter_readTypeWriteVrf_3;
  assign writeQueue_3_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_vd : 5'h0;
  assign writeQueue_3_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_groupCounter : _maskedWrite_out_3_bits_writeData_groupCounter;
  assign writeQueue_3_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_mask : _maskedWrite_out_3_bits_writeData_mask;
  assign writeQueue_3_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_data : _maskedWrite_out_3_bits_writeData_data;
  assign writeQueue_3_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_3 & _maskedWrite_out_3_bits_ffoByOther;
  wire [4:0]        exeResp_3_bits_vd_0 = instReg_vd + {1'h0, writeQueue_3_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_3_bits_offset_0 = writeQueue_3_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_3;
  wire              _dataNotInShifter_T_9 = exeResp_3_ready_0 & exeResp_3_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_3 = _dataNotInShifter_T_9 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_4 = waiteStageDeqFire & WillWriteLane[4];
  assign writeQueue_4_enq_valid = _maskedWrite_out_4_valid | dataNotInShifter_readTypeWriteVrf_4;
  assign writeQueue_4_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_vd : 5'h0;
  assign writeQueue_4_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_groupCounter : _maskedWrite_out_4_bits_writeData_groupCounter;
  assign writeQueue_4_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_mask : _maskedWrite_out_4_bits_writeData_mask;
  assign writeQueue_4_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_4 ? writeRequest_4_writeData_data : _maskedWrite_out_4_bits_writeData_data;
  assign writeQueue_4_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_4 & _maskedWrite_out_4_bits_ffoByOther;
  wire [4:0]        exeResp_4_bits_vd_0 = instReg_vd + {1'h0, writeQueue_4_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_4_bits_offset_0 = writeQueue_4_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_4;
  wire              _dataNotInShifter_T_12 = exeResp_4_ready_0 & exeResp_4_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_4 = _dataNotInShifter_T_12 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_5 = waiteStageDeqFire & WillWriteLane[5];
  assign writeQueue_5_enq_valid = _maskedWrite_out_5_valid | dataNotInShifter_readTypeWriteVrf_5;
  assign writeQueue_5_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_vd : 5'h0;
  assign writeQueue_5_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_groupCounter : _maskedWrite_out_5_bits_writeData_groupCounter;
  assign writeQueue_5_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_mask : _maskedWrite_out_5_bits_writeData_mask;
  assign writeQueue_5_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_5 ? writeRequest_5_writeData_data : _maskedWrite_out_5_bits_writeData_data;
  assign writeQueue_5_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_5 & _maskedWrite_out_5_bits_ffoByOther;
  wire [4:0]        exeResp_5_bits_vd_0 = instReg_vd + {1'h0, writeQueue_5_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_5_bits_offset_0 = writeQueue_5_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_5;
  wire              _dataNotInShifter_T_15 = exeResp_5_ready_0 & exeResp_5_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_5 = _dataNotInShifter_T_15 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_6 = waiteStageDeqFire & WillWriteLane[6];
  assign writeQueue_6_enq_valid = _maskedWrite_out_6_valid | dataNotInShifter_readTypeWriteVrf_6;
  assign writeQueue_6_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_vd : 5'h0;
  assign writeQueue_6_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_groupCounter : _maskedWrite_out_6_bits_writeData_groupCounter;
  assign writeQueue_6_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_mask : _maskedWrite_out_6_bits_writeData_mask;
  assign writeQueue_6_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_6 ? writeRequest_6_writeData_data : _maskedWrite_out_6_bits_writeData_data;
  assign writeQueue_6_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_6 & _maskedWrite_out_6_bits_ffoByOther;
  wire [4:0]        exeResp_6_bits_vd_0 = instReg_vd + {1'h0, writeQueue_6_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_6_bits_offset_0 = writeQueue_6_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_6;
  wire              _dataNotInShifter_T_18 = exeResp_6_ready_0 & exeResp_6_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_6 = _dataNotInShifter_T_18 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_7 = waiteStageDeqFire & WillWriteLane[7];
  assign writeQueue_7_enq_valid = _maskedWrite_out_7_valid | dataNotInShifter_readTypeWriteVrf_7;
  assign writeQueue_7_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_vd : 5'h0;
  assign writeQueue_7_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_groupCounter : _maskedWrite_out_7_bits_writeData_groupCounter;
  assign writeQueue_7_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_mask : _maskedWrite_out_7_bits_writeData_mask;
  assign writeQueue_7_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_7 ? writeRequest_7_writeData_data : _maskedWrite_out_7_bits_writeData_data;
  assign writeQueue_7_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_7 & _maskedWrite_out_7_bits_ffoByOther;
  wire [4:0]        exeResp_7_bits_vd_0 = instReg_vd + {1'h0, writeQueue_7_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_7_bits_offset_0 = writeQueue_7_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_7;
  wire              _dataNotInShifter_T_21 = exeResp_7_ready_0 & exeResp_7_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_7 = _dataNotInShifter_T_21 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_8 = waiteStageDeqFire & WillWriteLane[8];
  assign writeQueue_8_enq_valid = _maskedWrite_out_8_valid | dataNotInShifter_readTypeWriteVrf_8;
  assign writeQueue_8_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_vd : 5'h0;
  assign writeQueue_8_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_groupCounter : _maskedWrite_out_8_bits_writeData_groupCounter;
  assign writeQueue_8_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_mask : _maskedWrite_out_8_bits_writeData_mask;
  assign writeQueue_8_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_8 ? writeRequest_8_writeData_data : _maskedWrite_out_8_bits_writeData_data;
  assign writeQueue_8_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_8 & _maskedWrite_out_8_bits_ffoByOther;
  wire [4:0]        exeResp_8_bits_vd_0 = instReg_vd + {1'h0, writeQueue_8_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_8_bits_offset_0 = writeQueue_8_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_8;
  wire              _dataNotInShifter_T_24 = exeResp_8_ready_0 & exeResp_8_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_8 = _dataNotInShifter_T_24 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_9 = waiteStageDeqFire & WillWriteLane[9];
  assign writeQueue_9_enq_valid = _maskedWrite_out_9_valid | dataNotInShifter_readTypeWriteVrf_9;
  assign writeQueue_9_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_vd : 5'h0;
  assign writeQueue_9_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_groupCounter : _maskedWrite_out_9_bits_writeData_groupCounter;
  assign writeQueue_9_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_mask : _maskedWrite_out_9_bits_writeData_mask;
  assign writeQueue_9_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_9 ? writeRequest_9_writeData_data : _maskedWrite_out_9_bits_writeData_data;
  assign writeQueue_9_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_9 & _maskedWrite_out_9_bits_ffoByOther;
  wire [4:0]        exeResp_9_bits_vd_0 = instReg_vd + {1'h0, writeQueue_9_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_9_bits_offset_0 = writeQueue_9_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_9;
  wire              _dataNotInShifter_T_27 = exeResp_9_ready_0 & exeResp_9_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_9 = _dataNotInShifter_T_27 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_10 = waiteStageDeqFire & WillWriteLane[10];
  assign writeQueue_10_enq_valid = _maskedWrite_out_10_valid | dataNotInShifter_readTypeWriteVrf_10;
  assign writeQueue_10_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_vd : 5'h0;
  assign writeQueue_10_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_groupCounter : _maskedWrite_out_10_bits_writeData_groupCounter;
  assign writeQueue_10_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_mask : _maskedWrite_out_10_bits_writeData_mask;
  assign writeQueue_10_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_10 ? writeRequest_10_writeData_data : _maskedWrite_out_10_bits_writeData_data;
  assign writeQueue_10_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_10 & _maskedWrite_out_10_bits_ffoByOther;
  wire [4:0]        exeResp_10_bits_vd_0 = instReg_vd + {1'h0, writeQueue_10_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_10_bits_offset_0 = writeQueue_10_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_10;
  wire              _dataNotInShifter_T_30 = exeResp_10_ready_0 & exeResp_10_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_10 = _dataNotInShifter_T_30 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_11 = waiteStageDeqFire & WillWriteLane[11];
  assign writeQueue_11_enq_valid = _maskedWrite_out_11_valid | dataNotInShifter_readTypeWriteVrf_11;
  assign writeQueue_11_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_vd : 5'h0;
  assign writeQueue_11_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_groupCounter : _maskedWrite_out_11_bits_writeData_groupCounter;
  assign writeQueue_11_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_mask : _maskedWrite_out_11_bits_writeData_mask;
  assign writeQueue_11_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_11 ? writeRequest_11_writeData_data : _maskedWrite_out_11_bits_writeData_data;
  assign writeQueue_11_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_11 & _maskedWrite_out_11_bits_ffoByOther;
  wire [4:0]        exeResp_11_bits_vd_0 = instReg_vd + {1'h0, writeQueue_11_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_11_bits_offset_0 = writeQueue_11_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_11;
  wire              _dataNotInShifter_T_33 = exeResp_11_ready_0 & exeResp_11_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_11 = _dataNotInShifter_T_33 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_12 = waiteStageDeqFire & WillWriteLane[12];
  assign writeQueue_12_enq_valid = _maskedWrite_out_12_valid | dataNotInShifter_readTypeWriteVrf_12;
  assign writeQueue_12_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_vd : 5'h0;
  assign writeQueue_12_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_groupCounter : _maskedWrite_out_12_bits_writeData_groupCounter;
  assign writeQueue_12_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_mask : _maskedWrite_out_12_bits_writeData_mask;
  assign writeQueue_12_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_12 ? writeRequest_12_writeData_data : _maskedWrite_out_12_bits_writeData_data;
  assign writeQueue_12_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_12 & _maskedWrite_out_12_bits_ffoByOther;
  wire [4:0]        exeResp_12_bits_vd_0 = instReg_vd + {1'h0, writeQueue_12_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_12_bits_offset_0 = writeQueue_12_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_12;
  wire              _dataNotInShifter_T_36 = exeResp_12_ready_0 & exeResp_12_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_12 = _dataNotInShifter_T_36 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_13 = waiteStageDeqFire & WillWriteLane[13];
  assign writeQueue_13_enq_valid = _maskedWrite_out_13_valid | dataNotInShifter_readTypeWriteVrf_13;
  assign writeQueue_13_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_vd : 5'h0;
  assign writeQueue_13_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_groupCounter : _maskedWrite_out_13_bits_writeData_groupCounter;
  assign writeQueue_13_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_mask : _maskedWrite_out_13_bits_writeData_mask;
  assign writeQueue_13_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_13 ? writeRequest_13_writeData_data : _maskedWrite_out_13_bits_writeData_data;
  assign writeQueue_13_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_13 & _maskedWrite_out_13_bits_ffoByOther;
  wire [4:0]        exeResp_13_bits_vd_0 = instReg_vd + {1'h0, writeQueue_13_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_13_bits_offset_0 = writeQueue_13_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_13;
  wire              _dataNotInShifter_T_39 = exeResp_13_ready_0 & exeResp_13_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_13 = _dataNotInShifter_T_39 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_14 = waiteStageDeqFire & WillWriteLane[14];
  assign writeQueue_14_enq_valid = _maskedWrite_out_14_valid | dataNotInShifter_readTypeWriteVrf_14;
  assign writeQueue_14_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_vd : 5'h0;
  assign writeQueue_14_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_groupCounter : _maskedWrite_out_14_bits_writeData_groupCounter;
  assign writeQueue_14_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_mask : _maskedWrite_out_14_bits_writeData_mask;
  assign writeQueue_14_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_14 ? writeRequest_14_writeData_data : _maskedWrite_out_14_bits_writeData_data;
  assign writeQueue_14_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_14 & _maskedWrite_out_14_bits_ffoByOther;
  wire [4:0]        exeResp_14_bits_vd_0 = instReg_vd + {1'h0, writeQueue_14_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_14_bits_offset_0 = writeQueue_14_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_14;
  wire              _dataNotInShifter_T_42 = exeResp_14_ready_0 & exeResp_14_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_14 = _dataNotInShifter_T_42 ? 3'h1 : 3'h7;
  wire              dataNotInShifter_readTypeWriteVrf_15 = waiteStageDeqFire & WillWriteLane[15];
  assign writeQueue_15_enq_valid = _maskedWrite_out_15_valid | dataNotInShifter_readTypeWriteVrf_15;
  assign writeQueue_15_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_vd : 5'h0;
  assign writeQueue_15_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_groupCounter : _maskedWrite_out_15_bits_writeData_groupCounter;
  assign writeQueue_15_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_mask : _maskedWrite_out_15_bits_writeData_mask;
  assign writeQueue_15_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_15 ? writeRequest_15_writeData_data : _maskedWrite_out_15_bits_writeData_data;
  assign writeQueue_15_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_15 & _maskedWrite_out_15_bits_ffoByOther;
  wire [4:0]        exeResp_15_bits_vd_0 = instReg_vd + {1'h0, writeQueue_15_deq_bits_writeData_groupCounter[4:1]};
  wire              exeResp_15_bits_offset_0 = writeQueue_15_deq_bits_writeData_groupCounter[0];
  reg  [2:0]        dataNotInShifter_writeTokenCounter_15;
  wire              _dataNotInShifter_T_45 = exeResp_15_ready_0 & exeResp_15_valid_0;
  wire [2:0]        dataNotInShifter_writeTokenChange_15 = _dataNotInShifter_T_45 ? 3'h1 : 3'h7;
  wire              dataNotInShifter =
    dataNotInShifter_writeTokenCounter == 3'h0 & dataNotInShifter_writeTokenCounter_1 == 3'h0 & dataNotInShifter_writeTokenCounter_2 == 3'h0 & dataNotInShifter_writeTokenCounter_3 == 3'h0 & dataNotInShifter_writeTokenCounter_4 == 3'h0
    & dataNotInShifter_writeTokenCounter_5 == 3'h0 & dataNotInShifter_writeTokenCounter_6 == 3'h0 & dataNotInShifter_writeTokenCounter_7 == 3'h0 & dataNotInShifter_writeTokenCounter_8 == 3'h0 & dataNotInShifter_writeTokenCounter_9 == 3'h0
    & dataNotInShifter_writeTokenCounter_10 == 3'h0 & dataNotInShifter_writeTokenCounter_11 == 3'h0 & dataNotInShifter_writeTokenCounter_12 == 3'h0 & dataNotInShifter_writeTokenCounter_13 == 3'h0
    & dataNotInShifter_writeTokenCounter_14 == 3'h0 & dataNotInShifter_writeTokenCounter_15 == 3'h0;
  assign waiteStageDeqReady =
    (~(WillWriteLane[0]) | writeQueue_0_enq_ready) & (~(WillWriteLane[1]) | writeQueue_1_enq_ready) & (~(WillWriteLane[2]) | writeQueue_2_enq_ready) & (~(WillWriteLane[3]) | writeQueue_3_enq_ready)
    & (~(WillWriteLane[4]) | writeQueue_4_enq_ready) & (~(WillWriteLane[5]) | writeQueue_5_enq_ready) & (~(WillWriteLane[6]) | writeQueue_6_enq_ready) & (~(WillWriteLane[7]) | writeQueue_7_enq_ready)
    & (~(WillWriteLane[8]) | writeQueue_8_enq_ready) & (~(WillWriteLane[9]) | writeQueue_9_enq_ready) & (~(WillWriteLane[10]) | writeQueue_10_enq_ready) & (~(WillWriteLane[11]) | writeQueue_11_enq_ready)
    & (~(WillWriteLane[12]) | writeQueue_12_enq_ready) & (~(WillWriteLane[13]) | writeQueue_13_enq_ready) & (~(WillWriteLane[14]) | writeQueue_14_enq_ready) & (~(WillWriteLane[15]) | writeQueue_15_enq_ready);
  reg               waiteLastRequest;
  reg               waitQueueClear;
  wire              lastReportValid =
    waitQueueClear
    & ~(writeQueue_0_deq_valid | writeQueue_1_deq_valid | writeQueue_2_deq_valid | writeQueue_3_deq_valid | writeQueue_4_deq_valid | writeQueue_5_deq_valid | writeQueue_6_deq_valid | writeQueue_7_deq_valid | writeQueue_8_deq_valid
        | writeQueue_9_deq_valid | writeQueue_10_deq_valid | writeQueue_11_deq_valid | writeQueue_12_deq_valid | writeQueue_13_deq_valid | writeQueue_14_deq_valid | writeQueue_15_deq_valid) & dataNotInShifter;
  wire              executeStageInvalid = unitType[1] & ~compressUnitResultQueue_deq_valid & ~_compressUnit_stageValid | unitType[2] & _reduceUnit_in_ready | unitType[3];
  wire              executeStageClean = readType ? waiteStageDeqFire & waiteReadDataPipeReg_last : waiteLastRequest & _maskedWrite_stageClear & executeStageInvalid;
  wire              invalidEnq = instReq_valid & instReq_bits_vl == 11'h0 & ~enqMvRD;
  wire [7:0]        _lastReport_output = lastReportValid ? 8'h1 << instReg_instructionIndex : 8'h0;
  wire [31:0]       gatherData_bits_0 = readVS1Reg_dataValid ? readVS1Reg_data : 32'h0;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      gatherReadState <= 2'h0;
      gatherDatOffset <= 2'h0;
      gatherLane <= 4'h0;
      gatherOffset <= 1'h0;
      gatherGrowth <= 3'h0;
      instReg_instructionIndex <= 3'h0;
      instReg_decodeResult_orderReduce <= 1'h0;
      instReg_decodeResult_floatMul <= 1'h0;
      instReg_decodeResult_fpExecutionType <= 2'h0;
      instReg_decodeResult_float <= 1'h0;
      instReg_decodeResult_specialSlot <= 1'h0;
      instReg_decodeResult_topUop <= 5'h0;
      instReg_decodeResult_popCount <= 1'h0;
      instReg_decodeResult_ffo <= 1'h0;
      instReg_decodeResult_average <= 1'h0;
      instReg_decodeResult_reverse <= 1'h0;
      instReg_decodeResult_dontNeedExecuteInLane <= 1'h0;
      instReg_decodeResult_scheduler <= 1'h0;
      instReg_decodeResult_sReadVD <= 1'h0;
      instReg_decodeResult_vtype <= 1'h0;
      instReg_decodeResult_sWrite <= 1'h0;
      instReg_decodeResult_crossRead <= 1'h0;
      instReg_decodeResult_crossWrite <= 1'h0;
      instReg_decodeResult_maskUnit <= 1'h0;
      instReg_decodeResult_special <= 1'h0;
      instReg_decodeResult_saturate <= 1'h0;
      instReg_decodeResult_vwmacc <= 1'h0;
      instReg_decodeResult_readOnly <= 1'h0;
      instReg_decodeResult_maskSource <= 1'h0;
      instReg_decodeResult_maskDestination <= 1'h0;
      instReg_decodeResult_maskLogic <= 1'h0;
      instReg_decodeResult_uop <= 4'h0;
      instReg_decodeResult_iota <= 1'h0;
      instReg_decodeResult_mv <= 1'h0;
      instReg_decodeResult_extend <= 1'h0;
      instReg_decodeResult_unOrderWrite <= 1'h0;
      instReg_decodeResult_compress <= 1'h0;
      instReg_decodeResult_gather16 <= 1'h0;
      instReg_decodeResult_gather <= 1'h0;
      instReg_decodeResult_slid <= 1'h0;
      instReg_decodeResult_targetRd <= 1'h0;
      instReg_decodeResult_widenReduce <= 1'h0;
      instReg_decodeResult_red <= 1'h0;
      instReg_decodeResult_nr <= 1'h0;
      instReg_decodeResult_itype <= 1'h0;
      instReg_decodeResult_unsigned1 <= 1'h0;
      instReg_decodeResult_unsigned0 <= 1'h0;
      instReg_decodeResult_other <= 1'h0;
      instReg_decodeResult_multiCycle <= 1'h0;
      instReg_decodeResult_divider <= 1'h0;
      instReg_decodeResult_multiplier <= 1'h0;
      instReg_decodeResult_shift <= 1'h0;
      instReg_decodeResult_adder <= 1'h0;
      instReg_decodeResult_logic <= 1'h0;
      instReg_readFromScala <= 32'h0;
      instReg_sew <= 2'h0;
      instReg_vlmul <= 3'h0;
      instReg_maskType <= 1'h0;
      instReg_vxrm <= 3'h0;
      instReg_vs2 <= 5'h0;
      instReg_vs1 <= 5'h0;
      instReg_vd <= 5'h0;
      instReg_vl <= 11'h0;
      instVlValid <= 1'h0;
      readVS1Reg_dataValid <= 1'h0;
      readVS1Reg_requestSend <= 1'h0;
      readVS1Reg_sendToExecution <= 1'h0;
      readVS1Reg_data <= 32'h0;
      readVS1Reg_readIndex <= 4'h0;
      exeReqReg_0_valid <= 1'h0;
      exeReqReg_0_bits_source1 <= 32'h0;
      exeReqReg_0_bits_source2 <= 32'h0;
      exeReqReg_0_bits_index <= 3'h0;
      exeReqReg_0_bits_ffo <= 1'h0;
      exeReqReg_0_bits_fpReduceValid <= 1'h0;
      exeReqReg_1_valid <= 1'h0;
      exeReqReg_1_bits_source1 <= 32'h0;
      exeReqReg_1_bits_source2 <= 32'h0;
      exeReqReg_1_bits_index <= 3'h0;
      exeReqReg_1_bits_ffo <= 1'h0;
      exeReqReg_1_bits_fpReduceValid <= 1'h0;
      exeReqReg_2_valid <= 1'h0;
      exeReqReg_2_bits_source1 <= 32'h0;
      exeReqReg_2_bits_source2 <= 32'h0;
      exeReqReg_2_bits_index <= 3'h0;
      exeReqReg_2_bits_ffo <= 1'h0;
      exeReqReg_2_bits_fpReduceValid <= 1'h0;
      exeReqReg_3_valid <= 1'h0;
      exeReqReg_3_bits_source1 <= 32'h0;
      exeReqReg_3_bits_source2 <= 32'h0;
      exeReqReg_3_bits_index <= 3'h0;
      exeReqReg_3_bits_ffo <= 1'h0;
      exeReqReg_3_bits_fpReduceValid <= 1'h0;
      exeReqReg_4_valid <= 1'h0;
      exeReqReg_4_bits_source1 <= 32'h0;
      exeReqReg_4_bits_source2 <= 32'h0;
      exeReqReg_4_bits_index <= 3'h0;
      exeReqReg_4_bits_ffo <= 1'h0;
      exeReqReg_4_bits_fpReduceValid <= 1'h0;
      exeReqReg_5_valid <= 1'h0;
      exeReqReg_5_bits_source1 <= 32'h0;
      exeReqReg_5_bits_source2 <= 32'h0;
      exeReqReg_5_bits_index <= 3'h0;
      exeReqReg_5_bits_ffo <= 1'h0;
      exeReqReg_5_bits_fpReduceValid <= 1'h0;
      exeReqReg_6_valid <= 1'h0;
      exeReqReg_6_bits_source1 <= 32'h0;
      exeReqReg_6_bits_source2 <= 32'h0;
      exeReqReg_6_bits_index <= 3'h0;
      exeReqReg_6_bits_ffo <= 1'h0;
      exeReqReg_6_bits_fpReduceValid <= 1'h0;
      exeReqReg_7_valid <= 1'h0;
      exeReqReg_7_bits_source1 <= 32'h0;
      exeReqReg_7_bits_source2 <= 32'h0;
      exeReqReg_7_bits_index <= 3'h0;
      exeReqReg_7_bits_ffo <= 1'h0;
      exeReqReg_7_bits_fpReduceValid <= 1'h0;
      exeReqReg_8_valid <= 1'h0;
      exeReqReg_8_bits_source1 <= 32'h0;
      exeReqReg_8_bits_source2 <= 32'h0;
      exeReqReg_8_bits_index <= 3'h0;
      exeReqReg_8_bits_ffo <= 1'h0;
      exeReqReg_8_bits_fpReduceValid <= 1'h0;
      exeReqReg_9_valid <= 1'h0;
      exeReqReg_9_bits_source1 <= 32'h0;
      exeReqReg_9_bits_source2 <= 32'h0;
      exeReqReg_9_bits_index <= 3'h0;
      exeReqReg_9_bits_ffo <= 1'h0;
      exeReqReg_9_bits_fpReduceValid <= 1'h0;
      exeReqReg_10_valid <= 1'h0;
      exeReqReg_10_bits_source1 <= 32'h0;
      exeReqReg_10_bits_source2 <= 32'h0;
      exeReqReg_10_bits_index <= 3'h0;
      exeReqReg_10_bits_ffo <= 1'h0;
      exeReqReg_10_bits_fpReduceValid <= 1'h0;
      exeReqReg_11_valid <= 1'h0;
      exeReqReg_11_bits_source1 <= 32'h0;
      exeReqReg_11_bits_source2 <= 32'h0;
      exeReqReg_11_bits_index <= 3'h0;
      exeReqReg_11_bits_ffo <= 1'h0;
      exeReqReg_11_bits_fpReduceValid <= 1'h0;
      exeReqReg_12_valid <= 1'h0;
      exeReqReg_12_bits_source1 <= 32'h0;
      exeReqReg_12_bits_source2 <= 32'h0;
      exeReqReg_12_bits_index <= 3'h0;
      exeReqReg_12_bits_ffo <= 1'h0;
      exeReqReg_12_bits_fpReduceValid <= 1'h0;
      exeReqReg_13_valid <= 1'h0;
      exeReqReg_13_bits_source1 <= 32'h0;
      exeReqReg_13_bits_source2 <= 32'h0;
      exeReqReg_13_bits_index <= 3'h0;
      exeReqReg_13_bits_ffo <= 1'h0;
      exeReqReg_13_bits_fpReduceValid <= 1'h0;
      exeReqReg_14_valid <= 1'h0;
      exeReqReg_14_bits_source1 <= 32'h0;
      exeReqReg_14_bits_source2 <= 32'h0;
      exeReqReg_14_bits_index <= 3'h0;
      exeReqReg_14_bits_ffo <= 1'h0;
      exeReqReg_14_bits_fpReduceValid <= 1'h0;
      exeReqReg_15_valid <= 1'h0;
      exeReqReg_15_bits_source1 <= 32'h0;
      exeReqReg_15_bits_source2 <= 32'h0;
      exeReqReg_15_bits_index <= 3'h0;
      exeReqReg_15_bits_ffo <= 1'h0;
      exeReqReg_15_bits_fpReduceValid <= 1'h0;
      requestCounter <= 5'h0;
      executeIndex <= 2'h0;
      readIssueStageState_groupReadState <= 16'h0;
      readIssueStageState_needRead <= 16'h0;
      readIssueStageState_elementValid <= 16'h0;
      readIssueStageState_replaceVs1 <= 16'h0;
      readIssueStageState_readOffset <= 16'h0;
      readIssueStageState_accessLane_0 <= 4'h0;
      readIssueStageState_accessLane_1 <= 4'h0;
      readIssueStageState_accessLane_2 <= 4'h0;
      readIssueStageState_accessLane_3 <= 4'h0;
      readIssueStageState_accessLane_4 <= 4'h0;
      readIssueStageState_accessLane_5 <= 4'h0;
      readIssueStageState_accessLane_6 <= 4'h0;
      readIssueStageState_accessLane_7 <= 4'h0;
      readIssueStageState_accessLane_8 <= 4'h0;
      readIssueStageState_accessLane_9 <= 4'h0;
      readIssueStageState_accessLane_10 <= 4'h0;
      readIssueStageState_accessLane_11 <= 4'h0;
      readIssueStageState_accessLane_12 <= 4'h0;
      readIssueStageState_accessLane_13 <= 4'h0;
      readIssueStageState_accessLane_14 <= 4'h0;
      readIssueStageState_accessLane_15 <= 4'h0;
      readIssueStageState_vsGrowth_0 <= 3'h0;
      readIssueStageState_vsGrowth_1 <= 3'h0;
      readIssueStageState_vsGrowth_2 <= 3'h0;
      readIssueStageState_vsGrowth_3 <= 3'h0;
      readIssueStageState_vsGrowth_4 <= 3'h0;
      readIssueStageState_vsGrowth_5 <= 3'h0;
      readIssueStageState_vsGrowth_6 <= 3'h0;
      readIssueStageState_vsGrowth_7 <= 3'h0;
      readIssueStageState_vsGrowth_8 <= 3'h0;
      readIssueStageState_vsGrowth_9 <= 3'h0;
      readIssueStageState_vsGrowth_10 <= 3'h0;
      readIssueStageState_vsGrowth_11 <= 3'h0;
      readIssueStageState_vsGrowth_12 <= 3'h0;
      readIssueStageState_vsGrowth_13 <= 3'h0;
      readIssueStageState_vsGrowth_14 <= 3'h0;
      readIssueStageState_vsGrowth_15 <= 3'h0;
      readIssueStageState_executeGroup <= 7'h0;
      readIssueStageState_readDataOffset <= 32'h0;
      readIssueStageState_last <= 1'h0;
      readIssueStageValid <= 1'h0;
      tokenCheck_counter <= 4'h0;
      tokenCheck_counter_1 <= 4'h0;
      tokenCheck_counter_2 <= 4'h0;
      tokenCheck_counter_3 <= 4'h0;
      tokenCheck_counter_4 <= 4'h0;
      tokenCheck_counter_5 <= 4'h0;
      tokenCheck_counter_6 <= 4'h0;
      tokenCheck_counter_7 <= 4'h0;
      tokenCheck_counter_8 <= 4'h0;
      tokenCheck_counter_9 <= 4'h0;
      tokenCheck_counter_10 <= 4'h0;
      tokenCheck_counter_11 <= 4'h0;
      tokenCheck_counter_12 <= 4'h0;
      tokenCheck_counter_13 <= 4'h0;
      tokenCheck_counter_14 <= 4'h0;
      tokenCheck_counter_15 <= 4'h0;
      reorderQueueAllocate_counter <= 6'h0;
      reorderQueueAllocate_counterWillUpdate <= 6'h0;
      reorderQueueAllocate_counter_1 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_1 <= 6'h0;
      reorderQueueAllocate_counter_2 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_2 <= 6'h0;
      reorderQueueAllocate_counter_3 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_3 <= 6'h0;
      reorderQueueAllocate_counter_4 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_4 <= 6'h0;
      reorderQueueAllocate_counter_5 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_5 <= 6'h0;
      reorderQueueAllocate_counter_6 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_6 <= 6'h0;
      reorderQueueAllocate_counter_7 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_7 <= 6'h0;
      reorderQueueAllocate_counter_8 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_8 <= 6'h0;
      reorderQueueAllocate_counter_9 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_9 <= 6'h0;
      reorderQueueAllocate_counter_10 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_10 <= 6'h0;
      reorderQueueAllocate_counter_11 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_11 <= 6'h0;
      reorderQueueAllocate_counter_12 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_12 <= 6'h0;
      reorderQueueAllocate_counter_13 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_13 <= 6'h0;
      reorderQueueAllocate_counter_14 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_14 <= 6'h0;
      reorderQueueAllocate_counter_15 <= 6'h0;
      reorderQueueAllocate_counterWillUpdate_15 <= 6'h0;
      reorderStageValid <= 1'h0;
      reorderStageState_0 <= 5'h0;
      reorderStageState_1 <= 5'h0;
      reorderStageState_2 <= 5'h0;
      reorderStageState_3 <= 5'h0;
      reorderStageState_4 <= 5'h0;
      reorderStageState_5 <= 5'h0;
      reorderStageState_6 <= 5'h0;
      reorderStageState_7 <= 5'h0;
      reorderStageState_8 <= 5'h0;
      reorderStageState_9 <= 5'h0;
      reorderStageState_10 <= 5'h0;
      reorderStageState_11 <= 5'h0;
      reorderStageState_12 <= 5'h0;
      reorderStageState_13 <= 5'h0;
      reorderStageState_14 <= 5'h0;
      reorderStageState_15 <= 5'h0;
      reorderStageNeed_0 <= 5'h0;
      reorderStageNeed_1 <= 5'h0;
      reorderStageNeed_2 <= 5'h0;
      reorderStageNeed_3 <= 5'h0;
      reorderStageNeed_4 <= 5'h0;
      reorderStageNeed_5 <= 5'h0;
      reorderStageNeed_6 <= 5'h0;
      reorderStageNeed_7 <= 5'h0;
      reorderStageNeed_8 <= 5'h0;
      reorderStageNeed_9 <= 5'h0;
      reorderStageNeed_10 <= 5'h0;
      reorderStageNeed_11 <= 5'h0;
      reorderStageNeed_12 <= 5'h0;
      reorderStageNeed_13 <= 5'h0;
      reorderStageNeed_14 <= 5'h0;
      reorderStageNeed_15 <= 5'h0;
      waiteReadDataPipeReg_executeGroup <= 7'h0;
      waiteReadDataPipeReg_sourceValid <= 16'h0;
      waiteReadDataPipeReg_replaceVs1 <= 16'h0;
      waiteReadDataPipeReg_needRead <= 16'h0;
      waiteReadDataPipeReg_last <= 1'h0;
      waiteReadData_0 <= 32'h0;
      waiteReadData_1 <= 32'h0;
      waiteReadData_2 <= 32'h0;
      waiteReadData_3 <= 32'h0;
      waiteReadData_4 <= 32'h0;
      waiteReadData_5 <= 32'h0;
      waiteReadData_6 <= 32'h0;
      waiteReadData_7 <= 32'h0;
      waiteReadData_8 <= 32'h0;
      waiteReadData_9 <= 32'h0;
      waiteReadData_10 <= 32'h0;
      waiteReadData_11 <= 32'h0;
      waiteReadData_12 <= 32'h0;
      waiteReadData_13 <= 32'h0;
      waiteReadData_14 <= 32'h0;
      waiteReadData_15 <= 32'h0;
      waiteReadSate <= 16'h0;
      waiteReadStageValid <= 1'h0;
      dataNotInShifter_writeTokenCounter <= 3'h0;
      dataNotInShifter_writeTokenCounter_1 <= 3'h0;
      dataNotInShifter_writeTokenCounter_2 <= 3'h0;
      dataNotInShifter_writeTokenCounter_3 <= 3'h0;
      dataNotInShifter_writeTokenCounter_4 <= 3'h0;
      dataNotInShifter_writeTokenCounter_5 <= 3'h0;
      dataNotInShifter_writeTokenCounter_6 <= 3'h0;
      dataNotInShifter_writeTokenCounter_7 <= 3'h0;
      dataNotInShifter_writeTokenCounter_8 <= 3'h0;
      dataNotInShifter_writeTokenCounter_9 <= 3'h0;
      dataNotInShifter_writeTokenCounter_10 <= 3'h0;
      dataNotInShifter_writeTokenCounter_11 <= 3'h0;
      dataNotInShifter_writeTokenCounter_12 <= 3'h0;
      dataNotInShifter_writeTokenCounter_13 <= 3'h0;
      dataNotInShifter_writeTokenCounter_14 <= 3'h0;
      dataNotInShifter_writeTokenCounter_15 <= 3'h0;
      waiteLastRequest <= 1'h0;
      waitQueueClear <= 1'h0;
    end
    else begin
      automatic logic _GEN_106 = instReq_valid & (viotaReq | enqMvRD) | gatherRequestFire;
      automatic logic _GEN_107;
      automatic logic _GEN_108 = source1Change & viotaCounterAdd;
      _GEN_107 = instReq_valid | gatherRequestFire;
      if (v0UpdateVec_0_valid & ~v0UpdateVec_0_bits_offset)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & ~v0UpdateVec_1_bits_offset)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & ~v0UpdateVec_2_bits_offset)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & ~v0UpdateVec_3_bits_offset)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & ~v0UpdateVec_4_bits_offset)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & ~v0UpdateVec_5_bits_offset)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & ~v0UpdateVec_6_bits_offset)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & ~v0UpdateVec_7_bits_offset)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & ~v0UpdateVec_8_bits_offset)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & ~v0UpdateVec_9_bits_offset)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & ~v0UpdateVec_10_bits_offset)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & ~v0UpdateVec_11_bits_offset)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & ~v0UpdateVec_12_bits_offset)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & ~v0UpdateVec_13_bits_offset)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & ~v0UpdateVec_14_bits_offset)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & ~v0UpdateVec_15_bits_offset)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_15_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_4_valid & v0UpdateVec_4_bits_offset)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_4_bits_data;
      if (v0UpdateVec_5_valid & v0UpdateVec_5_bits_offset)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_5_bits_data;
      if (v0UpdateVec_6_valid & v0UpdateVec_6_bits_offset)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_6_bits_data;
      if (v0UpdateVec_7_valid & v0UpdateVec_7_bits_offset)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_7_bits_data;
      if (v0UpdateVec_8_valid & v0UpdateVec_8_bits_offset)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_8_bits_data;
      if (v0UpdateVec_9_valid & v0UpdateVec_9_bits_offset)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_9_bits_data;
      if (v0UpdateVec_10_valid & v0UpdateVec_10_bits_offset)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_10_bits_data;
      if (v0UpdateVec_11_valid & v0UpdateVec_11_bits_offset)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_11_bits_data;
      if (v0UpdateVec_12_valid & v0UpdateVec_12_bits_offset)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_12_bits_data;
      if (v0UpdateVec_13_valid & v0UpdateVec_13_bits_offset)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_13_bits_data;
      if (v0UpdateVec_14_valid & v0UpdateVec_14_bits_offset)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_14_bits_data;
      if (v0UpdateVec_15_valid & v0UpdateVec_15_bits_offset)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_15_bits_data;
      if (gatherData_ready_0 & gatherData_valid_0)
        gatherReadState <= 2'h0;
      else if (_tokenCheck_T & gatherSRead)
        gatherReadState <= 2'h2;
      else if (gatherRequestFire)
        gatherReadState <= {notNeedRead, 1'h1};
      else if (readTokenRelease_0 & gatherWaiteRead)
        gatherReadState <= 2'h3;
      if (gatherRequestFire) begin
        gatherDatOffset <= dataOffset;
        gatherLane <= accessLane;
        gatherOffset <= offset;
        gatherGrowth <= reallyGrowth;
      end
      if (_GEN_106 | instReq_valid)
        instReg_instructionIndex <= instReq_bits_instructionIndex;
      if (instReq_valid) begin
        instReg_decodeResult_orderReduce <= instReq_bits_decodeResult_orderReduce;
        instReg_decodeResult_floatMul <= instReq_bits_decodeResult_floatMul;
        instReg_decodeResult_fpExecutionType <= instReq_bits_decodeResult_fpExecutionType;
        instReg_decodeResult_float <= instReq_bits_decodeResult_float;
        instReg_decodeResult_specialSlot <= instReq_bits_decodeResult_specialSlot;
        instReg_decodeResult_topUop <= instReq_bits_decodeResult_topUop;
        instReg_decodeResult_popCount <= instReq_bits_decodeResult_popCount;
        instReg_decodeResult_ffo <= instReq_bits_decodeResult_ffo;
        instReg_decodeResult_average <= instReq_bits_decodeResult_average;
        instReg_decodeResult_reverse <= instReq_bits_decodeResult_reverse;
        instReg_decodeResult_dontNeedExecuteInLane <= instReq_bits_decodeResult_dontNeedExecuteInLane;
        instReg_decodeResult_scheduler <= instReq_bits_decodeResult_scheduler;
        instReg_decodeResult_sReadVD <= instReq_bits_decodeResult_sReadVD;
        instReg_decodeResult_vtype <= instReq_bits_decodeResult_vtype;
        instReg_decodeResult_sWrite <= instReq_bits_decodeResult_sWrite;
        instReg_decodeResult_crossRead <= instReq_bits_decodeResult_crossRead;
        instReg_decodeResult_crossWrite <= instReq_bits_decodeResult_crossWrite;
        instReg_decodeResult_maskUnit <= instReq_bits_decodeResult_maskUnit;
        instReg_decodeResult_special <= instReq_bits_decodeResult_special;
        instReg_decodeResult_saturate <= instReq_bits_decodeResult_saturate;
        instReg_decodeResult_vwmacc <= instReq_bits_decodeResult_vwmacc;
        instReg_decodeResult_readOnly <= instReq_bits_decodeResult_readOnly;
        instReg_decodeResult_maskSource <= instReq_bits_decodeResult_maskSource;
        instReg_decodeResult_maskDestination <= instReq_bits_decodeResult_maskDestination;
        instReg_decodeResult_maskLogic <= instReq_bits_decodeResult_maskLogic;
        instReg_decodeResult_uop <= instReq_bits_decodeResult_uop;
        instReg_decodeResult_iota <= instReq_bits_decodeResult_iota;
        instReg_decodeResult_mv <= instReq_bits_decodeResult_mv;
        instReg_decodeResult_extend <= instReq_bits_decodeResult_extend;
        instReg_decodeResult_unOrderWrite <= instReq_bits_decodeResult_unOrderWrite;
        instReg_decodeResult_compress <= instReq_bits_decodeResult_compress;
        instReg_decodeResult_gather16 <= instReq_bits_decodeResult_gather16;
        instReg_decodeResult_gather <= instReq_bits_decodeResult_gather;
        instReg_decodeResult_slid <= instReq_bits_decodeResult_slid;
        instReg_decodeResult_targetRd <= instReq_bits_decodeResult_targetRd;
        instReg_decodeResult_widenReduce <= instReq_bits_decodeResult_widenReduce;
        instReg_decodeResult_red <= instReq_bits_decodeResult_red;
        instReg_decodeResult_nr <= instReq_bits_decodeResult_nr;
        instReg_decodeResult_itype <= instReq_bits_decodeResult_itype;
        instReg_decodeResult_unsigned1 <= instReq_bits_decodeResult_unsigned1;
        instReg_decodeResult_unsigned0 <= instReq_bits_decodeResult_unsigned0;
        instReg_decodeResult_other <= instReq_bits_decodeResult_other;
        instReg_decodeResult_multiCycle <= instReq_bits_decodeResult_multiCycle;
        instReg_decodeResult_divider <= instReq_bits_decodeResult_divider;
        instReg_decodeResult_multiplier <= instReq_bits_decodeResult_multiplier;
        instReg_decodeResult_shift <= instReq_bits_decodeResult_shift;
        instReg_decodeResult_adder <= instReq_bits_decodeResult_adder;
        instReg_decodeResult_logic <= instReq_bits_decodeResult_logic;
        instReg_readFromScala <= instReq_bits_readFromScala;
        instReg_sew <= instReq_bits_sew;
        instReg_vlmul <= instReq_bits_vlmul;
        instReg_maskType <= instReq_bits_maskType;
        instReg_vxrm <= instReq_bits_vxrm;
        instReg_vs2 <= instReq_bits_vs2;
        instReg_vd <= instReq_bits_vd;
        instReg_vl <= instReq_bits_vl;
      end
      if (_GEN_106)
        instReg_vs1 <= instReq_bits_vs2;
      else if (instReq_valid)
        instReg_vs1 <= instReq_bits_vs1;
      if (|{instReq_valid, _lastReport_output})
        instVlValid <= ((|instReq_bits_vl) | enqMvRD) & instReq_valid;
      readVS1Reg_dataValid <= ~_GEN_108 & (readTokenRelease_0 | ~_GEN_107 & readVS1Reg_dataValid);
      readVS1Reg_requestSend <= ~_GEN_108 & (_tokenCheck_T | ~_GEN_107 & readVS1Reg_requestSend);
      readVS1Reg_sendToExecution <= _view__firstGroup_T_1 | viotaCounterAdd | ~_GEN_107 & readVS1Reg_sendToExecution;
      if (readTokenRelease_0) begin
        readVS1Reg_data <= readData_readDataQueue_deq_bits;
        waiteReadData_0 <= readData_readDataQueue_deq_bits;
      end
      if (_GEN_108)
        readVS1Reg_readIndex <= readVS1Reg_readIndex + 4'h1;
      else if (_GEN_107)
        readVS1Reg_readIndex <= 4'h0;
      if (tokenIO_0_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_0_valid <= tokenIO_0_maskRequestRelease_0 & ~viota;
      if (tokenIO_0_maskRequestRelease_0) begin
        exeReqReg_0_bits_source1 <= exeRequestQueue_0_deq_bits_source1;
        exeReqReg_0_bits_source2 <= exeRequestQueue_0_deq_bits_source2;
        exeReqReg_0_bits_index <= exeRequestQueue_0_deq_bits_index;
        exeReqReg_0_bits_ffo <= exeRequestQueue_0_deq_bits_ffo;
        exeReqReg_0_bits_fpReduceValid <= exeRequestQueue_0_deq_bits_fpReduceValid;
      end
      if (tokenIO_1_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_1_valid <= tokenIO_1_maskRequestRelease_0 & ~viota;
      if (tokenIO_1_maskRequestRelease_0) begin
        exeReqReg_1_bits_source1 <= exeRequestQueue_1_deq_bits_source1;
        exeReqReg_1_bits_source2 <= exeRequestQueue_1_deq_bits_source2;
        exeReqReg_1_bits_index <= exeRequestQueue_1_deq_bits_index;
        exeReqReg_1_bits_ffo <= exeRequestQueue_1_deq_bits_ffo;
        exeReqReg_1_bits_fpReduceValid <= exeRequestQueue_1_deq_bits_fpReduceValid;
      end
      if (tokenIO_2_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_2_valid <= tokenIO_2_maskRequestRelease_0 & ~viota;
      if (tokenIO_2_maskRequestRelease_0) begin
        exeReqReg_2_bits_source1 <= exeRequestQueue_2_deq_bits_source1;
        exeReqReg_2_bits_source2 <= exeRequestQueue_2_deq_bits_source2;
        exeReqReg_2_bits_index <= exeRequestQueue_2_deq_bits_index;
        exeReqReg_2_bits_ffo <= exeRequestQueue_2_deq_bits_ffo;
        exeReqReg_2_bits_fpReduceValid <= exeRequestQueue_2_deq_bits_fpReduceValid;
      end
      if (tokenIO_3_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_3_valid <= tokenIO_3_maskRequestRelease_0 & ~viota;
      if (tokenIO_3_maskRequestRelease_0) begin
        exeReqReg_3_bits_source1 <= exeRequestQueue_3_deq_bits_source1;
        exeReqReg_3_bits_source2 <= exeRequestQueue_3_deq_bits_source2;
        exeReqReg_3_bits_index <= exeRequestQueue_3_deq_bits_index;
        exeReqReg_3_bits_ffo <= exeRequestQueue_3_deq_bits_ffo;
        exeReqReg_3_bits_fpReduceValid <= exeRequestQueue_3_deq_bits_fpReduceValid;
      end
      if (tokenIO_4_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_4_valid <= tokenIO_4_maskRequestRelease_0 & ~viota;
      if (tokenIO_4_maskRequestRelease_0) begin
        exeReqReg_4_bits_source1 <= exeRequestQueue_4_deq_bits_source1;
        exeReqReg_4_bits_source2 <= exeRequestQueue_4_deq_bits_source2;
        exeReqReg_4_bits_index <= exeRequestQueue_4_deq_bits_index;
        exeReqReg_4_bits_ffo <= exeRequestQueue_4_deq_bits_ffo;
        exeReqReg_4_bits_fpReduceValid <= exeRequestQueue_4_deq_bits_fpReduceValid;
      end
      if (tokenIO_5_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_5_valid <= tokenIO_5_maskRequestRelease_0 & ~viota;
      if (tokenIO_5_maskRequestRelease_0) begin
        exeReqReg_5_bits_source1 <= exeRequestQueue_5_deq_bits_source1;
        exeReqReg_5_bits_source2 <= exeRequestQueue_5_deq_bits_source2;
        exeReqReg_5_bits_index <= exeRequestQueue_5_deq_bits_index;
        exeReqReg_5_bits_ffo <= exeRequestQueue_5_deq_bits_ffo;
        exeReqReg_5_bits_fpReduceValid <= exeRequestQueue_5_deq_bits_fpReduceValid;
      end
      if (tokenIO_6_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_6_valid <= tokenIO_6_maskRequestRelease_0 & ~viota;
      if (tokenIO_6_maskRequestRelease_0) begin
        exeReqReg_6_bits_source1 <= exeRequestQueue_6_deq_bits_source1;
        exeReqReg_6_bits_source2 <= exeRequestQueue_6_deq_bits_source2;
        exeReqReg_6_bits_index <= exeRequestQueue_6_deq_bits_index;
        exeReqReg_6_bits_ffo <= exeRequestQueue_6_deq_bits_ffo;
        exeReqReg_6_bits_fpReduceValid <= exeRequestQueue_6_deq_bits_fpReduceValid;
      end
      if (tokenIO_7_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_7_valid <= tokenIO_7_maskRequestRelease_0 & ~viota;
      if (tokenIO_7_maskRequestRelease_0) begin
        exeReqReg_7_bits_source1 <= exeRequestQueue_7_deq_bits_source1;
        exeReqReg_7_bits_source2 <= exeRequestQueue_7_deq_bits_source2;
        exeReqReg_7_bits_index <= exeRequestQueue_7_deq_bits_index;
        exeReqReg_7_bits_ffo <= exeRequestQueue_7_deq_bits_ffo;
        exeReqReg_7_bits_fpReduceValid <= exeRequestQueue_7_deq_bits_fpReduceValid;
      end
      if (tokenIO_8_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_8_valid <= tokenIO_8_maskRequestRelease_0 & ~viota;
      if (tokenIO_8_maskRequestRelease_0) begin
        exeReqReg_8_bits_source1 <= exeRequestQueue_8_deq_bits_source1;
        exeReqReg_8_bits_source2 <= exeRequestQueue_8_deq_bits_source2;
        exeReqReg_8_bits_index <= exeRequestQueue_8_deq_bits_index;
        exeReqReg_8_bits_ffo <= exeRequestQueue_8_deq_bits_ffo;
        exeReqReg_8_bits_fpReduceValid <= exeRequestQueue_8_deq_bits_fpReduceValid;
      end
      if (tokenIO_9_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_9_valid <= tokenIO_9_maskRequestRelease_0 & ~viota;
      if (tokenIO_9_maskRequestRelease_0) begin
        exeReqReg_9_bits_source1 <= exeRequestQueue_9_deq_bits_source1;
        exeReqReg_9_bits_source2 <= exeRequestQueue_9_deq_bits_source2;
        exeReqReg_9_bits_index <= exeRequestQueue_9_deq_bits_index;
        exeReqReg_9_bits_ffo <= exeRequestQueue_9_deq_bits_ffo;
        exeReqReg_9_bits_fpReduceValid <= exeRequestQueue_9_deq_bits_fpReduceValid;
      end
      if (tokenIO_10_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_10_valid <= tokenIO_10_maskRequestRelease_0 & ~viota;
      if (tokenIO_10_maskRequestRelease_0) begin
        exeReqReg_10_bits_source1 <= exeRequestQueue_10_deq_bits_source1;
        exeReqReg_10_bits_source2 <= exeRequestQueue_10_deq_bits_source2;
        exeReqReg_10_bits_index <= exeRequestQueue_10_deq_bits_index;
        exeReqReg_10_bits_ffo <= exeRequestQueue_10_deq_bits_ffo;
        exeReqReg_10_bits_fpReduceValid <= exeRequestQueue_10_deq_bits_fpReduceValid;
      end
      if (tokenIO_11_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_11_valid <= tokenIO_11_maskRequestRelease_0 & ~viota;
      if (tokenIO_11_maskRequestRelease_0) begin
        exeReqReg_11_bits_source1 <= exeRequestQueue_11_deq_bits_source1;
        exeReqReg_11_bits_source2 <= exeRequestQueue_11_deq_bits_source2;
        exeReqReg_11_bits_index <= exeRequestQueue_11_deq_bits_index;
        exeReqReg_11_bits_ffo <= exeRequestQueue_11_deq_bits_ffo;
        exeReqReg_11_bits_fpReduceValid <= exeRequestQueue_11_deq_bits_fpReduceValid;
      end
      if (tokenIO_12_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_12_valid <= tokenIO_12_maskRequestRelease_0 & ~viota;
      if (tokenIO_12_maskRequestRelease_0) begin
        exeReqReg_12_bits_source1 <= exeRequestQueue_12_deq_bits_source1;
        exeReqReg_12_bits_source2 <= exeRequestQueue_12_deq_bits_source2;
        exeReqReg_12_bits_index <= exeRequestQueue_12_deq_bits_index;
        exeReqReg_12_bits_ffo <= exeRequestQueue_12_deq_bits_ffo;
        exeReqReg_12_bits_fpReduceValid <= exeRequestQueue_12_deq_bits_fpReduceValid;
      end
      if (tokenIO_13_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_13_valid <= tokenIO_13_maskRequestRelease_0 & ~viota;
      if (tokenIO_13_maskRequestRelease_0) begin
        exeReqReg_13_bits_source1 <= exeRequestQueue_13_deq_bits_source1;
        exeReqReg_13_bits_source2 <= exeRequestQueue_13_deq_bits_source2;
        exeReqReg_13_bits_index <= exeRequestQueue_13_deq_bits_index;
        exeReqReg_13_bits_ffo <= exeRequestQueue_13_deq_bits_ffo;
        exeReqReg_13_bits_fpReduceValid <= exeRequestQueue_13_deq_bits_fpReduceValid;
      end
      if (tokenIO_14_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_14_valid <= tokenIO_14_maskRequestRelease_0 & ~viota;
      if (tokenIO_14_maskRequestRelease_0) begin
        exeReqReg_14_bits_source1 <= exeRequestQueue_14_deq_bits_source1;
        exeReqReg_14_bits_source2 <= exeRequestQueue_14_deq_bits_source2;
        exeReqReg_14_bits_index <= exeRequestQueue_14_deq_bits_index;
        exeReqReg_14_bits_ffo <= exeRequestQueue_14_deq_bits_ffo;
        exeReqReg_14_bits_fpReduceValid <= exeRequestQueue_14_deq_bits_fpReduceValid;
      end
      if (tokenIO_15_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_15_valid <= tokenIO_15_maskRequestRelease_0 & ~viota;
      if (tokenIO_15_maskRequestRelease_0) begin
        exeReqReg_15_bits_source1 <= exeRequestQueue_15_deq_bits_source1;
        exeReqReg_15_bits_source2 <= exeRequestQueue_15_deq_bits_source2;
        exeReqReg_15_bits_index <= exeRequestQueue_15_deq_bits_index;
        exeReqReg_15_bits_ffo <= exeRequestQueue_15_deq_bits_ffo;
        exeReqReg_15_bits_fpReduceValid <= exeRequestQueue_15_deq_bits_fpReduceValid;
      end
      if (instReq_valid | groupCounterAdd)
        requestCounter <= instReq_valid ? 5'h0 : requestCounter + 5'h1;
      if (requestStageDeq & anyDataValid)
        executeIndex <= executeIndex + executeIndexGrowth[1:0];
      if (readIssueStageEnq) begin
        readIssueStageState_groupReadState <= 16'h0;
        readIssueStageState_needRead <= _GEN_90 ? _slideAddressGen_indexDeq_bits_needRead : ~notReadSelect;
        readIssueStageState_elementValid <= _GEN_90 ? _slideAddressGen_indexDeq_bits_elementValid : elementValidSelect;
        readIssueStageState_replaceVs1 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_replaceVs1 : 16'h0;
        readIssueStageState_readOffset <= _GEN_90 ? _slideAddressGen_indexDeq_bits_readOffset : offsetSelect;
        readIssueStageState_accessLane_0 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_0 : accessLaneSelect[3:0];
        readIssueStageState_accessLane_1 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_1 : accessLaneSelect[7:4];
        readIssueStageState_accessLane_2 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_2 : accessLaneSelect[11:8];
        readIssueStageState_accessLane_3 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_3 : accessLaneSelect[15:12];
        readIssueStageState_accessLane_4 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_4 : accessLaneSelect[19:16];
        readIssueStageState_accessLane_5 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_5 : accessLaneSelect[23:20];
        readIssueStageState_accessLane_6 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_6 : accessLaneSelect[27:24];
        readIssueStageState_accessLane_7 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_7 : accessLaneSelect[31:28];
        readIssueStageState_accessLane_8 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_8 : accessLaneSelect[35:32];
        readIssueStageState_accessLane_9 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_9 : accessLaneSelect[39:36];
        readIssueStageState_accessLane_10 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_10 : accessLaneSelect[43:40];
        readIssueStageState_accessLane_11 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_11 : accessLaneSelect[47:44];
        readIssueStageState_accessLane_12 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_12 : accessLaneSelect[51:48];
        readIssueStageState_accessLane_13 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_13 : accessLaneSelect[55:52];
        readIssueStageState_accessLane_14 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_14 : accessLaneSelect[59:56];
        readIssueStageState_accessLane_15 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_accessLane_15 : accessLaneSelect[63:60];
        readIssueStageState_vsGrowth_0 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_0 : growthSelect[2:0];
        readIssueStageState_vsGrowth_1 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_1 : growthSelect[5:3];
        readIssueStageState_vsGrowth_2 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_2 : growthSelect[8:6];
        readIssueStageState_vsGrowth_3 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_3 : growthSelect[11:9];
        readIssueStageState_vsGrowth_4 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_4 : growthSelect[14:12];
        readIssueStageState_vsGrowth_5 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_5 : growthSelect[17:15];
        readIssueStageState_vsGrowth_6 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_6 : growthSelect[20:18];
        readIssueStageState_vsGrowth_7 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_7 : growthSelect[23:21];
        readIssueStageState_vsGrowth_8 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_8 : growthSelect[26:24];
        readIssueStageState_vsGrowth_9 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_9 : growthSelect[29:27];
        readIssueStageState_vsGrowth_10 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_10 : growthSelect[32:30];
        readIssueStageState_vsGrowth_11 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_11 : growthSelect[35:33];
        readIssueStageState_vsGrowth_12 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_12 : growthSelect[38:36];
        readIssueStageState_vsGrowth_13 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_13 : growthSelect[41:39];
        readIssueStageState_vsGrowth_14 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_14 : growthSelect[44:42];
        readIssueStageState_vsGrowth_15 <= _GEN_90 ? _slideAddressGen_indexDeq_bits_vsGrowth_15 : growthSelect[47:45];
        readIssueStageState_executeGroup <= _GEN_90 ? _slideAddressGen_indexDeq_bits_executeGroup : executeGroup;
        readIssueStageState_readDataOffset <= _GEN_90 ? _slideAddressGen_indexDeq_bits_readDataOffset : dataOffsetSelect;
        readIssueStageState_last <= _GEN_90 ? _slideAddressGen_indexDeq_bits_last : isVlBoundary;
      end
      else if (anyReadFire)
        readIssueStageState_groupReadState <= readStateUpdate;
      if (readTypeRequestDeq ^ readIssueStageEnq)
        readIssueStageValid <= readIssueStageEnq;
      if (_tokenCheck_T ^ readTokenRelease_0)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (pipeReadFire_1 ^ readTokenRelease_1)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (pipeReadFire_2 ^ readTokenRelease_2)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (pipeReadFire_3 ^ readTokenRelease_3)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (pipeReadFire_4 ^ readTokenRelease_4)
        tokenCheck_counter_4 <= tokenCheck_counter_4 + tokenCheck_counterChange_4;
      if (pipeReadFire_5 ^ readTokenRelease_5)
        tokenCheck_counter_5 <= tokenCheck_counter_5 + tokenCheck_counterChange_5;
      if (pipeReadFire_6 ^ readTokenRelease_6)
        tokenCheck_counter_6 <= tokenCheck_counter_6 + tokenCheck_counterChange_6;
      if (pipeReadFire_7 ^ readTokenRelease_7)
        tokenCheck_counter_7 <= tokenCheck_counter_7 + tokenCheck_counterChange_7;
      if (pipeReadFire_8 ^ readTokenRelease_8)
        tokenCheck_counter_8 <= tokenCheck_counter_8 + tokenCheck_counterChange_8;
      if (pipeReadFire_9 ^ readTokenRelease_9)
        tokenCheck_counter_9 <= tokenCheck_counter_9 + tokenCheck_counterChange_9;
      if (pipeReadFire_10 ^ readTokenRelease_10)
        tokenCheck_counter_10 <= tokenCheck_counter_10 + tokenCheck_counterChange_10;
      if (pipeReadFire_11 ^ readTokenRelease_11)
        tokenCheck_counter_11 <= tokenCheck_counter_11 + tokenCheck_counterChange_11;
      if (pipeReadFire_12 ^ readTokenRelease_12)
        tokenCheck_counter_12 <= tokenCheck_counter_12 + tokenCheck_counterChange_12;
      if (pipeReadFire_13 ^ readTokenRelease_13)
        tokenCheck_counter_13 <= tokenCheck_counter_13 + tokenCheck_counterChange_13;
      if (pipeReadFire_14 ^ readTokenRelease_14)
        tokenCheck_counter_14 <= tokenCheck_counter_14 + tokenCheck_counterChange_14;
      if (pipeReadFire_15 ^ readTokenRelease_15)
        tokenCheck_counter_15 <= tokenCheck_counter_15 + tokenCheck_counterChange_15;
      if (reorderQueueAllocate_release | readIssueStageEnq) begin
        reorderQueueAllocate_counter <= reorderQueueAllocate_counterUpdate;
        reorderQueueAllocate_counterWillUpdate <= reorderQueueAllocate_counterUpdate + 6'h10;
      end
      if (reorderQueueAllocate_release_1 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_1 <= reorderQueueAllocate_counterUpdate_1;
        reorderQueueAllocate_counterWillUpdate_1 <= reorderQueueAllocate_counterUpdate_1 + 6'h10;
      end
      if (reorderQueueAllocate_release_2 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_2 <= reorderQueueAllocate_counterUpdate_2;
        reorderQueueAllocate_counterWillUpdate_2 <= reorderQueueAllocate_counterUpdate_2 + 6'h10;
      end
      if (reorderQueueAllocate_release_3 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_3 <= reorderQueueAllocate_counterUpdate_3;
        reorderQueueAllocate_counterWillUpdate_3 <= reorderQueueAllocate_counterUpdate_3 + 6'h10;
      end
      if (reorderQueueAllocate_release_4 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_4 <= reorderQueueAllocate_counterUpdate_4;
        reorderQueueAllocate_counterWillUpdate_4 <= reorderQueueAllocate_counterUpdate_4 + 6'h10;
      end
      if (reorderQueueAllocate_release_5 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_5 <= reorderQueueAllocate_counterUpdate_5;
        reorderQueueAllocate_counterWillUpdate_5 <= reorderQueueAllocate_counterUpdate_5 + 6'h10;
      end
      if (reorderQueueAllocate_release_6 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_6 <= reorderQueueAllocate_counterUpdate_6;
        reorderQueueAllocate_counterWillUpdate_6 <= reorderQueueAllocate_counterUpdate_6 + 6'h10;
      end
      if (reorderQueueAllocate_release_7 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_7 <= reorderQueueAllocate_counterUpdate_7;
        reorderQueueAllocate_counterWillUpdate_7 <= reorderQueueAllocate_counterUpdate_7 + 6'h10;
      end
      if (reorderQueueAllocate_release_8 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_8 <= reorderQueueAllocate_counterUpdate_8;
        reorderQueueAllocate_counterWillUpdate_8 <= reorderQueueAllocate_counterUpdate_8 + 6'h10;
      end
      if (reorderQueueAllocate_release_9 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_9 <= reorderQueueAllocate_counterUpdate_9;
        reorderQueueAllocate_counterWillUpdate_9 <= reorderQueueAllocate_counterUpdate_9 + 6'h10;
      end
      if (reorderQueueAllocate_release_10 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_10 <= reorderQueueAllocate_counterUpdate_10;
        reorderQueueAllocate_counterWillUpdate_10 <= reorderQueueAllocate_counterUpdate_10 + 6'h10;
      end
      if (reorderQueueAllocate_release_11 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_11 <= reorderQueueAllocate_counterUpdate_11;
        reorderQueueAllocate_counterWillUpdate_11 <= reorderQueueAllocate_counterUpdate_11 + 6'h10;
      end
      if (reorderQueueAllocate_release_12 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_12 <= reorderQueueAllocate_counterUpdate_12;
        reorderQueueAllocate_counterWillUpdate_12 <= reorderQueueAllocate_counterUpdate_12 + 6'h10;
      end
      if (reorderQueueAllocate_release_13 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_13 <= reorderQueueAllocate_counterUpdate_13;
        reorderQueueAllocate_counterWillUpdate_13 <= reorderQueueAllocate_counterUpdate_13 + 6'h10;
      end
      if (reorderQueueAllocate_release_14 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_14 <= reorderQueueAllocate_counterUpdate_14;
        reorderQueueAllocate_counterWillUpdate_14 <= reorderQueueAllocate_counterUpdate_14 + 6'h10;
      end
      if (reorderQueueAllocate_release_15 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_15 <= reorderQueueAllocate_counterUpdate_15;
        reorderQueueAllocate_counterWillUpdate_15 <= reorderQueueAllocate_counterUpdate_15 + 6'h10;
      end
      if (reorderStageEnqFire ^ reorderStageDeqFire)
        reorderStageValid <= reorderStageEnqFire;
      if (_write1HPipe_0_T & readType)
        reorderStageState_0 <= reorderStageState_0 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_0 <= 5'h0;
      if (_write1HPipe_1_T & readType)
        reorderStageState_1 <= reorderStageState_1 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_1 <= 5'h0;
      if (_write1HPipe_2_T & readType)
        reorderStageState_2 <= reorderStageState_2 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_2 <= 5'h0;
      if (_write1HPipe_3_T & readType)
        reorderStageState_3 <= reorderStageState_3 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_3 <= 5'h0;
      if (_write1HPipe_4_T & readType)
        reorderStageState_4 <= reorderStageState_4 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_4 <= 5'h0;
      if (_write1HPipe_5_T & readType)
        reorderStageState_5 <= reorderStageState_5 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_5 <= 5'h0;
      if (_write1HPipe_6_T & readType)
        reorderStageState_6 <= reorderStageState_6 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_6 <= 5'h0;
      if (_write1HPipe_7_T & readType)
        reorderStageState_7 <= reorderStageState_7 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_7 <= 5'h0;
      if (_write1HPipe_8_T & readType)
        reorderStageState_8 <= reorderStageState_8 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_8 <= 5'h0;
      if (_write1HPipe_9_T & readType)
        reorderStageState_9 <= reorderStageState_9 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_9 <= 5'h0;
      if (_write1HPipe_10_T & readType)
        reorderStageState_10 <= reorderStageState_10 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_10 <= 5'h0;
      if (_write1HPipe_11_T & readType)
        reorderStageState_11 <= reorderStageState_11 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_11 <= 5'h0;
      if (_write1HPipe_12_T & readType)
        reorderStageState_12 <= reorderStageState_12 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_12 <= 5'h0;
      if (_write1HPipe_13_T & readType)
        reorderStageState_13 <= reorderStageState_13 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_13 <= 5'h0;
      if (_write1HPipe_14_T & readType)
        reorderStageState_14 <= reorderStageState_14 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_14 <= 5'h0;
      if (_write1HPipe_15_T & readType)
        reorderStageState_15 <= reorderStageState_15 + 5'h1;
      else if (reorderStageEnqFire)
        reorderStageState_15 <= 5'h0;
      if (reorderStageEnqFire) begin
        reorderStageNeed_0 <= accessCountQueue_deq_bits_0;
        reorderStageNeed_1 <= accessCountQueue_deq_bits_1;
        reorderStageNeed_2 <= accessCountQueue_deq_bits_2;
        reorderStageNeed_3 <= accessCountQueue_deq_bits_3;
        reorderStageNeed_4 <= accessCountQueue_deq_bits_4;
        reorderStageNeed_5 <= accessCountQueue_deq_bits_5;
        reorderStageNeed_6 <= accessCountQueue_deq_bits_6;
        reorderStageNeed_7 <= accessCountQueue_deq_bits_7;
        reorderStageNeed_8 <= accessCountQueue_deq_bits_8;
        reorderStageNeed_9 <= accessCountQueue_deq_bits_9;
        reorderStageNeed_10 <= accessCountQueue_deq_bits_10;
        reorderStageNeed_11 <= accessCountQueue_deq_bits_11;
        reorderStageNeed_12 <= accessCountQueue_deq_bits_12;
        reorderStageNeed_13 <= accessCountQueue_deq_bits_13;
        reorderStageNeed_14 <= accessCountQueue_deq_bits_14;
        reorderStageNeed_15 <= accessCountQueue_deq_bits_15;
      end
      if (waiteStageEnqFire) begin
        waiteReadDataPipeReg_executeGroup <= readWaitQueue_deq_bits_executeGroup;
        waiteReadDataPipeReg_sourceValid <= readWaitQueue_deq_bits_sourceValid;
        waiteReadDataPipeReg_replaceVs1 <= readWaitQueue_deq_bits_replaceVs1;
        waiteReadDataPipeReg_needRead <= readWaitQueue_deq_bits_needRead;
        waiteReadDataPipeReg_last <= readWaitQueue_deq_bits_last;
      end
      if (readTokenRelease_1)
        waiteReadData_1 <= readData_readDataQueue_1_deq_bits;
      if (readTokenRelease_2)
        waiteReadData_2 <= readData_readDataQueue_2_deq_bits;
      if (readTokenRelease_3)
        waiteReadData_3 <= readData_readDataQueue_3_deq_bits;
      if (readTokenRelease_4)
        waiteReadData_4 <= readData_readDataQueue_4_deq_bits;
      if (readTokenRelease_5)
        waiteReadData_5 <= readData_readDataQueue_5_deq_bits;
      if (readTokenRelease_6)
        waiteReadData_6 <= readData_readDataQueue_6_deq_bits;
      if (readTokenRelease_7)
        waiteReadData_7 <= readData_readDataQueue_7_deq_bits;
      if (readTokenRelease_8)
        waiteReadData_8 <= readData_readDataQueue_8_deq_bits;
      if (readTokenRelease_9)
        waiteReadData_9 <= readData_readDataQueue_9_deq_bits;
      if (readTokenRelease_10)
        waiteReadData_10 <= readData_readDataQueue_10_deq_bits;
      if (readTokenRelease_11)
        waiteReadData_11 <= readData_readDataQueue_11_deq_bits;
      if (readTokenRelease_12)
        waiteReadData_12 <= readData_readDataQueue_12_deq_bits;
      if (readTokenRelease_13)
        waiteReadData_13 <= readData_readDataQueue_13_deq_bits;
      if (readTokenRelease_14)
        waiteReadData_14 <= readData_readDataQueue_14_deq_bits;
      if (readTokenRelease_15)
        waiteReadData_15 <= readData_readDataQueue_15_deq_bits;
      if (waiteStageEnqFire & (|readResultValid))
        waiteReadSate <= readResultValid;
      else if (|readResultValid)
        waiteReadSate <= waiteReadSate | readResultValid;
      else if (waiteStageEnqFire)
        waiteReadSate <= 16'h0;
      if (waiteStageDeqFire ^ waiteStageEnqFire)
        waiteReadStageValid <= waiteStageEnqFire;
      if (_dataNotInShifter_T ^ writeRelease_0)
        dataNotInShifter_writeTokenCounter <= dataNotInShifter_writeTokenCounter + dataNotInShifter_writeTokenChange;
      if (_dataNotInShifter_T_3 ^ writeRelease_1)
        dataNotInShifter_writeTokenCounter_1 <= dataNotInShifter_writeTokenCounter_1 + dataNotInShifter_writeTokenChange_1;
      if (_dataNotInShifter_T_6 ^ writeRelease_2)
        dataNotInShifter_writeTokenCounter_2 <= dataNotInShifter_writeTokenCounter_2 + dataNotInShifter_writeTokenChange_2;
      if (_dataNotInShifter_T_9 ^ writeRelease_3)
        dataNotInShifter_writeTokenCounter_3 <= dataNotInShifter_writeTokenCounter_3 + dataNotInShifter_writeTokenChange_3;
      if (_dataNotInShifter_T_12 ^ writeRelease_4)
        dataNotInShifter_writeTokenCounter_4 <= dataNotInShifter_writeTokenCounter_4 + dataNotInShifter_writeTokenChange_4;
      if (_dataNotInShifter_T_15 ^ writeRelease_5)
        dataNotInShifter_writeTokenCounter_5 <= dataNotInShifter_writeTokenCounter_5 + dataNotInShifter_writeTokenChange_5;
      if (_dataNotInShifter_T_18 ^ writeRelease_6)
        dataNotInShifter_writeTokenCounter_6 <= dataNotInShifter_writeTokenCounter_6 + dataNotInShifter_writeTokenChange_6;
      if (_dataNotInShifter_T_21 ^ writeRelease_7)
        dataNotInShifter_writeTokenCounter_7 <= dataNotInShifter_writeTokenCounter_7 + dataNotInShifter_writeTokenChange_7;
      if (_dataNotInShifter_T_24 ^ writeRelease_8)
        dataNotInShifter_writeTokenCounter_8 <= dataNotInShifter_writeTokenCounter_8 + dataNotInShifter_writeTokenChange_8;
      if (_dataNotInShifter_T_27 ^ writeRelease_9)
        dataNotInShifter_writeTokenCounter_9 <= dataNotInShifter_writeTokenCounter_9 + dataNotInShifter_writeTokenChange_9;
      if (_dataNotInShifter_T_30 ^ writeRelease_10)
        dataNotInShifter_writeTokenCounter_10 <= dataNotInShifter_writeTokenCounter_10 + dataNotInShifter_writeTokenChange_10;
      if (_dataNotInShifter_T_33 ^ writeRelease_11)
        dataNotInShifter_writeTokenCounter_11 <= dataNotInShifter_writeTokenCounter_11 + dataNotInShifter_writeTokenChange_11;
      if (_dataNotInShifter_T_36 ^ writeRelease_12)
        dataNotInShifter_writeTokenCounter_12 <= dataNotInShifter_writeTokenCounter_12 + dataNotInShifter_writeTokenChange_12;
      if (_dataNotInShifter_T_39 ^ writeRelease_13)
        dataNotInShifter_writeTokenCounter_13 <= dataNotInShifter_writeTokenCounter_13 + dataNotInShifter_writeTokenChange_13;
      if (_dataNotInShifter_T_42 ^ writeRelease_14)
        dataNotInShifter_writeTokenCounter_14 <= dataNotInShifter_writeTokenCounter_14 + dataNotInShifter_writeTokenChange_14;
      if (_dataNotInShifter_T_45 ^ writeRelease_15)
        dataNotInShifter_writeTokenCounter_15 <= dataNotInShifter_writeTokenCounter_15 + dataNotInShifter_writeTokenChange_15;
      waiteLastRequest <= ~readType & requestStageDeq & lastGroup | ~lastReportValid & waiteLastRequest;
      waitQueueClear <= executeStageClean | invalidEnq | ~lastReportValid & waitQueueClear;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:113];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h72; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[7'h0];
        v0_1 = _RANDOM[7'h1];
        v0_2 = _RANDOM[7'h2];
        v0_3 = _RANDOM[7'h3];
        v0_4 = _RANDOM[7'h4];
        v0_5 = _RANDOM[7'h5];
        v0_6 = _RANDOM[7'h6];
        v0_7 = _RANDOM[7'h7];
        v0_8 = _RANDOM[7'h8];
        v0_9 = _RANDOM[7'h9];
        v0_10 = _RANDOM[7'hA];
        v0_11 = _RANDOM[7'hB];
        v0_12 = _RANDOM[7'hC];
        v0_13 = _RANDOM[7'hD];
        v0_14 = _RANDOM[7'hE];
        v0_15 = _RANDOM[7'hF];
        v0_16 = _RANDOM[7'h10];
        v0_17 = _RANDOM[7'h11];
        v0_18 = _RANDOM[7'h12];
        v0_19 = _RANDOM[7'h13];
        v0_20 = _RANDOM[7'h14];
        v0_21 = _RANDOM[7'h15];
        v0_22 = _RANDOM[7'h16];
        v0_23 = _RANDOM[7'h17];
        v0_24 = _RANDOM[7'h18];
        v0_25 = _RANDOM[7'h19];
        v0_26 = _RANDOM[7'h1A];
        v0_27 = _RANDOM[7'h1B];
        v0_28 = _RANDOM[7'h1C];
        v0_29 = _RANDOM[7'h1D];
        v0_30 = _RANDOM[7'h1E];
        v0_31 = _RANDOM[7'h1F];
        gatherReadState = _RANDOM[7'h20][1:0];
        gatherDatOffset = _RANDOM[7'h20][3:2];
        gatherLane = _RANDOM[7'h20][7:4];
        gatherOffset = _RANDOM[7'h20][8];
        gatherGrowth = _RANDOM[7'h20][11:9];
        instReg_instructionIndex = _RANDOM[7'h20][14:12];
        instReg_decodeResult_orderReduce = _RANDOM[7'h20][15];
        instReg_decodeResult_floatMul = _RANDOM[7'h20][16];
        instReg_decodeResult_fpExecutionType = _RANDOM[7'h20][18:17];
        instReg_decodeResult_float = _RANDOM[7'h20][19];
        instReg_decodeResult_specialSlot = _RANDOM[7'h20][20];
        instReg_decodeResult_topUop = _RANDOM[7'h20][25:21];
        instReg_decodeResult_popCount = _RANDOM[7'h20][26];
        instReg_decodeResult_ffo = _RANDOM[7'h20][27];
        instReg_decodeResult_average = _RANDOM[7'h20][28];
        instReg_decodeResult_reverse = _RANDOM[7'h20][29];
        instReg_decodeResult_dontNeedExecuteInLane = _RANDOM[7'h20][30];
        instReg_decodeResult_scheduler = _RANDOM[7'h20][31];
        instReg_decodeResult_sReadVD = _RANDOM[7'h21][0];
        instReg_decodeResult_vtype = _RANDOM[7'h21][1];
        instReg_decodeResult_sWrite = _RANDOM[7'h21][2];
        instReg_decodeResult_crossRead = _RANDOM[7'h21][3];
        instReg_decodeResult_crossWrite = _RANDOM[7'h21][4];
        instReg_decodeResult_maskUnit = _RANDOM[7'h21][5];
        instReg_decodeResult_special = _RANDOM[7'h21][6];
        instReg_decodeResult_saturate = _RANDOM[7'h21][7];
        instReg_decodeResult_vwmacc = _RANDOM[7'h21][8];
        instReg_decodeResult_readOnly = _RANDOM[7'h21][9];
        instReg_decodeResult_maskSource = _RANDOM[7'h21][10];
        instReg_decodeResult_maskDestination = _RANDOM[7'h21][11];
        instReg_decodeResult_maskLogic = _RANDOM[7'h21][12];
        instReg_decodeResult_uop = _RANDOM[7'h21][16:13];
        instReg_decodeResult_iota = _RANDOM[7'h21][17];
        instReg_decodeResult_mv = _RANDOM[7'h21][18];
        instReg_decodeResult_extend = _RANDOM[7'h21][19];
        instReg_decodeResult_unOrderWrite = _RANDOM[7'h21][20];
        instReg_decodeResult_compress = _RANDOM[7'h21][21];
        instReg_decodeResult_gather16 = _RANDOM[7'h21][22];
        instReg_decodeResult_gather = _RANDOM[7'h21][23];
        instReg_decodeResult_slid = _RANDOM[7'h21][24];
        instReg_decodeResult_targetRd = _RANDOM[7'h21][25];
        instReg_decodeResult_widenReduce = _RANDOM[7'h21][26];
        instReg_decodeResult_red = _RANDOM[7'h21][27];
        instReg_decodeResult_nr = _RANDOM[7'h21][28];
        instReg_decodeResult_itype = _RANDOM[7'h21][29];
        instReg_decodeResult_unsigned1 = _RANDOM[7'h21][30];
        instReg_decodeResult_unsigned0 = _RANDOM[7'h21][31];
        instReg_decodeResult_other = _RANDOM[7'h22][0];
        instReg_decodeResult_multiCycle = _RANDOM[7'h22][1];
        instReg_decodeResult_divider = _RANDOM[7'h22][2];
        instReg_decodeResult_multiplier = _RANDOM[7'h22][3];
        instReg_decodeResult_shift = _RANDOM[7'h22][4];
        instReg_decodeResult_adder = _RANDOM[7'h22][5];
        instReg_decodeResult_logic = _RANDOM[7'h22][6];
        instReg_readFromScala = {_RANDOM[7'h22][31:7], _RANDOM[7'h23][6:0]};
        instReg_sew = _RANDOM[7'h23][8:7];
        instReg_vlmul = _RANDOM[7'h23][11:9];
        instReg_maskType = _RANDOM[7'h23][12];
        instReg_vxrm = _RANDOM[7'h23][15:13];
        instReg_vs2 = _RANDOM[7'h23][20:16];
        instReg_vs1 = _RANDOM[7'h23][25:21];
        instReg_vd = _RANDOM[7'h23][30:26];
        instReg_vl = {_RANDOM[7'h23][31], _RANDOM[7'h24][9:0]};
        instVlValid = _RANDOM[7'h24][10];
        readVS1Reg_dataValid = _RANDOM[7'h24][11];
        readVS1Reg_requestSend = _RANDOM[7'h24][12];
        readVS1Reg_sendToExecution = _RANDOM[7'h24][13];
        readVS1Reg_data = {_RANDOM[7'h24][31:14], _RANDOM[7'h25][13:0]};
        readVS1Reg_readIndex = _RANDOM[7'h25][17:14];
        exeReqReg_0_valid = _RANDOM[7'h26][2];
        exeReqReg_0_bits_source1 = {_RANDOM[7'h26][31:3], _RANDOM[7'h27][2:0]};
        exeReqReg_0_bits_source2 = {_RANDOM[7'h27][31:3], _RANDOM[7'h28][2:0]};
        exeReqReg_0_bits_index = _RANDOM[7'h28][5:3];
        exeReqReg_0_bits_ffo = _RANDOM[7'h28][6];
        exeReqReg_0_bits_fpReduceValid = _RANDOM[7'h28][7];
        exeReqReg_1_valid = _RANDOM[7'h28][8];
        exeReqReg_1_bits_source1 = {_RANDOM[7'h28][31:9], _RANDOM[7'h29][8:0]};
        exeReqReg_1_bits_source2 = {_RANDOM[7'h29][31:9], _RANDOM[7'h2A][8:0]};
        exeReqReg_1_bits_index = _RANDOM[7'h2A][11:9];
        exeReqReg_1_bits_ffo = _RANDOM[7'h2A][12];
        exeReqReg_1_bits_fpReduceValid = _RANDOM[7'h2A][13];
        exeReqReg_2_valid = _RANDOM[7'h2A][14];
        exeReqReg_2_bits_source1 = {_RANDOM[7'h2A][31:15], _RANDOM[7'h2B][14:0]};
        exeReqReg_2_bits_source2 = {_RANDOM[7'h2B][31:15], _RANDOM[7'h2C][14:0]};
        exeReqReg_2_bits_index = _RANDOM[7'h2C][17:15];
        exeReqReg_2_bits_ffo = _RANDOM[7'h2C][18];
        exeReqReg_2_bits_fpReduceValid = _RANDOM[7'h2C][19];
        exeReqReg_3_valid = _RANDOM[7'h2C][20];
        exeReqReg_3_bits_source1 = {_RANDOM[7'h2C][31:21], _RANDOM[7'h2D][20:0]};
        exeReqReg_3_bits_source2 = {_RANDOM[7'h2D][31:21], _RANDOM[7'h2E][20:0]};
        exeReqReg_3_bits_index = _RANDOM[7'h2E][23:21];
        exeReqReg_3_bits_ffo = _RANDOM[7'h2E][24];
        exeReqReg_3_bits_fpReduceValid = _RANDOM[7'h2E][25];
        exeReqReg_4_valid = _RANDOM[7'h2E][26];
        exeReqReg_4_bits_source1 = {_RANDOM[7'h2E][31:27], _RANDOM[7'h2F][26:0]};
        exeReqReg_4_bits_source2 = {_RANDOM[7'h2F][31:27], _RANDOM[7'h30][26:0]};
        exeReqReg_4_bits_index = _RANDOM[7'h30][29:27];
        exeReqReg_4_bits_ffo = _RANDOM[7'h30][30];
        exeReqReg_4_bits_fpReduceValid = _RANDOM[7'h30][31];
        exeReqReg_5_valid = _RANDOM[7'h31][0];
        exeReqReg_5_bits_source1 = {_RANDOM[7'h31][31:1], _RANDOM[7'h32][0]};
        exeReqReg_5_bits_source2 = {_RANDOM[7'h32][31:1], _RANDOM[7'h33][0]};
        exeReqReg_5_bits_index = _RANDOM[7'h33][3:1];
        exeReqReg_5_bits_ffo = _RANDOM[7'h33][4];
        exeReqReg_5_bits_fpReduceValid = _RANDOM[7'h33][5];
        exeReqReg_6_valid = _RANDOM[7'h33][6];
        exeReqReg_6_bits_source1 = {_RANDOM[7'h33][31:7], _RANDOM[7'h34][6:0]};
        exeReqReg_6_bits_source2 = {_RANDOM[7'h34][31:7], _RANDOM[7'h35][6:0]};
        exeReqReg_6_bits_index = _RANDOM[7'h35][9:7];
        exeReqReg_6_bits_ffo = _RANDOM[7'h35][10];
        exeReqReg_6_bits_fpReduceValid = _RANDOM[7'h35][11];
        exeReqReg_7_valid = _RANDOM[7'h35][12];
        exeReqReg_7_bits_source1 = {_RANDOM[7'h35][31:13], _RANDOM[7'h36][12:0]};
        exeReqReg_7_bits_source2 = {_RANDOM[7'h36][31:13], _RANDOM[7'h37][12:0]};
        exeReqReg_7_bits_index = _RANDOM[7'h37][15:13];
        exeReqReg_7_bits_ffo = _RANDOM[7'h37][16];
        exeReqReg_7_bits_fpReduceValid = _RANDOM[7'h37][17];
        exeReqReg_8_valid = _RANDOM[7'h37][18];
        exeReqReg_8_bits_source1 = {_RANDOM[7'h37][31:19], _RANDOM[7'h38][18:0]};
        exeReqReg_8_bits_source2 = {_RANDOM[7'h38][31:19], _RANDOM[7'h39][18:0]};
        exeReqReg_8_bits_index = _RANDOM[7'h39][21:19];
        exeReqReg_8_bits_ffo = _RANDOM[7'h39][22];
        exeReqReg_8_bits_fpReduceValid = _RANDOM[7'h39][23];
        exeReqReg_9_valid = _RANDOM[7'h39][24];
        exeReqReg_9_bits_source1 = {_RANDOM[7'h39][31:25], _RANDOM[7'h3A][24:0]};
        exeReqReg_9_bits_source2 = {_RANDOM[7'h3A][31:25], _RANDOM[7'h3B][24:0]};
        exeReqReg_9_bits_index = _RANDOM[7'h3B][27:25];
        exeReqReg_9_bits_ffo = _RANDOM[7'h3B][28];
        exeReqReg_9_bits_fpReduceValid = _RANDOM[7'h3B][29];
        exeReqReg_10_valid = _RANDOM[7'h3B][30];
        exeReqReg_10_bits_source1 = {_RANDOM[7'h3B][31], _RANDOM[7'h3C][30:0]};
        exeReqReg_10_bits_source2 = {_RANDOM[7'h3C][31], _RANDOM[7'h3D][30:0]};
        exeReqReg_10_bits_index = {_RANDOM[7'h3D][31], _RANDOM[7'h3E][1:0]};
        exeReqReg_10_bits_ffo = _RANDOM[7'h3E][2];
        exeReqReg_10_bits_fpReduceValid = _RANDOM[7'h3E][3];
        exeReqReg_11_valid = _RANDOM[7'h3E][4];
        exeReqReg_11_bits_source1 = {_RANDOM[7'h3E][31:5], _RANDOM[7'h3F][4:0]};
        exeReqReg_11_bits_source2 = {_RANDOM[7'h3F][31:5], _RANDOM[7'h40][4:0]};
        exeReqReg_11_bits_index = _RANDOM[7'h40][7:5];
        exeReqReg_11_bits_ffo = _RANDOM[7'h40][8];
        exeReqReg_11_bits_fpReduceValid = _RANDOM[7'h40][9];
        exeReqReg_12_valid = _RANDOM[7'h40][10];
        exeReqReg_12_bits_source1 = {_RANDOM[7'h40][31:11], _RANDOM[7'h41][10:0]};
        exeReqReg_12_bits_source2 = {_RANDOM[7'h41][31:11], _RANDOM[7'h42][10:0]};
        exeReqReg_12_bits_index = _RANDOM[7'h42][13:11];
        exeReqReg_12_bits_ffo = _RANDOM[7'h42][14];
        exeReqReg_12_bits_fpReduceValid = _RANDOM[7'h42][15];
        exeReqReg_13_valid = _RANDOM[7'h42][16];
        exeReqReg_13_bits_source1 = {_RANDOM[7'h42][31:17], _RANDOM[7'h43][16:0]};
        exeReqReg_13_bits_source2 = {_RANDOM[7'h43][31:17], _RANDOM[7'h44][16:0]};
        exeReqReg_13_bits_index = _RANDOM[7'h44][19:17];
        exeReqReg_13_bits_ffo = _RANDOM[7'h44][20];
        exeReqReg_13_bits_fpReduceValid = _RANDOM[7'h44][21];
        exeReqReg_14_valid = _RANDOM[7'h44][22];
        exeReqReg_14_bits_source1 = {_RANDOM[7'h44][31:23], _RANDOM[7'h45][22:0]};
        exeReqReg_14_bits_source2 = {_RANDOM[7'h45][31:23], _RANDOM[7'h46][22:0]};
        exeReqReg_14_bits_index = _RANDOM[7'h46][25:23];
        exeReqReg_14_bits_ffo = _RANDOM[7'h46][26];
        exeReqReg_14_bits_fpReduceValid = _RANDOM[7'h46][27];
        exeReqReg_15_valid = _RANDOM[7'h46][28];
        exeReqReg_15_bits_source1 = {_RANDOM[7'h46][31:29], _RANDOM[7'h47][28:0]};
        exeReqReg_15_bits_source2 = {_RANDOM[7'h47][31:29], _RANDOM[7'h48][28:0]};
        exeReqReg_15_bits_index = _RANDOM[7'h48][31:29];
        exeReqReg_15_bits_ffo = _RANDOM[7'h49][0];
        exeReqReg_15_bits_fpReduceValid = _RANDOM[7'h49][1];
        requestCounter = _RANDOM[7'h49][6:2];
        executeIndex = _RANDOM[7'h49][8:7];
        readIssueStageState_groupReadState = _RANDOM[7'h49][24:9];
        readIssueStageState_needRead = {_RANDOM[7'h49][31:25], _RANDOM[7'h4A][8:0]};
        readIssueStageState_elementValid = _RANDOM[7'h4A][24:9];
        readIssueStageState_replaceVs1 = {_RANDOM[7'h4A][31:25], _RANDOM[7'h4B][8:0]};
        readIssueStageState_readOffset = _RANDOM[7'h4B][24:9];
        readIssueStageState_accessLane_0 = _RANDOM[7'h4B][28:25];
        readIssueStageState_accessLane_1 = {_RANDOM[7'h4B][31:29], _RANDOM[7'h4C][0]};
        readIssueStageState_accessLane_2 = _RANDOM[7'h4C][4:1];
        readIssueStageState_accessLane_3 = _RANDOM[7'h4C][8:5];
        readIssueStageState_accessLane_4 = _RANDOM[7'h4C][12:9];
        readIssueStageState_accessLane_5 = _RANDOM[7'h4C][16:13];
        readIssueStageState_accessLane_6 = _RANDOM[7'h4C][20:17];
        readIssueStageState_accessLane_7 = _RANDOM[7'h4C][24:21];
        readIssueStageState_accessLane_8 = _RANDOM[7'h4C][28:25];
        readIssueStageState_accessLane_9 = {_RANDOM[7'h4C][31:29], _RANDOM[7'h4D][0]};
        readIssueStageState_accessLane_10 = _RANDOM[7'h4D][4:1];
        readIssueStageState_accessLane_11 = _RANDOM[7'h4D][8:5];
        readIssueStageState_accessLane_12 = _RANDOM[7'h4D][12:9];
        readIssueStageState_accessLane_13 = _RANDOM[7'h4D][16:13];
        readIssueStageState_accessLane_14 = _RANDOM[7'h4D][20:17];
        readIssueStageState_accessLane_15 = _RANDOM[7'h4D][24:21];
        readIssueStageState_vsGrowth_0 = _RANDOM[7'h4D][27:25];
        readIssueStageState_vsGrowth_1 = _RANDOM[7'h4D][30:28];
        readIssueStageState_vsGrowth_2 = {_RANDOM[7'h4D][31], _RANDOM[7'h4E][1:0]};
        readIssueStageState_vsGrowth_3 = _RANDOM[7'h4E][4:2];
        readIssueStageState_vsGrowth_4 = _RANDOM[7'h4E][7:5];
        readIssueStageState_vsGrowth_5 = _RANDOM[7'h4E][10:8];
        readIssueStageState_vsGrowth_6 = _RANDOM[7'h4E][13:11];
        readIssueStageState_vsGrowth_7 = _RANDOM[7'h4E][16:14];
        readIssueStageState_vsGrowth_8 = _RANDOM[7'h4E][19:17];
        readIssueStageState_vsGrowth_9 = _RANDOM[7'h4E][22:20];
        readIssueStageState_vsGrowth_10 = _RANDOM[7'h4E][25:23];
        readIssueStageState_vsGrowth_11 = _RANDOM[7'h4E][28:26];
        readIssueStageState_vsGrowth_12 = _RANDOM[7'h4E][31:29];
        readIssueStageState_vsGrowth_13 = _RANDOM[7'h4F][2:0];
        readIssueStageState_vsGrowth_14 = _RANDOM[7'h4F][5:3];
        readIssueStageState_vsGrowth_15 = _RANDOM[7'h4F][8:6];
        readIssueStageState_executeGroup = _RANDOM[7'h4F][15:9];
        readIssueStageState_readDataOffset = {_RANDOM[7'h4F][31:16], _RANDOM[7'h50][15:0]};
        readIssueStageState_last = _RANDOM[7'h50][16];
        readIssueStageValid = _RANDOM[7'h50][17];
        tokenCheck_counter = _RANDOM[7'h50][21:18];
        tokenCheck_counter_1 = _RANDOM[7'h50][25:22];
        tokenCheck_counter_2 = _RANDOM[7'h50][29:26];
        tokenCheck_counter_3 = {_RANDOM[7'h50][31:30], _RANDOM[7'h51][1:0]};
        tokenCheck_counter_4 = _RANDOM[7'h51][5:2];
        tokenCheck_counter_5 = _RANDOM[7'h51][9:6];
        tokenCheck_counter_6 = _RANDOM[7'h51][13:10];
        tokenCheck_counter_7 = _RANDOM[7'h51][17:14];
        tokenCheck_counter_8 = _RANDOM[7'h51][21:18];
        tokenCheck_counter_9 = _RANDOM[7'h51][25:22];
        tokenCheck_counter_10 = _RANDOM[7'h51][29:26];
        tokenCheck_counter_11 = {_RANDOM[7'h51][31:30], _RANDOM[7'h52][1:0]};
        tokenCheck_counter_12 = _RANDOM[7'h52][5:2];
        tokenCheck_counter_13 = _RANDOM[7'h52][9:6];
        tokenCheck_counter_14 = _RANDOM[7'h52][13:10];
        tokenCheck_counter_15 = _RANDOM[7'h52][17:14];
        reorderQueueAllocate_counter = _RANDOM[7'h52][23:18];
        reorderQueueAllocate_counterWillUpdate = _RANDOM[7'h52][29:24];
        reorderQueueAllocate_counter_1 = {_RANDOM[7'h52][31:30], _RANDOM[7'h53][3:0]};
        reorderQueueAllocate_counterWillUpdate_1 = _RANDOM[7'h53][9:4];
        reorderQueueAllocate_counter_2 = _RANDOM[7'h53][15:10];
        reorderQueueAllocate_counterWillUpdate_2 = _RANDOM[7'h53][21:16];
        reorderQueueAllocate_counter_3 = _RANDOM[7'h53][27:22];
        reorderQueueAllocate_counterWillUpdate_3 = {_RANDOM[7'h53][31:28], _RANDOM[7'h54][1:0]};
        reorderQueueAllocate_counter_4 = _RANDOM[7'h54][7:2];
        reorderQueueAllocate_counterWillUpdate_4 = _RANDOM[7'h54][13:8];
        reorderQueueAllocate_counter_5 = _RANDOM[7'h54][19:14];
        reorderQueueAllocate_counterWillUpdate_5 = _RANDOM[7'h54][25:20];
        reorderQueueAllocate_counter_6 = _RANDOM[7'h54][31:26];
        reorderQueueAllocate_counterWillUpdate_6 = _RANDOM[7'h55][5:0];
        reorderQueueAllocate_counter_7 = _RANDOM[7'h55][11:6];
        reorderQueueAllocate_counterWillUpdate_7 = _RANDOM[7'h55][17:12];
        reorderQueueAllocate_counter_8 = _RANDOM[7'h55][23:18];
        reorderQueueAllocate_counterWillUpdate_8 = _RANDOM[7'h55][29:24];
        reorderQueueAllocate_counter_9 = {_RANDOM[7'h55][31:30], _RANDOM[7'h56][3:0]};
        reorderQueueAllocate_counterWillUpdate_9 = _RANDOM[7'h56][9:4];
        reorderQueueAllocate_counter_10 = _RANDOM[7'h56][15:10];
        reorderQueueAllocate_counterWillUpdate_10 = _RANDOM[7'h56][21:16];
        reorderQueueAllocate_counter_11 = _RANDOM[7'h56][27:22];
        reorderQueueAllocate_counterWillUpdate_11 = {_RANDOM[7'h56][31:28], _RANDOM[7'h57][1:0]};
        reorderQueueAllocate_counter_12 = _RANDOM[7'h57][7:2];
        reorderQueueAllocate_counterWillUpdate_12 = _RANDOM[7'h57][13:8];
        reorderQueueAllocate_counter_13 = _RANDOM[7'h57][19:14];
        reorderQueueAllocate_counterWillUpdate_13 = _RANDOM[7'h57][25:20];
        reorderQueueAllocate_counter_14 = _RANDOM[7'h57][31:26];
        reorderQueueAllocate_counterWillUpdate_14 = _RANDOM[7'h58][5:0];
        reorderQueueAllocate_counter_15 = _RANDOM[7'h58][11:6];
        reorderQueueAllocate_counterWillUpdate_15 = _RANDOM[7'h58][17:12];
        reorderStageValid = _RANDOM[7'h58][18];
        reorderStageState_0 = _RANDOM[7'h58][23:19];
        reorderStageState_1 = _RANDOM[7'h58][28:24];
        reorderStageState_2 = {_RANDOM[7'h58][31:29], _RANDOM[7'h59][1:0]};
        reorderStageState_3 = _RANDOM[7'h59][6:2];
        reorderStageState_4 = _RANDOM[7'h59][11:7];
        reorderStageState_5 = _RANDOM[7'h59][16:12];
        reorderStageState_6 = _RANDOM[7'h59][21:17];
        reorderStageState_7 = _RANDOM[7'h59][26:22];
        reorderStageState_8 = _RANDOM[7'h59][31:27];
        reorderStageState_9 = _RANDOM[7'h5A][4:0];
        reorderStageState_10 = _RANDOM[7'h5A][9:5];
        reorderStageState_11 = _RANDOM[7'h5A][14:10];
        reorderStageState_12 = _RANDOM[7'h5A][19:15];
        reorderStageState_13 = _RANDOM[7'h5A][24:20];
        reorderStageState_14 = _RANDOM[7'h5A][29:25];
        reorderStageState_15 = {_RANDOM[7'h5A][31:30], _RANDOM[7'h5B][2:0]};
        reorderStageNeed_0 = _RANDOM[7'h5B][7:3];
        reorderStageNeed_1 = _RANDOM[7'h5B][12:8];
        reorderStageNeed_2 = _RANDOM[7'h5B][17:13];
        reorderStageNeed_3 = _RANDOM[7'h5B][22:18];
        reorderStageNeed_4 = _RANDOM[7'h5B][27:23];
        reorderStageNeed_5 = {_RANDOM[7'h5B][31:28], _RANDOM[7'h5C][0]};
        reorderStageNeed_6 = _RANDOM[7'h5C][5:1];
        reorderStageNeed_7 = _RANDOM[7'h5C][10:6];
        reorderStageNeed_8 = _RANDOM[7'h5C][15:11];
        reorderStageNeed_9 = _RANDOM[7'h5C][20:16];
        reorderStageNeed_10 = _RANDOM[7'h5C][25:21];
        reorderStageNeed_11 = _RANDOM[7'h5C][30:26];
        reorderStageNeed_12 = {_RANDOM[7'h5C][31], _RANDOM[7'h5D][3:0]};
        reorderStageNeed_13 = _RANDOM[7'h5D][8:4];
        reorderStageNeed_14 = _RANDOM[7'h5D][13:9];
        reorderStageNeed_15 = _RANDOM[7'h5D][18:14];
        waiteReadDataPipeReg_executeGroup = _RANDOM[7'h5D][25:19];
        waiteReadDataPipeReg_sourceValid = {_RANDOM[7'h5D][31:26], _RANDOM[7'h5E][9:0]};
        waiteReadDataPipeReg_replaceVs1 = _RANDOM[7'h5E][25:10];
        waiteReadDataPipeReg_needRead = {_RANDOM[7'h5E][31:26], _RANDOM[7'h5F][9:0]};
        waiteReadDataPipeReg_last = _RANDOM[7'h5F][10];
        waiteReadData_0 = {_RANDOM[7'h5F][31:11], _RANDOM[7'h60][10:0]};
        waiteReadData_1 = {_RANDOM[7'h60][31:11], _RANDOM[7'h61][10:0]};
        waiteReadData_2 = {_RANDOM[7'h61][31:11], _RANDOM[7'h62][10:0]};
        waiteReadData_3 = {_RANDOM[7'h62][31:11], _RANDOM[7'h63][10:0]};
        waiteReadData_4 = {_RANDOM[7'h63][31:11], _RANDOM[7'h64][10:0]};
        waiteReadData_5 = {_RANDOM[7'h64][31:11], _RANDOM[7'h65][10:0]};
        waiteReadData_6 = {_RANDOM[7'h65][31:11], _RANDOM[7'h66][10:0]};
        waiteReadData_7 = {_RANDOM[7'h66][31:11], _RANDOM[7'h67][10:0]};
        waiteReadData_8 = {_RANDOM[7'h67][31:11], _RANDOM[7'h68][10:0]};
        waiteReadData_9 = {_RANDOM[7'h68][31:11], _RANDOM[7'h69][10:0]};
        waiteReadData_10 = {_RANDOM[7'h69][31:11], _RANDOM[7'h6A][10:0]};
        waiteReadData_11 = {_RANDOM[7'h6A][31:11], _RANDOM[7'h6B][10:0]};
        waiteReadData_12 = {_RANDOM[7'h6B][31:11], _RANDOM[7'h6C][10:0]};
        waiteReadData_13 = {_RANDOM[7'h6C][31:11], _RANDOM[7'h6D][10:0]};
        waiteReadData_14 = {_RANDOM[7'h6D][31:11], _RANDOM[7'h6E][10:0]};
        waiteReadData_15 = {_RANDOM[7'h6E][31:11], _RANDOM[7'h6F][10:0]};
        waiteReadSate = _RANDOM[7'h6F][26:11];
        waiteReadStageValid = _RANDOM[7'h6F][27];
        dataNotInShifter_writeTokenCounter = _RANDOM[7'h6F][30:28];
        dataNotInShifter_writeTokenCounter_1 = {_RANDOM[7'h6F][31], _RANDOM[7'h70][1:0]};
        dataNotInShifter_writeTokenCounter_2 = _RANDOM[7'h70][4:2];
        dataNotInShifter_writeTokenCounter_3 = _RANDOM[7'h70][7:5];
        dataNotInShifter_writeTokenCounter_4 = _RANDOM[7'h70][10:8];
        dataNotInShifter_writeTokenCounter_5 = _RANDOM[7'h70][13:11];
        dataNotInShifter_writeTokenCounter_6 = _RANDOM[7'h70][16:14];
        dataNotInShifter_writeTokenCounter_7 = _RANDOM[7'h70][19:17];
        dataNotInShifter_writeTokenCounter_8 = _RANDOM[7'h70][22:20];
        dataNotInShifter_writeTokenCounter_9 = _RANDOM[7'h70][25:23];
        dataNotInShifter_writeTokenCounter_10 = _RANDOM[7'h70][28:26];
        dataNotInShifter_writeTokenCounter_11 = _RANDOM[7'h70][31:29];
        dataNotInShifter_writeTokenCounter_12 = _RANDOM[7'h71][2:0];
        dataNotInShifter_writeTokenCounter_13 = _RANDOM[7'h71][5:3];
        dataNotInShifter_writeTokenCounter_14 = _RANDOM[7'h71][8:6];
        dataNotInShifter_writeTokenCounter_15 = _RANDOM[7'h71][11:9];
        waiteLastRequest = _RANDOM[7'h71][12];
        waitQueueClear = _RANDOM[7'h71][13];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire              exeRequestQueue_0_empty;
  assign exeRequestQueue_0_empty = _exeRequestQueue_queue_fifo_empty;
  wire              exeRequestQueue_0_full;
  assign exeRequestQueue_0_full = _exeRequestQueue_queue_fifo_full;
  wire              exeRequestQueue_1_empty;
  assign exeRequestQueue_1_empty = _exeRequestQueue_queue_fifo_1_empty;
  wire              exeRequestQueue_1_full;
  assign exeRequestQueue_1_full = _exeRequestQueue_queue_fifo_1_full;
  wire              exeRequestQueue_2_empty;
  assign exeRequestQueue_2_empty = _exeRequestQueue_queue_fifo_2_empty;
  wire              exeRequestQueue_2_full;
  assign exeRequestQueue_2_full = _exeRequestQueue_queue_fifo_2_full;
  wire              exeRequestQueue_3_empty;
  assign exeRequestQueue_3_empty = _exeRequestQueue_queue_fifo_3_empty;
  wire              exeRequestQueue_3_full;
  assign exeRequestQueue_3_full = _exeRequestQueue_queue_fifo_3_full;
  wire              exeRequestQueue_4_empty;
  assign exeRequestQueue_4_empty = _exeRequestQueue_queue_fifo_4_empty;
  wire              exeRequestQueue_4_full;
  assign exeRequestQueue_4_full = _exeRequestQueue_queue_fifo_4_full;
  wire              exeRequestQueue_5_empty;
  assign exeRequestQueue_5_empty = _exeRequestQueue_queue_fifo_5_empty;
  wire              exeRequestQueue_5_full;
  assign exeRequestQueue_5_full = _exeRequestQueue_queue_fifo_5_full;
  wire              exeRequestQueue_6_empty;
  assign exeRequestQueue_6_empty = _exeRequestQueue_queue_fifo_6_empty;
  wire              exeRequestQueue_6_full;
  assign exeRequestQueue_6_full = _exeRequestQueue_queue_fifo_6_full;
  wire              exeRequestQueue_7_empty;
  assign exeRequestQueue_7_empty = _exeRequestQueue_queue_fifo_7_empty;
  wire              exeRequestQueue_7_full;
  assign exeRequestQueue_7_full = _exeRequestQueue_queue_fifo_7_full;
  wire              exeRequestQueue_8_empty;
  assign exeRequestQueue_8_empty = _exeRequestQueue_queue_fifo_8_empty;
  wire              exeRequestQueue_8_full;
  assign exeRequestQueue_8_full = _exeRequestQueue_queue_fifo_8_full;
  wire              exeRequestQueue_9_empty;
  assign exeRequestQueue_9_empty = _exeRequestQueue_queue_fifo_9_empty;
  wire              exeRequestQueue_9_full;
  assign exeRequestQueue_9_full = _exeRequestQueue_queue_fifo_9_full;
  wire              exeRequestQueue_10_empty;
  assign exeRequestQueue_10_empty = _exeRequestQueue_queue_fifo_10_empty;
  wire              exeRequestQueue_10_full;
  assign exeRequestQueue_10_full = _exeRequestQueue_queue_fifo_10_full;
  wire              exeRequestQueue_11_empty;
  assign exeRequestQueue_11_empty = _exeRequestQueue_queue_fifo_11_empty;
  wire              exeRequestQueue_11_full;
  assign exeRequestQueue_11_full = _exeRequestQueue_queue_fifo_11_full;
  wire              exeRequestQueue_12_empty;
  assign exeRequestQueue_12_empty = _exeRequestQueue_queue_fifo_12_empty;
  wire              exeRequestQueue_12_full;
  assign exeRequestQueue_12_full = _exeRequestQueue_queue_fifo_12_full;
  wire              exeRequestQueue_13_empty;
  assign exeRequestQueue_13_empty = _exeRequestQueue_queue_fifo_13_empty;
  wire              exeRequestQueue_13_full;
  assign exeRequestQueue_13_full = _exeRequestQueue_queue_fifo_13_full;
  wire              exeRequestQueue_14_empty;
  assign exeRequestQueue_14_empty = _exeRequestQueue_queue_fifo_14_empty;
  wire              exeRequestQueue_14_full;
  assign exeRequestQueue_14_full = _exeRequestQueue_queue_fifo_14_full;
  wire              exeRequestQueue_15_empty;
  assign exeRequestQueue_15_empty = _exeRequestQueue_queue_fifo_15_empty;
  wire              exeRequestQueue_15_full;
  assign exeRequestQueue_15_full = _exeRequestQueue_queue_fifo_15_full;
  wire              accessCountQueue_empty;
  assign accessCountQueue_empty = _accessCountQueue_fifo_empty;
  wire              accessCountQueue_full;
  assign accessCountQueue_full = _accessCountQueue_fifo_full;
  wire              readWaitQueue_empty;
  assign readWaitQueue_empty = _readWaitQueue_fifo_empty;
  wire              readWaitQueue_full;
  assign readWaitQueue_full = _readWaitQueue_fifo_full;
  assign compressUnitResultQueue_empty = _compressUnitResultQueue_fifo_empty;
  wire              compressUnitResultQueue_full;
  assign compressUnitResultQueue_full = _compressUnitResultQueue_fifo_full;
  wire              reorderQueueVec_0_empty;
  assign reorderQueueVec_0_empty = _reorderQueueVec_fifo_empty;
  wire              reorderQueueVec_0_full;
  assign reorderQueueVec_0_full = _reorderQueueVec_fifo_full;
  wire              reorderQueueVec_1_empty;
  assign reorderQueueVec_1_empty = _reorderQueueVec_fifo_1_empty;
  wire              reorderQueueVec_1_full;
  assign reorderQueueVec_1_full = _reorderQueueVec_fifo_1_full;
  wire              reorderQueueVec_2_empty;
  assign reorderQueueVec_2_empty = _reorderQueueVec_fifo_2_empty;
  wire              reorderQueueVec_2_full;
  assign reorderQueueVec_2_full = _reorderQueueVec_fifo_2_full;
  wire              reorderQueueVec_3_empty;
  assign reorderQueueVec_3_empty = _reorderQueueVec_fifo_3_empty;
  wire              reorderQueueVec_3_full;
  assign reorderQueueVec_3_full = _reorderQueueVec_fifo_3_full;
  wire              reorderQueueVec_4_empty;
  assign reorderQueueVec_4_empty = _reorderQueueVec_fifo_4_empty;
  wire              reorderQueueVec_4_full;
  assign reorderQueueVec_4_full = _reorderQueueVec_fifo_4_full;
  wire              reorderQueueVec_5_empty;
  assign reorderQueueVec_5_empty = _reorderQueueVec_fifo_5_empty;
  wire              reorderQueueVec_5_full;
  assign reorderQueueVec_5_full = _reorderQueueVec_fifo_5_full;
  wire              reorderQueueVec_6_empty;
  assign reorderQueueVec_6_empty = _reorderQueueVec_fifo_6_empty;
  wire              reorderQueueVec_6_full;
  assign reorderQueueVec_6_full = _reorderQueueVec_fifo_6_full;
  wire              reorderQueueVec_7_empty;
  assign reorderQueueVec_7_empty = _reorderQueueVec_fifo_7_empty;
  wire              reorderQueueVec_7_full;
  assign reorderQueueVec_7_full = _reorderQueueVec_fifo_7_full;
  wire              reorderQueueVec_8_empty;
  assign reorderQueueVec_8_empty = _reorderQueueVec_fifo_8_empty;
  wire              reorderQueueVec_8_full;
  assign reorderQueueVec_8_full = _reorderQueueVec_fifo_8_full;
  wire              reorderQueueVec_9_empty;
  assign reorderQueueVec_9_empty = _reorderQueueVec_fifo_9_empty;
  wire              reorderQueueVec_9_full;
  assign reorderQueueVec_9_full = _reorderQueueVec_fifo_9_full;
  wire              reorderQueueVec_10_empty;
  assign reorderQueueVec_10_empty = _reorderQueueVec_fifo_10_empty;
  wire              reorderQueueVec_10_full;
  assign reorderQueueVec_10_full = _reorderQueueVec_fifo_10_full;
  wire              reorderQueueVec_11_empty;
  assign reorderQueueVec_11_empty = _reorderQueueVec_fifo_11_empty;
  wire              reorderQueueVec_11_full;
  assign reorderQueueVec_11_full = _reorderQueueVec_fifo_11_full;
  wire              reorderQueueVec_12_empty;
  assign reorderQueueVec_12_empty = _reorderQueueVec_fifo_12_empty;
  wire              reorderQueueVec_12_full;
  assign reorderQueueVec_12_full = _reorderQueueVec_fifo_12_full;
  wire              reorderQueueVec_13_empty;
  assign reorderQueueVec_13_empty = _reorderQueueVec_fifo_13_empty;
  wire              reorderQueueVec_13_full;
  assign reorderQueueVec_13_full = _reorderQueueVec_fifo_13_full;
  wire              reorderQueueVec_14_empty;
  assign reorderQueueVec_14_empty = _reorderQueueVec_fifo_14_empty;
  wire              reorderQueueVec_14_full;
  assign reorderQueueVec_14_full = _reorderQueueVec_fifo_14_full;
  wire              reorderQueueVec_15_empty;
  assign reorderQueueVec_15_empty = _reorderQueueVec_fifo_15_empty;
  wire              reorderQueueVec_15_full;
  assign reorderQueueVec_15_full = _reorderQueueVec_fifo_15_full;
  wire              readMessageQueue_empty;
  assign readMessageQueue_empty = _readMessageQueue_fifo_empty;
  wire              readMessageQueue_full;
  assign readMessageQueue_full = _readMessageQueue_fifo_full;
  wire              readMessageQueue_1_empty;
  assign readMessageQueue_1_empty = _readMessageQueue_fifo_1_empty;
  wire              readMessageQueue_1_full;
  assign readMessageQueue_1_full = _readMessageQueue_fifo_1_full;
  wire              readMessageQueue_2_empty;
  assign readMessageQueue_2_empty = _readMessageQueue_fifo_2_empty;
  wire              readMessageQueue_2_full;
  assign readMessageQueue_2_full = _readMessageQueue_fifo_2_full;
  wire              readMessageQueue_3_empty;
  assign readMessageQueue_3_empty = _readMessageQueue_fifo_3_empty;
  wire              readMessageQueue_3_full;
  assign readMessageQueue_3_full = _readMessageQueue_fifo_3_full;
  wire              readMessageQueue_4_empty;
  assign readMessageQueue_4_empty = _readMessageQueue_fifo_4_empty;
  wire              readMessageQueue_4_full;
  assign readMessageQueue_4_full = _readMessageQueue_fifo_4_full;
  wire              readMessageQueue_5_empty;
  assign readMessageQueue_5_empty = _readMessageQueue_fifo_5_empty;
  wire              readMessageQueue_5_full;
  assign readMessageQueue_5_full = _readMessageQueue_fifo_5_full;
  wire              readMessageQueue_6_empty;
  assign readMessageQueue_6_empty = _readMessageQueue_fifo_6_empty;
  wire              readMessageQueue_6_full;
  assign readMessageQueue_6_full = _readMessageQueue_fifo_6_full;
  wire              readMessageQueue_7_empty;
  assign readMessageQueue_7_empty = _readMessageQueue_fifo_7_empty;
  wire              readMessageQueue_7_full;
  assign readMessageQueue_7_full = _readMessageQueue_fifo_7_full;
  wire              readMessageQueue_8_empty;
  assign readMessageQueue_8_empty = _readMessageQueue_fifo_8_empty;
  wire              readMessageQueue_8_full;
  assign readMessageQueue_8_full = _readMessageQueue_fifo_8_full;
  wire              readMessageQueue_9_empty;
  assign readMessageQueue_9_empty = _readMessageQueue_fifo_9_empty;
  wire              readMessageQueue_9_full;
  assign readMessageQueue_9_full = _readMessageQueue_fifo_9_full;
  wire              readMessageQueue_10_empty;
  assign readMessageQueue_10_empty = _readMessageQueue_fifo_10_empty;
  wire              readMessageQueue_10_full;
  assign readMessageQueue_10_full = _readMessageQueue_fifo_10_full;
  wire              readMessageQueue_11_empty;
  assign readMessageQueue_11_empty = _readMessageQueue_fifo_11_empty;
  wire              readMessageQueue_11_full;
  assign readMessageQueue_11_full = _readMessageQueue_fifo_11_full;
  wire              readMessageQueue_12_empty;
  assign readMessageQueue_12_empty = _readMessageQueue_fifo_12_empty;
  wire              readMessageQueue_12_full;
  assign readMessageQueue_12_full = _readMessageQueue_fifo_12_full;
  wire              readMessageQueue_13_empty;
  assign readMessageQueue_13_empty = _readMessageQueue_fifo_13_empty;
  wire              readMessageQueue_13_full;
  assign readMessageQueue_13_full = _readMessageQueue_fifo_13_full;
  wire              readMessageQueue_14_empty;
  assign readMessageQueue_14_empty = _readMessageQueue_fifo_14_empty;
  wire              readMessageQueue_14_full;
  assign readMessageQueue_14_full = _readMessageQueue_fifo_14_full;
  wire              readMessageQueue_15_empty;
  assign readMessageQueue_15_empty = _readMessageQueue_fifo_15_empty;
  wire              readMessageQueue_15_full;
  assign readMessageQueue_15_full = _readMessageQueue_fifo_15_full;
  wire              readData_readDataQueue_empty;
  assign readData_readDataQueue_empty = _readData_readDataQueue_fifo_empty;
  wire              readData_readDataQueue_full;
  assign readData_readDataQueue_full = _readData_readDataQueue_fifo_full;
  wire              readData_readDataQueue_1_empty;
  assign readData_readDataQueue_1_empty = _readData_readDataQueue_fifo_1_empty;
  wire              readData_readDataQueue_1_full;
  assign readData_readDataQueue_1_full = _readData_readDataQueue_fifo_1_full;
  wire              readData_readDataQueue_2_empty;
  assign readData_readDataQueue_2_empty = _readData_readDataQueue_fifo_2_empty;
  wire              readData_readDataQueue_2_full;
  assign readData_readDataQueue_2_full = _readData_readDataQueue_fifo_2_full;
  wire              readData_readDataQueue_3_empty;
  assign readData_readDataQueue_3_empty = _readData_readDataQueue_fifo_3_empty;
  wire              readData_readDataQueue_3_full;
  assign readData_readDataQueue_3_full = _readData_readDataQueue_fifo_3_full;
  wire              readData_readDataQueue_4_empty;
  assign readData_readDataQueue_4_empty = _readData_readDataQueue_fifo_4_empty;
  wire              readData_readDataQueue_4_full;
  assign readData_readDataQueue_4_full = _readData_readDataQueue_fifo_4_full;
  wire              readData_readDataQueue_5_empty;
  assign readData_readDataQueue_5_empty = _readData_readDataQueue_fifo_5_empty;
  wire              readData_readDataQueue_5_full;
  assign readData_readDataQueue_5_full = _readData_readDataQueue_fifo_5_full;
  wire              readData_readDataQueue_6_empty;
  assign readData_readDataQueue_6_empty = _readData_readDataQueue_fifo_6_empty;
  wire              readData_readDataQueue_6_full;
  assign readData_readDataQueue_6_full = _readData_readDataQueue_fifo_6_full;
  wire              readData_readDataQueue_7_empty;
  assign readData_readDataQueue_7_empty = _readData_readDataQueue_fifo_7_empty;
  wire              readData_readDataQueue_7_full;
  assign readData_readDataQueue_7_full = _readData_readDataQueue_fifo_7_full;
  wire              readData_readDataQueue_8_empty;
  assign readData_readDataQueue_8_empty = _readData_readDataQueue_fifo_8_empty;
  wire              readData_readDataQueue_8_full;
  assign readData_readDataQueue_8_full = _readData_readDataQueue_fifo_8_full;
  wire              readData_readDataQueue_9_empty;
  assign readData_readDataQueue_9_empty = _readData_readDataQueue_fifo_9_empty;
  wire              readData_readDataQueue_9_full;
  assign readData_readDataQueue_9_full = _readData_readDataQueue_fifo_9_full;
  wire              readData_readDataQueue_10_empty;
  assign readData_readDataQueue_10_empty = _readData_readDataQueue_fifo_10_empty;
  wire              readData_readDataQueue_10_full;
  assign readData_readDataQueue_10_full = _readData_readDataQueue_fifo_10_full;
  wire              readData_readDataQueue_11_empty;
  assign readData_readDataQueue_11_empty = _readData_readDataQueue_fifo_11_empty;
  wire              readData_readDataQueue_11_full;
  assign readData_readDataQueue_11_full = _readData_readDataQueue_fifo_11_full;
  wire              readData_readDataQueue_12_empty;
  assign readData_readDataQueue_12_empty = _readData_readDataQueue_fifo_12_empty;
  wire              readData_readDataQueue_12_full;
  assign readData_readDataQueue_12_full = _readData_readDataQueue_fifo_12_full;
  wire              readData_readDataQueue_13_empty;
  assign readData_readDataQueue_13_empty = _readData_readDataQueue_fifo_13_empty;
  wire              readData_readDataQueue_13_full;
  assign readData_readDataQueue_13_full = _readData_readDataQueue_fifo_13_full;
  wire              readData_readDataQueue_14_empty;
  assign readData_readDataQueue_14_empty = _readData_readDataQueue_fifo_14_empty;
  wire              readData_readDataQueue_14_full;
  assign readData_readDataQueue_14_full = _readData_readDataQueue_fifo_14_full;
  wire              readData_readDataQueue_15_empty;
  assign readData_readDataQueue_15_empty = _readData_readDataQueue_fifo_15_empty;
  wire              readData_readDataQueue_15_full;
  assign readData_readDataQueue_15_full = _readData_readDataQueue_fifo_15_full;
  assign compressUnitResultQueue_enq_valid = _compressUnit_out_compressValid;
  assign compressUnitResultQueue_enq_bits_compressValid = _compressUnit_out_compressValid;
  wire              writeQueue_0_empty;
  assign writeQueue_0_empty = _writeQueue_fifo_empty;
  wire              writeQueue_0_full;
  assign writeQueue_0_full = _writeQueue_fifo_full;
  wire              writeQueue_1_empty;
  assign writeQueue_1_empty = _writeQueue_fifo_1_empty;
  wire              writeQueue_1_full;
  assign writeQueue_1_full = _writeQueue_fifo_1_full;
  wire              writeQueue_2_empty;
  assign writeQueue_2_empty = _writeQueue_fifo_2_empty;
  wire              writeQueue_2_full;
  assign writeQueue_2_full = _writeQueue_fifo_2_full;
  wire              writeQueue_3_empty;
  assign writeQueue_3_empty = _writeQueue_fifo_3_empty;
  wire              writeQueue_3_full;
  assign writeQueue_3_full = _writeQueue_fifo_3_full;
  wire              writeQueue_4_empty;
  assign writeQueue_4_empty = _writeQueue_fifo_4_empty;
  wire              writeQueue_4_full;
  assign writeQueue_4_full = _writeQueue_fifo_4_full;
  wire              writeQueue_5_empty;
  assign writeQueue_5_empty = _writeQueue_fifo_5_empty;
  wire              writeQueue_5_full;
  assign writeQueue_5_full = _writeQueue_fifo_5_full;
  wire              writeQueue_6_empty;
  assign writeQueue_6_empty = _writeQueue_fifo_6_empty;
  wire              writeQueue_6_full;
  assign writeQueue_6_full = _writeQueue_fifo_6_full;
  wire              writeQueue_7_empty;
  assign writeQueue_7_empty = _writeQueue_fifo_7_empty;
  wire              writeQueue_7_full;
  assign writeQueue_7_full = _writeQueue_fifo_7_full;
  wire              writeQueue_8_empty;
  assign writeQueue_8_empty = _writeQueue_fifo_8_empty;
  wire              writeQueue_8_full;
  assign writeQueue_8_full = _writeQueue_fifo_8_full;
  wire              writeQueue_9_empty;
  assign writeQueue_9_empty = _writeQueue_fifo_9_empty;
  wire              writeQueue_9_full;
  assign writeQueue_9_full = _writeQueue_fifo_9_full;
  wire              writeQueue_10_empty;
  assign writeQueue_10_empty = _writeQueue_fifo_10_empty;
  wire              writeQueue_10_full;
  assign writeQueue_10_full = _writeQueue_fifo_10_full;
  wire              writeQueue_11_empty;
  assign writeQueue_11_empty = _writeQueue_fifo_11_empty;
  wire              writeQueue_11_full;
  assign writeQueue_11_full = _writeQueue_fifo_11_full;
  wire              writeQueue_12_empty;
  assign writeQueue_12_empty = _writeQueue_fifo_12_empty;
  wire              writeQueue_12_full;
  assign writeQueue_12_full = _writeQueue_fifo_12_full;
  wire              writeQueue_13_empty;
  assign writeQueue_13_empty = _writeQueue_fifo_13_empty;
  wire              writeQueue_13_full;
  assign writeQueue_13_full = _writeQueue_fifo_13_full;
  wire              writeQueue_14_empty;
  assign writeQueue_14_empty = _writeQueue_fifo_14_empty;
  wire              writeQueue_14_full;
  assign writeQueue_14_full = _writeQueue_fifo_14_full;
  wire              writeQueue_15_empty;
  assign writeQueue_15_empty = _writeQueue_fifo_15_empty;
  wire              writeQueue_15_full;
  assign writeQueue_15_full = _writeQueue_fifo_15_full;
  BitLevelMaskWrite maskedWrite (
    .clock                              (clock),
    .reset                              (reset),
    .needWAR                            (maskDestinationType),
    .vd                                 (instReg_vd),
    .in_0_ready                         (_maskedWrite_in_0_ready),
    .in_0_valid                         (unitType[2] ? _reduceUnit_out_valid : executeValid & maskFilter),
    .in_0_bits_data                     (unitType[2] ? _reduceUnit_out_bits_data : executeResult[31:0]),
    .in_0_bits_bitMask                  (currentMaskGroupForDestination[31:0]),
    .in_0_bits_mask                     (unitType[2] ? _reduceUnit_out_bits_mask : executeWriteByteMask[3:0]),
    .in_0_bits_groupCounter             (unitType[2] ? 5'h0 : executeDeqGroupCounter[4:0]),
    .in_0_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[0] & ffo),
    .in_1_ready                         (_maskedWrite_in_1_ready),
    .in_1_valid                         (executeValid & maskFilter_1),
    .in_1_bits_data                     (executeResult[63:32]),
    .in_1_bits_bitMask                  (currentMaskGroupForDestination[63:32]),
    .in_1_bits_mask                     (executeWriteByteMask[7:4]),
    .in_1_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_1_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[1] & ffo),
    .in_2_ready                         (_maskedWrite_in_2_ready),
    .in_2_valid                         (executeValid & maskFilter_2),
    .in_2_bits_data                     (executeResult[95:64]),
    .in_2_bits_bitMask                  (currentMaskGroupForDestination[95:64]),
    .in_2_bits_mask                     (executeWriteByteMask[11:8]),
    .in_2_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_2_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[2] & ffo),
    .in_3_ready                         (_maskedWrite_in_3_ready),
    .in_3_valid                         (executeValid & maskFilter_3),
    .in_3_bits_data                     (executeResult[127:96]),
    .in_3_bits_bitMask                  (currentMaskGroupForDestination[127:96]),
    .in_3_bits_mask                     (executeWriteByteMask[15:12]),
    .in_3_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_3_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[3] & ffo),
    .in_4_ready                         (_maskedWrite_in_4_ready),
    .in_4_valid                         (executeValid & maskFilter_4),
    .in_4_bits_data                     (executeResult[159:128]),
    .in_4_bits_bitMask                  (currentMaskGroupForDestination[159:128]),
    .in_4_bits_mask                     (executeWriteByteMask[19:16]),
    .in_4_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_4_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[4] & ffo),
    .in_5_ready                         (_maskedWrite_in_5_ready),
    .in_5_valid                         (executeValid & maskFilter_5),
    .in_5_bits_data                     (executeResult[191:160]),
    .in_5_bits_bitMask                  (currentMaskGroupForDestination[191:160]),
    .in_5_bits_mask                     (executeWriteByteMask[23:20]),
    .in_5_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_5_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[5] & ffo),
    .in_6_ready                         (_maskedWrite_in_6_ready),
    .in_6_valid                         (executeValid & maskFilter_6),
    .in_6_bits_data                     (executeResult[223:192]),
    .in_6_bits_bitMask                  (currentMaskGroupForDestination[223:192]),
    .in_6_bits_mask                     (executeWriteByteMask[27:24]),
    .in_6_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_6_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[6] & ffo),
    .in_7_ready                         (_maskedWrite_in_7_ready),
    .in_7_valid                         (executeValid & maskFilter_7),
    .in_7_bits_data                     (executeResult[255:224]),
    .in_7_bits_bitMask                  (currentMaskGroupForDestination[255:224]),
    .in_7_bits_mask                     (executeWriteByteMask[31:28]),
    .in_7_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_7_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[7] & ffo),
    .in_8_ready                         (_maskedWrite_in_8_ready),
    .in_8_valid                         (executeValid & maskFilter_8),
    .in_8_bits_data                     (executeResult[287:256]),
    .in_8_bits_bitMask                  (currentMaskGroupForDestination[287:256]),
    .in_8_bits_mask                     (executeWriteByteMask[35:32]),
    .in_8_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_8_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[8] & ffo),
    .in_9_ready                         (_maskedWrite_in_9_ready),
    .in_9_valid                         (executeValid & maskFilter_9),
    .in_9_bits_data                     (executeResult[319:288]),
    .in_9_bits_bitMask                  (currentMaskGroupForDestination[319:288]),
    .in_9_bits_mask                     (executeWriteByteMask[39:36]),
    .in_9_bits_groupCounter             (executeDeqGroupCounter[4:0]),
    .in_9_bits_ffoByOther               (compressUnitResultQueue_deq_bits_ffoOutput[9] & ffo),
    .in_10_ready                        (_maskedWrite_in_10_ready),
    .in_10_valid                        (executeValid & maskFilter_10),
    .in_10_bits_data                    (executeResult[351:320]),
    .in_10_bits_bitMask                 (currentMaskGroupForDestination[351:320]),
    .in_10_bits_mask                    (executeWriteByteMask[43:40]),
    .in_10_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_10_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[10] & ffo),
    .in_11_ready                        (_maskedWrite_in_11_ready),
    .in_11_valid                        (executeValid & maskFilter_11),
    .in_11_bits_data                    (executeResult[383:352]),
    .in_11_bits_bitMask                 (currentMaskGroupForDestination[383:352]),
    .in_11_bits_mask                    (executeWriteByteMask[47:44]),
    .in_11_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_11_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[11] & ffo),
    .in_12_ready                        (_maskedWrite_in_12_ready),
    .in_12_valid                        (executeValid & maskFilter_12),
    .in_12_bits_data                    (executeResult[415:384]),
    .in_12_bits_bitMask                 (currentMaskGroupForDestination[415:384]),
    .in_12_bits_mask                    (executeWriteByteMask[51:48]),
    .in_12_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_12_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[12] & ffo),
    .in_13_ready                        (_maskedWrite_in_13_ready),
    .in_13_valid                        (executeValid & maskFilter_13),
    .in_13_bits_data                    (executeResult[447:416]),
    .in_13_bits_bitMask                 (currentMaskGroupForDestination[447:416]),
    .in_13_bits_mask                    (executeWriteByteMask[55:52]),
    .in_13_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_13_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[13] & ffo),
    .in_14_ready                        (_maskedWrite_in_14_ready),
    .in_14_valid                        (executeValid & maskFilter_14),
    .in_14_bits_data                    (executeResult[479:448]),
    .in_14_bits_bitMask                 (currentMaskGroupForDestination[479:448]),
    .in_14_bits_mask                    (executeWriteByteMask[59:56]),
    .in_14_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_14_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[14] & ffo),
    .in_15_ready                        (_maskedWrite_in_15_ready),
    .in_15_valid                        (executeValid & maskFilter_15),
    .in_15_bits_data                    (executeResult[511:480]),
    .in_15_bits_bitMask                 (currentMaskGroupForDestination[511:480]),
    .in_15_bits_mask                    (executeWriteByteMask[63:60]),
    .in_15_bits_groupCounter            (executeDeqGroupCounter[4:0]),
    .in_15_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[15] & ffo),
    .out_0_ready                        (writeQueue_0_enq_ready),
    .out_0_valid                        (_maskedWrite_out_0_valid),
    .out_0_bits_ffoByOther              (_maskedWrite_out_0_bits_ffoByOther),
    .out_0_bits_writeData_data          (_maskedWrite_out_0_bits_writeData_data),
    .out_0_bits_writeData_mask          (_maskedWrite_out_0_bits_writeData_mask),
    .out_0_bits_writeData_groupCounter  (_maskedWrite_out_0_bits_writeData_groupCounter),
    .out_1_ready                        (writeQueue_1_enq_ready),
    .out_1_valid                        (_maskedWrite_out_1_valid),
    .out_1_bits_ffoByOther              (_maskedWrite_out_1_bits_ffoByOther),
    .out_1_bits_writeData_data          (_maskedWrite_out_1_bits_writeData_data),
    .out_1_bits_writeData_mask          (_maskedWrite_out_1_bits_writeData_mask),
    .out_1_bits_writeData_groupCounter  (_maskedWrite_out_1_bits_writeData_groupCounter),
    .out_2_ready                        (writeQueue_2_enq_ready),
    .out_2_valid                        (_maskedWrite_out_2_valid),
    .out_2_bits_ffoByOther              (_maskedWrite_out_2_bits_ffoByOther),
    .out_2_bits_writeData_data          (_maskedWrite_out_2_bits_writeData_data),
    .out_2_bits_writeData_mask          (_maskedWrite_out_2_bits_writeData_mask),
    .out_2_bits_writeData_groupCounter  (_maskedWrite_out_2_bits_writeData_groupCounter),
    .out_3_ready                        (writeQueue_3_enq_ready),
    .out_3_valid                        (_maskedWrite_out_3_valid),
    .out_3_bits_ffoByOther              (_maskedWrite_out_3_bits_ffoByOther),
    .out_3_bits_writeData_data          (_maskedWrite_out_3_bits_writeData_data),
    .out_3_bits_writeData_mask          (_maskedWrite_out_3_bits_writeData_mask),
    .out_3_bits_writeData_groupCounter  (_maskedWrite_out_3_bits_writeData_groupCounter),
    .out_4_ready                        (writeQueue_4_enq_ready),
    .out_4_valid                        (_maskedWrite_out_4_valid),
    .out_4_bits_ffoByOther              (_maskedWrite_out_4_bits_ffoByOther),
    .out_4_bits_writeData_data          (_maskedWrite_out_4_bits_writeData_data),
    .out_4_bits_writeData_mask          (_maskedWrite_out_4_bits_writeData_mask),
    .out_4_bits_writeData_groupCounter  (_maskedWrite_out_4_bits_writeData_groupCounter),
    .out_5_ready                        (writeQueue_5_enq_ready),
    .out_5_valid                        (_maskedWrite_out_5_valid),
    .out_5_bits_ffoByOther              (_maskedWrite_out_5_bits_ffoByOther),
    .out_5_bits_writeData_data          (_maskedWrite_out_5_bits_writeData_data),
    .out_5_bits_writeData_mask          (_maskedWrite_out_5_bits_writeData_mask),
    .out_5_bits_writeData_groupCounter  (_maskedWrite_out_5_bits_writeData_groupCounter),
    .out_6_ready                        (writeQueue_6_enq_ready),
    .out_6_valid                        (_maskedWrite_out_6_valid),
    .out_6_bits_ffoByOther              (_maskedWrite_out_6_bits_ffoByOther),
    .out_6_bits_writeData_data          (_maskedWrite_out_6_bits_writeData_data),
    .out_6_bits_writeData_mask          (_maskedWrite_out_6_bits_writeData_mask),
    .out_6_bits_writeData_groupCounter  (_maskedWrite_out_6_bits_writeData_groupCounter),
    .out_7_ready                        (writeQueue_7_enq_ready),
    .out_7_valid                        (_maskedWrite_out_7_valid),
    .out_7_bits_ffoByOther              (_maskedWrite_out_7_bits_ffoByOther),
    .out_7_bits_writeData_data          (_maskedWrite_out_7_bits_writeData_data),
    .out_7_bits_writeData_mask          (_maskedWrite_out_7_bits_writeData_mask),
    .out_7_bits_writeData_groupCounter  (_maskedWrite_out_7_bits_writeData_groupCounter),
    .out_8_ready                        (writeQueue_8_enq_ready),
    .out_8_valid                        (_maskedWrite_out_8_valid),
    .out_8_bits_ffoByOther              (_maskedWrite_out_8_bits_ffoByOther),
    .out_8_bits_writeData_data          (_maskedWrite_out_8_bits_writeData_data),
    .out_8_bits_writeData_mask          (_maskedWrite_out_8_bits_writeData_mask),
    .out_8_bits_writeData_groupCounter  (_maskedWrite_out_8_bits_writeData_groupCounter),
    .out_9_ready                        (writeQueue_9_enq_ready),
    .out_9_valid                        (_maskedWrite_out_9_valid),
    .out_9_bits_ffoByOther              (_maskedWrite_out_9_bits_ffoByOther),
    .out_9_bits_writeData_data          (_maskedWrite_out_9_bits_writeData_data),
    .out_9_bits_writeData_mask          (_maskedWrite_out_9_bits_writeData_mask),
    .out_9_bits_writeData_groupCounter  (_maskedWrite_out_9_bits_writeData_groupCounter),
    .out_10_ready                       (writeQueue_10_enq_ready),
    .out_10_valid                       (_maskedWrite_out_10_valid),
    .out_10_bits_ffoByOther             (_maskedWrite_out_10_bits_ffoByOther),
    .out_10_bits_writeData_data         (_maskedWrite_out_10_bits_writeData_data),
    .out_10_bits_writeData_mask         (_maskedWrite_out_10_bits_writeData_mask),
    .out_10_bits_writeData_groupCounter (_maskedWrite_out_10_bits_writeData_groupCounter),
    .out_11_ready                       (writeQueue_11_enq_ready),
    .out_11_valid                       (_maskedWrite_out_11_valid),
    .out_11_bits_ffoByOther             (_maskedWrite_out_11_bits_ffoByOther),
    .out_11_bits_writeData_data         (_maskedWrite_out_11_bits_writeData_data),
    .out_11_bits_writeData_mask         (_maskedWrite_out_11_bits_writeData_mask),
    .out_11_bits_writeData_groupCounter (_maskedWrite_out_11_bits_writeData_groupCounter),
    .out_12_ready                       (writeQueue_12_enq_ready),
    .out_12_valid                       (_maskedWrite_out_12_valid),
    .out_12_bits_ffoByOther             (_maskedWrite_out_12_bits_ffoByOther),
    .out_12_bits_writeData_data         (_maskedWrite_out_12_bits_writeData_data),
    .out_12_bits_writeData_mask         (_maskedWrite_out_12_bits_writeData_mask),
    .out_12_bits_writeData_groupCounter (_maskedWrite_out_12_bits_writeData_groupCounter),
    .out_13_ready                       (writeQueue_13_enq_ready),
    .out_13_valid                       (_maskedWrite_out_13_valid),
    .out_13_bits_ffoByOther             (_maskedWrite_out_13_bits_ffoByOther),
    .out_13_bits_writeData_data         (_maskedWrite_out_13_bits_writeData_data),
    .out_13_bits_writeData_mask         (_maskedWrite_out_13_bits_writeData_mask),
    .out_13_bits_writeData_groupCounter (_maskedWrite_out_13_bits_writeData_groupCounter),
    .out_14_ready                       (writeQueue_14_enq_ready),
    .out_14_valid                       (_maskedWrite_out_14_valid),
    .out_14_bits_ffoByOther             (_maskedWrite_out_14_bits_ffoByOther),
    .out_14_bits_writeData_data         (_maskedWrite_out_14_bits_writeData_data),
    .out_14_bits_writeData_mask         (_maskedWrite_out_14_bits_writeData_mask),
    .out_14_bits_writeData_groupCounter (_maskedWrite_out_14_bits_writeData_groupCounter),
    .out_15_ready                       (writeQueue_15_enq_ready),
    .out_15_valid                       (_maskedWrite_out_15_valid),
    .out_15_bits_ffoByOther             (_maskedWrite_out_15_bits_ffoByOther),
    .out_15_bits_writeData_data         (_maskedWrite_out_15_bits_writeData_data),
    .out_15_bits_writeData_mask         (_maskedWrite_out_15_bits_writeData_mask),
    .out_15_bits_writeData_groupCounter (_maskedWrite_out_15_bits_writeData_groupCounter),
    .readChannel_0_ready                (readChannel_0_ready_0),
    .readChannel_0_valid                (_maskedWrite_readChannel_0_valid),
    .readChannel_0_bits_vs              (_maskedWrite_readChannel_0_bits_vs),
    .readChannel_0_bits_offset          (_maskedWrite_readChannel_0_bits_offset),
    .readChannel_1_ready                (readChannel_1_ready_0),
    .readChannel_1_valid                (_maskedWrite_readChannel_1_valid),
    .readChannel_1_bits_vs              (_maskedWrite_readChannel_1_bits_vs),
    .readChannel_1_bits_offset          (_maskedWrite_readChannel_1_bits_offset),
    .readChannel_2_ready                (readChannel_2_ready_0),
    .readChannel_2_valid                (_maskedWrite_readChannel_2_valid),
    .readChannel_2_bits_vs              (_maskedWrite_readChannel_2_bits_vs),
    .readChannel_2_bits_offset          (_maskedWrite_readChannel_2_bits_offset),
    .readChannel_3_ready                (readChannel_3_ready_0),
    .readChannel_3_valid                (_maskedWrite_readChannel_3_valid),
    .readChannel_3_bits_vs              (_maskedWrite_readChannel_3_bits_vs),
    .readChannel_3_bits_offset          (_maskedWrite_readChannel_3_bits_offset),
    .readChannel_4_ready                (readChannel_4_ready_0),
    .readChannel_4_valid                (_maskedWrite_readChannel_4_valid),
    .readChannel_4_bits_vs              (_maskedWrite_readChannel_4_bits_vs),
    .readChannel_4_bits_offset          (_maskedWrite_readChannel_4_bits_offset),
    .readChannel_5_ready                (readChannel_5_ready_0),
    .readChannel_5_valid                (_maskedWrite_readChannel_5_valid),
    .readChannel_5_bits_vs              (_maskedWrite_readChannel_5_bits_vs),
    .readChannel_5_bits_offset          (_maskedWrite_readChannel_5_bits_offset),
    .readChannel_6_ready                (readChannel_6_ready_0),
    .readChannel_6_valid                (_maskedWrite_readChannel_6_valid),
    .readChannel_6_bits_vs              (_maskedWrite_readChannel_6_bits_vs),
    .readChannel_6_bits_offset          (_maskedWrite_readChannel_6_bits_offset),
    .readChannel_7_ready                (readChannel_7_ready_0),
    .readChannel_7_valid                (_maskedWrite_readChannel_7_valid),
    .readChannel_7_bits_vs              (_maskedWrite_readChannel_7_bits_vs),
    .readChannel_7_bits_offset          (_maskedWrite_readChannel_7_bits_offset),
    .readChannel_8_ready                (readChannel_8_ready_0),
    .readChannel_8_valid                (_maskedWrite_readChannel_8_valid),
    .readChannel_8_bits_vs              (_maskedWrite_readChannel_8_bits_vs),
    .readChannel_8_bits_offset          (_maskedWrite_readChannel_8_bits_offset),
    .readChannel_9_ready                (readChannel_9_ready_0),
    .readChannel_9_valid                (_maskedWrite_readChannel_9_valid),
    .readChannel_9_bits_vs              (_maskedWrite_readChannel_9_bits_vs),
    .readChannel_9_bits_offset          (_maskedWrite_readChannel_9_bits_offset),
    .readChannel_10_ready               (readChannel_10_ready_0),
    .readChannel_10_valid               (_maskedWrite_readChannel_10_valid),
    .readChannel_10_bits_vs             (_maskedWrite_readChannel_10_bits_vs),
    .readChannel_10_bits_offset         (_maskedWrite_readChannel_10_bits_offset),
    .readChannel_11_ready               (readChannel_11_ready_0),
    .readChannel_11_valid               (_maskedWrite_readChannel_11_valid),
    .readChannel_11_bits_vs             (_maskedWrite_readChannel_11_bits_vs),
    .readChannel_11_bits_offset         (_maskedWrite_readChannel_11_bits_offset),
    .readChannel_12_ready               (readChannel_12_ready_0),
    .readChannel_12_valid               (_maskedWrite_readChannel_12_valid),
    .readChannel_12_bits_vs             (_maskedWrite_readChannel_12_bits_vs),
    .readChannel_12_bits_offset         (_maskedWrite_readChannel_12_bits_offset),
    .readChannel_13_ready               (readChannel_13_ready_0),
    .readChannel_13_valid               (_maskedWrite_readChannel_13_valid),
    .readChannel_13_bits_vs             (_maskedWrite_readChannel_13_bits_vs),
    .readChannel_13_bits_offset         (_maskedWrite_readChannel_13_bits_offset),
    .readChannel_14_ready               (readChannel_14_ready_0),
    .readChannel_14_valid               (_maskedWrite_readChannel_14_valid),
    .readChannel_14_bits_vs             (_maskedWrite_readChannel_14_bits_vs),
    .readChannel_14_bits_offset         (_maskedWrite_readChannel_14_bits_offset),
    .readChannel_15_ready               (readChannel_15_ready_0),
    .readChannel_15_valid               (_maskedWrite_readChannel_15_valid),
    .readChannel_15_bits_vs             (_maskedWrite_readChannel_15_bits_vs),
    .readChannel_15_bits_offset         (_maskedWrite_readChannel_15_bits_offset),
    .readResult_0_valid                 (readResult_0_valid),
    .readResult_0_bits                  (readResult_0_bits),
    .readResult_1_valid                 (readResult_1_valid),
    .readResult_1_bits                  (readResult_1_bits),
    .readResult_2_valid                 (readResult_2_valid),
    .readResult_2_bits                  (readResult_2_bits),
    .readResult_3_valid                 (readResult_3_valid),
    .readResult_3_bits                  (readResult_3_bits),
    .readResult_4_valid                 (readResult_4_valid),
    .readResult_4_bits                  (readResult_4_bits),
    .readResult_5_valid                 (readResult_5_valid),
    .readResult_5_bits                  (readResult_5_bits),
    .readResult_6_valid                 (readResult_6_valid),
    .readResult_6_bits                  (readResult_6_bits),
    .readResult_7_valid                 (readResult_7_valid),
    .readResult_7_bits                  (readResult_7_bits),
    .readResult_8_valid                 (readResult_8_valid),
    .readResult_8_bits                  (readResult_8_bits),
    .readResult_9_valid                 (readResult_9_valid),
    .readResult_9_bits                  (readResult_9_bits),
    .readResult_10_valid                (readResult_10_valid),
    .readResult_10_bits                 (readResult_10_bits),
    .readResult_11_valid                (readResult_11_valid),
    .readResult_11_bits                 (readResult_11_bits),
    .readResult_12_valid                (readResult_12_valid),
    .readResult_12_bits                 (readResult_12_bits),
    .readResult_13_valid                (readResult_13_valid),
    .readResult_13_bits                 (readResult_13_bits),
    .readResult_14_valid                (readResult_14_valid),
    .readResult_14_bits                 (readResult_14_bits),
    .readResult_15_valid                (readResult_15_valid),
    .readResult_15_bits                 (readResult_15_bits),
    .stageClear                         (_maskedWrite_stageClear)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_0_enq_ready & exeRequestQueue_0_enq_valid & ~(_exeRequestQueue_queue_fifo_empty & exeRequestQueue_0_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_0_deq_ready & ~_exeRequestQueue_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn),
    .empty        (_exeRequestQueue_queue_fifo_empty),
    .almost_empty (exeRequestQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_0_almostFull),
    .full         (_exeRequestQueue_queue_fifo_full),
    .error        (_exeRequestQueue_queue_fifo_error),
    .data_out     (_exeRequestQueue_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_1_enq_ready & exeRequestQueue_1_enq_valid & ~(_exeRequestQueue_queue_fifo_1_empty & exeRequestQueue_1_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_1_deq_ready & ~_exeRequestQueue_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_1),
    .empty        (_exeRequestQueue_queue_fifo_1_empty),
    .almost_empty (exeRequestQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_1_almostFull),
    .full         (_exeRequestQueue_queue_fifo_1_full),
    .error        (_exeRequestQueue_queue_fifo_1_error),
    .data_out     (_exeRequestQueue_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_2_enq_ready & exeRequestQueue_2_enq_valid & ~(_exeRequestQueue_queue_fifo_2_empty & exeRequestQueue_2_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_2_deq_ready & ~_exeRequestQueue_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_2),
    .empty        (_exeRequestQueue_queue_fifo_2_empty),
    .almost_empty (exeRequestQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_2_almostFull),
    .full         (_exeRequestQueue_queue_fifo_2_full),
    .error        (_exeRequestQueue_queue_fifo_2_error),
    .data_out     (_exeRequestQueue_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_3_enq_ready & exeRequestQueue_3_enq_valid & ~(_exeRequestQueue_queue_fifo_3_empty & exeRequestQueue_3_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_3_deq_ready & ~_exeRequestQueue_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_3),
    .empty        (_exeRequestQueue_queue_fifo_3_empty),
    .almost_empty (exeRequestQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_3_almostFull),
    .full         (_exeRequestQueue_queue_fifo_3_full),
    .error        (_exeRequestQueue_queue_fifo_3_error),
    .data_out     (_exeRequestQueue_queue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_4_enq_ready & exeRequestQueue_4_enq_valid & ~(_exeRequestQueue_queue_fifo_4_empty & exeRequestQueue_4_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_4_deq_ready & ~_exeRequestQueue_queue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_4),
    .empty        (_exeRequestQueue_queue_fifo_4_empty),
    .almost_empty (exeRequestQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_4_almostFull),
    .full         (_exeRequestQueue_queue_fifo_4_full),
    .error        (_exeRequestQueue_queue_fifo_4_error),
    .data_out     (_exeRequestQueue_queue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_5_enq_ready & exeRequestQueue_5_enq_valid & ~(_exeRequestQueue_queue_fifo_5_empty & exeRequestQueue_5_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_5_deq_ready & ~_exeRequestQueue_queue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_5),
    .empty        (_exeRequestQueue_queue_fifo_5_empty),
    .almost_empty (exeRequestQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_5_almostFull),
    .full         (_exeRequestQueue_queue_fifo_5_full),
    .error        (_exeRequestQueue_queue_fifo_5_error),
    .data_out     (_exeRequestQueue_queue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_6_enq_ready & exeRequestQueue_6_enq_valid & ~(_exeRequestQueue_queue_fifo_6_empty & exeRequestQueue_6_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_6_deq_ready & ~_exeRequestQueue_queue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_6),
    .empty        (_exeRequestQueue_queue_fifo_6_empty),
    .almost_empty (exeRequestQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_6_almostFull),
    .full         (_exeRequestQueue_queue_fifo_6_full),
    .error        (_exeRequestQueue_queue_fifo_6_error),
    .data_out     (_exeRequestQueue_queue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_7_enq_ready & exeRequestQueue_7_enq_valid & ~(_exeRequestQueue_queue_fifo_7_empty & exeRequestQueue_7_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_7_deq_ready & ~_exeRequestQueue_queue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_7),
    .empty        (_exeRequestQueue_queue_fifo_7_empty),
    .almost_empty (exeRequestQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_7_almostFull),
    .full         (_exeRequestQueue_queue_fifo_7_full),
    .error        (_exeRequestQueue_queue_fifo_7_error),
    .data_out     (_exeRequestQueue_queue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_8_enq_ready & exeRequestQueue_8_enq_valid & ~(_exeRequestQueue_queue_fifo_8_empty & exeRequestQueue_8_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_8_deq_ready & ~_exeRequestQueue_queue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_8),
    .empty        (_exeRequestQueue_queue_fifo_8_empty),
    .almost_empty (exeRequestQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_8_almostFull),
    .full         (_exeRequestQueue_queue_fifo_8_full),
    .error        (_exeRequestQueue_queue_fifo_8_error),
    .data_out     (_exeRequestQueue_queue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_9_enq_ready & exeRequestQueue_9_enq_valid & ~(_exeRequestQueue_queue_fifo_9_empty & exeRequestQueue_9_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_9_deq_ready & ~_exeRequestQueue_queue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_9),
    .empty        (_exeRequestQueue_queue_fifo_9_empty),
    .almost_empty (exeRequestQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_9_almostFull),
    .full         (_exeRequestQueue_queue_fifo_9_full),
    .error        (_exeRequestQueue_queue_fifo_9_error),
    .data_out     (_exeRequestQueue_queue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_10_enq_ready & exeRequestQueue_10_enq_valid & ~(_exeRequestQueue_queue_fifo_10_empty & exeRequestQueue_10_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_10_deq_ready & ~_exeRequestQueue_queue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_10),
    .empty        (_exeRequestQueue_queue_fifo_10_empty),
    .almost_empty (exeRequestQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_10_almostFull),
    .full         (_exeRequestQueue_queue_fifo_10_full),
    .error        (_exeRequestQueue_queue_fifo_10_error),
    .data_out     (_exeRequestQueue_queue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_11_enq_ready & exeRequestQueue_11_enq_valid & ~(_exeRequestQueue_queue_fifo_11_empty & exeRequestQueue_11_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_11_deq_ready & ~_exeRequestQueue_queue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_11),
    .empty        (_exeRequestQueue_queue_fifo_11_empty),
    .almost_empty (exeRequestQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_11_almostFull),
    .full         (_exeRequestQueue_queue_fifo_11_full),
    .error        (_exeRequestQueue_queue_fifo_11_error),
    .data_out     (_exeRequestQueue_queue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_12_enq_ready & exeRequestQueue_12_enq_valid & ~(_exeRequestQueue_queue_fifo_12_empty & exeRequestQueue_12_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_12_deq_ready & ~_exeRequestQueue_queue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_12),
    .empty        (_exeRequestQueue_queue_fifo_12_empty),
    .almost_empty (exeRequestQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_12_almostFull),
    .full         (_exeRequestQueue_queue_fifo_12_full),
    .error        (_exeRequestQueue_queue_fifo_12_error),
    .data_out     (_exeRequestQueue_queue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_13_enq_ready & exeRequestQueue_13_enq_valid & ~(_exeRequestQueue_queue_fifo_13_empty & exeRequestQueue_13_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_13_deq_ready & ~_exeRequestQueue_queue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_13),
    .empty        (_exeRequestQueue_queue_fifo_13_empty),
    .almost_empty (exeRequestQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_13_almostFull),
    .full         (_exeRequestQueue_queue_fifo_13_full),
    .error        (_exeRequestQueue_queue_fifo_13_error),
    .data_out     (_exeRequestQueue_queue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_14_enq_ready & exeRequestQueue_14_enq_valid & ~(_exeRequestQueue_queue_fifo_14_empty & exeRequestQueue_14_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_14_deq_ready & ~_exeRequestQueue_queue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_14),
    .empty        (_exeRequestQueue_queue_fifo_14_empty),
    .almost_empty (exeRequestQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_14_almostFull),
    .full         (_exeRequestQueue_queue_fifo_14_full),
    .error        (_exeRequestQueue_queue_fifo_14_error),
    .data_out     (_exeRequestQueue_queue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(69)
  ) exeRequestQueue_queue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_15_enq_ready & exeRequestQueue_15_enq_valid & ~(_exeRequestQueue_queue_fifo_15_empty & exeRequestQueue_15_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_15_deq_ready & ~_exeRequestQueue_queue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_15),
    .empty        (_exeRequestQueue_queue_fifo_15_empty),
    .almost_empty (exeRequestQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_15_almostFull),
    .full         (_exeRequestQueue_queue_fifo_15_full),
    .error        (_exeRequestQueue_queue_fifo_15_error),
    .data_out     (_exeRequestQueue_queue_fifo_15_data_out)
  );
  SlideIndexGen slideAddressGen (
    .clock                              (clock),
    .reset                              (reset),
    .newInstruction                     (instReq_valid & (|instReq_bits_vl)),
    .instructionReq_decodeResult_topUop (instReg_decodeResult_topUop),
    .instructionReq_readFromScala       (instReg_readFromScala),
    .instructionReq_sew                 (instReg_sew),
    .instructionReq_vlmul               (instReg_vlmul),
    .instructionReq_maskType            (instReg_maskType),
    .instructionReq_vl                  (instReg_vl),
    .indexDeq_ready                     (slideAddressGen_indexDeq_ready),
    .indexDeq_valid                     (_slideAddressGen_indexDeq_valid),
    .indexDeq_bits_needRead             (_slideAddressGen_indexDeq_bits_needRead),
    .indexDeq_bits_elementValid         (_slideAddressGen_indexDeq_bits_elementValid),
    .indexDeq_bits_replaceVs1           (_slideAddressGen_indexDeq_bits_replaceVs1),
    .indexDeq_bits_readOffset           (_slideAddressGen_indexDeq_bits_readOffset),
    .indexDeq_bits_accessLane_0         (_slideAddressGen_indexDeq_bits_accessLane_0),
    .indexDeq_bits_accessLane_1         (_slideAddressGen_indexDeq_bits_accessLane_1),
    .indexDeq_bits_accessLane_2         (_slideAddressGen_indexDeq_bits_accessLane_2),
    .indexDeq_bits_accessLane_3         (_slideAddressGen_indexDeq_bits_accessLane_3),
    .indexDeq_bits_accessLane_4         (_slideAddressGen_indexDeq_bits_accessLane_4),
    .indexDeq_bits_accessLane_5         (_slideAddressGen_indexDeq_bits_accessLane_5),
    .indexDeq_bits_accessLane_6         (_slideAddressGen_indexDeq_bits_accessLane_6),
    .indexDeq_bits_accessLane_7         (_slideAddressGen_indexDeq_bits_accessLane_7),
    .indexDeq_bits_accessLane_8         (_slideAddressGen_indexDeq_bits_accessLane_8),
    .indexDeq_bits_accessLane_9         (_slideAddressGen_indexDeq_bits_accessLane_9),
    .indexDeq_bits_accessLane_10        (_slideAddressGen_indexDeq_bits_accessLane_10),
    .indexDeq_bits_accessLane_11        (_slideAddressGen_indexDeq_bits_accessLane_11),
    .indexDeq_bits_accessLane_12        (_slideAddressGen_indexDeq_bits_accessLane_12),
    .indexDeq_bits_accessLane_13        (_slideAddressGen_indexDeq_bits_accessLane_13),
    .indexDeq_bits_accessLane_14        (_slideAddressGen_indexDeq_bits_accessLane_14),
    .indexDeq_bits_accessLane_15        (_slideAddressGen_indexDeq_bits_accessLane_15),
    .indexDeq_bits_vsGrowth_0           (_slideAddressGen_indexDeq_bits_vsGrowth_0),
    .indexDeq_bits_vsGrowth_1           (_slideAddressGen_indexDeq_bits_vsGrowth_1),
    .indexDeq_bits_vsGrowth_2           (_slideAddressGen_indexDeq_bits_vsGrowth_2),
    .indexDeq_bits_vsGrowth_3           (_slideAddressGen_indexDeq_bits_vsGrowth_3),
    .indexDeq_bits_vsGrowth_4           (_slideAddressGen_indexDeq_bits_vsGrowth_4),
    .indexDeq_bits_vsGrowth_5           (_slideAddressGen_indexDeq_bits_vsGrowth_5),
    .indexDeq_bits_vsGrowth_6           (_slideAddressGen_indexDeq_bits_vsGrowth_6),
    .indexDeq_bits_vsGrowth_7           (_slideAddressGen_indexDeq_bits_vsGrowth_7),
    .indexDeq_bits_vsGrowth_8           (_slideAddressGen_indexDeq_bits_vsGrowth_8),
    .indexDeq_bits_vsGrowth_9           (_slideAddressGen_indexDeq_bits_vsGrowth_9),
    .indexDeq_bits_vsGrowth_10          (_slideAddressGen_indexDeq_bits_vsGrowth_10),
    .indexDeq_bits_vsGrowth_11          (_slideAddressGen_indexDeq_bits_vsGrowth_11),
    .indexDeq_bits_vsGrowth_12          (_slideAddressGen_indexDeq_bits_vsGrowth_12),
    .indexDeq_bits_vsGrowth_13          (_slideAddressGen_indexDeq_bits_vsGrowth_13),
    .indexDeq_bits_vsGrowth_14          (_slideAddressGen_indexDeq_bits_vsGrowth_14),
    .indexDeq_bits_vsGrowth_15          (_slideAddressGen_indexDeq_bits_vsGrowth_15),
    .indexDeq_bits_executeGroup         (_slideAddressGen_indexDeq_bits_executeGroup),
    .indexDeq_bits_readDataOffset       (_slideAddressGen_indexDeq_bits_readDataOffset),
    .indexDeq_bits_last                 (_slideAddressGen_indexDeq_bits_last),
    .slideGroupOut                      (_slideAddressGen_slideGroupOut),
    .slideMaskInput                     (_GEN_40[_slideAddressGen_slideGroupOut[5:0]])
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(80)
  ) accessCountQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(accessCountQueue_enq_ready & accessCountQueue_enq_valid)),
    .pop_req_n    (~(accessCountQueue_deq_ready & ~_accessCountQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (accessCountQueue_dataIn),
    .empty        (_accessCountQueue_fifo_empty),
    .almost_empty (accessCountQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (accessCountQueue_almostFull),
    .full         (_accessCountQueue_fifo_full),
    .error        (_accessCountQueue_fifo_error),
    .data_out     (_accessCountQueue_fifo_data_out)
  );
  MaskUnitReadCrossBar readCrossBar (
    .input_0_ready             (_readCrossBar_input_0_ready),
    .input_0_valid             (readCrossBar_input_0_valid),
    .input_0_bits_vs           (selectExecuteReq_0_bits_vs),
    .input_0_bits_offset       (selectExecuteReq_0_bits_offset),
    .input_0_bits_readLane     (selectExecuteReq_0_bits_readLane),
    .input_0_bits_dataOffset   (selectExecuteReq_0_bits_dataOffset),
    .input_1_ready             (_readCrossBar_input_1_ready),
    .input_1_valid             (readCrossBar_input_1_valid),
    .input_1_bits_vs           (selectExecuteReq_1_bits_vs),
    .input_1_bits_offset       (selectExecuteReq_1_bits_offset),
    .input_1_bits_readLane     (selectExecuteReq_1_bits_readLane),
    .input_1_bits_dataOffset   (selectExecuteReq_1_bits_dataOffset),
    .input_2_ready             (_readCrossBar_input_2_ready),
    .input_2_valid             (readCrossBar_input_2_valid),
    .input_2_bits_vs           (selectExecuteReq_2_bits_vs),
    .input_2_bits_offset       (selectExecuteReq_2_bits_offset),
    .input_2_bits_readLane     (selectExecuteReq_2_bits_readLane),
    .input_2_bits_dataOffset   (selectExecuteReq_2_bits_dataOffset),
    .input_3_ready             (_readCrossBar_input_3_ready),
    .input_3_valid             (readCrossBar_input_3_valid),
    .input_3_bits_vs           (selectExecuteReq_3_bits_vs),
    .input_3_bits_offset       (selectExecuteReq_3_bits_offset),
    .input_3_bits_readLane     (selectExecuteReq_3_bits_readLane),
    .input_3_bits_dataOffset   (selectExecuteReq_3_bits_dataOffset),
    .input_4_ready             (_readCrossBar_input_4_ready),
    .input_4_valid             (readCrossBar_input_4_valid),
    .input_4_bits_vs           (selectExecuteReq_4_bits_vs),
    .input_4_bits_offset       (selectExecuteReq_4_bits_offset),
    .input_4_bits_readLane     (selectExecuteReq_4_bits_readLane),
    .input_4_bits_dataOffset   (selectExecuteReq_4_bits_dataOffset),
    .input_5_ready             (_readCrossBar_input_5_ready),
    .input_5_valid             (readCrossBar_input_5_valid),
    .input_5_bits_vs           (selectExecuteReq_5_bits_vs),
    .input_5_bits_offset       (selectExecuteReq_5_bits_offset),
    .input_5_bits_readLane     (selectExecuteReq_5_bits_readLane),
    .input_5_bits_dataOffset   (selectExecuteReq_5_bits_dataOffset),
    .input_6_ready             (_readCrossBar_input_6_ready),
    .input_6_valid             (readCrossBar_input_6_valid),
    .input_6_bits_vs           (selectExecuteReq_6_bits_vs),
    .input_6_bits_offset       (selectExecuteReq_6_bits_offset),
    .input_6_bits_readLane     (selectExecuteReq_6_bits_readLane),
    .input_6_bits_dataOffset   (selectExecuteReq_6_bits_dataOffset),
    .input_7_ready             (_readCrossBar_input_7_ready),
    .input_7_valid             (readCrossBar_input_7_valid),
    .input_7_bits_vs           (selectExecuteReq_7_bits_vs),
    .input_7_bits_offset       (selectExecuteReq_7_bits_offset),
    .input_7_bits_readLane     (selectExecuteReq_7_bits_readLane),
    .input_7_bits_dataOffset   (selectExecuteReq_7_bits_dataOffset),
    .input_8_ready             (_readCrossBar_input_8_ready),
    .input_8_valid             (readCrossBar_input_8_valid),
    .input_8_bits_vs           (selectExecuteReq_8_bits_vs),
    .input_8_bits_offset       (selectExecuteReq_8_bits_offset),
    .input_8_bits_readLane     (selectExecuteReq_8_bits_readLane),
    .input_8_bits_dataOffset   (selectExecuteReq_8_bits_dataOffset),
    .input_9_ready             (_readCrossBar_input_9_ready),
    .input_9_valid             (readCrossBar_input_9_valid),
    .input_9_bits_vs           (selectExecuteReq_9_bits_vs),
    .input_9_bits_offset       (selectExecuteReq_9_bits_offset),
    .input_9_bits_readLane     (selectExecuteReq_9_bits_readLane),
    .input_9_bits_dataOffset   (selectExecuteReq_9_bits_dataOffset),
    .input_10_ready            (_readCrossBar_input_10_ready),
    .input_10_valid            (readCrossBar_input_10_valid),
    .input_10_bits_vs          (selectExecuteReq_10_bits_vs),
    .input_10_bits_offset      (selectExecuteReq_10_bits_offset),
    .input_10_bits_readLane    (selectExecuteReq_10_bits_readLane),
    .input_10_bits_dataOffset  (selectExecuteReq_10_bits_dataOffset),
    .input_11_ready            (_readCrossBar_input_11_ready),
    .input_11_valid            (readCrossBar_input_11_valid),
    .input_11_bits_vs          (selectExecuteReq_11_bits_vs),
    .input_11_bits_offset      (selectExecuteReq_11_bits_offset),
    .input_11_bits_readLane    (selectExecuteReq_11_bits_readLane),
    .input_11_bits_dataOffset  (selectExecuteReq_11_bits_dataOffset),
    .input_12_ready            (_readCrossBar_input_12_ready),
    .input_12_valid            (readCrossBar_input_12_valid),
    .input_12_bits_vs          (selectExecuteReq_12_bits_vs),
    .input_12_bits_offset      (selectExecuteReq_12_bits_offset),
    .input_12_bits_readLane    (selectExecuteReq_12_bits_readLane),
    .input_12_bits_dataOffset  (selectExecuteReq_12_bits_dataOffset),
    .input_13_ready            (_readCrossBar_input_13_ready),
    .input_13_valid            (readCrossBar_input_13_valid),
    .input_13_bits_vs          (selectExecuteReq_13_bits_vs),
    .input_13_bits_offset      (selectExecuteReq_13_bits_offset),
    .input_13_bits_readLane    (selectExecuteReq_13_bits_readLane),
    .input_13_bits_dataOffset  (selectExecuteReq_13_bits_dataOffset),
    .input_14_ready            (_readCrossBar_input_14_ready),
    .input_14_valid            (readCrossBar_input_14_valid),
    .input_14_bits_vs          (selectExecuteReq_14_bits_vs),
    .input_14_bits_offset      (selectExecuteReq_14_bits_offset),
    .input_14_bits_readLane    (selectExecuteReq_14_bits_readLane),
    .input_14_bits_dataOffset  (selectExecuteReq_14_bits_dataOffset),
    .input_15_ready            (_readCrossBar_input_15_ready),
    .input_15_valid            (readCrossBar_input_15_valid),
    .input_15_bits_vs          (selectExecuteReq_15_bits_vs),
    .input_15_bits_offset      (selectExecuteReq_15_bits_offset),
    .input_15_bits_readLane    (selectExecuteReq_15_bits_readLane),
    .input_15_bits_dataOffset  (selectExecuteReq_15_bits_dataOffset),
    .output_0_ready            (readChannel_0_ready_0 & readMessageQueue_enq_ready),
    .output_0_valid            (_readCrossBar_output_0_valid),
    .output_0_bits_vs          (_readCrossBar_output_0_bits_vs),
    .output_0_bits_offset      (_readCrossBar_output_0_bits_offset),
    .output_0_bits_writeIndex  (_readCrossBar_output_0_bits_writeIndex),
    .output_0_bits_dataOffset  (readMessageQueue_enq_bits_dataOffset),
    .output_1_ready            (readChannel_1_ready_0 & readMessageQueue_1_enq_ready),
    .output_1_valid            (_readCrossBar_output_1_valid),
    .output_1_bits_vs          (_readCrossBar_output_1_bits_vs),
    .output_1_bits_offset      (_readCrossBar_output_1_bits_offset),
    .output_1_bits_writeIndex  (_readCrossBar_output_1_bits_writeIndex),
    .output_1_bits_dataOffset  (readMessageQueue_1_enq_bits_dataOffset),
    .output_2_ready            (readChannel_2_ready_0 & readMessageQueue_2_enq_ready),
    .output_2_valid            (_readCrossBar_output_2_valid),
    .output_2_bits_vs          (_readCrossBar_output_2_bits_vs),
    .output_2_bits_offset      (_readCrossBar_output_2_bits_offset),
    .output_2_bits_writeIndex  (_readCrossBar_output_2_bits_writeIndex),
    .output_2_bits_dataOffset  (readMessageQueue_2_enq_bits_dataOffset),
    .output_3_ready            (readChannel_3_ready_0 & readMessageQueue_3_enq_ready),
    .output_3_valid            (_readCrossBar_output_3_valid),
    .output_3_bits_vs          (_readCrossBar_output_3_bits_vs),
    .output_3_bits_offset      (_readCrossBar_output_3_bits_offset),
    .output_3_bits_writeIndex  (_readCrossBar_output_3_bits_writeIndex),
    .output_3_bits_dataOffset  (readMessageQueue_3_enq_bits_dataOffset),
    .output_4_ready            (readChannel_4_ready_0 & readMessageQueue_4_enq_ready),
    .output_4_valid            (_readCrossBar_output_4_valid),
    .output_4_bits_vs          (_readCrossBar_output_4_bits_vs),
    .output_4_bits_offset      (_readCrossBar_output_4_bits_offset),
    .output_4_bits_writeIndex  (_readCrossBar_output_4_bits_writeIndex),
    .output_4_bits_dataOffset  (readMessageQueue_4_enq_bits_dataOffset),
    .output_5_ready            (readChannel_5_ready_0 & readMessageQueue_5_enq_ready),
    .output_5_valid            (_readCrossBar_output_5_valid),
    .output_5_bits_vs          (_readCrossBar_output_5_bits_vs),
    .output_5_bits_offset      (_readCrossBar_output_5_bits_offset),
    .output_5_bits_writeIndex  (_readCrossBar_output_5_bits_writeIndex),
    .output_5_bits_dataOffset  (readMessageQueue_5_enq_bits_dataOffset),
    .output_6_ready            (readChannel_6_ready_0 & readMessageQueue_6_enq_ready),
    .output_6_valid            (_readCrossBar_output_6_valid),
    .output_6_bits_vs          (_readCrossBar_output_6_bits_vs),
    .output_6_bits_offset      (_readCrossBar_output_6_bits_offset),
    .output_6_bits_writeIndex  (_readCrossBar_output_6_bits_writeIndex),
    .output_6_bits_dataOffset  (readMessageQueue_6_enq_bits_dataOffset),
    .output_7_ready            (readChannel_7_ready_0 & readMessageQueue_7_enq_ready),
    .output_7_valid            (_readCrossBar_output_7_valid),
    .output_7_bits_vs          (_readCrossBar_output_7_bits_vs),
    .output_7_bits_offset      (_readCrossBar_output_7_bits_offset),
    .output_7_bits_writeIndex  (_readCrossBar_output_7_bits_writeIndex),
    .output_7_bits_dataOffset  (readMessageQueue_7_enq_bits_dataOffset),
    .output_8_ready            (readChannel_8_ready_0 & readMessageQueue_8_enq_ready),
    .output_8_valid            (_readCrossBar_output_8_valid),
    .output_8_bits_vs          (_readCrossBar_output_8_bits_vs),
    .output_8_bits_offset      (_readCrossBar_output_8_bits_offset),
    .output_8_bits_writeIndex  (_readCrossBar_output_8_bits_writeIndex),
    .output_8_bits_dataOffset  (readMessageQueue_8_enq_bits_dataOffset),
    .output_9_ready            (readChannel_9_ready_0 & readMessageQueue_9_enq_ready),
    .output_9_valid            (_readCrossBar_output_9_valid),
    .output_9_bits_vs          (_readCrossBar_output_9_bits_vs),
    .output_9_bits_offset      (_readCrossBar_output_9_bits_offset),
    .output_9_bits_writeIndex  (_readCrossBar_output_9_bits_writeIndex),
    .output_9_bits_dataOffset  (readMessageQueue_9_enq_bits_dataOffset),
    .output_10_ready           (readChannel_10_ready_0 & readMessageQueue_10_enq_ready),
    .output_10_valid           (_readCrossBar_output_10_valid),
    .output_10_bits_vs         (_readCrossBar_output_10_bits_vs),
    .output_10_bits_offset     (_readCrossBar_output_10_bits_offset),
    .output_10_bits_writeIndex (_readCrossBar_output_10_bits_writeIndex),
    .output_10_bits_dataOffset (readMessageQueue_10_enq_bits_dataOffset),
    .output_11_ready           (readChannel_11_ready_0 & readMessageQueue_11_enq_ready),
    .output_11_valid           (_readCrossBar_output_11_valid),
    .output_11_bits_vs         (_readCrossBar_output_11_bits_vs),
    .output_11_bits_offset     (_readCrossBar_output_11_bits_offset),
    .output_11_bits_writeIndex (_readCrossBar_output_11_bits_writeIndex),
    .output_11_bits_dataOffset (readMessageQueue_11_enq_bits_dataOffset),
    .output_12_ready           (readChannel_12_ready_0 & readMessageQueue_12_enq_ready),
    .output_12_valid           (_readCrossBar_output_12_valid),
    .output_12_bits_vs         (_readCrossBar_output_12_bits_vs),
    .output_12_bits_offset     (_readCrossBar_output_12_bits_offset),
    .output_12_bits_writeIndex (_readCrossBar_output_12_bits_writeIndex),
    .output_12_bits_dataOffset (readMessageQueue_12_enq_bits_dataOffset),
    .output_13_ready           (readChannel_13_ready_0 & readMessageQueue_13_enq_ready),
    .output_13_valid           (_readCrossBar_output_13_valid),
    .output_13_bits_vs         (_readCrossBar_output_13_bits_vs),
    .output_13_bits_offset     (_readCrossBar_output_13_bits_offset),
    .output_13_bits_writeIndex (_readCrossBar_output_13_bits_writeIndex),
    .output_13_bits_dataOffset (readMessageQueue_13_enq_bits_dataOffset),
    .output_14_ready           (readChannel_14_ready_0 & readMessageQueue_14_enq_ready),
    .output_14_valid           (_readCrossBar_output_14_valid),
    .output_14_bits_vs         (_readCrossBar_output_14_bits_vs),
    .output_14_bits_offset     (_readCrossBar_output_14_bits_offset),
    .output_14_bits_writeIndex (_readCrossBar_output_14_bits_writeIndex),
    .output_14_bits_dataOffset (readMessageQueue_14_enq_bits_dataOffset),
    .output_15_ready           (readChannel_15_ready_0 & readMessageQueue_15_enq_ready),
    .output_15_valid           (_readCrossBar_output_15_valid),
    .output_15_bits_vs         (_readCrossBar_output_15_bits_vs),
    .output_15_bits_offset     (_readCrossBar_output_15_bits_offset),
    .output_15_bits_writeIndex (_readCrossBar_output_15_bits_writeIndex),
    .output_15_bits_dataOffset (readMessageQueue_15_enq_bits_dataOffset)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(56)
  ) readWaitQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readWaitQueue_enq_ready & readWaitQueue_enq_valid)),
    .pop_req_n    (~(readWaitQueue_deq_ready & ~_readWaitQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readWaitQueue_dataIn),
    .empty        (_readWaitQueue_fifo_empty),
    .almost_empty (readWaitQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readWaitQueue_almostFull),
    .full         (_readWaitQueue_fifo_full),
    .error        (_readWaitQueue_fifo_error),
    .data_out     (_readWaitQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(598)
  ) compressUnitResultQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(compressUnitResultQueue_enq_ready & compressUnitResultQueue_enq_valid & ~(_compressUnitResultQueue_fifo_empty & compressUnitResultQueue_deq_ready))),
    .pop_req_n    (~(compressUnitResultQueue_deq_ready & ~_compressUnitResultQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (compressUnitResultQueue_dataIn),
    .empty        (_compressUnitResultQueue_fifo_empty),
    .almost_empty (compressUnitResultQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (compressUnitResultQueue_almostFull),
    .full         (_compressUnitResultQueue_fifo_full),
    .error        (_compressUnitResultQueue_fifo_error),
    .data_out     (_compressUnitResultQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_0_enq_ready & reorderQueueVec_0_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_0_deq_ready & ~_reorderQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn),
    .empty        (_reorderQueueVec_fifo_empty),
    .almost_empty (reorderQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_0_almostFull),
    .full         (_reorderQueueVec_fifo_full),
    .error        (_reorderQueueVec_fifo_error),
    .data_out     (_reorderQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_1_enq_ready & reorderQueueVec_1_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_1_deq_ready & ~_reorderQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_1),
    .empty        (_reorderQueueVec_fifo_1_empty),
    .almost_empty (reorderQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_1_almostFull),
    .full         (_reorderQueueVec_fifo_1_full),
    .error        (_reorderQueueVec_fifo_1_error),
    .data_out     (_reorderQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_2_enq_ready & reorderQueueVec_2_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_2_deq_ready & ~_reorderQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_2),
    .empty        (_reorderQueueVec_fifo_2_empty),
    .almost_empty (reorderQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_2_almostFull),
    .full         (_reorderQueueVec_fifo_2_full),
    .error        (_reorderQueueVec_fifo_2_error),
    .data_out     (_reorderQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_3_enq_ready & reorderQueueVec_3_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_3_deq_ready & ~_reorderQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_3),
    .empty        (_reorderQueueVec_fifo_3_empty),
    .almost_empty (reorderQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_3_almostFull),
    .full         (_reorderQueueVec_fifo_3_full),
    .error        (_reorderQueueVec_fifo_3_error),
    .data_out     (_reorderQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_4_enq_ready & reorderQueueVec_4_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_4_deq_ready & ~_reorderQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_4),
    .empty        (_reorderQueueVec_fifo_4_empty),
    .almost_empty (reorderQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_4_almostFull),
    .full         (_reorderQueueVec_fifo_4_full),
    .error        (_reorderQueueVec_fifo_4_error),
    .data_out     (_reorderQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_5_enq_ready & reorderQueueVec_5_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_5_deq_ready & ~_reorderQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_5),
    .empty        (_reorderQueueVec_fifo_5_empty),
    .almost_empty (reorderQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_5_almostFull),
    .full         (_reorderQueueVec_fifo_5_full),
    .error        (_reorderQueueVec_fifo_5_error),
    .data_out     (_reorderQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_6_enq_ready & reorderQueueVec_6_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_6_deq_ready & ~_reorderQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_6),
    .empty        (_reorderQueueVec_fifo_6_empty),
    .almost_empty (reorderQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_6_almostFull),
    .full         (_reorderQueueVec_fifo_6_full),
    .error        (_reorderQueueVec_fifo_6_error),
    .data_out     (_reorderQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_7_enq_ready & reorderQueueVec_7_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_7_deq_ready & ~_reorderQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_7),
    .empty        (_reorderQueueVec_fifo_7_empty),
    .almost_empty (reorderQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_7_almostFull),
    .full         (_reorderQueueVec_fifo_7_full),
    .error        (_reorderQueueVec_fifo_7_error),
    .data_out     (_reorderQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_8_enq_ready & reorderQueueVec_8_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_8_deq_ready & ~_reorderQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_8),
    .empty        (_reorderQueueVec_fifo_8_empty),
    .almost_empty (reorderQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_8_almostFull),
    .full         (_reorderQueueVec_fifo_8_full),
    .error        (_reorderQueueVec_fifo_8_error),
    .data_out     (_reorderQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_9_enq_ready & reorderQueueVec_9_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_9_deq_ready & ~_reorderQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_9),
    .empty        (_reorderQueueVec_fifo_9_empty),
    .almost_empty (reorderQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_9_almostFull),
    .full         (_reorderQueueVec_fifo_9_full),
    .error        (_reorderQueueVec_fifo_9_error),
    .data_out     (_reorderQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_10_enq_ready & reorderQueueVec_10_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_10_deq_ready & ~_reorderQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_10),
    .empty        (_reorderQueueVec_fifo_10_empty),
    .almost_empty (reorderQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_10_almostFull),
    .full         (_reorderQueueVec_fifo_10_full),
    .error        (_reorderQueueVec_fifo_10_error),
    .data_out     (_reorderQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_11_enq_ready & reorderQueueVec_11_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_11_deq_ready & ~_reorderQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_11),
    .empty        (_reorderQueueVec_fifo_11_empty),
    .almost_empty (reorderQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_11_almostFull),
    .full         (_reorderQueueVec_fifo_11_full),
    .error        (_reorderQueueVec_fifo_11_error),
    .data_out     (_reorderQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_12_enq_ready & reorderQueueVec_12_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_12_deq_ready & ~_reorderQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_12),
    .empty        (_reorderQueueVec_fifo_12_empty),
    .almost_empty (reorderQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_12_almostFull),
    .full         (_reorderQueueVec_fifo_12_full),
    .error        (_reorderQueueVec_fifo_12_error),
    .data_out     (_reorderQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_13_enq_ready & reorderQueueVec_13_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_13_deq_ready & ~_reorderQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_13),
    .empty        (_reorderQueueVec_fifo_13_empty),
    .almost_empty (reorderQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_13_almostFull),
    .full         (_reorderQueueVec_fifo_13_full),
    .error        (_reorderQueueVec_fifo_13_error),
    .data_out     (_reorderQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_14_enq_ready & reorderQueueVec_14_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_14_deq_ready & ~_reorderQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_14),
    .empty        (_reorderQueueVec_fifo_14_empty),
    .almost_empty (reorderQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_14_almostFull),
    .full         (_reorderQueueVec_fifo_14_full),
    .error        (_reorderQueueVec_fifo_14_error),
    .data_out     (_reorderQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(48)
  ) reorderQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_15_enq_ready & reorderQueueVec_15_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_15_deq_ready & ~_reorderQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_15),
    .empty        (_reorderQueueVec_fifo_15_empty),
    .almost_empty (reorderQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_15_almostFull),
    .full         (_reorderQueueVec_fifo_15_full),
    .error        (_reorderQueueVec_fifo_15_error),
    .data_out     (_reorderQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_enq_ready & readMessageQueue_enq_valid)),
    .pop_req_n    (~(readMessageQueue_deq_ready & ~_readMessageQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn),
    .empty        (_readMessageQueue_fifo_empty),
    .almost_empty (readMessageQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_almostFull),
    .full         (_readMessageQueue_fifo_full),
    .error        (_readMessageQueue_fifo_error),
    .data_out     (_readMessageQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_1_enq_ready & readMessageQueue_1_enq_valid)),
    .pop_req_n    (~(readMessageQueue_1_deq_ready & ~_readMessageQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_1),
    .empty        (_readMessageQueue_fifo_1_empty),
    .almost_empty (readMessageQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_1_almostFull),
    .full         (_readMessageQueue_fifo_1_full),
    .error        (_readMessageQueue_fifo_1_error),
    .data_out     (_readMessageQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_2_enq_ready & readMessageQueue_2_enq_valid)),
    .pop_req_n    (~(readMessageQueue_2_deq_ready & ~_readMessageQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_2),
    .empty        (_readMessageQueue_fifo_2_empty),
    .almost_empty (readMessageQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_2_almostFull),
    .full         (_readMessageQueue_fifo_2_full),
    .error        (_readMessageQueue_fifo_2_error),
    .data_out     (_readMessageQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_3_enq_ready & readMessageQueue_3_enq_valid)),
    .pop_req_n    (~(readMessageQueue_3_deq_ready & ~_readMessageQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_3),
    .empty        (_readMessageQueue_fifo_3_empty),
    .almost_empty (readMessageQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_3_almostFull),
    .full         (_readMessageQueue_fifo_3_full),
    .error        (_readMessageQueue_fifo_3_error),
    .data_out     (_readMessageQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_4_enq_ready & readMessageQueue_4_enq_valid)),
    .pop_req_n    (~(readMessageQueue_4_deq_ready & ~_readMessageQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_4),
    .empty        (_readMessageQueue_fifo_4_empty),
    .almost_empty (readMessageQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_4_almostFull),
    .full         (_readMessageQueue_fifo_4_full),
    .error        (_readMessageQueue_fifo_4_error),
    .data_out     (_readMessageQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_5_enq_ready & readMessageQueue_5_enq_valid)),
    .pop_req_n    (~(readMessageQueue_5_deq_ready & ~_readMessageQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_5),
    .empty        (_readMessageQueue_fifo_5_empty),
    .almost_empty (readMessageQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_5_almostFull),
    .full         (_readMessageQueue_fifo_5_full),
    .error        (_readMessageQueue_fifo_5_error),
    .data_out     (_readMessageQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_6_enq_ready & readMessageQueue_6_enq_valid)),
    .pop_req_n    (~(readMessageQueue_6_deq_ready & ~_readMessageQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_6),
    .empty        (_readMessageQueue_fifo_6_empty),
    .almost_empty (readMessageQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_6_almostFull),
    .full         (_readMessageQueue_fifo_6_full),
    .error        (_readMessageQueue_fifo_6_error),
    .data_out     (_readMessageQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_7_enq_ready & readMessageQueue_7_enq_valid)),
    .pop_req_n    (~(readMessageQueue_7_deq_ready & ~_readMessageQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_7),
    .empty        (_readMessageQueue_fifo_7_empty),
    .almost_empty (readMessageQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_7_almostFull),
    .full         (_readMessageQueue_fifo_7_full),
    .error        (_readMessageQueue_fifo_7_error),
    .data_out     (_readMessageQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_8_enq_ready & readMessageQueue_8_enq_valid)),
    .pop_req_n    (~(readMessageQueue_8_deq_ready & ~_readMessageQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_8),
    .empty        (_readMessageQueue_fifo_8_empty),
    .almost_empty (readMessageQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_8_almostFull),
    .full         (_readMessageQueue_fifo_8_full),
    .error        (_readMessageQueue_fifo_8_error),
    .data_out     (_readMessageQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_9_enq_ready & readMessageQueue_9_enq_valid)),
    .pop_req_n    (~(readMessageQueue_9_deq_ready & ~_readMessageQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_9),
    .empty        (_readMessageQueue_fifo_9_empty),
    .almost_empty (readMessageQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_9_almostFull),
    .full         (_readMessageQueue_fifo_9_full),
    .error        (_readMessageQueue_fifo_9_error),
    .data_out     (_readMessageQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_10_enq_ready & readMessageQueue_10_enq_valid)),
    .pop_req_n    (~(readMessageQueue_10_deq_ready & ~_readMessageQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_10),
    .empty        (_readMessageQueue_fifo_10_empty),
    .almost_empty (readMessageQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_10_almostFull),
    .full         (_readMessageQueue_fifo_10_full),
    .error        (_readMessageQueue_fifo_10_error),
    .data_out     (_readMessageQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_11_enq_ready & readMessageQueue_11_enq_valid)),
    .pop_req_n    (~(readMessageQueue_11_deq_ready & ~_readMessageQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_11),
    .empty        (_readMessageQueue_fifo_11_empty),
    .almost_empty (readMessageQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_11_almostFull),
    .full         (_readMessageQueue_fifo_11_full),
    .error        (_readMessageQueue_fifo_11_error),
    .data_out     (_readMessageQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_12_enq_ready & readMessageQueue_12_enq_valid)),
    .pop_req_n    (~(readMessageQueue_12_deq_ready & ~_readMessageQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_12),
    .empty        (_readMessageQueue_fifo_12_empty),
    .almost_empty (readMessageQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_12_almostFull),
    .full         (_readMessageQueue_fifo_12_full),
    .error        (_readMessageQueue_fifo_12_error),
    .data_out     (_readMessageQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_13_enq_ready & readMessageQueue_13_enq_valid)),
    .pop_req_n    (~(readMessageQueue_13_deq_ready & ~_readMessageQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_13),
    .empty        (_readMessageQueue_fifo_13_empty),
    .almost_empty (readMessageQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_13_almostFull),
    .full         (_readMessageQueue_fifo_13_full),
    .error        (_readMessageQueue_fifo_13_error),
    .data_out     (_readMessageQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_14_enq_ready & readMessageQueue_14_enq_valid)),
    .pop_req_n    (~(readMessageQueue_14_deq_ready & ~_readMessageQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_14),
    .empty        (_readMessageQueue_fifo_14_empty),
    .almost_empty (readMessageQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_14_almostFull),
    .full         (_readMessageQueue_fifo_14_full),
    .error        (_readMessageQueue_fifo_14_error),
    .data_out     (_readMessageQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(18)
  ) readMessageQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_15_enq_ready & readMessageQueue_15_enq_valid)),
    .pop_req_n    (~(readMessageQueue_15_deq_ready & ~_readMessageQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_15),
    .empty        (_readMessageQueue_fifo_15_empty),
    .almost_empty (readMessageQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_15_almostFull),
    .full         (_readMessageQueue_fifo_15_full),
    .error        (_readMessageQueue_fifo_15_error),
    .data_out     (_readMessageQueue_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_enq_ready & readData_readDataQueue_enq_valid & ~(_readData_readDataQueue_fifo_empty & readData_readDataQueue_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_deq_ready & ~_readData_readDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_enq_bits),
    .empty        (_readData_readDataQueue_fifo_empty),
    .almost_empty (readData_readDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_almostFull),
    .full         (_readData_readDataQueue_fifo_full),
    .error        (_readData_readDataQueue_fifo_error),
    .data_out     (_readData_readDataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_1_enq_ready & readData_readDataQueue_1_enq_valid & ~(_readData_readDataQueue_fifo_1_empty & readData_readDataQueue_1_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_1_deq_ready & ~_readData_readDataQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_1_enq_bits),
    .empty        (_readData_readDataQueue_fifo_1_empty),
    .almost_empty (readData_readDataQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_1_almostFull),
    .full         (_readData_readDataQueue_fifo_1_full),
    .error        (_readData_readDataQueue_fifo_1_error),
    .data_out     (_readData_readDataQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_2_enq_ready & readData_readDataQueue_2_enq_valid & ~(_readData_readDataQueue_fifo_2_empty & readData_readDataQueue_2_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_2_deq_ready & ~_readData_readDataQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_2_enq_bits),
    .empty        (_readData_readDataQueue_fifo_2_empty),
    .almost_empty (readData_readDataQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_2_almostFull),
    .full         (_readData_readDataQueue_fifo_2_full),
    .error        (_readData_readDataQueue_fifo_2_error),
    .data_out     (_readData_readDataQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_3_enq_ready & readData_readDataQueue_3_enq_valid & ~(_readData_readDataQueue_fifo_3_empty & readData_readDataQueue_3_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_3_deq_ready & ~_readData_readDataQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_3_enq_bits),
    .empty        (_readData_readDataQueue_fifo_3_empty),
    .almost_empty (readData_readDataQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_3_almostFull),
    .full         (_readData_readDataQueue_fifo_3_full),
    .error        (_readData_readDataQueue_fifo_3_error),
    .data_out     (_readData_readDataQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_4_enq_ready & readData_readDataQueue_4_enq_valid & ~(_readData_readDataQueue_fifo_4_empty & readData_readDataQueue_4_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_4_deq_ready & ~_readData_readDataQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_4_enq_bits),
    .empty        (_readData_readDataQueue_fifo_4_empty),
    .almost_empty (readData_readDataQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_4_almostFull),
    .full         (_readData_readDataQueue_fifo_4_full),
    .error        (_readData_readDataQueue_fifo_4_error),
    .data_out     (_readData_readDataQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_5_enq_ready & readData_readDataQueue_5_enq_valid & ~(_readData_readDataQueue_fifo_5_empty & readData_readDataQueue_5_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_5_deq_ready & ~_readData_readDataQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_5_enq_bits),
    .empty        (_readData_readDataQueue_fifo_5_empty),
    .almost_empty (readData_readDataQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_5_almostFull),
    .full         (_readData_readDataQueue_fifo_5_full),
    .error        (_readData_readDataQueue_fifo_5_error),
    .data_out     (_readData_readDataQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_6_enq_ready & readData_readDataQueue_6_enq_valid & ~(_readData_readDataQueue_fifo_6_empty & readData_readDataQueue_6_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_6_deq_ready & ~_readData_readDataQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_6_enq_bits),
    .empty        (_readData_readDataQueue_fifo_6_empty),
    .almost_empty (readData_readDataQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_6_almostFull),
    .full         (_readData_readDataQueue_fifo_6_full),
    .error        (_readData_readDataQueue_fifo_6_error),
    .data_out     (_readData_readDataQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_7_enq_ready & readData_readDataQueue_7_enq_valid & ~(_readData_readDataQueue_fifo_7_empty & readData_readDataQueue_7_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_7_deq_ready & ~_readData_readDataQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_7_enq_bits),
    .empty        (_readData_readDataQueue_fifo_7_empty),
    .almost_empty (readData_readDataQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_7_almostFull),
    .full         (_readData_readDataQueue_fifo_7_full),
    .error        (_readData_readDataQueue_fifo_7_error),
    .data_out     (_readData_readDataQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_8_enq_ready & readData_readDataQueue_8_enq_valid & ~(_readData_readDataQueue_fifo_8_empty & readData_readDataQueue_8_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_8_deq_ready & ~_readData_readDataQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_8_enq_bits),
    .empty        (_readData_readDataQueue_fifo_8_empty),
    .almost_empty (readData_readDataQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_8_almostFull),
    .full         (_readData_readDataQueue_fifo_8_full),
    .error        (_readData_readDataQueue_fifo_8_error),
    .data_out     (_readData_readDataQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_9_enq_ready & readData_readDataQueue_9_enq_valid & ~(_readData_readDataQueue_fifo_9_empty & readData_readDataQueue_9_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_9_deq_ready & ~_readData_readDataQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_9_enq_bits),
    .empty        (_readData_readDataQueue_fifo_9_empty),
    .almost_empty (readData_readDataQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_9_almostFull),
    .full         (_readData_readDataQueue_fifo_9_full),
    .error        (_readData_readDataQueue_fifo_9_error),
    .data_out     (_readData_readDataQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_10_enq_ready & readData_readDataQueue_10_enq_valid & ~(_readData_readDataQueue_fifo_10_empty & readData_readDataQueue_10_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_10_deq_ready & ~_readData_readDataQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_10_enq_bits),
    .empty        (_readData_readDataQueue_fifo_10_empty),
    .almost_empty (readData_readDataQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_10_almostFull),
    .full         (_readData_readDataQueue_fifo_10_full),
    .error        (_readData_readDataQueue_fifo_10_error),
    .data_out     (_readData_readDataQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_11_enq_ready & readData_readDataQueue_11_enq_valid & ~(_readData_readDataQueue_fifo_11_empty & readData_readDataQueue_11_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_11_deq_ready & ~_readData_readDataQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_11_enq_bits),
    .empty        (_readData_readDataQueue_fifo_11_empty),
    .almost_empty (readData_readDataQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_11_almostFull),
    .full         (_readData_readDataQueue_fifo_11_full),
    .error        (_readData_readDataQueue_fifo_11_error),
    .data_out     (_readData_readDataQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_12_enq_ready & readData_readDataQueue_12_enq_valid & ~(_readData_readDataQueue_fifo_12_empty & readData_readDataQueue_12_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_12_deq_ready & ~_readData_readDataQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_12_enq_bits),
    .empty        (_readData_readDataQueue_fifo_12_empty),
    .almost_empty (readData_readDataQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_12_almostFull),
    .full         (_readData_readDataQueue_fifo_12_full),
    .error        (_readData_readDataQueue_fifo_12_error),
    .data_out     (_readData_readDataQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_13_enq_ready & readData_readDataQueue_13_enq_valid & ~(_readData_readDataQueue_fifo_13_empty & readData_readDataQueue_13_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_13_deq_ready & ~_readData_readDataQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_13_enq_bits),
    .empty        (_readData_readDataQueue_fifo_13_empty),
    .almost_empty (readData_readDataQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_13_almostFull),
    .full         (_readData_readDataQueue_fifo_13_full),
    .error        (_readData_readDataQueue_fifo_13_error),
    .data_out     (_readData_readDataQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_14_enq_ready & readData_readDataQueue_14_enq_valid & ~(_readData_readDataQueue_fifo_14_empty & readData_readDataQueue_14_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_14_deq_ready & ~_readData_readDataQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_14_enq_bits),
    .empty        (_readData_readDataQueue_fifo_14_empty),
    .almost_empty (readData_readDataQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_14_almostFull),
    .full         (_readData_readDataQueue_fifo_14_full),
    .error        (_readData_readDataQueue_fifo_14_error),
    .data_out     (_readData_readDataQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_15_enq_ready & readData_readDataQueue_15_enq_valid & ~(_readData_readDataQueue_fifo_15_empty & readData_readDataQueue_15_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_15_deq_ready & ~_readData_readDataQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_15_enq_bits),
    .empty        (_readData_readDataQueue_fifo_15_empty),
    .almost_empty (readData_readDataQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_15_almostFull),
    .full         (_readData_readDataQueue_fifo_15_full),
    .error        (_readData_readDataQueue_fifo_15_error),
    .data_out     (_readData_readDataQueue_fifo_15_data_out)
  );
  MaskCompress compressUnit (
    .clock                  (clock),
    .reset                  (reset),
    .in_valid               (viotaCounterAdd),
    .in_bits_maskType       (instReg_maskType),
    .in_bits_eew            (instReg_sew),
    .in_bits_uop            (instReg_decodeResult_topUop[2:0]),
    .in_bits_readFromScalar (instReg_readFromScala),
    .in_bits_source1        (source1Select),
    .in_bits_mask           (executeElementMask[31:0]),
    .in_bits_source2        (source2),
    .in_bits_pipeData       (source1),
    .in_bits_groupCounter   (requestCounter),
    .in_bits_ffoInput       ({view__in_bits_ffoInput_hi, view__in_bits_ffoInput_lo}),
    .in_bits_validInput     ({view__in_bits_validInput_hi, view__in_bits_validInput_lo}),
    .in_bits_lastCompress   (lastGroup),
    .out_data               (compressUnitResultQueue_enq_bits_data),
    .out_mask               (compressUnitResultQueue_enq_bits_mask),
    .out_groupCounter       (compressUnitResultQueue_enq_bits_groupCounter),
    .out_ffoOutput          (compressUnitResultQueue_enq_bits_ffoOutput),
    .out_compressValid      (_compressUnit_out_compressValid),
    .newInstruction         (instReq_valid),
    .ffoInstruction         (&(instReq_bits_decodeResult_topUop[2:1])),
    .writeData              (_compressUnit_writeData),
    .stageValid             (_compressUnit_stageValid)
  );
  MaskReduce reduceUnit (
    .clock                 (clock),
    .reset                 (reset),
    .in_ready              (_reduceUnit_in_ready),
    .in_valid              (reduceUnit_in_valid),
    .in_bits_maskType      (instReg_maskType),
    .in_bits_eew           (instReg_sew),
    .in_bits_uop           (instReg_decodeResult_topUop[2:0]),
    .in_bits_readVS1       (readVS1Reg_data),
    .in_bits_source2       (source2),
    .in_bits_sourceValid   ({view__in_bits_sourceValid_hi, view__in_bits_sourceValid_lo}),
    .in_bits_lastGroup     (lastGroup),
    .in_bits_vxrm          (instReg_vxrm),
    .in_bits_aluUop        (instReg_decodeResult_uop),
    .in_bits_sign          (~instReg_decodeResult_unsigned1),
    .in_bits_fpSourceValid ({view__in_bits_fpSourceValid_hi, view__in_bits_fpSourceValid_lo}),
    .out_valid             (_reduceUnit_out_valid),
    .out_bits_data         (_reduceUnit_out_bits_data),
    .out_bits_mask         (_reduceUnit_out_bits_mask),
    .firstGroup            (~readVS1Reg_sendToExecution & _view__firstGroup_T_1),
    .newInstruction        (instReq_valid),
    .validInst             (|instReg_vl),
    .pop                   (instReg_decodeResult_popCount)
  );
  MaskExtend extendUnit (
    .in_eew          (instReg_sew),
    .in_uop          (instReg_decodeResult_topUop[2:0]),
    .in_source2      (source2),
    .in_groupCounter (extendGroupCount[4:0]),
    .out             (_extendUnit_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_0_enq_ready & writeQueue_0_enq_valid)),
    .pop_req_n    (~(writeQueue_0_deq_ready & ~_writeQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn),
    .empty        (_writeQueue_fifo_empty),
    .almost_empty (writeQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_0_almostFull),
    .full         (_writeQueue_fifo_full),
    .error        (_writeQueue_fifo_error),
    .data_out     (_writeQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_1_enq_ready & writeQueue_1_enq_valid)),
    .pop_req_n    (~(writeQueue_1_deq_ready & ~_writeQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_1),
    .empty        (_writeQueue_fifo_1_empty),
    .almost_empty (writeQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_1_almostFull),
    .full         (_writeQueue_fifo_1_full),
    .error        (_writeQueue_fifo_1_error),
    .data_out     (_writeQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_2_enq_ready & writeQueue_2_enq_valid)),
    .pop_req_n    (~(writeQueue_2_deq_ready & ~_writeQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_2),
    .empty        (_writeQueue_fifo_2_empty),
    .almost_empty (writeQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_2_almostFull),
    .full         (_writeQueue_fifo_2_full),
    .error        (_writeQueue_fifo_2_error),
    .data_out     (_writeQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_3_enq_ready & writeQueue_3_enq_valid)),
    .pop_req_n    (~(writeQueue_3_deq_ready & ~_writeQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_3),
    .empty        (_writeQueue_fifo_3_empty),
    .almost_empty (writeQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_3_almostFull),
    .full         (_writeQueue_fifo_3_full),
    .error        (_writeQueue_fifo_3_error),
    .data_out     (_writeQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_4_enq_ready & writeQueue_4_enq_valid)),
    .pop_req_n    (~(writeQueue_4_deq_ready & ~_writeQueue_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_4),
    .empty        (_writeQueue_fifo_4_empty),
    .almost_empty (writeQueue_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_4_almostFull),
    .full         (_writeQueue_fifo_4_full),
    .error        (_writeQueue_fifo_4_error),
    .data_out     (_writeQueue_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_5_enq_ready & writeQueue_5_enq_valid)),
    .pop_req_n    (~(writeQueue_5_deq_ready & ~_writeQueue_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_5),
    .empty        (_writeQueue_fifo_5_empty),
    .almost_empty (writeQueue_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_5_almostFull),
    .full         (_writeQueue_fifo_5_full),
    .error        (_writeQueue_fifo_5_error),
    .data_out     (_writeQueue_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_6_enq_ready & writeQueue_6_enq_valid)),
    .pop_req_n    (~(writeQueue_6_deq_ready & ~_writeQueue_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_6),
    .empty        (_writeQueue_fifo_6_empty),
    .almost_empty (writeQueue_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_6_almostFull),
    .full         (_writeQueue_fifo_6_full),
    .error        (_writeQueue_fifo_6_error),
    .data_out     (_writeQueue_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_7_enq_ready & writeQueue_7_enq_valid)),
    .pop_req_n    (~(writeQueue_7_deq_ready & ~_writeQueue_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_7),
    .empty        (_writeQueue_fifo_7_empty),
    .almost_empty (writeQueue_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_7_almostFull),
    .full         (_writeQueue_fifo_7_full),
    .error        (_writeQueue_fifo_7_error),
    .data_out     (_writeQueue_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_8_enq_ready & writeQueue_8_enq_valid)),
    .pop_req_n    (~(writeQueue_8_deq_ready & ~_writeQueue_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_8),
    .empty        (_writeQueue_fifo_8_empty),
    .almost_empty (writeQueue_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_8_almostFull),
    .full         (_writeQueue_fifo_8_full),
    .error        (_writeQueue_fifo_8_error),
    .data_out     (_writeQueue_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_9_enq_ready & writeQueue_9_enq_valid)),
    .pop_req_n    (~(writeQueue_9_deq_ready & ~_writeQueue_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_9),
    .empty        (_writeQueue_fifo_9_empty),
    .almost_empty (writeQueue_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_9_almostFull),
    .full         (_writeQueue_fifo_9_full),
    .error        (_writeQueue_fifo_9_error),
    .data_out     (_writeQueue_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_10_enq_ready & writeQueue_10_enq_valid)),
    .pop_req_n    (~(writeQueue_10_deq_ready & ~_writeQueue_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_10),
    .empty        (_writeQueue_fifo_10_empty),
    .almost_empty (writeQueue_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_10_almostFull),
    .full         (_writeQueue_fifo_10_full),
    .error        (_writeQueue_fifo_10_error),
    .data_out     (_writeQueue_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_11_enq_ready & writeQueue_11_enq_valid)),
    .pop_req_n    (~(writeQueue_11_deq_ready & ~_writeQueue_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_11),
    .empty        (_writeQueue_fifo_11_empty),
    .almost_empty (writeQueue_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_11_almostFull),
    .full         (_writeQueue_fifo_11_full),
    .error        (_writeQueue_fifo_11_error),
    .data_out     (_writeQueue_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_12_enq_ready & writeQueue_12_enq_valid)),
    .pop_req_n    (~(writeQueue_12_deq_ready & ~_writeQueue_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_12),
    .empty        (_writeQueue_fifo_12_empty),
    .almost_empty (writeQueue_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_12_almostFull),
    .full         (_writeQueue_fifo_12_full),
    .error        (_writeQueue_fifo_12_error),
    .data_out     (_writeQueue_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_13_enq_ready & writeQueue_13_enq_valid)),
    .pop_req_n    (~(writeQueue_13_deq_ready & ~_writeQueue_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_13),
    .empty        (_writeQueue_fifo_13_empty),
    .almost_empty (writeQueue_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_13_almostFull),
    .full         (_writeQueue_fifo_13_full),
    .error        (_writeQueue_fifo_13_error),
    .data_out     (_writeQueue_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_14_enq_ready & writeQueue_14_enq_valid)),
    .pop_req_n    (~(writeQueue_14_deq_ready & ~_writeQueue_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_14),
    .empty        (_writeQueue_fifo_14_empty),
    .almost_empty (writeQueue_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_14_almostFull),
    .full         (_writeQueue_fifo_14_full),
    .error        (_writeQueue_fifo_14_error),
    .data_out     (_writeQueue_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(50)
  ) writeQueue_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_15_enq_ready & writeQueue_15_enq_valid)),
    .pop_req_n    (~(writeQueue_15_deq_ready & ~_writeQueue_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_15),
    .empty        (_writeQueue_fifo_15_empty),
    .almost_empty (writeQueue_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_15_almostFull),
    .full         (_writeQueue_fifo_15_full),
    .error        (_writeQueue_fifo_15_error),
    .data_out     (_writeQueue_fifo_15_data_out)
  );
  assign exeResp_0_valid = exeResp_0_valid_0;
  assign exeResp_0_bits_vd = exeResp_0_bits_vd_0;
  assign exeResp_0_bits_offset = exeResp_0_bits_offset_0;
  assign exeResp_0_bits_mask = exeResp_0_bits_mask_0;
  assign exeResp_0_bits_data = exeResp_0_bits_data_0;
  assign exeResp_0_bits_instructionIndex = exeResp_0_bits_instructionIndex_0;
  assign exeResp_1_valid = exeResp_1_valid_0;
  assign exeResp_1_bits_vd = exeResp_1_bits_vd_0;
  assign exeResp_1_bits_offset = exeResp_1_bits_offset_0;
  assign exeResp_1_bits_mask = exeResp_1_bits_mask_0;
  assign exeResp_1_bits_data = exeResp_1_bits_data_0;
  assign exeResp_1_bits_instructionIndex = exeResp_1_bits_instructionIndex_0;
  assign exeResp_2_valid = exeResp_2_valid_0;
  assign exeResp_2_bits_vd = exeResp_2_bits_vd_0;
  assign exeResp_2_bits_offset = exeResp_2_bits_offset_0;
  assign exeResp_2_bits_mask = exeResp_2_bits_mask_0;
  assign exeResp_2_bits_data = exeResp_2_bits_data_0;
  assign exeResp_2_bits_instructionIndex = exeResp_2_bits_instructionIndex_0;
  assign exeResp_3_valid = exeResp_3_valid_0;
  assign exeResp_3_bits_vd = exeResp_3_bits_vd_0;
  assign exeResp_3_bits_offset = exeResp_3_bits_offset_0;
  assign exeResp_3_bits_mask = exeResp_3_bits_mask_0;
  assign exeResp_3_bits_data = exeResp_3_bits_data_0;
  assign exeResp_3_bits_instructionIndex = exeResp_3_bits_instructionIndex_0;
  assign exeResp_4_valid = exeResp_4_valid_0;
  assign exeResp_4_bits_vd = exeResp_4_bits_vd_0;
  assign exeResp_4_bits_offset = exeResp_4_bits_offset_0;
  assign exeResp_4_bits_mask = exeResp_4_bits_mask_0;
  assign exeResp_4_bits_data = exeResp_4_bits_data_0;
  assign exeResp_4_bits_instructionIndex = exeResp_4_bits_instructionIndex_0;
  assign exeResp_5_valid = exeResp_5_valid_0;
  assign exeResp_5_bits_vd = exeResp_5_bits_vd_0;
  assign exeResp_5_bits_offset = exeResp_5_bits_offset_0;
  assign exeResp_5_bits_mask = exeResp_5_bits_mask_0;
  assign exeResp_5_bits_data = exeResp_5_bits_data_0;
  assign exeResp_5_bits_instructionIndex = exeResp_5_bits_instructionIndex_0;
  assign exeResp_6_valid = exeResp_6_valid_0;
  assign exeResp_6_bits_vd = exeResp_6_bits_vd_0;
  assign exeResp_6_bits_offset = exeResp_6_bits_offset_0;
  assign exeResp_6_bits_mask = exeResp_6_bits_mask_0;
  assign exeResp_6_bits_data = exeResp_6_bits_data_0;
  assign exeResp_6_bits_instructionIndex = exeResp_6_bits_instructionIndex_0;
  assign exeResp_7_valid = exeResp_7_valid_0;
  assign exeResp_7_bits_vd = exeResp_7_bits_vd_0;
  assign exeResp_7_bits_offset = exeResp_7_bits_offset_0;
  assign exeResp_7_bits_mask = exeResp_7_bits_mask_0;
  assign exeResp_7_bits_data = exeResp_7_bits_data_0;
  assign exeResp_7_bits_instructionIndex = exeResp_7_bits_instructionIndex_0;
  assign exeResp_8_valid = exeResp_8_valid_0;
  assign exeResp_8_bits_vd = exeResp_8_bits_vd_0;
  assign exeResp_8_bits_offset = exeResp_8_bits_offset_0;
  assign exeResp_8_bits_mask = exeResp_8_bits_mask_0;
  assign exeResp_8_bits_data = exeResp_8_bits_data_0;
  assign exeResp_8_bits_instructionIndex = exeResp_8_bits_instructionIndex_0;
  assign exeResp_9_valid = exeResp_9_valid_0;
  assign exeResp_9_bits_vd = exeResp_9_bits_vd_0;
  assign exeResp_9_bits_offset = exeResp_9_bits_offset_0;
  assign exeResp_9_bits_mask = exeResp_9_bits_mask_0;
  assign exeResp_9_bits_data = exeResp_9_bits_data_0;
  assign exeResp_9_bits_instructionIndex = exeResp_9_bits_instructionIndex_0;
  assign exeResp_10_valid = exeResp_10_valid_0;
  assign exeResp_10_bits_vd = exeResp_10_bits_vd_0;
  assign exeResp_10_bits_offset = exeResp_10_bits_offset_0;
  assign exeResp_10_bits_mask = exeResp_10_bits_mask_0;
  assign exeResp_10_bits_data = exeResp_10_bits_data_0;
  assign exeResp_10_bits_instructionIndex = exeResp_10_bits_instructionIndex_0;
  assign exeResp_11_valid = exeResp_11_valid_0;
  assign exeResp_11_bits_vd = exeResp_11_bits_vd_0;
  assign exeResp_11_bits_offset = exeResp_11_bits_offset_0;
  assign exeResp_11_bits_mask = exeResp_11_bits_mask_0;
  assign exeResp_11_bits_data = exeResp_11_bits_data_0;
  assign exeResp_11_bits_instructionIndex = exeResp_11_bits_instructionIndex_0;
  assign exeResp_12_valid = exeResp_12_valid_0;
  assign exeResp_12_bits_vd = exeResp_12_bits_vd_0;
  assign exeResp_12_bits_offset = exeResp_12_bits_offset_0;
  assign exeResp_12_bits_mask = exeResp_12_bits_mask_0;
  assign exeResp_12_bits_data = exeResp_12_bits_data_0;
  assign exeResp_12_bits_instructionIndex = exeResp_12_bits_instructionIndex_0;
  assign exeResp_13_valid = exeResp_13_valid_0;
  assign exeResp_13_bits_vd = exeResp_13_bits_vd_0;
  assign exeResp_13_bits_offset = exeResp_13_bits_offset_0;
  assign exeResp_13_bits_mask = exeResp_13_bits_mask_0;
  assign exeResp_13_bits_data = exeResp_13_bits_data_0;
  assign exeResp_13_bits_instructionIndex = exeResp_13_bits_instructionIndex_0;
  assign exeResp_14_valid = exeResp_14_valid_0;
  assign exeResp_14_bits_vd = exeResp_14_bits_vd_0;
  assign exeResp_14_bits_offset = exeResp_14_bits_offset_0;
  assign exeResp_14_bits_mask = exeResp_14_bits_mask_0;
  assign exeResp_14_bits_data = exeResp_14_bits_data_0;
  assign exeResp_14_bits_instructionIndex = exeResp_14_bits_instructionIndex_0;
  assign exeResp_15_valid = exeResp_15_valid_0;
  assign exeResp_15_bits_vd = exeResp_15_bits_vd_0;
  assign exeResp_15_bits_offset = exeResp_15_bits_offset_0;
  assign exeResp_15_bits_mask = exeResp_15_bits_mask_0;
  assign exeResp_15_bits_data = exeResp_15_bits_data_0;
  assign exeResp_15_bits_instructionIndex = exeResp_15_bits_instructionIndex_0;
  assign tokenIO_0_maskRequestRelease = tokenIO_0_maskRequestRelease_0;
  assign tokenIO_1_maskRequestRelease = tokenIO_1_maskRequestRelease_0;
  assign tokenIO_2_maskRequestRelease = tokenIO_2_maskRequestRelease_0;
  assign tokenIO_3_maskRequestRelease = tokenIO_3_maskRequestRelease_0;
  assign tokenIO_4_maskRequestRelease = tokenIO_4_maskRequestRelease_0;
  assign tokenIO_5_maskRequestRelease = tokenIO_5_maskRequestRelease_0;
  assign tokenIO_6_maskRequestRelease = tokenIO_6_maskRequestRelease_0;
  assign tokenIO_7_maskRequestRelease = tokenIO_7_maskRequestRelease_0;
  assign tokenIO_8_maskRequestRelease = tokenIO_8_maskRequestRelease_0;
  assign tokenIO_9_maskRequestRelease = tokenIO_9_maskRequestRelease_0;
  assign tokenIO_10_maskRequestRelease = tokenIO_10_maskRequestRelease_0;
  assign tokenIO_11_maskRequestRelease = tokenIO_11_maskRequestRelease_0;
  assign tokenIO_12_maskRequestRelease = tokenIO_12_maskRequestRelease_0;
  assign tokenIO_13_maskRequestRelease = tokenIO_13_maskRequestRelease_0;
  assign tokenIO_14_maskRequestRelease = tokenIO_14_maskRequestRelease_0;
  assign tokenIO_15_maskRequestRelease = tokenIO_15_maskRequestRelease_0;
  assign readChannel_0_valid = readChannel_0_valid_0;
  assign readChannel_0_bits_vs = readChannel_0_bits_vs_0;
  assign readChannel_0_bits_offset = readChannel_0_bits_offset_0;
  assign readChannel_0_bits_instructionIndex = readChannel_0_bits_instructionIndex_0;
  assign readChannel_1_valid = readChannel_1_valid_0;
  assign readChannel_1_bits_vs = readChannel_1_bits_vs_0;
  assign readChannel_1_bits_offset = readChannel_1_bits_offset_0;
  assign readChannel_1_bits_instructionIndex = readChannel_1_bits_instructionIndex_0;
  assign readChannel_2_valid = readChannel_2_valid_0;
  assign readChannel_2_bits_vs = readChannel_2_bits_vs_0;
  assign readChannel_2_bits_offset = readChannel_2_bits_offset_0;
  assign readChannel_2_bits_instructionIndex = readChannel_2_bits_instructionIndex_0;
  assign readChannel_3_valid = readChannel_3_valid_0;
  assign readChannel_3_bits_vs = readChannel_3_bits_vs_0;
  assign readChannel_3_bits_offset = readChannel_3_bits_offset_0;
  assign readChannel_3_bits_instructionIndex = readChannel_3_bits_instructionIndex_0;
  assign readChannel_4_valid = readChannel_4_valid_0;
  assign readChannel_4_bits_vs = readChannel_4_bits_vs_0;
  assign readChannel_4_bits_offset = readChannel_4_bits_offset_0;
  assign readChannel_4_bits_instructionIndex = readChannel_4_bits_instructionIndex_0;
  assign readChannel_5_valid = readChannel_5_valid_0;
  assign readChannel_5_bits_vs = readChannel_5_bits_vs_0;
  assign readChannel_5_bits_offset = readChannel_5_bits_offset_0;
  assign readChannel_5_bits_instructionIndex = readChannel_5_bits_instructionIndex_0;
  assign readChannel_6_valid = readChannel_6_valid_0;
  assign readChannel_6_bits_vs = readChannel_6_bits_vs_0;
  assign readChannel_6_bits_offset = readChannel_6_bits_offset_0;
  assign readChannel_6_bits_instructionIndex = readChannel_6_bits_instructionIndex_0;
  assign readChannel_7_valid = readChannel_7_valid_0;
  assign readChannel_7_bits_vs = readChannel_7_bits_vs_0;
  assign readChannel_7_bits_offset = readChannel_7_bits_offset_0;
  assign readChannel_7_bits_instructionIndex = readChannel_7_bits_instructionIndex_0;
  assign readChannel_8_valid = readChannel_8_valid_0;
  assign readChannel_8_bits_vs = readChannel_8_bits_vs_0;
  assign readChannel_8_bits_offset = readChannel_8_bits_offset_0;
  assign readChannel_8_bits_instructionIndex = readChannel_8_bits_instructionIndex_0;
  assign readChannel_9_valid = readChannel_9_valid_0;
  assign readChannel_9_bits_vs = readChannel_9_bits_vs_0;
  assign readChannel_9_bits_offset = readChannel_9_bits_offset_0;
  assign readChannel_9_bits_instructionIndex = readChannel_9_bits_instructionIndex_0;
  assign readChannel_10_valid = readChannel_10_valid_0;
  assign readChannel_10_bits_vs = readChannel_10_bits_vs_0;
  assign readChannel_10_bits_offset = readChannel_10_bits_offset_0;
  assign readChannel_10_bits_instructionIndex = readChannel_10_bits_instructionIndex_0;
  assign readChannel_11_valid = readChannel_11_valid_0;
  assign readChannel_11_bits_vs = readChannel_11_bits_vs_0;
  assign readChannel_11_bits_offset = readChannel_11_bits_offset_0;
  assign readChannel_11_bits_instructionIndex = readChannel_11_bits_instructionIndex_0;
  assign readChannel_12_valid = readChannel_12_valid_0;
  assign readChannel_12_bits_vs = readChannel_12_bits_vs_0;
  assign readChannel_12_bits_offset = readChannel_12_bits_offset_0;
  assign readChannel_12_bits_instructionIndex = readChannel_12_bits_instructionIndex_0;
  assign readChannel_13_valid = readChannel_13_valid_0;
  assign readChannel_13_bits_vs = readChannel_13_bits_vs_0;
  assign readChannel_13_bits_offset = readChannel_13_bits_offset_0;
  assign readChannel_13_bits_instructionIndex = readChannel_13_bits_instructionIndex_0;
  assign readChannel_14_valid = readChannel_14_valid_0;
  assign readChannel_14_bits_vs = readChannel_14_bits_vs_0;
  assign readChannel_14_bits_offset = readChannel_14_bits_offset_0;
  assign readChannel_14_bits_instructionIndex = readChannel_14_bits_instructionIndex_0;
  assign readChannel_15_valid = readChannel_15_valid_0;
  assign readChannel_15_bits_vs = readChannel_15_bits_vs_0;
  assign readChannel_15_bits_offset = readChannel_15_bits_offset_0;
  assign readChannel_15_bits_instructionIndex = readChannel_15_bits_instructionIndex_0;
  assign lastReport = _lastReport_output;
  assign laneMaskInput_0 = laneMaskSelect_0[0] ? v0SelectBySew[63:32] : v0SelectBySew[31:0];
  assign laneMaskInput_1 = laneMaskSelect_1[0] ? v0SelectBySew_1[63:32] : v0SelectBySew_1[31:0];
  assign laneMaskInput_2 = laneMaskSelect_2[0] ? v0SelectBySew_2[63:32] : v0SelectBySew_2[31:0];
  assign laneMaskInput_3 = laneMaskSelect_3[0] ? v0SelectBySew_3[63:32] : v0SelectBySew_3[31:0];
  assign laneMaskInput_4 = laneMaskSelect_4[0] ? v0SelectBySew_4[63:32] : v0SelectBySew_4[31:0];
  assign laneMaskInput_5 = laneMaskSelect_5[0] ? v0SelectBySew_5[63:32] : v0SelectBySew_5[31:0];
  assign laneMaskInput_6 = laneMaskSelect_6[0] ? v0SelectBySew_6[63:32] : v0SelectBySew_6[31:0];
  assign laneMaskInput_7 = laneMaskSelect_7[0] ? v0SelectBySew_7[63:32] : v0SelectBySew_7[31:0];
  assign laneMaskInput_8 = laneMaskSelect_8[0] ? v0SelectBySew_8[63:32] : v0SelectBySew_8[31:0];
  assign laneMaskInput_9 = laneMaskSelect_9[0] ? v0SelectBySew_9[63:32] : v0SelectBySew_9[31:0];
  assign laneMaskInput_10 = laneMaskSelect_10[0] ? v0SelectBySew_10[63:32] : v0SelectBySew_10[31:0];
  assign laneMaskInput_11 = laneMaskSelect_11[0] ? v0SelectBySew_11[63:32] : v0SelectBySew_11[31:0];
  assign laneMaskInput_12 = laneMaskSelect_12[0] ? v0SelectBySew_12[63:32] : v0SelectBySew_12[31:0];
  assign laneMaskInput_13 = laneMaskSelect_13[0] ? v0SelectBySew_13[63:32] : v0SelectBySew_13[31:0];
  assign laneMaskInput_14 = laneMaskSelect_14[0] ? v0SelectBySew_14[63:32] : v0SelectBySew_14[31:0];
  assign laneMaskInput_15 = laneMaskSelect_15[0] ? v0SelectBySew_15[63:32] : v0SelectBySew_15[31:0];
  assign writeRDData = instReg_decodeResult_popCount ? _reduceUnit_out_bits_data : _compressUnit_writeData;
  assign gatherData_valid = gatherData_valid_0;
  assign gatherData_bits = gatherData_bits_0;
endmodule

