
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LoadUnit(
  input          clock,
                 reset,
                 lsuRequest_valid,
  input  [2:0]   lsuRequest_bits_instructionInformation_nf,
  input          lsuRequest_bits_instructionInformation_mew,
  input  [1:0]   lsuRequest_bits_instructionInformation_mop,
  input  [4:0]   lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]   lsuRequest_bits_instructionInformation_eew,
  input  [4:0]   lsuRequest_bits_instructionInformation_vs3,
  input          lsuRequest_bits_instructionInformation_isStore,
                 lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  lsuRequest_bits_rs1Data,
                 lsuRequest_bits_rs2Data,
  input  [2:0]   lsuRequest_bits_instructionIndex,
  input  [11:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
  input  [15:0]  maskInput,
  output         maskSelect_valid,
  output [6:0]   maskSelect_bits,
  input          addressConflict,
                 memRequest_ready,
  output         memRequest_valid,
  output [7:0]   memRequest_bits_src,
  output [31:0]  memRequest_bits_address,
  output         memResponse_ready,
  input          memResponse_valid,
  input  [127:0] memResponse_bits_data,
  input  [7:0]   memResponse_bits_index,
  output         status_idle,
                 status_last,
  output [2:0]   status_instructionIndex,
  output         status_changeMaskGroup,
  output [31:0]  status_startAddress,
                 status_endAddress,
  input          vrfWritePort_0_ready,
  output         vrfWritePort_0_valid,
  output [4:0]   vrfWritePort_0_bits_vd,
  output [3:0]   vrfWritePort_0_bits_offset,
                 vrfWritePort_0_bits_mask,
  output [31:0]  vrfWritePort_0_bits_data,
  output [2:0]   vrfWritePort_0_bits_instructionIndex,
  input          vrfWritePort_1_ready,
  output         vrfWritePort_1_valid,
  output [4:0]   vrfWritePort_1_bits_vd,
  output [3:0]   vrfWritePort_1_bits_offset,
                 vrfWritePort_1_bits_mask,
  output [31:0]  vrfWritePort_1_bits_data,
  output [2:0]   vrfWritePort_1_bits_instructionIndex,
  input          vrfWritePort_2_ready,
  output         vrfWritePort_2_valid,
  output [4:0]   vrfWritePort_2_bits_vd,
  output [3:0]   vrfWritePort_2_bits_offset,
                 vrfWritePort_2_bits_mask,
  output [31:0]  vrfWritePort_2_bits_data,
  output [2:0]   vrfWritePort_2_bits_instructionIndex,
  input          vrfWritePort_3_ready,
  output         vrfWritePort_3_valid,
  output [4:0]   vrfWritePort_3_bits_vd,
  output [3:0]   vrfWritePort_3_bits_offset,
                 vrfWritePort_3_bits_mask,
  output [31:0]  vrfWritePort_3_bits_data,
  output [2:0]   vrfWritePort_3_bits_instructionIndex
);

  wire          memRequest_ready_0 = memRequest_ready;
  wire          memResponse_valid_0 = memResponse_valid;
  wire [127:0]  memResponse_bits_data_0 = memResponse_bits_data;
  wire [7:0]    memResponse_bits_index_0 = memResponse_bits_index;
  wire          vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire          vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire          vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire          vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire [511:0]  hi = 512'h0;
  wire [511:0]  hi_1 = 512'h0;
  wire [511:0]  hi_2 = 512'h0;
  wire [511:0]  hi_3 = 512'h0;
  wire [511:0]  hi_8 = 512'h0;
  wire [511:0]  hi_9 = 512'h0;
  wire [511:0]  hi_10 = 512'h0;
  wire [511:0]  hi_11 = 512'h0;
  wire [511:0]  hi_16 = 512'h0;
  wire [511:0]  hi_17 = 512'h0;
  wire [511:0]  hi_18 = 512'h0;
  wire [511:0]  hi_19 = 512'h0;
  wire [255:0]  lo_hi = 256'h0;
  wire [255:0]  hi_lo = 256'h0;
  wire [255:0]  hi_hi = 256'h0;
  wire [255:0]  lo_hi_1 = 256'h0;
  wire [255:0]  hi_lo_1 = 256'h0;
  wire [255:0]  hi_hi_1 = 256'h0;
  wire [255:0]  hi_lo_2 = 256'h0;
  wire [255:0]  hi_hi_2 = 256'h0;
  wire [255:0]  hi_lo_3 = 256'h0;
  wire [255:0]  hi_hi_3 = 256'h0;
  wire [255:0]  hi_hi_4 = 256'h0;
  wire [255:0]  hi_hi_5 = 256'h0;
  wire [255:0]  lo_hi_8 = 256'h0;
  wire [255:0]  hi_lo_8 = 256'h0;
  wire [255:0]  hi_hi_8 = 256'h0;
  wire [255:0]  lo_hi_9 = 256'h0;
  wire [255:0]  hi_lo_9 = 256'h0;
  wire [255:0]  hi_hi_9 = 256'h0;
  wire [255:0]  hi_lo_10 = 256'h0;
  wire [255:0]  hi_hi_10 = 256'h0;
  wire [255:0]  hi_lo_11 = 256'h0;
  wire [255:0]  hi_hi_11 = 256'h0;
  wire [255:0]  hi_hi_12 = 256'h0;
  wire [255:0]  hi_hi_13 = 256'h0;
  wire [255:0]  lo_hi_16 = 256'h0;
  wire [255:0]  hi_lo_16 = 256'h0;
  wire [255:0]  hi_hi_16 = 256'h0;
  wire [255:0]  lo_hi_17 = 256'h0;
  wire [255:0]  hi_lo_17 = 256'h0;
  wire [255:0]  hi_hi_17 = 256'h0;
  wire [255:0]  hi_lo_18 = 256'h0;
  wire [255:0]  hi_hi_18 = 256'h0;
  wire [255:0]  hi_lo_19 = 256'h0;
  wire [255:0]  hi_hi_19 = 256'h0;
  wire [255:0]  hi_hi_20 = 256'h0;
  wire [255:0]  hi_hi_21 = 256'h0;
  wire [127:0]  res_1 = 128'h0;
  wire [127:0]  res_2 = 128'h0;
  wire [127:0]  res_3 = 128'h0;
  wire [127:0]  res_4 = 128'h0;
  wire [127:0]  res_5 = 128'h0;
  wire [127:0]  res_6 = 128'h0;
  wire [127:0]  res_7 = 128'h0;
  wire [127:0]  res_10 = 128'h0;
  wire [127:0]  res_11 = 128'h0;
  wire [127:0]  res_12 = 128'h0;
  wire [127:0]  res_13 = 128'h0;
  wire [127:0]  res_14 = 128'h0;
  wire [127:0]  res_15 = 128'h0;
  wire [127:0]  res_19 = 128'h0;
  wire [127:0]  res_20 = 128'h0;
  wire [127:0]  res_21 = 128'h0;
  wire [127:0]  res_22 = 128'h0;
  wire [127:0]  res_23 = 128'h0;
  wire [127:0]  res_28 = 128'h0;
  wire [127:0]  res_29 = 128'h0;
  wire [127:0]  res_30 = 128'h0;
  wire [127:0]  res_31 = 128'h0;
  wire [127:0]  res_37 = 128'h0;
  wire [127:0]  res_38 = 128'h0;
  wire [127:0]  res_39 = 128'h0;
  wire [127:0]  res_46 = 128'h0;
  wire [127:0]  res_47 = 128'h0;
  wire [127:0]  res_55 = 128'h0;
  wire [127:0]  res_65 = 128'h0;
  wire [127:0]  res_66 = 128'h0;
  wire [127:0]  res_67 = 128'h0;
  wire [127:0]  res_68 = 128'h0;
  wire [127:0]  res_69 = 128'h0;
  wire [127:0]  res_70 = 128'h0;
  wire [127:0]  res_71 = 128'h0;
  wire [127:0]  res_74 = 128'h0;
  wire [127:0]  res_75 = 128'h0;
  wire [127:0]  res_76 = 128'h0;
  wire [127:0]  res_77 = 128'h0;
  wire [127:0]  res_78 = 128'h0;
  wire [127:0]  res_79 = 128'h0;
  wire [127:0]  res_83 = 128'h0;
  wire [127:0]  res_84 = 128'h0;
  wire [127:0]  res_85 = 128'h0;
  wire [127:0]  res_86 = 128'h0;
  wire [127:0]  res_87 = 128'h0;
  wire [127:0]  res_92 = 128'h0;
  wire [127:0]  res_93 = 128'h0;
  wire [127:0]  res_94 = 128'h0;
  wire [127:0]  res_95 = 128'h0;
  wire [127:0]  res_101 = 128'h0;
  wire [127:0]  res_102 = 128'h0;
  wire [127:0]  res_103 = 128'h0;
  wire [127:0]  res_110 = 128'h0;
  wire [127:0]  res_111 = 128'h0;
  wire [127:0]  res_119 = 128'h0;
  wire [127:0]  res_129 = 128'h0;
  wire [127:0]  res_130 = 128'h0;
  wire [127:0]  res_131 = 128'h0;
  wire [127:0]  res_132 = 128'h0;
  wire [127:0]  res_133 = 128'h0;
  wire [127:0]  res_134 = 128'h0;
  wire [127:0]  res_135 = 128'h0;
  wire [127:0]  res_138 = 128'h0;
  wire [127:0]  res_139 = 128'h0;
  wire [127:0]  res_140 = 128'h0;
  wire [127:0]  res_141 = 128'h0;
  wire [127:0]  res_142 = 128'h0;
  wire [127:0]  res_143 = 128'h0;
  wire [127:0]  res_147 = 128'h0;
  wire [127:0]  res_148 = 128'h0;
  wire [127:0]  res_149 = 128'h0;
  wire [127:0]  res_150 = 128'h0;
  wire [127:0]  res_151 = 128'h0;
  wire [127:0]  res_156 = 128'h0;
  wire [127:0]  res_157 = 128'h0;
  wire [127:0]  res_158 = 128'h0;
  wire [127:0]  res_159 = 128'h0;
  wire [127:0]  res_165 = 128'h0;
  wire [127:0]  res_166 = 128'h0;
  wire [127:0]  res_167 = 128'h0;
  wire [127:0]  res_174 = 128'h0;
  wire [127:0]  res_175 = 128'h0;
  wire [127:0]  res_183 = 128'h0;
  wire          vrfWritePort_0_bits_last = 1'h0;
  wire          vrfWritePort_1_bits_last = 1'h0;
  wire          vrfWritePort_2_bits_last = 1'h0;
  wire          vrfWritePort_3_bits_last = 1'h0;
  wire [31:0]   requestAddress;
  wire          unalignedEnqueueReady;
  reg  [2:0]    lsuRequestReg_instructionInformation_nf;
  reg           lsuRequestReg_instructionInformation_mew;
  reg  [1:0]    lsuRequestReg_instructionInformation_mop;
  reg  [4:0]    lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]    lsuRequestReg_instructionInformation_eew;
  reg  [4:0]    lsuRequestReg_instructionInformation_vs3;
  reg           lsuRequestReg_instructionInformation_isStore;
  reg           lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]   lsuRequestReg_rs1Data;
  reg  [31:0]   lsuRequestReg_rs2Data;
  reg  [2:0]    lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_0_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_1_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_2_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_3_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [11:0]   csrInterfaceReg_vl;
  reg  [11:0]   csrInterfaceReg_vStart;
  reg  [2:0]    csrInterfaceReg_vlmul;
  reg  [1:0]    csrInterfaceReg_vSew;
  reg  [1:0]    csrInterfaceReg_vxrm;
  reg           csrInterfaceReg_vta;
  reg           csrInterfaceReg_vma;
  reg           requestFireNext;
  reg  [1:0]    dataEEW;
  wire [3:0]    _dataEEWOH_T = 4'h1 << dataEEW;
  wire [2:0]    dataEEWOH = _dataEEWOH_T[2:0];
  wire          isMaskType = lsuRequest_valid ? lsuRequest_bits_instructionInformation_maskedLoadStore : lsuRequestReg_instructionInformation_maskedLoadStore;
  wire [15:0]   maskAmend = isMaskType ? maskInput : 16'hFFFF;
  reg  [15:0]   maskReg;
  wire [15:0]   _lastMaskAmend_T_1 = 16'h1 << csrInterface_vl[3:0];
  wire [13:0]   _GEN = _lastMaskAmend_T_1[14:1] | _lastMaskAmend_T_1[15:2];
  wire [12:0]   _GEN_0 = _GEN[12:0] | {_lastMaskAmend_T_1[15], _GEN[13:2]};
  wire [10:0]   _GEN_1 = _GEN_0[10:0] | {_lastMaskAmend_T_1[15], _GEN[13], _GEN_0[12:4]};
  wire [14:0]   lastMaskAmend = {_lastMaskAmend_T_1[15], _GEN[13], _GEN_0[12:11], _GEN_1[10:7], _GEN_1[6:0] | {_lastMaskAmend_T_1[15], _GEN[13], _GEN_0[12:11], _GEN_1[10:8]}};
  reg           needAmend;
  reg  [14:0]   lastMaskAmendReg;
  wire [1:0]    countEndForGroup = {1'h0, dataEEWOH[1]} | {2{dataEEWOH[2]}};
  reg  [6:0]    maskGroupCounter;
  wire [6:0]    nextMaskGroup = maskGroupCounter + 7'h1;
  reg  [1:0]    maskCounterInGroup;
  wire [1:0]    nextMaskCount = maskCounterInGroup + 2'h1;
  wire          isLastDataGroup = maskCounterInGroup == countEndForGroup;
  wire [6:0]    _maskSelect_bits_output = lsuRequest_valid ? 7'h0 : nextMaskGroup;
  reg  [15:0]   maskForGroup;
  reg           isLastMaskGroup;
  wire [15:0]   maskWire = maskReg & (needAmend & isLastMaskGroup ? {1'h0, lastMaskAmendReg} : 16'hFFFF);
  wire [3:0]    maskForGroupWire_lo_lo_lo = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]    maskForGroupWire_lo_lo = {maskForGroupWire_lo_lo_hi, maskForGroupWire_lo_lo_lo};
  wire [3:0]    maskForGroupWire_lo_hi_lo = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]    maskForGroupWire_lo_hi = {maskForGroupWire_lo_hi_hi, maskForGroupWire_lo_hi_lo};
  wire [15:0]   maskForGroupWire_lo = {maskForGroupWire_lo_hi, maskForGroupWire_lo_lo};
  wire [3:0]    maskForGroupWire_hi_lo_lo = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]    maskForGroupWire_hi_lo = {maskForGroupWire_hi_lo_hi, maskForGroupWire_hi_lo_lo};
  wire [3:0]    maskForGroupWire_hi_hi_lo = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]    maskForGroupWire_hi_hi = {maskForGroupWire_hi_hi_hi, maskForGroupWire_hi_hi_lo};
  wire [15:0]   maskForGroupWire_hi = {maskForGroupWire_hi_hi, maskForGroupWire_hi_lo};
  wire [3:0]    maskForGroupWire_lo_lo_lo_1 = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi_1 = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]    maskForGroupWire_lo_lo_1 = {maskForGroupWire_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_hi_lo_1 = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi_1 = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]    maskForGroupWire_lo_hi_1 = {maskForGroupWire_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_1};
  wire [15:0]   maskForGroupWire_lo_1 = {maskForGroupWire_lo_hi_1, maskForGroupWire_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_lo_lo_1 = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi_1 = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]    maskForGroupWire_hi_lo_1 = {maskForGroupWire_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_hi_lo_1 = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi_1 = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]    maskForGroupWire_hi_hi_1 = {maskForGroupWire_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_1};
  wire [15:0]   maskForGroupWire_hi_1 = {maskForGroupWire_hi_hi_1, maskForGroupWire_hi_lo_1};
  wire [3:0]    _maskForGroupWire_T_69 = 4'h1 << maskCounterInGroup;
  wire [7:0]    maskForGroupWire_lo_lo_lo_2 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_2 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_2 = {maskForGroupWire_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_hi_lo_2 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_2 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_hi_2 = {maskForGroupWire_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_2};
  wire [31:0]   maskForGroupWire_lo_2 = {maskForGroupWire_lo_hi_2, maskForGroupWire_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_lo_lo_2 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_2 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_hi_lo_2 = {maskForGroupWire_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_hi_lo_2 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_2 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_hi_hi_2 = {maskForGroupWire_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_2};
  wire [31:0]   maskForGroupWire_hi_2 = {maskForGroupWire_hi_hi_2, maskForGroupWire_hi_lo_2};
  wire [7:0]    maskForGroupWire_lo_lo_lo_3 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_3 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_3 = {maskForGroupWire_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_hi_lo_3 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_3 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_hi_3 = {maskForGroupWire_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_3};
  wire [31:0]   maskForGroupWire_lo_3 = {maskForGroupWire_lo_hi_3, maskForGroupWire_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_lo_lo_3 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_3 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_hi_lo_3 = {maskForGroupWire_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_hi_lo_3 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_3 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_hi_hi_3 = {maskForGroupWire_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_3};
  wire [31:0]   maskForGroupWire_hi_3 = {maskForGroupWire_hi_hi_3, maskForGroupWire_hi_lo_3};
  wire [7:0]    maskForGroupWire_lo_lo_lo_4 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_4 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_4 = {maskForGroupWire_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_hi_lo_4 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_4 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_hi_4 = {maskForGroupWire_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_4};
  wire [31:0]   maskForGroupWire_lo_4 = {maskForGroupWire_lo_hi_4, maskForGroupWire_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_lo_lo_4 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_4 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_hi_lo_4 = {maskForGroupWire_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_hi_lo_4 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_4 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_hi_hi_4 = {maskForGroupWire_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_4};
  wire [31:0]   maskForGroupWire_hi_4 = {maskForGroupWire_hi_hi_4, maskForGroupWire_hi_lo_4};
  wire [7:0]    maskForGroupWire_lo_lo_lo_5 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_5 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_5 = {maskForGroupWire_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_hi_lo_5 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_5 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_hi_5 = {maskForGroupWire_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_5};
  wire [31:0]   maskForGroupWire_lo_5 = {maskForGroupWire_lo_hi_5, maskForGroupWire_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_lo_lo_5 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_5 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_hi_lo_5 = {maskForGroupWire_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_hi_lo_5 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_5 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_hi_hi_5 = {maskForGroupWire_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_5};
  wire [31:0]   maskForGroupWire_hi_5 = {maskForGroupWire_hi_hi_5, maskForGroupWire_hi_lo_5};
  wire [15:0]   maskForGroupWire =
    (dataEEWOH[0] ? maskWire : 16'h0) | (dataEEWOH[1] ? (maskCounterInGroup[0] ? maskForGroupWire_hi : maskForGroupWire_lo_1) : 16'h0)
    | (dataEEWOH[2]
         ? (_maskForGroupWire_T_69[0] ? maskForGroupWire_lo_2[15:0] : 16'h0) | (_maskForGroupWire_T_69[1] ? maskForGroupWire_lo_3[31:16] : 16'h0) | (_maskForGroupWire_T_69[2] ? maskForGroupWire_hi_4[15:0] : 16'h0)
           | (_maskForGroupWire_T_69[3] ? maskForGroupWire_hi_5[31:16] : 16'h0)
         : 16'h0);
  wire [1:0]    initSendState_lo = maskForGroupWire[1:0];
  wire [1:0]    initSendState_hi = maskForGroupWire[3:2];
  wire          initSendState_0 = |{initSendState_hi, initSendState_lo};
  wire [1:0]    initSendState_lo_1 = maskForGroupWire[5:4];
  wire [1:0]    initSendState_hi_1 = maskForGroupWire[7:6];
  wire          initSendState_1 = |{initSendState_hi_1, initSendState_lo_1};
  wire [1:0]    initSendState_lo_2 = maskForGroupWire[9:8];
  wire [1:0]    initSendState_hi_2 = maskForGroupWire[11:10];
  wire          initSendState_2 = |{initSendState_hi_2, initSendState_lo_2};
  wire [1:0]    initSendState_lo_3 = maskForGroupWire[13:12];
  wire [1:0]    initSendState_hi_3 = maskForGroupWire[15:14];
  wire          initSendState_3 = |{initSendState_hi_3, initSendState_lo_3};
  reg  [127:0]  accessData_0;
  reg  [127:0]  accessData_1;
  reg  [127:0]  accessData_2;
  reg  [127:0]  accessData_3;
  reg  [127:0]  accessData_4;
  reg  [127:0]  accessData_5;
  reg  [127:0]  accessData_6;
  reg  [127:0]  accessData_7;
  reg  [2:0]    accessPtr;
  reg           accessState_0;
  reg           accessState_1;
  reg           accessState_2;
  reg           accessState_3;
  wire          accessStateUpdate_0;
  wire          accessStateUpdate_1;
  wire [1:0]    accessStateCheck_lo = {accessStateUpdate_1, accessStateUpdate_0};
  wire          accessStateUpdate_2;
  wire          accessStateUpdate_3;
  wire [1:0]    accessStateCheck_hi = {accessStateUpdate_3, accessStateUpdate_2};
  wire          accessStateCheck = {accessStateCheck_hi, accessStateCheck_lo} == 4'h0;
  reg  [6:0]    dataGroup;
  reg  [127:0]  dataBuffer_0;
  reg  [127:0]  dataBuffer_1;
  reg  [127:0]  dataBuffer_2;
  reg  [127:0]  dataBuffer_3;
  reg  [127:0]  dataBuffer_4;
  reg  [127:0]  dataBuffer_5;
  reg  [127:0]  dataBuffer_6;
  reg  [127:0]  dataBuffer_7;
  reg  [7:0]    bufferBaseCacheLineIndex;
  reg  [2:0]    cacheLineIndexInBuffer;
  wire [3:0]    initOffset = lsuRequestReg_rs1Data[3:0];
  wire          invalidInstruction = csrInterface_vl == 12'h0;
  reg           invalidInstructionNext;
  wire          wholeType = lsuRequest_bits_instructionInformation_lumop[3];
  wire [2:0]    nfCorrection = wholeType ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [3:0]    segmentInstructionIndexInterval;
  wire [18:0]   bytePerInstruction = {3'h0, {12'h0, {1'h0, nfCorrection} + 4'h1} * {4'h0, csrInterface_vl}} << lsuRequest_bits_instructionInformation_eew;
  wire [18:0]   accessMemSize = bytePerInstruction + {15'h0, lsuRequest_bits_rs1Data[3:0]};
  wire [14:0]   lastCacheLineIndex = accessMemSize[18:4] - {14'h0, accessMemSize[3:0] == 4'h0};
  wire [14:0]   lastWriteVrfIndex = bytePerInstruction[18:4] - {14'h0, bytePerInstruction[3:0] == 4'h0};
  reg  [14:0]   lastWriteVrfIndexReg;
  reg           lastCacheNeedPush;
  reg  [14:0]   cacheLineNumberReg;
  wire          memRequest_valid_0;
  wire          _lastCacheRequest_T = memRequest_ready_0 & memRequest_valid_0;
  reg  [7:0]    cacheLineIndex;
  wire [7:0]    memRequest_bits_src_0 = cacheLineIndex;
  wire [7:0]    nextCacheLineIndex = cacheLineIndex + 8'h1;
  wire          validInstruction = ~invalidInstruction & lsuRequest_valid;
  wire          lastRequest = cacheLineNumberReg == {7'h0, cacheLineIndex};
  reg           sendRequest;
  assign requestAddress = {lsuRequestReg_rs1Data[31:4] + {20'h0, cacheLineIndex}, 4'h0};
  wire [31:0]   memRequest_bits_address_0 = requestAddress;
  reg           writeReadyReg;
  assign memRequest_valid_0 = sendRequest & ~addressConflict;
  wire          memResponse_ready_0;
  wire          unalignedEnqueueFire = memResponse_ready_0 & memResponse_valid_0;
  wire          anyLastCacheLineAck = unalignedEnqueueFire & {7'h0, memResponse_bits_index_0} == cacheLineNumberReg;
  wire          alignedDequeueValid;
  wire [127:0]  alignedDequeue_bits_data_lo_40;
  reg           unalignedCacheLine_valid;
  reg  [127:0]  unalignedCacheLine_bits_data;
  reg  [7:0]    unalignedCacheLine_bits_index;
  wire [7:0]    alignedDequeue_bits_index = unalignedCacheLine_bits_index;
  wire          alignedDequeue_ready;
  assign unalignedEnqueueReady = alignedDequeue_ready | ~unalignedCacheLine_valid;
  assign memResponse_ready_0 = unalignedEnqueueReady;
  wire [7:0]    nextIndex = unalignedCacheLine_valid ? unalignedCacheLine_bits_index + 8'h1 : 8'h0;
  assign alignedDequeueValid = unalignedCacheLine_valid & (memResponse_valid_0 | {7'h0, unalignedCacheLine_bits_index} == cacheLineNumberReg & lastCacheNeedPush);
  wire          alignedDequeue_valid = alignedDequeueValid;
  wire          _bufferTailFire_T = alignedDequeue_ready & alignedDequeue_valid;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo = {unalignedCacheLine_bits_data[8], unalignedCacheLine_bits_data[0]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi = {unalignedCacheLine_bits_data[24], unalignedCacheLine_bits_data[16]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo = {alignedDequeue_bits_data_lo_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo = {unalignedCacheLine_bits_data[40], unalignedCacheLine_bits_data[32]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi = {unalignedCacheLine_bits_data[56], unalignedCacheLine_bits_data[48]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi = {alignedDequeue_bits_data_lo_lo_hi_hi, alignedDequeue_bits_data_lo_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_lo = {alignedDequeue_bits_data_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo = {unalignedCacheLine_bits_data[72], unalignedCacheLine_bits_data[64]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi = {unalignedCacheLine_bits_data[88], unalignedCacheLine_bits_data[80]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo = {alignedDequeue_bits_data_lo_hi_lo_hi, alignedDequeue_bits_data_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo = {unalignedCacheLine_bits_data[104], unalignedCacheLine_bits_data[96]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi = {unalignedCacheLine_bits_data[120], unalignedCacheLine_bits_data[112]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi = {alignedDequeue_bits_data_lo_hi_hi_hi, alignedDequeue_bits_data_lo_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_hi = {alignedDequeue_bits_data_lo_hi_hi, alignedDequeue_bits_data_lo_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_lo = {alignedDequeue_bits_data_lo_hi, alignedDequeue_bits_data_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo = {memResponse_bits_data_0[8], memResponse_bits_data_0[0]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi = {memResponse_bits_data_0[24], memResponse_bits_data_0[16]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo = {alignedDequeue_bits_data_hi_lo_lo_hi, alignedDequeue_bits_data_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo = {memResponse_bits_data_0[40], memResponse_bits_data_0[32]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi = {memResponse_bits_data_0[56], memResponse_bits_data_0[48]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi = {alignedDequeue_bits_data_hi_lo_hi_hi, alignedDequeue_bits_data_hi_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_lo = {alignedDequeue_bits_data_hi_lo_hi, alignedDequeue_bits_data_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo = {memResponse_bits_data_0[72], memResponse_bits_data_0[64]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi = {memResponse_bits_data_0[88], memResponse_bits_data_0[80]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo = {alignedDequeue_bits_data_hi_hi_lo_hi, alignedDequeue_bits_data_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo = {memResponse_bits_data_0[104], memResponse_bits_data_0[96]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi = {memResponse_bits_data_0[120], memResponse_bits_data_0[112]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi = {alignedDequeue_bits_data_hi_hi_hi_hi, alignedDequeue_bits_data_hi_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_hi = {alignedDequeue_bits_data_hi_hi_hi, alignedDequeue_bits_data_hi_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_hi = {alignedDequeue_bits_data_hi_hi, alignedDequeue_bits_data_hi_lo};
  wire [31:0]   _GEN_2 = {28'h0, initOffset};
  wire [31:0]   _alignedDequeue_bits_data_T_258 = {alignedDequeue_bits_data_hi, alignedDequeue_bits_data_lo} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_1 = {unalignedCacheLine_bits_data[9], unalignedCacheLine_bits_data[1]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_1 = {unalignedCacheLine_bits_data[25], unalignedCacheLine_bits_data[17]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_1 = {unalignedCacheLine_bits_data[41], unalignedCacheLine_bits_data[33]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_1 = {unalignedCacheLine_bits_data[57], unalignedCacheLine_bits_data[49]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_1 = {alignedDequeue_bits_data_lo_lo_hi_hi_1, alignedDequeue_bits_data_lo_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_1 = {unalignedCacheLine_bits_data[73], unalignedCacheLine_bits_data[65]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_1 = {unalignedCacheLine_bits_data[89], unalignedCacheLine_bits_data[81]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_1 = {alignedDequeue_bits_data_lo_hi_lo_hi_1, alignedDequeue_bits_data_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_1 = {unalignedCacheLine_bits_data[105], unalignedCacheLine_bits_data[97]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_1 = {unalignedCacheLine_bits_data[121], unalignedCacheLine_bits_data[113]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_hi_1, alignedDequeue_bits_data_lo_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_1, alignedDequeue_bits_data_lo_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_lo_1 = {alignedDequeue_bits_data_lo_hi_1, alignedDequeue_bits_data_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_1 = {memResponse_bits_data_0[9], memResponse_bits_data_0[1]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_1 = {memResponse_bits_data_0[25], memResponse_bits_data_0[17]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_1 = {alignedDequeue_bits_data_hi_lo_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_1 = {memResponse_bits_data_0[41], memResponse_bits_data_0[33]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_1 = {memResponse_bits_data_0[57], memResponse_bits_data_0[49]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_1 = {alignedDequeue_bits_data_hi_lo_hi_hi_1, alignedDequeue_bits_data_hi_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_1 = {alignedDequeue_bits_data_hi_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_1 = {memResponse_bits_data_0[73], memResponse_bits_data_0[65]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_1 = {memResponse_bits_data_0[89], memResponse_bits_data_0[81]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_1 = {alignedDequeue_bits_data_hi_hi_lo_hi_1, alignedDequeue_bits_data_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_1 = {memResponse_bits_data_0[105], memResponse_bits_data_0[97]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_1 = {memResponse_bits_data_0[121], memResponse_bits_data_0[113]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_hi_1 = {alignedDequeue_bits_data_hi_hi_1, alignedDequeue_bits_data_hi_lo_1};
  wire [31:0]   _alignedDequeue_bits_data_T_292 = {alignedDequeue_bits_data_hi_1, alignedDequeue_bits_data_lo_1} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_2 = {unalignedCacheLine_bits_data[10], unalignedCacheLine_bits_data[2]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_2 = {unalignedCacheLine_bits_data[26], unalignedCacheLine_bits_data[18]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_2 = {unalignedCacheLine_bits_data[42], unalignedCacheLine_bits_data[34]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_2 = {unalignedCacheLine_bits_data[58], unalignedCacheLine_bits_data[50]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_2 = {alignedDequeue_bits_data_lo_lo_hi_hi_2, alignedDequeue_bits_data_lo_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_2 = {unalignedCacheLine_bits_data[74], unalignedCacheLine_bits_data[66]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_2 = {unalignedCacheLine_bits_data[90], unalignedCacheLine_bits_data[82]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_2 = {alignedDequeue_bits_data_lo_hi_lo_hi_2, alignedDequeue_bits_data_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_2 = {unalignedCacheLine_bits_data[106], unalignedCacheLine_bits_data[98]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_2 = {unalignedCacheLine_bits_data[122], unalignedCacheLine_bits_data[114]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_hi_2, alignedDequeue_bits_data_lo_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_2, alignedDequeue_bits_data_lo_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_lo_2 = {alignedDequeue_bits_data_lo_hi_2, alignedDequeue_bits_data_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_2 = {memResponse_bits_data_0[10], memResponse_bits_data_0[2]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_2 = {memResponse_bits_data_0[26], memResponse_bits_data_0[18]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_2 = {alignedDequeue_bits_data_hi_lo_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_2 = {memResponse_bits_data_0[42], memResponse_bits_data_0[34]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_2 = {memResponse_bits_data_0[58], memResponse_bits_data_0[50]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_2 = {alignedDequeue_bits_data_hi_lo_hi_hi_2, alignedDequeue_bits_data_hi_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_2 = {alignedDequeue_bits_data_hi_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_2 = {memResponse_bits_data_0[74], memResponse_bits_data_0[66]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_2 = {memResponse_bits_data_0[90], memResponse_bits_data_0[82]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_2 = {alignedDequeue_bits_data_hi_hi_lo_hi_2, alignedDequeue_bits_data_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_2 = {memResponse_bits_data_0[106], memResponse_bits_data_0[98]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_2 = {memResponse_bits_data_0[122], memResponse_bits_data_0[114]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_hi_2 = {alignedDequeue_bits_data_hi_hi_2, alignedDequeue_bits_data_hi_lo_2};
  wire [31:0]   _alignedDequeue_bits_data_T_326 = {alignedDequeue_bits_data_hi_2, alignedDequeue_bits_data_lo_2} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_3 = {unalignedCacheLine_bits_data[11], unalignedCacheLine_bits_data[3]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_3 = {unalignedCacheLine_bits_data[27], unalignedCacheLine_bits_data[19]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_3 = {unalignedCacheLine_bits_data[43], unalignedCacheLine_bits_data[35]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_3 = {unalignedCacheLine_bits_data[59], unalignedCacheLine_bits_data[51]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_3 = {alignedDequeue_bits_data_lo_lo_hi_hi_3, alignedDequeue_bits_data_lo_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_3 = {unalignedCacheLine_bits_data[75], unalignedCacheLine_bits_data[67]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_3 = {unalignedCacheLine_bits_data[91], unalignedCacheLine_bits_data[83]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_3 = {alignedDequeue_bits_data_lo_hi_lo_hi_3, alignedDequeue_bits_data_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_3 = {unalignedCacheLine_bits_data[107], unalignedCacheLine_bits_data[99]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_3 = {unalignedCacheLine_bits_data[123], unalignedCacheLine_bits_data[115]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_hi_3, alignedDequeue_bits_data_lo_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_3, alignedDequeue_bits_data_lo_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_lo_3 = {alignedDequeue_bits_data_lo_hi_3, alignedDequeue_bits_data_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_3 = {memResponse_bits_data_0[11], memResponse_bits_data_0[3]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_3 = {memResponse_bits_data_0[27], memResponse_bits_data_0[19]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_3 = {alignedDequeue_bits_data_hi_lo_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_3 = {memResponse_bits_data_0[43], memResponse_bits_data_0[35]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_3 = {memResponse_bits_data_0[59], memResponse_bits_data_0[51]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_3 = {alignedDequeue_bits_data_hi_lo_hi_hi_3, alignedDequeue_bits_data_hi_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_3 = {alignedDequeue_bits_data_hi_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_3 = {memResponse_bits_data_0[75], memResponse_bits_data_0[67]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_3 = {memResponse_bits_data_0[91], memResponse_bits_data_0[83]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_3 = {alignedDequeue_bits_data_hi_hi_lo_hi_3, alignedDequeue_bits_data_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_3 = {memResponse_bits_data_0[107], memResponse_bits_data_0[99]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_3 = {memResponse_bits_data_0[123], memResponse_bits_data_0[115]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_hi_3 = {alignedDequeue_bits_data_hi_hi_3, alignedDequeue_bits_data_hi_lo_3};
  wire [31:0]   _alignedDequeue_bits_data_T_360 = {alignedDequeue_bits_data_hi_3, alignedDequeue_bits_data_lo_3} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_4 = {unalignedCacheLine_bits_data[12], unalignedCacheLine_bits_data[4]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_4 = {unalignedCacheLine_bits_data[28], unalignedCacheLine_bits_data[20]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_4 = {unalignedCacheLine_bits_data[44], unalignedCacheLine_bits_data[36]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_4 = {unalignedCacheLine_bits_data[60], unalignedCacheLine_bits_data[52]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_4 = {alignedDequeue_bits_data_lo_lo_hi_hi_4, alignedDequeue_bits_data_lo_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_4 = {unalignedCacheLine_bits_data[76], unalignedCacheLine_bits_data[68]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_4 = {unalignedCacheLine_bits_data[92], unalignedCacheLine_bits_data[84]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_4 = {alignedDequeue_bits_data_lo_hi_lo_hi_4, alignedDequeue_bits_data_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_4 = {unalignedCacheLine_bits_data[108], unalignedCacheLine_bits_data[100]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_4 = {unalignedCacheLine_bits_data[124], unalignedCacheLine_bits_data[116]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_hi_4, alignedDequeue_bits_data_lo_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_4, alignedDequeue_bits_data_lo_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_lo_4 = {alignedDequeue_bits_data_lo_hi_4, alignedDequeue_bits_data_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_4 = {memResponse_bits_data_0[12], memResponse_bits_data_0[4]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_4 = {memResponse_bits_data_0[28], memResponse_bits_data_0[20]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_4 = {alignedDequeue_bits_data_hi_lo_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_4 = {memResponse_bits_data_0[44], memResponse_bits_data_0[36]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_4 = {memResponse_bits_data_0[60], memResponse_bits_data_0[52]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_4 = {alignedDequeue_bits_data_hi_lo_hi_hi_4, alignedDequeue_bits_data_hi_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_4 = {alignedDequeue_bits_data_hi_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_4 = {memResponse_bits_data_0[76], memResponse_bits_data_0[68]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_4 = {memResponse_bits_data_0[92], memResponse_bits_data_0[84]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_4 = {alignedDequeue_bits_data_hi_hi_lo_hi_4, alignedDequeue_bits_data_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_4 = {memResponse_bits_data_0[108], memResponse_bits_data_0[100]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_4 = {memResponse_bits_data_0[124], memResponse_bits_data_0[116]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_hi_4 = {alignedDequeue_bits_data_hi_hi_4, alignedDequeue_bits_data_hi_lo_4};
  wire [31:0]   _alignedDequeue_bits_data_T_394 = {alignedDequeue_bits_data_hi_4, alignedDequeue_bits_data_lo_4} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_5 = {unalignedCacheLine_bits_data[13], unalignedCacheLine_bits_data[5]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_5 = {unalignedCacheLine_bits_data[29], unalignedCacheLine_bits_data[21]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_5 = {unalignedCacheLine_bits_data[45], unalignedCacheLine_bits_data[37]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_5 = {unalignedCacheLine_bits_data[61], unalignedCacheLine_bits_data[53]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_5 = {alignedDequeue_bits_data_lo_lo_hi_hi_5, alignedDequeue_bits_data_lo_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_5 = {unalignedCacheLine_bits_data[77], unalignedCacheLine_bits_data[69]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_5 = {unalignedCacheLine_bits_data[93], unalignedCacheLine_bits_data[85]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_5 = {alignedDequeue_bits_data_lo_hi_lo_hi_5, alignedDequeue_bits_data_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_5 = {unalignedCacheLine_bits_data[109], unalignedCacheLine_bits_data[101]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_5 = {unalignedCacheLine_bits_data[125], unalignedCacheLine_bits_data[117]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_hi_5, alignedDequeue_bits_data_lo_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_5, alignedDequeue_bits_data_lo_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_lo_5 = {alignedDequeue_bits_data_lo_hi_5, alignedDequeue_bits_data_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_5 = {memResponse_bits_data_0[13], memResponse_bits_data_0[5]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_5 = {memResponse_bits_data_0[29], memResponse_bits_data_0[21]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_5 = {alignedDequeue_bits_data_hi_lo_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_5 = {memResponse_bits_data_0[45], memResponse_bits_data_0[37]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_5 = {memResponse_bits_data_0[61], memResponse_bits_data_0[53]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_5 = {alignedDequeue_bits_data_hi_lo_hi_hi_5, alignedDequeue_bits_data_hi_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_5 = {alignedDequeue_bits_data_hi_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_5 = {memResponse_bits_data_0[77], memResponse_bits_data_0[69]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_5 = {memResponse_bits_data_0[93], memResponse_bits_data_0[85]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_5 = {alignedDequeue_bits_data_hi_hi_lo_hi_5, alignedDequeue_bits_data_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_5 = {memResponse_bits_data_0[109], memResponse_bits_data_0[101]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_5 = {memResponse_bits_data_0[125], memResponse_bits_data_0[117]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_hi_5 = {alignedDequeue_bits_data_hi_hi_5, alignedDequeue_bits_data_hi_lo_5};
  wire [31:0]   _alignedDequeue_bits_data_T_428 = {alignedDequeue_bits_data_hi_5, alignedDequeue_bits_data_lo_5} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_6 = {unalignedCacheLine_bits_data[14], unalignedCacheLine_bits_data[6]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_6 = {unalignedCacheLine_bits_data[30], unalignedCacheLine_bits_data[22]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_6 = {unalignedCacheLine_bits_data[46], unalignedCacheLine_bits_data[38]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_6 = {unalignedCacheLine_bits_data[62], unalignedCacheLine_bits_data[54]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_6 = {alignedDequeue_bits_data_lo_lo_hi_hi_6, alignedDequeue_bits_data_lo_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_6 = {unalignedCacheLine_bits_data[78], unalignedCacheLine_bits_data[70]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_6 = {unalignedCacheLine_bits_data[94], unalignedCacheLine_bits_data[86]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_6 = {alignedDequeue_bits_data_lo_hi_lo_hi_6, alignedDequeue_bits_data_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_6 = {unalignedCacheLine_bits_data[110], unalignedCacheLine_bits_data[102]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_6 = {unalignedCacheLine_bits_data[126], unalignedCacheLine_bits_data[118]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_hi_6, alignedDequeue_bits_data_lo_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_6, alignedDequeue_bits_data_lo_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_lo_6 = {alignedDequeue_bits_data_lo_hi_6, alignedDequeue_bits_data_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_6 = {memResponse_bits_data_0[14], memResponse_bits_data_0[6]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_6 = {memResponse_bits_data_0[30], memResponse_bits_data_0[22]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_6 = {alignedDequeue_bits_data_hi_lo_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_6 = {memResponse_bits_data_0[46], memResponse_bits_data_0[38]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_6 = {memResponse_bits_data_0[62], memResponse_bits_data_0[54]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_6 = {alignedDequeue_bits_data_hi_lo_hi_hi_6, alignedDequeue_bits_data_hi_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_6 = {alignedDequeue_bits_data_hi_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_6 = {memResponse_bits_data_0[78], memResponse_bits_data_0[70]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_6 = {memResponse_bits_data_0[94], memResponse_bits_data_0[86]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_6 = {alignedDequeue_bits_data_hi_hi_lo_hi_6, alignedDequeue_bits_data_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_6 = {memResponse_bits_data_0[110], memResponse_bits_data_0[102]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_6 = {memResponse_bits_data_0[126], memResponse_bits_data_0[118]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_hi_6 = {alignedDequeue_bits_data_hi_hi_6, alignedDequeue_bits_data_hi_lo_6};
  wire [31:0]   _alignedDequeue_bits_data_T_462 = {alignedDequeue_bits_data_hi_6, alignedDequeue_bits_data_lo_6} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_7 = {unalignedCacheLine_bits_data[15], unalignedCacheLine_bits_data[7]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_7 = {unalignedCacheLine_bits_data[31], unalignedCacheLine_bits_data[23]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_7 = {unalignedCacheLine_bits_data[47], unalignedCacheLine_bits_data[39]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_7 = {unalignedCacheLine_bits_data[63], unalignedCacheLine_bits_data[55]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_7 = {alignedDequeue_bits_data_lo_lo_hi_hi_7, alignedDequeue_bits_data_lo_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_7 = {unalignedCacheLine_bits_data[79], unalignedCacheLine_bits_data[71]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_7 = {unalignedCacheLine_bits_data[95], unalignedCacheLine_bits_data[87]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_7 = {alignedDequeue_bits_data_lo_hi_lo_hi_7, alignedDequeue_bits_data_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_7 = {unalignedCacheLine_bits_data[111], unalignedCacheLine_bits_data[103]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_7 = {unalignedCacheLine_bits_data[127], unalignedCacheLine_bits_data[119]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_hi_7, alignedDequeue_bits_data_lo_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_7, alignedDequeue_bits_data_lo_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_lo_7 = {alignedDequeue_bits_data_lo_hi_7, alignedDequeue_bits_data_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_7 = {memResponse_bits_data_0[15], memResponse_bits_data_0[7]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_7 = {memResponse_bits_data_0[31], memResponse_bits_data_0[23]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_7 = {alignedDequeue_bits_data_hi_lo_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_7 = {memResponse_bits_data_0[47], memResponse_bits_data_0[39]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_7 = {memResponse_bits_data_0[63], memResponse_bits_data_0[55]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_7 = {alignedDequeue_bits_data_hi_lo_hi_hi_7, alignedDequeue_bits_data_hi_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_7 = {alignedDequeue_bits_data_hi_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_7 = {memResponse_bits_data_0[79], memResponse_bits_data_0[71]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_7 = {memResponse_bits_data_0[95], memResponse_bits_data_0[87]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_7 = {alignedDequeue_bits_data_hi_hi_lo_hi_7, alignedDequeue_bits_data_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_7 = {memResponse_bits_data_0[111], memResponse_bits_data_0[103]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_7 = {memResponse_bits_data_0[127], memResponse_bits_data_0[119]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_hi_7 = {alignedDequeue_bits_data_hi_hi_7, alignedDequeue_bits_data_hi_lo_7};
  wire [31:0]   _alignedDequeue_bits_data_T_496 = {alignedDequeue_bits_data_hi_7, alignedDequeue_bits_data_lo_7} >> _GEN_2;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_8 = {_alignedDequeue_bits_data_T_292[0], _alignedDequeue_bits_data_T_258[0]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_8 = {_alignedDequeue_bits_data_T_360[0], _alignedDequeue_bits_data_T_326[0]};
  wire [3:0]    alignedDequeue_bits_data_lo_8 = {alignedDequeue_bits_data_lo_hi_8, alignedDequeue_bits_data_lo_lo_8};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_8 = {_alignedDequeue_bits_data_T_428[0], _alignedDequeue_bits_data_T_394[0]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_8 = {_alignedDequeue_bits_data_T_496[0], _alignedDequeue_bits_data_T_462[0]};
  wire [3:0]    alignedDequeue_bits_data_hi_8 = {alignedDequeue_bits_data_hi_hi_8, alignedDequeue_bits_data_hi_lo_8};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_9 = {_alignedDequeue_bits_data_T_292[1], _alignedDequeue_bits_data_T_258[1]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_9 = {_alignedDequeue_bits_data_T_360[1], _alignedDequeue_bits_data_T_326[1]};
  wire [3:0]    alignedDequeue_bits_data_lo_9 = {alignedDequeue_bits_data_lo_hi_9, alignedDequeue_bits_data_lo_lo_9};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_9 = {_alignedDequeue_bits_data_T_428[1], _alignedDequeue_bits_data_T_394[1]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_9 = {_alignedDequeue_bits_data_T_496[1], _alignedDequeue_bits_data_T_462[1]};
  wire [3:0]    alignedDequeue_bits_data_hi_9 = {alignedDequeue_bits_data_hi_hi_9, alignedDequeue_bits_data_hi_lo_9};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_10 = {_alignedDequeue_bits_data_T_292[2], _alignedDequeue_bits_data_T_258[2]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_10 = {_alignedDequeue_bits_data_T_360[2], _alignedDequeue_bits_data_T_326[2]};
  wire [3:0]    alignedDequeue_bits_data_lo_10 = {alignedDequeue_bits_data_lo_hi_10, alignedDequeue_bits_data_lo_lo_10};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_10 = {_alignedDequeue_bits_data_T_428[2], _alignedDequeue_bits_data_T_394[2]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_10 = {_alignedDequeue_bits_data_T_496[2], _alignedDequeue_bits_data_T_462[2]};
  wire [3:0]    alignedDequeue_bits_data_hi_10 = {alignedDequeue_bits_data_hi_hi_10, alignedDequeue_bits_data_hi_lo_10};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_11 = {_alignedDequeue_bits_data_T_292[3], _alignedDequeue_bits_data_T_258[3]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_11 = {_alignedDequeue_bits_data_T_360[3], _alignedDequeue_bits_data_T_326[3]};
  wire [3:0]    alignedDequeue_bits_data_lo_11 = {alignedDequeue_bits_data_lo_hi_11, alignedDequeue_bits_data_lo_lo_11};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_11 = {_alignedDequeue_bits_data_T_428[3], _alignedDequeue_bits_data_T_394[3]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_11 = {_alignedDequeue_bits_data_T_496[3], _alignedDequeue_bits_data_T_462[3]};
  wire [3:0]    alignedDequeue_bits_data_hi_11 = {alignedDequeue_bits_data_hi_hi_11, alignedDequeue_bits_data_hi_lo_11};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_12 = {_alignedDequeue_bits_data_T_292[4], _alignedDequeue_bits_data_T_258[4]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_12 = {_alignedDequeue_bits_data_T_360[4], _alignedDequeue_bits_data_T_326[4]};
  wire [3:0]    alignedDequeue_bits_data_lo_12 = {alignedDequeue_bits_data_lo_hi_12, alignedDequeue_bits_data_lo_lo_12};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_12 = {_alignedDequeue_bits_data_T_428[4], _alignedDequeue_bits_data_T_394[4]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_12 = {_alignedDequeue_bits_data_T_496[4], _alignedDequeue_bits_data_T_462[4]};
  wire [3:0]    alignedDequeue_bits_data_hi_12 = {alignedDequeue_bits_data_hi_hi_12, alignedDequeue_bits_data_hi_lo_12};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_13 = {_alignedDequeue_bits_data_T_292[5], _alignedDequeue_bits_data_T_258[5]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_13 = {_alignedDequeue_bits_data_T_360[5], _alignedDequeue_bits_data_T_326[5]};
  wire [3:0]    alignedDequeue_bits_data_lo_13 = {alignedDequeue_bits_data_lo_hi_13, alignedDequeue_bits_data_lo_lo_13};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_13 = {_alignedDequeue_bits_data_T_428[5], _alignedDequeue_bits_data_T_394[5]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_13 = {_alignedDequeue_bits_data_T_496[5], _alignedDequeue_bits_data_T_462[5]};
  wire [3:0]    alignedDequeue_bits_data_hi_13 = {alignedDequeue_bits_data_hi_hi_13, alignedDequeue_bits_data_hi_lo_13};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_14 = {_alignedDequeue_bits_data_T_292[6], _alignedDequeue_bits_data_T_258[6]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_14 = {_alignedDequeue_bits_data_T_360[6], _alignedDequeue_bits_data_T_326[6]};
  wire [3:0]    alignedDequeue_bits_data_lo_14 = {alignedDequeue_bits_data_lo_hi_14, alignedDequeue_bits_data_lo_lo_14};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_14 = {_alignedDequeue_bits_data_T_428[6], _alignedDequeue_bits_data_T_394[6]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_14 = {_alignedDequeue_bits_data_T_496[6], _alignedDequeue_bits_data_T_462[6]};
  wire [3:0]    alignedDequeue_bits_data_hi_14 = {alignedDequeue_bits_data_hi_hi_14, alignedDequeue_bits_data_hi_lo_14};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_15 = {_alignedDequeue_bits_data_T_292[7], _alignedDequeue_bits_data_T_258[7]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_15 = {_alignedDequeue_bits_data_T_360[7], _alignedDequeue_bits_data_T_326[7]};
  wire [3:0]    alignedDequeue_bits_data_lo_15 = {alignedDequeue_bits_data_lo_hi_15, alignedDequeue_bits_data_lo_lo_15};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_15 = {_alignedDequeue_bits_data_T_428[7], _alignedDequeue_bits_data_T_394[7]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_15 = {_alignedDequeue_bits_data_T_496[7], _alignedDequeue_bits_data_T_462[7]};
  wire [3:0]    alignedDequeue_bits_data_hi_15 = {alignedDequeue_bits_data_hi_hi_15, alignedDequeue_bits_data_hi_lo_15};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_16 = {_alignedDequeue_bits_data_T_292[8], _alignedDequeue_bits_data_T_258[8]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_16 = {_alignedDequeue_bits_data_T_360[8], _alignedDequeue_bits_data_T_326[8]};
  wire [3:0]    alignedDequeue_bits_data_lo_16 = {alignedDequeue_bits_data_lo_hi_16, alignedDequeue_bits_data_lo_lo_16};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_16 = {_alignedDequeue_bits_data_T_428[8], _alignedDequeue_bits_data_T_394[8]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_16 = {_alignedDequeue_bits_data_T_496[8], _alignedDequeue_bits_data_T_462[8]};
  wire [3:0]    alignedDequeue_bits_data_hi_16 = {alignedDequeue_bits_data_hi_hi_16, alignedDequeue_bits_data_hi_lo_16};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_17 = {_alignedDequeue_bits_data_T_292[9], _alignedDequeue_bits_data_T_258[9]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_17 = {_alignedDequeue_bits_data_T_360[9], _alignedDequeue_bits_data_T_326[9]};
  wire [3:0]    alignedDequeue_bits_data_lo_17 = {alignedDequeue_bits_data_lo_hi_17, alignedDequeue_bits_data_lo_lo_17};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_17 = {_alignedDequeue_bits_data_T_428[9], _alignedDequeue_bits_data_T_394[9]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_17 = {_alignedDequeue_bits_data_T_496[9], _alignedDequeue_bits_data_T_462[9]};
  wire [3:0]    alignedDequeue_bits_data_hi_17 = {alignedDequeue_bits_data_hi_hi_17, alignedDequeue_bits_data_hi_lo_17};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_18 = {_alignedDequeue_bits_data_T_292[10], _alignedDequeue_bits_data_T_258[10]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_18 = {_alignedDequeue_bits_data_T_360[10], _alignedDequeue_bits_data_T_326[10]};
  wire [3:0]    alignedDequeue_bits_data_lo_18 = {alignedDequeue_bits_data_lo_hi_18, alignedDequeue_bits_data_lo_lo_18};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_18 = {_alignedDequeue_bits_data_T_428[10], _alignedDequeue_bits_data_T_394[10]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_18 = {_alignedDequeue_bits_data_T_496[10], _alignedDequeue_bits_data_T_462[10]};
  wire [3:0]    alignedDequeue_bits_data_hi_18 = {alignedDequeue_bits_data_hi_hi_18, alignedDequeue_bits_data_hi_lo_18};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_19 = {_alignedDequeue_bits_data_T_292[11], _alignedDequeue_bits_data_T_258[11]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_19 = {_alignedDequeue_bits_data_T_360[11], _alignedDequeue_bits_data_T_326[11]};
  wire [3:0]    alignedDequeue_bits_data_lo_19 = {alignedDequeue_bits_data_lo_hi_19, alignedDequeue_bits_data_lo_lo_19};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_19 = {_alignedDequeue_bits_data_T_428[11], _alignedDequeue_bits_data_T_394[11]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_19 = {_alignedDequeue_bits_data_T_496[11], _alignedDequeue_bits_data_T_462[11]};
  wire [3:0]    alignedDequeue_bits_data_hi_19 = {alignedDequeue_bits_data_hi_hi_19, alignedDequeue_bits_data_hi_lo_19};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_20 = {_alignedDequeue_bits_data_T_292[12], _alignedDequeue_bits_data_T_258[12]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_20 = {_alignedDequeue_bits_data_T_360[12], _alignedDequeue_bits_data_T_326[12]};
  wire [3:0]    alignedDequeue_bits_data_lo_20 = {alignedDequeue_bits_data_lo_hi_20, alignedDequeue_bits_data_lo_lo_20};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_20 = {_alignedDequeue_bits_data_T_428[12], _alignedDequeue_bits_data_T_394[12]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_20 = {_alignedDequeue_bits_data_T_496[12], _alignedDequeue_bits_data_T_462[12]};
  wire [3:0]    alignedDequeue_bits_data_hi_20 = {alignedDequeue_bits_data_hi_hi_20, alignedDequeue_bits_data_hi_lo_20};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_21 = {_alignedDequeue_bits_data_T_292[13], _alignedDequeue_bits_data_T_258[13]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_21 = {_alignedDequeue_bits_data_T_360[13], _alignedDequeue_bits_data_T_326[13]};
  wire [3:0]    alignedDequeue_bits_data_lo_21 = {alignedDequeue_bits_data_lo_hi_21, alignedDequeue_bits_data_lo_lo_21};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_21 = {_alignedDequeue_bits_data_T_428[13], _alignedDequeue_bits_data_T_394[13]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_21 = {_alignedDequeue_bits_data_T_496[13], _alignedDequeue_bits_data_T_462[13]};
  wire [3:0]    alignedDequeue_bits_data_hi_21 = {alignedDequeue_bits_data_hi_hi_21, alignedDequeue_bits_data_hi_lo_21};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_22 = {_alignedDequeue_bits_data_T_292[14], _alignedDequeue_bits_data_T_258[14]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_22 = {_alignedDequeue_bits_data_T_360[14], _alignedDequeue_bits_data_T_326[14]};
  wire [3:0]    alignedDequeue_bits_data_lo_22 = {alignedDequeue_bits_data_lo_hi_22, alignedDequeue_bits_data_lo_lo_22};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_22 = {_alignedDequeue_bits_data_T_428[14], _alignedDequeue_bits_data_T_394[14]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_22 = {_alignedDequeue_bits_data_T_496[14], _alignedDequeue_bits_data_T_462[14]};
  wire [3:0]    alignedDequeue_bits_data_hi_22 = {alignedDequeue_bits_data_hi_hi_22, alignedDequeue_bits_data_hi_lo_22};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_23 = {_alignedDequeue_bits_data_T_292[15], _alignedDequeue_bits_data_T_258[15]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_23 = {_alignedDequeue_bits_data_T_360[15], _alignedDequeue_bits_data_T_326[15]};
  wire [3:0]    alignedDequeue_bits_data_lo_23 = {alignedDequeue_bits_data_lo_hi_23, alignedDequeue_bits_data_lo_lo_23};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_23 = {_alignedDequeue_bits_data_T_428[15], _alignedDequeue_bits_data_T_394[15]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_23 = {_alignedDequeue_bits_data_T_496[15], _alignedDequeue_bits_data_T_462[15]};
  wire [3:0]    alignedDequeue_bits_data_hi_23 = {alignedDequeue_bits_data_hi_hi_23, alignedDequeue_bits_data_hi_lo_23};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_24 = {_alignedDequeue_bits_data_T_292[16], _alignedDequeue_bits_data_T_258[16]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_24 = {_alignedDequeue_bits_data_T_360[16], _alignedDequeue_bits_data_T_326[16]};
  wire [3:0]    alignedDequeue_bits_data_lo_24 = {alignedDequeue_bits_data_lo_hi_24, alignedDequeue_bits_data_lo_lo_24};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_24 = {_alignedDequeue_bits_data_T_428[16], _alignedDequeue_bits_data_T_394[16]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_24 = {_alignedDequeue_bits_data_T_496[16], _alignedDequeue_bits_data_T_462[16]};
  wire [3:0]    alignedDequeue_bits_data_hi_24 = {alignedDequeue_bits_data_hi_hi_24, alignedDequeue_bits_data_hi_lo_24};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_25 = {_alignedDequeue_bits_data_T_292[17], _alignedDequeue_bits_data_T_258[17]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_25 = {_alignedDequeue_bits_data_T_360[17], _alignedDequeue_bits_data_T_326[17]};
  wire [3:0]    alignedDequeue_bits_data_lo_25 = {alignedDequeue_bits_data_lo_hi_25, alignedDequeue_bits_data_lo_lo_25};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_25 = {_alignedDequeue_bits_data_T_428[17], _alignedDequeue_bits_data_T_394[17]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_25 = {_alignedDequeue_bits_data_T_496[17], _alignedDequeue_bits_data_T_462[17]};
  wire [3:0]    alignedDequeue_bits_data_hi_25 = {alignedDequeue_bits_data_hi_hi_25, alignedDequeue_bits_data_hi_lo_25};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_26 = {_alignedDequeue_bits_data_T_292[18], _alignedDequeue_bits_data_T_258[18]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_26 = {_alignedDequeue_bits_data_T_360[18], _alignedDequeue_bits_data_T_326[18]};
  wire [3:0]    alignedDequeue_bits_data_lo_26 = {alignedDequeue_bits_data_lo_hi_26, alignedDequeue_bits_data_lo_lo_26};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_26 = {_alignedDequeue_bits_data_T_428[18], _alignedDequeue_bits_data_T_394[18]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_26 = {_alignedDequeue_bits_data_T_496[18], _alignedDequeue_bits_data_T_462[18]};
  wire [3:0]    alignedDequeue_bits_data_hi_26 = {alignedDequeue_bits_data_hi_hi_26, alignedDequeue_bits_data_hi_lo_26};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_27 = {_alignedDequeue_bits_data_T_292[19], _alignedDequeue_bits_data_T_258[19]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_27 = {_alignedDequeue_bits_data_T_360[19], _alignedDequeue_bits_data_T_326[19]};
  wire [3:0]    alignedDequeue_bits_data_lo_27 = {alignedDequeue_bits_data_lo_hi_27, alignedDequeue_bits_data_lo_lo_27};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_27 = {_alignedDequeue_bits_data_T_428[19], _alignedDequeue_bits_data_T_394[19]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_27 = {_alignedDequeue_bits_data_T_496[19], _alignedDequeue_bits_data_T_462[19]};
  wire [3:0]    alignedDequeue_bits_data_hi_27 = {alignedDequeue_bits_data_hi_hi_27, alignedDequeue_bits_data_hi_lo_27};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_28 = {_alignedDequeue_bits_data_T_292[20], _alignedDequeue_bits_data_T_258[20]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_28 = {_alignedDequeue_bits_data_T_360[20], _alignedDequeue_bits_data_T_326[20]};
  wire [3:0]    alignedDequeue_bits_data_lo_28 = {alignedDequeue_bits_data_lo_hi_28, alignedDequeue_bits_data_lo_lo_28};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_28 = {_alignedDequeue_bits_data_T_428[20], _alignedDequeue_bits_data_T_394[20]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_28 = {_alignedDequeue_bits_data_T_496[20], _alignedDequeue_bits_data_T_462[20]};
  wire [3:0]    alignedDequeue_bits_data_hi_28 = {alignedDequeue_bits_data_hi_hi_28, alignedDequeue_bits_data_hi_lo_28};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_29 = {_alignedDequeue_bits_data_T_292[21], _alignedDequeue_bits_data_T_258[21]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_29 = {_alignedDequeue_bits_data_T_360[21], _alignedDequeue_bits_data_T_326[21]};
  wire [3:0]    alignedDequeue_bits_data_lo_29 = {alignedDequeue_bits_data_lo_hi_29, alignedDequeue_bits_data_lo_lo_29};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_29 = {_alignedDequeue_bits_data_T_428[21], _alignedDequeue_bits_data_T_394[21]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_29 = {_alignedDequeue_bits_data_T_496[21], _alignedDequeue_bits_data_T_462[21]};
  wire [3:0]    alignedDequeue_bits_data_hi_29 = {alignedDequeue_bits_data_hi_hi_29, alignedDequeue_bits_data_hi_lo_29};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_30 = {_alignedDequeue_bits_data_T_292[22], _alignedDequeue_bits_data_T_258[22]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_30 = {_alignedDequeue_bits_data_T_360[22], _alignedDequeue_bits_data_T_326[22]};
  wire [3:0]    alignedDequeue_bits_data_lo_30 = {alignedDequeue_bits_data_lo_hi_30, alignedDequeue_bits_data_lo_lo_30};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_30 = {_alignedDequeue_bits_data_T_428[22], _alignedDequeue_bits_data_T_394[22]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_30 = {_alignedDequeue_bits_data_T_496[22], _alignedDequeue_bits_data_T_462[22]};
  wire [3:0]    alignedDequeue_bits_data_hi_30 = {alignedDequeue_bits_data_hi_hi_30, alignedDequeue_bits_data_hi_lo_30};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_31 = {_alignedDequeue_bits_data_T_292[23], _alignedDequeue_bits_data_T_258[23]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_31 = {_alignedDequeue_bits_data_T_360[23], _alignedDequeue_bits_data_T_326[23]};
  wire [3:0]    alignedDequeue_bits_data_lo_31 = {alignedDequeue_bits_data_lo_hi_31, alignedDequeue_bits_data_lo_lo_31};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_31 = {_alignedDequeue_bits_data_T_428[23], _alignedDequeue_bits_data_T_394[23]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_31 = {_alignedDequeue_bits_data_T_496[23], _alignedDequeue_bits_data_T_462[23]};
  wire [3:0]    alignedDequeue_bits_data_hi_31 = {alignedDequeue_bits_data_hi_hi_31, alignedDequeue_bits_data_hi_lo_31};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_32 = {_alignedDequeue_bits_data_T_292[24], _alignedDequeue_bits_data_T_258[24]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_32 = {_alignedDequeue_bits_data_T_360[24], _alignedDequeue_bits_data_T_326[24]};
  wire [3:0]    alignedDequeue_bits_data_lo_32 = {alignedDequeue_bits_data_lo_hi_32, alignedDequeue_bits_data_lo_lo_32};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_32 = {_alignedDequeue_bits_data_T_428[24], _alignedDequeue_bits_data_T_394[24]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_32 = {_alignedDequeue_bits_data_T_496[24], _alignedDequeue_bits_data_T_462[24]};
  wire [3:0]    alignedDequeue_bits_data_hi_32 = {alignedDequeue_bits_data_hi_hi_32, alignedDequeue_bits_data_hi_lo_32};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_33 = {_alignedDequeue_bits_data_T_292[25], _alignedDequeue_bits_data_T_258[25]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_33 = {_alignedDequeue_bits_data_T_360[25], _alignedDequeue_bits_data_T_326[25]};
  wire [3:0]    alignedDequeue_bits_data_lo_33 = {alignedDequeue_bits_data_lo_hi_33, alignedDequeue_bits_data_lo_lo_33};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_33 = {_alignedDequeue_bits_data_T_428[25], _alignedDequeue_bits_data_T_394[25]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_33 = {_alignedDequeue_bits_data_T_496[25], _alignedDequeue_bits_data_T_462[25]};
  wire [3:0]    alignedDequeue_bits_data_hi_33 = {alignedDequeue_bits_data_hi_hi_33, alignedDequeue_bits_data_hi_lo_33};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_34 = {_alignedDequeue_bits_data_T_292[26], _alignedDequeue_bits_data_T_258[26]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_34 = {_alignedDequeue_bits_data_T_360[26], _alignedDequeue_bits_data_T_326[26]};
  wire [3:0]    alignedDequeue_bits_data_lo_34 = {alignedDequeue_bits_data_lo_hi_34, alignedDequeue_bits_data_lo_lo_34};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_34 = {_alignedDequeue_bits_data_T_428[26], _alignedDequeue_bits_data_T_394[26]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_34 = {_alignedDequeue_bits_data_T_496[26], _alignedDequeue_bits_data_T_462[26]};
  wire [3:0]    alignedDequeue_bits_data_hi_34 = {alignedDequeue_bits_data_hi_hi_34, alignedDequeue_bits_data_hi_lo_34};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_35 = {_alignedDequeue_bits_data_T_292[27], _alignedDequeue_bits_data_T_258[27]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_35 = {_alignedDequeue_bits_data_T_360[27], _alignedDequeue_bits_data_T_326[27]};
  wire [3:0]    alignedDequeue_bits_data_lo_35 = {alignedDequeue_bits_data_lo_hi_35, alignedDequeue_bits_data_lo_lo_35};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_35 = {_alignedDequeue_bits_data_T_428[27], _alignedDequeue_bits_data_T_394[27]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_35 = {_alignedDequeue_bits_data_T_496[27], _alignedDequeue_bits_data_T_462[27]};
  wire [3:0]    alignedDequeue_bits_data_hi_35 = {alignedDequeue_bits_data_hi_hi_35, alignedDequeue_bits_data_hi_lo_35};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_36 = {_alignedDequeue_bits_data_T_292[28], _alignedDequeue_bits_data_T_258[28]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_36 = {_alignedDequeue_bits_data_T_360[28], _alignedDequeue_bits_data_T_326[28]};
  wire [3:0]    alignedDequeue_bits_data_lo_36 = {alignedDequeue_bits_data_lo_hi_36, alignedDequeue_bits_data_lo_lo_36};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_36 = {_alignedDequeue_bits_data_T_428[28], _alignedDequeue_bits_data_T_394[28]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_36 = {_alignedDequeue_bits_data_T_496[28], _alignedDequeue_bits_data_T_462[28]};
  wire [3:0]    alignedDequeue_bits_data_hi_36 = {alignedDequeue_bits_data_hi_hi_36, alignedDequeue_bits_data_hi_lo_36};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_37 = {_alignedDequeue_bits_data_T_292[29], _alignedDequeue_bits_data_T_258[29]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_37 = {_alignedDequeue_bits_data_T_360[29], _alignedDequeue_bits_data_T_326[29]};
  wire [3:0]    alignedDequeue_bits_data_lo_37 = {alignedDequeue_bits_data_lo_hi_37, alignedDequeue_bits_data_lo_lo_37};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_37 = {_alignedDequeue_bits_data_T_428[29], _alignedDequeue_bits_data_T_394[29]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_37 = {_alignedDequeue_bits_data_T_496[29], _alignedDequeue_bits_data_T_462[29]};
  wire [3:0]    alignedDequeue_bits_data_hi_37 = {alignedDequeue_bits_data_hi_hi_37, alignedDequeue_bits_data_hi_lo_37};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_38 = {_alignedDequeue_bits_data_T_292[30], _alignedDequeue_bits_data_T_258[30]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_38 = {_alignedDequeue_bits_data_T_360[30], _alignedDequeue_bits_data_T_326[30]};
  wire [3:0]    alignedDequeue_bits_data_lo_38 = {alignedDequeue_bits_data_lo_hi_38, alignedDequeue_bits_data_lo_lo_38};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_38 = {_alignedDequeue_bits_data_T_428[30], _alignedDequeue_bits_data_T_394[30]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_38 = {_alignedDequeue_bits_data_T_496[30], _alignedDequeue_bits_data_T_462[30]};
  wire [3:0]    alignedDequeue_bits_data_hi_38 = {alignedDequeue_bits_data_hi_hi_38, alignedDequeue_bits_data_hi_lo_38};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_39 = {_alignedDequeue_bits_data_T_292[31], _alignedDequeue_bits_data_T_258[31]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_39 = {_alignedDequeue_bits_data_T_360[31], _alignedDequeue_bits_data_T_326[31]};
  wire [3:0]    alignedDequeue_bits_data_lo_39 = {alignedDequeue_bits_data_lo_hi_39, alignedDequeue_bits_data_lo_lo_39};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_39 = {_alignedDequeue_bits_data_T_428[31], _alignedDequeue_bits_data_T_394[31]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_39 = {_alignedDequeue_bits_data_T_496[31], _alignedDequeue_bits_data_T_462[31]};
  wire [3:0]    alignedDequeue_bits_data_hi_39 = {alignedDequeue_bits_data_hi_hi_39, alignedDequeue_bits_data_hi_lo_39};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_9, alignedDequeue_bits_data_lo_9, alignedDequeue_bits_data_hi_8, alignedDequeue_bits_data_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_11, alignedDequeue_bits_data_lo_11, alignedDequeue_bits_data_hi_10, alignedDequeue_bits_data_lo_10};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_lo_8 = {alignedDequeue_bits_data_lo_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_13, alignedDequeue_bits_data_lo_13, alignedDequeue_bits_data_hi_12, alignedDequeue_bits_data_lo_12};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_15, alignedDequeue_bits_data_lo_15, alignedDequeue_bits_data_hi_14, alignedDequeue_bits_data_lo_14};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_hi_8 = {alignedDequeue_bits_data_lo_lo_hi_hi_8, alignedDequeue_bits_data_lo_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_lo_40 = {alignedDequeue_bits_data_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_17, alignedDequeue_bits_data_lo_17, alignedDequeue_bits_data_hi_16, alignedDequeue_bits_data_lo_16};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_19, alignedDequeue_bits_data_lo_19, alignedDequeue_bits_data_hi_18, alignedDequeue_bits_data_lo_18};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_lo_8 = {alignedDequeue_bits_data_lo_hi_lo_hi_8, alignedDequeue_bits_data_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_21, alignedDequeue_bits_data_lo_21, alignedDequeue_bits_data_hi_20, alignedDequeue_bits_data_lo_20};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_23, alignedDequeue_bits_data_lo_23, alignedDequeue_bits_data_hi_22, alignedDequeue_bits_data_lo_22};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_hi_8 = {alignedDequeue_bits_data_lo_hi_hi_hi_8, alignedDequeue_bits_data_lo_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_hi_40 = {alignedDequeue_bits_data_lo_hi_hi_8, alignedDequeue_bits_data_lo_hi_lo_8};
  assign alignedDequeue_bits_data_lo_40 = {alignedDequeue_bits_data_lo_hi_40, alignedDequeue_bits_data_lo_lo_40};
  wire [127:0]  alignedDequeue_bits_data = alignedDequeue_bits_data_lo_40;
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_25, alignedDequeue_bits_data_lo_25, alignedDequeue_bits_data_hi_24, alignedDequeue_bits_data_lo_24};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_27, alignedDequeue_bits_data_lo_27, alignedDequeue_bits_data_hi_26, alignedDequeue_bits_data_lo_26};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_lo_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_29, alignedDequeue_bits_data_lo_29, alignedDequeue_bits_data_hi_28, alignedDequeue_bits_data_lo_28};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_31, alignedDequeue_bits_data_lo_31, alignedDequeue_bits_data_hi_30, alignedDequeue_bits_data_lo_30};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_lo_hi_hi_8, alignedDequeue_bits_data_hi_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_lo_40 = {alignedDequeue_bits_data_hi_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_33, alignedDequeue_bits_data_lo_33, alignedDequeue_bits_data_hi_32, alignedDequeue_bits_data_lo_32};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_35, alignedDequeue_bits_data_lo_35, alignedDequeue_bits_data_hi_34, alignedDequeue_bits_data_lo_34};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_hi_lo_hi_8, alignedDequeue_bits_data_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_37, alignedDequeue_bits_data_lo_37, alignedDequeue_bits_data_hi_36, alignedDequeue_bits_data_lo_36};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_39, alignedDequeue_bits_data_lo_39, alignedDequeue_bits_data_hi_38, alignedDequeue_bits_data_lo_38};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_hi_40 = {alignedDequeue_bits_data_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_hi_40 = {alignedDequeue_bits_data_hi_hi_40, alignedDequeue_bits_data_hi_lo_40};
  reg           bufferFull;
  wire          bufferTailFire;
  wire          bufferDequeueValid = bufferFull | bufferTailFire;
  wire          writeStageReady;
  wire          bufferDequeueReady;
  wire          bufferDequeueFire = bufferDequeueReady & bufferDequeueValid;
  assign alignedDequeue_ready = ~bufferFull;
  wire [7:0]    bufferEnqueueSelect = _bufferTailFire_T ? 8'h1 << cacheLineIndexInBuffer : 8'h0;
  wire [127:0]  dataBufferUpdate_0 = bufferEnqueueSelect[0] ? alignedDequeue_bits_data : dataBuffer_0;
  wire [127:0]  dataBufferUpdate_1 = bufferEnqueueSelect[1] ? alignedDequeue_bits_data : dataBuffer_1;
  wire [127:0]  dataBufferUpdate_2 = bufferEnqueueSelect[2] ? alignedDequeue_bits_data : dataBuffer_2;
  wire [127:0]  dataBufferUpdate_3 = bufferEnqueueSelect[3] ? alignedDequeue_bits_data : dataBuffer_3;
  wire [127:0]  dataBufferUpdate_4 = bufferEnqueueSelect[4] ? alignedDequeue_bits_data : dataBuffer_4;
  wire [127:0]  dataBufferUpdate_5 = bufferEnqueueSelect[5] ? alignedDequeue_bits_data : dataBuffer_5;
  wire [127:0]  dataBufferUpdate_6 = bufferEnqueueSelect[6] ? alignedDequeue_bits_data : dataBuffer_6;
  wire [127:0]  dataBufferUpdate_7 = bufferEnqueueSelect[7] ? alignedDequeue_bits_data : dataBuffer_7;
  wire [127:0]  dataSelect_0 = bufferFull ? dataBuffer_0 : dataBufferUpdate_0;
  wire [127:0]  dataSelect_1 = bufferFull ? dataBuffer_1 : dataBufferUpdate_1;
  wire [127:0]  dataSelect_2 = bufferFull ? dataBuffer_2 : dataBufferUpdate_2;
  wire [127:0]  dataSelect_3 = bufferFull ? dataBuffer_3 : dataBufferUpdate_3;
  wire [127:0]  dataSelect_4 = bufferFull ? dataBuffer_4 : dataBufferUpdate_4;
  wire [127:0]  dataSelect_5 = bufferFull ? dataBuffer_5 : dataBufferUpdate_5;
  wire [127:0]  dataSelect_6 = bufferFull ? dataBuffer_6 : dataBufferUpdate_6;
  wire [127:0]  dataSelect_7 = bufferFull ? dataBuffer_7 : dataBufferUpdate_7;
  wire          lastCacheLineForThisGroup = cacheLineIndexInBuffer == lsuRequestReg_instructionInformation_nf;
  wire          lastCacheLineForInst = {7'h0, alignedDequeue_bits_index} == lastWriteVrfIndexReg;
  assign bufferTailFire = _bufferTailFire_T & (lastCacheLineForThisGroup | lastCacheLineForInst);
  reg           waitForFirstDataGroup;
  wire          lastPtr = accessPtr == 3'h0;
  assign writeStageReady = lastPtr & accessStateCheck;
  assign bufferDequeueReady = writeStageReady;
  wire          _maskSelect_valid_output = bufferDequeueFire & isLastDataGroup;
  wire [255:0]  _GEN_3 = {dataSelect_1, dataSelect_0};
  wire [255:0]  dataGroup_lo_lo;
  assign dataGroup_lo_lo = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1;
  assign dataGroup_lo_lo_1 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_2;
  assign dataGroup_lo_lo_2 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_3;
  assign dataGroup_lo_lo_3 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_4;
  assign dataGroup_lo_lo_4 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_5;
  assign dataGroup_lo_lo_5 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_6;
  assign dataGroup_lo_lo_6 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_7;
  assign dataGroup_lo_lo_7 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_8;
  assign dataGroup_lo_lo_8 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_9;
  assign dataGroup_lo_lo_9 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_10;
  assign dataGroup_lo_lo_10 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_11;
  assign dataGroup_lo_lo_11 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_12;
  assign dataGroup_lo_lo_12 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_13;
  assign dataGroup_lo_lo_13 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_14;
  assign dataGroup_lo_lo_14 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_15;
  assign dataGroup_lo_lo_15 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_16;
  assign dataGroup_lo_lo_16 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_17;
  assign dataGroup_lo_lo_17 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_18;
  assign dataGroup_lo_lo_18 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_19;
  assign dataGroup_lo_lo_19 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_20;
  assign dataGroup_lo_lo_20 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_21;
  assign dataGroup_lo_lo_21 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_22;
  assign dataGroup_lo_lo_22 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_23;
  assign dataGroup_lo_lo_23 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_24;
  assign dataGroup_lo_lo_24 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_25;
  assign dataGroup_lo_lo_25 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_26;
  assign dataGroup_lo_lo_26 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_27;
  assign dataGroup_lo_lo_27 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_28;
  assign dataGroup_lo_lo_28 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_29;
  assign dataGroup_lo_lo_29 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_30;
  assign dataGroup_lo_lo_30 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_31;
  assign dataGroup_lo_lo_31 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_32;
  assign dataGroup_lo_lo_32 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_33;
  assign dataGroup_lo_lo_33 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_34;
  assign dataGroup_lo_lo_34 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_35;
  assign dataGroup_lo_lo_35 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_36;
  assign dataGroup_lo_lo_36 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_37;
  assign dataGroup_lo_lo_37 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_38;
  assign dataGroup_lo_lo_38 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_39;
  assign dataGroup_lo_lo_39 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_40;
  assign dataGroup_lo_lo_40 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_41;
  assign dataGroup_lo_lo_41 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_42;
  assign dataGroup_lo_lo_42 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_43;
  assign dataGroup_lo_lo_43 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_44;
  assign dataGroup_lo_lo_44 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_45;
  assign dataGroup_lo_lo_45 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_46;
  assign dataGroup_lo_lo_46 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_47;
  assign dataGroup_lo_lo_47 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_48;
  assign dataGroup_lo_lo_48 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_49;
  assign dataGroup_lo_lo_49 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_50;
  assign dataGroup_lo_lo_50 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_51;
  assign dataGroup_lo_lo_51 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_52;
  assign dataGroup_lo_lo_52 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_53;
  assign dataGroup_lo_lo_53 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_54;
  assign dataGroup_lo_lo_54 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_55;
  assign dataGroup_lo_lo_55 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_56;
  assign dataGroup_lo_lo_56 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_57;
  assign dataGroup_lo_lo_57 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_58;
  assign dataGroup_lo_lo_58 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_59;
  assign dataGroup_lo_lo_59 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_60;
  assign dataGroup_lo_lo_60 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_61;
  assign dataGroup_lo_lo_61 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_62;
  assign dataGroup_lo_lo_62 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_63;
  assign dataGroup_lo_lo_63 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_64;
  assign dataGroup_lo_lo_64 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_65;
  assign dataGroup_lo_lo_65 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_66;
  assign dataGroup_lo_lo_66 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_67;
  assign dataGroup_lo_lo_67 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_68;
  assign dataGroup_lo_lo_68 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_69;
  assign dataGroup_lo_lo_69 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_70;
  assign dataGroup_lo_lo_70 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_71;
  assign dataGroup_lo_lo_71 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_72;
  assign dataGroup_lo_lo_72 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_73;
  assign dataGroup_lo_lo_73 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_74;
  assign dataGroup_lo_lo_74 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_75;
  assign dataGroup_lo_lo_75 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_76;
  assign dataGroup_lo_lo_76 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_77;
  assign dataGroup_lo_lo_77 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_78;
  assign dataGroup_lo_lo_78 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_79;
  assign dataGroup_lo_lo_79 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_80;
  assign dataGroup_lo_lo_80 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_81;
  assign dataGroup_lo_lo_81 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_82;
  assign dataGroup_lo_lo_82 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_83;
  assign dataGroup_lo_lo_83 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_84;
  assign dataGroup_lo_lo_84 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_85;
  assign dataGroup_lo_lo_85 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_86;
  assign dataGroup_lo_lo_86 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_87;
  assign dataGroup_lo_lo_87 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_88;
  assign dataGroup_lo_lo_88 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_89;
  assign dataGroup_lo_lo_89 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_90;
  assign dataGroup_lo_lo_90 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_91;
  assign dataGroup_lo_lo_91 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_92;
  assign dataGroup_lo_lo_92 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_93;
  assign dataGroup_lo_lo_93 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_94;
  assign dataGroup_lo_lo_94 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_95;
  assign dataGroup_lo_lo_95 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_96;
  assign dataGroup_lo_lo_96 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_97;
  assign dataGroup_lo_lo_97 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_98;
  assign dataGroup_lo_lo_98 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_99;
  assign dataGroup_lo_lo_99 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_100;
  assign dataGroup_lo_lo_100 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_101;
  assign dataGroup_lo_lo_101 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_102;
  assign dataGroup_lo_lo_102 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_103;
  assign dataGroup_lo_lo_103 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_104;
  assign dataGroup_lo_lo_104 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_105;
  assign dataGroup_lo_lo_105 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_106;
  assign dataGroup_lo_lo_106 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_107;
  assign dataGroup_lo_lo_107 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_108;
  assign dataGroup_lo_lo_108 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_109;
  assign dataGroup_lo_lo_109 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_110;
  assign dataGroup_lo_lo_110 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_111;
  assign dataGroup_lo_lo_111 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_112;
  assign dataGroup_lo_lo_112 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_113;
  assign dataGroup_lo_lo_113 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_114;
  assign dataGroup_lo_lo_114 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_115;
  assign dataGroup_lo_lo_115 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_116;
  assign dataGroup_lo_lo_116 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_117;
  assign dataGroup_lo_lo_117 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_118;
  assign dataGroup_lo_lo_118 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_119;
  assign dataGroup_lo_lo_119 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_120;
  assign dataGroup_lo_lo_120 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_121;
  assign dataGroup_lo_lo_121 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_122;
  assign dataGroup_lo_lo_122 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_123;
  assign dataGroup_lo_lo_123 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_124;
  assign dataGroup_lo_lo_124 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_125;
  assign dataGroup_lo_lo_125 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_126;
  assign dataGroup_lo_lo_126 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_127;
  assign dataGroup_lo_lo_127 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_128;
  assign dataGroup_lo_lo_128 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_129;
  assign dataGroup_lo_lo_129 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_130;
  assign dataGroup_lo_lo_130 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_131;
  assign dataGroup_lo_lo_131 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_132;
  assign dataGroup_lo_lo_132 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_133;
  assign dataGroup_lo_lo_133 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_134;
  assign dataGroup_lo_lo_134 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_135;
  assign dataGroup_lo_lo_135 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_136;
  assign dataGroup_lo_lo_136 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_137;
  assign dataGroup_lo_lo_137 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_138;
  assign dataGroup_lo_lo_138 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_139;
  assign dataGroup_lo_lo_139 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_140;
  assign dataGroup_lo_lo_140 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_141;
  assign dataGroup_lo_lo_141 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_142;
  assign dataGroup_lo_lo_142 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_143;
  assign dataGroup_lo_lo_143 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_144;
  assign dataGroup_lo_lo_144 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_145;
  assign dataGroup_lo_lo_145 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_146;
  assign dataGroup_lo_lo_146 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_147;
  assign dataGroup_lo_lo_147 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_148;
  assign dataGroup_lo_lo_148 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_149;
  assign dataGroup_lo_lo_149 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_150;
  assign dataGroup_lo_lo_150 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_151;
  assign dataGroup_lo_lo_151 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_152;
  assign dataGroup_lo_lo_152 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_153;
  assign dataGroup_lo_lo_153 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_154;
  assign dataGroup_lo_lo_154 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_155;
  assign dataGroup_lo_lo_155 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_156;
  assign dataGroup_lo_lo_156 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_157;
  assign dataGroup_lo_lo_157 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_158;
  assign dataGroup_lo_lo_158 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_159;
  assign dataGroup_lo_lo_159 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_160;
  assign dataGroup_lo_lo_160 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_161;
  assign dataGroup_lo_lo_161 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_162;
  assign dataGroup_lo_lo_162 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_163;
  assign dataGroup_lo_lo_163 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_164;
  assign dataGroup_lo_lo_164 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_165;
  assign dataGroup_lo_lo_165 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_166;
  assign dataGroup_lo_lo_166 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_167;
  assign dataGroup_lo_lo_167 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_168;
  assign dataGroup_lo_lo_168 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_169;
  assign dataGroup_lo_lo_169 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_170;
  assign dataGroup_lo_lo_170 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_171;
  assign dataGroup_lo_lo_171 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_172;
  assign dataGroup_lo_lo_172 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_173;
  assign dataGroup_lo_lo_173 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_174;
  assign dataGroup_lo_lo_174 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_175;
  assign dataGroup_lo_lo_175 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_176;
  assign dataGroup_lo_lo_176 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_177;
  assign dataGroup_lo_lo_177 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_178;
  assign dataGroup_lo_lo_178 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_179;
  assign dataGroup_lo_lo_179 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_180;
  assign dataGroup_lo_lo_180 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_181;
  assign dataGroup_lo_lo_181 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_182;
  assign dataGroup_lo_lo_182 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_183;
  assign dataGroup_lo_lo_183 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_184;
  assign dataGroup_lo_lo_184 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_185;
  assign dataGroup_lo_lo_185 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_186;
  assign dataGroup_lo_lo_186 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_187;
  assign dataGroup_lo_lo_187 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_188;
  assign dataGroup_lo_lo_188 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_189;
  assign dataGroup_lo_lo_189 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_190;
  assign dataGroup_lo_lo_190 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_191;
  assign dataGroup_lo_lo_191 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_192;
  assign dataGroup_lo_lo_192 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_193;
  assign dataGroup_lo_lo_193 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_194;
  assign dataGroup_lo_lo_194 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_195;
  assign dataGroup_lo_lo_195 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_196;
  assign dataGroup_lo_lo_196 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_197;
  assign dataGroup_lo_lo_197 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_198;
  assign dataGroup_lo_lo_198 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_199;
  assign dataGroup_lo_lo_199 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_200;
  assign dataGroup_lo_lo_200 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_201;
  assign dataGroup_lo_lo_201 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_202;
  assign dataGroup_lo_lo_202 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_203;
  assign dataGroup_lo_lo_203 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_204;
  assign dataGroup_lo_lo_204 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_205;
  assign dataGroup_lo_lo_205 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_206;
  assign dataGroup_lo_lo_206 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_207;
  assign dataGroup_lo_lo_207 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_208;
  assign dataGroup_lo_lo_208 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_209;
  assign dataGroup_lo_lo_209 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_210;
  assign dataGroup_lo_lo_210 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_211;
  assign dataGroup_lo_lo_211 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_212;
  assign dataGroup_lo_lo_212 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_213;
  assign dataGroup_lo_lo_213 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_214;
  assign dataGroup_lo_lo_214 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_215;
  assign dataGroup_lo_lo_215 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_216;
  assign dataGroup_lo_lo_216 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_217;
  assign dataGroup_lo_lo_217 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_218;
  assign dataGroup_lo_lo_218 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_219;
  assign dataGroup_lo_lo_219 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_220;
  assign dataGroup_lo_lo_220 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_221;
  assign dataGroup_lo_lo_221 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_222;
  assign dataGroup_lo_lo_222 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_223;
  assign dataGroup_lo_lo_223 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_224;
  assign dataGroup_lo_lo_224 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_225;
  assign dataGroup_lo_lo_225 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_226;
  assign dataGroup_lo_lo_226 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_227;
  assign dataGroup_lo_lo_227 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_228;
  assign dataGroup_lo_lo_228 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_229;
  assign dataGroup_lo_lo_229 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_230;
  assign dataGroup_lo_lo_230 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_231;
  assign dataGroup_lo_lo_231 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_232;
  assign dataGroup_lo_lo_232 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_233;
  assign dataGroup_lo_lo_233 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_234;
  assign dataGroup_lo_lo_234 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_235;
  assign dataGroup_lo_lo_235 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_236;
  assign dataGroup_lo_lo_236 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_237;
  assign dataGroup_lo_lo_237 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_238;
  assign dataGroup_lo_lo_238 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_239;
  assign dataGroup_lo_lo_239 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_240;
  assign dataGroup_lo_lo_240 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_241;
  assign dataGroup_lo_lo_241 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_242;
  assign dataGroup_lo_lo_242 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_243;
  assign dataGroup_lo_lo_243 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_244;
  assign dataGroup_lo_lo_244 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_245;
  assign dataGroup_lo_lo_245 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_246;
  assign dataGroup_lo_lo_246 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_247;
  assign dataGroup_lo_lo_247 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_248;
  assign dataGroup_lo_lo_248 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_249;
  assign dataGroup_lo_lo_249 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_250;
  assign dataGroup_lo_lo_250 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_251;
  assign dataGroup_lo_lo_251 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_252;
  assign dataGroup_lo_lo_252 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_253;
  assign dataGroup_lo_lo_253 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_254;
  assign dataGroup_lo_lo_254 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_255;
  assign dataGroup_lo_lo_255 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_256;
  assign dataGroup_lo_lo_256 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_257;
  assign dataGroup_lo_lo_257 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_258;
  assign dataGroup_lo_lo_258 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_259;
  assign dataGroup_lo_lo_259 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_260;
  assign dataGroup_lo_lo_260 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_261;
  assign dataGroup_lo_lo_261 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_262;
  assign dataGroup_lo_lo_262 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_263;
  assign dataGroup_lo_lo_263 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_264;
  assign dataGroup_lo_lo_264 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_265;
  assign dataGroup_lo_lo_265 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_266;
  assign dataGroup_lo_lo_266 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_267;
  assign dataGroup_lo_lo_267 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_268;
  assign dataGroup_lo_lo_268 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_269;
  assign dataGroup_lo_lo_269 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_270;
  assign dataGroup_lo_lo_270 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_271;
  assign dataGroup_lo_lo_271 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_272;
  assign dataGroup_lo_lo_272 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_273;
  assign dataGroup_lo_lo_273 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_274;
  assign dataGroup_lo_lo_274 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_275;
  assign dataGroup_lo_lo_275 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_276;
  assign dataGroup_lo_lo_276 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_277;
  assign dataGroup_lo_lo_277 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_278;
  assign dataGroup_lo_lo_278 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_279;
  assign dataGroup_lo_lo_279 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_280;
  assign dataGroup_lo_lo_280 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_281;
  assign dataGroup_lo_lo_281 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_282;
  assign dataGroup_lo_lo_282 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_283;
  assign dataGroup_lo_lo_283 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_284;
  assign dataGroup_lo_lo_284 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_285;
  assign dataGroup_lo_lo_285 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_286;
  assign dataGroup_lo_lo_286 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_287;
  assign dataGroup_lo_lo_287 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_288;
  assign dataGroup_lo_lo_288 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_289;
  assign dataGroup_lo_lo_289 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_290;
  assign dataGroup_lo_lo_290 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_291;
  assign dataGroup_lo_lo_291 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_292;
  assign dataGroup_lo_lo_292 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_293;
  assign dataGroup_lo_lo_293 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_294;
  assign dataGroup_lo_lo_294 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_295;
  assign dataGroup_lo_lo_295 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_296;
  assign dataGroup_lo_lo_296 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_297;
  assign dataGroup_lo_lo_297 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_298;
  assign dataGroup_lo_lo_298 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_299;
  assign dataGroup_lo_lo_299 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_300;
  assign dataGroup_lo_lo_300 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_301;
  assign dataGroup_lo_lo_301 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_302;
  assign dataGroup_lo_lo_302 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_303;
  assign dataGroup_lo_lo_303 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_304;
  assign dataGroup_lo_lo_304 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_305;
  assign dataGroup_lo_lo_305 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_306;
  assign dataGroup_lo_lo_306 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_307;
  assign dataGroup_lo_lo_307 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_308;
  assign dataGroup_lo_lo_308 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_309;
  assign dataGroup_lo_lo_309 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_310;
  assign dataGroup_lo_lo_310 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_311;
  assign dataGroup_lo_lo_311 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_312;
  assign dataGroup_lo_lo_312 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_313;
  assign dataGroup_lo_lo_313 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_314;
  assign dataGroup_lo_lo_314 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_315;
  assign dataGroup_lo_lo_315 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_316;
  assign dataGroup_lo_lo_316 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_317;
  assign dataGroup_lo_lo_317 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_318;
  assign dataGroup_lo_lo_318 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_319;
  assign dataGroup_lo_lo_319 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_320;
  assign dataGroup_lo_lo_320 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_321;
  assign dataGroup_lo_lo_321 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_322;
  assign dataGroup_lo_lo_322 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_323;
  assign dataGroup_lo_lo_323 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_324;
  assign dataGroup_lo_lo_324 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_325;
  assign dataGroup_lo_lo_325 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_326;
  assign dataGroup_lo_lo_326 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_327;
  assign dataGroup_lo_lo_327 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_328;
  assign dataGroup_lo_lo_328 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_329;
  assign dataGroup_lo_lo_329 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_330;
  assign dataGroup_lo_lo_330 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_331;
  assign dataGroup_lo_lo_331 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_332;
  assign dataGroup_lo_lo_332 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_333;
  assign dataGroup_lo_lo_333 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_334;
  assign dataGroup_lo_lo_334 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_335;
  assign dataGroup_lo_lo_335 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_336;
  assign dataGroup_lo_lo_336 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_337;
  assign dataGroup_lo_lo_337 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_338;
  assign dataGroup_lo_lo_338 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_339;
  assign dataGroup_lo_lo_339 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_340;
  assign dataGroup_lo_lo_340 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_341;
  assign dataGroup_lo_lo_341 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_342;
  assign dataGroup_lo_lo_342 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_343;
  assign dataGroup_lo_lo_343 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_344;
  assign dataGroup_lo_lo_344 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_345;
  assign dataGroup_lo_lo_345 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_346;
  assign dataGroup_lo_lo_346 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_347;
  assign dataGroup_lo_lo_347 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_348;
  assign dataGroup_lo_lo_348 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_349;
  assign dataGroup_lo_lo_349 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_350;
  assign dataGroup_lo_lo_350 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_351;
  assign dataGroup_lo_lo_351 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_352;
  assign dataGroup_lo_lo_352 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_353;
  assign dataGroup_lo_lo_353 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_354;
  assign dataGroup_lo_lo_354 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_355;
  assign dataGroup_lo_lo_355 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_356;
  assign dataGroup_lo_lo_356 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_357;
  assign dataGroup_lo_lo_357 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_358;
  assign dataGroup_lo_lo_358 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_359;
  assign dataGroup_lo_lo_359 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_360;
  assign dataGroup_lo_lo_360 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_361;
  assign dataGroup_lo_lo_361 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_362;
  assign dataGroup_lo_lo_362 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_363;
  assign dataGroup_lo_lo_363 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_364;
  assign dataGroup_lo_lo_364 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_365;
  assign dataGroup_lo_lo_365 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_366;
  assign dataGroup_lo_lo_366 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_367;
  assign dataGroup_lo_lo_367 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_368;
  assign dataGroup_lo_lo_368 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_369;
  assign dataGroup_lo_lo_369 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_370;
  assign dataGroup_lo_lo_370 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_371;
  assign dataGroup_lo_lo_371 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_372;
  assign dataGroup_lo_lo_372 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_373;
  assign dataGroup_lo_lo_373 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_374;
  assign dataGroup_lo_lo_374 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_375;
  assign dataGroup_lo_lo_375 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_376;
  assign dataGroup_lo_lo_376 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_377;
  assign dataGroup_lo_lo_377 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_378;
  assign dataGroup_lo_lo_378 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_379;
  assign dataGroup_lo_lo_379 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_380;
  assign dataGroup_lo_lo_380 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_381;
  assign dataGroup_lo_lo_381 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_382;
  assign dataGroup_lo_lo_382 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_383;
  assign dataGroup_lo_lo_383 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_384;
  assign dataGroup_lo_lo_384 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_385;
  assign dataGroup_lo_lo_385 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_386;
  assign dataGroup_lo_lo_386 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_387;
  assign dataGroup_lo_lo_387 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_388;
  assign dataGroup_lo_lo_388 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_389;
  assign dataGroup_lo_lo_389 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_390;
  assign dataGroup_lo_lo_390 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_391;
  assign dataGroup_lo_lo_391 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_392;
  assign dataGroup_lo_lo_392 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_393;
  assign dataGroup_lo_lo_393 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_394;
  assign dataGroup_lo_lo_394 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_395;
  assign dataGroup_lo_lo_395 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_396;
  assign dataGroup_lo_lo_396 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_397;
  assign dataGroup_lo_lo_397 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_398;
  assign dataGroup_lo_lo_398 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_399;
  assign dataGroup_lo_lo_399 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_400;
  assign dataGroup_lo_lo_400 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_401;
  assign dataGroup_lo_lo_401 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_402;
  assign dataGroup_lo_lo_402 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_403;
  assign dataGroup_lo_lo_403 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_404;
  assign dataGroup_lo_lo_404 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_405;
  assign dataGroup_lo_lo_405 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_406;
  assign dataGroup_lo_lo_406 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_407;
  assign dataGroup_lo_lo_407 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_408;
  assign dataGroup_lo_lo_408 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_409;
  assign dataGroup_lo_lo_409 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_410;
  assign dataGroup_lo_lo_410 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_411;
  assign dataGroup_lo_lo_411 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_412;
  assign dataGroup_lo_lo_412 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_413;
  assign dataGroup_lo_lo_413 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_414;
  assign dataGroup_lo_lo_414 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_415;
  assign dataGroup_lo_lo_415 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_416;
  assign dataGroup_lo_lo_416 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_417;
  assign dataGroup_lo_lo_417 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_418;
  assign dataGroup_lo_lo_418 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_419;
  assign dataGroup_lo_lo_419 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_420;
  assign dataGroup_lo_lo_420 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_421;
  assign dataGroup_lo_lo_421 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_422;
  assign dataGroup_lo_lo_422 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_423;
  assign dataGroup_lo_lo_423 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_424;
  assign dataGroup_lo_lo_424 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_425;
  assign dataGroup_lo_lo_425 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_426;
  assign dataGroup_lo_lo_426 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_427;
  assign dataGroup_lo_lo_427 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_428;
  assign dataGroup_lo_lo_428 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_429;
  assign dataGroup_lo_lo_429 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_430;
  assign dataGroup_lo_lo_430 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_431;
  assign dataGroup_lo_lo_431 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_432;
  assign dataGroup_lo_lo_432 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_433;
  assign dataGroup_lo_lo_433 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_434;
  assign dataGroup_lo_lo_434 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_435;
  assign dataGroup_lo_lo_435 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_436;
  assign dataGroup_lo_lo_436 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_437;
  assign dataGroup_lo_lo_437 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_438;
  assign dataGroup_lo_lo_438 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_439;
  assign dataGroup_lo_lo_439 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_440;
  assign dataGroup_lo_lo_440 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_441;
  assign dataGroup_lo_lo_441 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_442;
  assign dataGroup_lo_lo_442 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_443;
  assign dataGroup_lo_lo_443 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_444;
  assign dataGroup_lo_lo_444 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_445;
  assign dataGroup_lo_lo_445 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_446;
  assign dataGroup_lo_lo_446 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_447;
  assign dataGroup_lo_lo_447 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_448;
  assign dataGroup_lo_lo_448 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_449;
  assign dataGroup_lo_lo_449 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_450;
  assign dataGroup_lo_lo_450 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_451;
  assign dataGroup_lo_lo_451 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_452;
  assign dataGroup_lo_lo_452 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_453;
  assign dataGroup_lo_lo_453 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_454;
  assign dataGroup_lo_lo_454 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_455;
  assign dataGroup_lo_lo_455 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_456;
  assign dataGroup_lo_lo_456 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_457;
  assign dataGroup_lo_lo_457 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_458;
  assign dataGroup_lo_lo_458 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_459;
  assign dataGroup_lo_lo_459 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_460;
  assign dataGroup_lo_lo_460 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_461;
  assign dataGroup_lo_lo_461 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_462;
  assign dataGroup_lo_lo_462 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_463;
  assign dataGroup_lo_lo_463 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_464;
  assign dataGroup_lo_lo_464 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_465;
  assign dataGroup_lo_lo_465 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_466;
  assign dataGroup_lo_lo_466 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_467;
  assign dataGroup_lo_lo_467 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_468;
  assign dataGroup_lo_lo_468 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_469;
  assign dataGroup_lo_lo_469 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_470;
  assign dataGroup_lo_lo_470 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_471;
  assign dataGroup_lo_lo_471 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_472;
  assign dataGroup_lo_lo_472 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_473;
  assign dataGroup_lo_lo_473 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_474;
  assign dataGroup_lo_lo_474 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_475;
  assign dataGroup_lo_lo_475 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_476;
  assign dataGroup_lo_lo_476 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_477;
  assign dataGroup_lo_lo_477 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_478;
  assign dataGroup_lo_lo_478 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_479;
  assign dataGroup_lo_lo_479 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_480;
  assign dataGroup_lo_lo_480 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_481;
  assign dataGroup_lo_lo_481 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_482;
  assign dataGroup_lo_lo_482 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_483;
  assign dataGroup_lo_lo_483 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_484;
  assign dataGroup_lo_lo_484 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_485;
  assign dataGroup_lo_lo_485 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_486;
  assign dataGroup_lo_lo_486 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_487;
  assign dataGroup_lo_lo_487 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_488;
  assign dataGroup_lo_lo_488 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_489;
  assign dataGroup_lo_lo_489 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_490;
  assign dataGroup_lo_lo_490 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_491;
  assign dataGroup_lo_lo_491 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_492;
  assign dataGroup_lo_lo_492 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_493;
  assign dataGroup_lo_lo_493 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_494;
  assign dataGroup_lo_lo_494 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_495;
  assign dataGroup_lo_lo_495 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_496;
  assign dataGroup_lo_lo_496 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_497;
  assign dataGroup_lo_lo_497 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_498;
  assign dataGroup_lo_lo_498 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_499;
  assign dataGroup_lo_lo_499 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_500;
  assign dataGroup_lo_lo_500 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_501;
  assign dataGroup_lo_lo_501 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_502;
  assign dataGroup_lo_lo_502 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_503;
  assign dataGroup_lo_lo_503 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_504;
  assign dataGroup_lo_lo_504 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_505;
  assign dataGroup_lo_lo_505 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_506;
  assign dataGroup_lo_lo_506 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_507;
  assign dataGroup_lo_lo_507 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_508;
  assign dataGroup_lo_lo_508 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_509;
  assign dataGroup_lo_lo_509 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_510;
  assign dataGroup_lo_lo_510 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_511;
  assign dataGroup_lo_lo_511 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_512;
  assign dataGroup_lo_lo_512 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_513;
  assign dataGroup_lo_lo_513 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_514;
  assign dataGroup_lo_lo_514 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_515;
  assign dataGroup_lo_lo_515 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_516;
  assign dataGroup_lo_lo_516 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_517;
  assign dataGroup_lo_lo_517 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_518;
  assign dataGroup_lo_lo_518 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_519;
  assign dataGroup_lo_lo_519 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_520;
  assign dataGroup_lo_lo_520 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_521;
  assign dataGroup_lo_lo_521 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_522;
  assign dataGroup_lo_lo_522 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_523;
  assign dataGroup_lo_lo_523 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_524;
  assign dataGroup_lo_lo_524 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_525;
  assign dataGroup_lo_lo_525 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_526;
  assign dataGroup_lo_lo_526 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_527;
  assign dataGroup_lo_lo_527 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_528;
  assign dataGroup_lo_lo_528 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_529;
  assign dataGroup_lo_lo_529 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_530;
  assign dataGroup_lo_lo_530 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_531;
  assign dataGroup_lo_lo_531 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_532;
  assign dataGroup_lo_lo_532 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_533;
  assign dataGroup_lo_lo_533 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_534;
  assign dataGroup_lo_lo_534 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_535;
  assign dataGroup_lo_lo_535 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_536;
  assign dataGroup_lo_lo_536 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_537;
  assign dataGroup_lo_lo_537 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_538;
  assign dataGroup_lo_lo_538 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_539;
  assign dataGroup_lo_lo_539 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_540;
  assign dataGroup_lo_lo_540 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_541;
  assign dataGroup_lo_lo_541 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_542;
  assign dataGroup_lo_lo_542 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_543;
  assign dataGroup_lo_lo_543 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_544;
  assign dataGroup_lo_lo_544 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_545;
  assign dataGroup_lo_lo_545 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_546;
  assign dataGroup_lo_lo_546 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_547;
  assign dataGroup_lo_lo_547 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_548;
  assign dataGroup_lo_lo_548 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_549;
  assign dataGroup_lo_lo_549 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_550;
  assign dataGroup_lo_lo_550 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_551;
  assign dataGroup_lo_lo_551 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_552;
  assign dataGroup_lo_lo_552 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_553;
  assign dataGroup_lo_lo_553 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_554;
  assign dataGroup_lo_lo_554 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_555;
  assign dataGroup_lo_lo_555 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_556;
  assign dataGroup_lo_lo_556 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_557;
  assign dataGroup_lo_lo_557 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_558;
  assign dataGroup_lo_lo_558 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_559;
  assign dataGroup_lo_lo_559 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_560;
  assign dataGroup_lo_lo_560 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_561;
  assign dataGroup_lo_lo_561 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_562;
  assign dataGroup_lo_lo_562 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_563;
  assign dataGroup_lo_lo_563 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_564;
  assign dataGroup_lo_lo_564 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_565;
  assign dataGroup_lo_lo_565 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_566;
  assign dataGroup_lo_lo_566 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_567;
  assign dataGroup_lo_lo_567 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_568;
  assign dataGroup_lo_lo_568 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_569;
  assign dataGroup_lo_lo_569 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_570;
  assign dataGroup_lo_lo_570 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_571;
  assign dataGroup_lo_lo_571 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_572;
  assign dataGroup_lo_lo_572 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_573;
  assign dataGroup_lo_lo_573 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_574;
  assign dataGroup_lo_lo_574 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_575;
  assign dataGroup_lo_lo_575 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_576;
  assign dataGroup_lo_lo_576 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_577;
  assign dataGroup_lo_lo_577 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_578;
  assign dataGroup_lo_lo_578 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_579;
  assign dataGroup_lo_lo_579 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_580;
  assign dataGroup_lo_lo_580 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_581;
  assign dataGroup_lo_lo_581 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_582;
  assign dataGroup_lo_lo_582 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_583;
  assign dataGroup_lo_lo_583 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_584;
  assign dataGroup_lo_lo_584 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_585;
  assign dataGroup_lo_lo_585 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_586;
  assign dataGroup_lo_lo_586 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_587;
  assign dataGroup_lo_lo_587 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_588;
  assign dataGroup_lo_lo_588 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_589;
  assign dataGroup_lo_lo_589 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_590;
  assign dataGroup_lo_lo_590 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_591;
  assign dataGroup_lo_lo_591 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_592;
  assign dataGroup_lo_lo_592 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_593;
  assign dataGroup_lo_lo_593 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_594;
  assign dataGroup_lo_lo_594 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_595;
  assign dataGroup_lo_lo_595 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_596;
  assign dataGroup_lo_lo_596 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_597;
  assign dataGroup_lo_lo_597 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_598;
  assign dataGroup_lo_lo_598 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_599;
  assign dataGroup_lo_lo_599 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_600;
  assign dataGroup_lo_lo_600 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_601;
  assign dataGroup_lo_lo_601 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_602;
  assign dataGroup_lo_lo_602 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_603;
  assign dataGroup_lo_lo_603 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_604;
  assign dataGroup_lo_lo_604 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_605;
  assign dataGroup_lo_lo_605 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_606;
  assign dataGroup_lo_lo_606 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_607;
  assign dataGroup_lo_lo_607 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_608;
  assign dataGroup_lo_lo_608 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_609;
  assign dataGroup_lo_lo_609 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_610;
  assign dataGroup_lo_lo_610 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_611;
  assign dataGroup_lo_lo_611 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_612;
  assign dataGroup_lo_lo_612 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_613;
  assign dataGroup_lo_lo_613 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_614;
  assign dataGroup_lo_lo_614 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_615;
  assign dataGroup_lo_lo_615 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_616;
  assign dataGroup_lo_lo_616 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_617;
  assign dataGroup_lo_lo_617 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_618;
  assign dataGroup_lo_lo_618 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_619;
  assign dataGroup_lo_lo_619 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_620;
  assign dataGroup_lo_lo_620 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_621;
  assign dataGroup_lo_lo_621 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_622;
  assign dataGroup_lo_lo_622 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_623;
  assign dataGroup_lo_lo_623 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_624;
  assign dataGroup_lo_lo_624 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_625;
  assign dataGroup_lo_lo_625 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_626;
  assign dataGroup_lo_lo_626 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_627;
  assign dataGroup_lo_lo_627 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_628;
  assign dataGroup_lo_lo_628 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_629;
  assign dataGroup_lo_lo_629 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_630;
  assign dataGroup_lo_lo_630 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_631;
  assign dataGroup_lo_lo_631 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_632;
  assign dataGroup_lo_lo_632 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_633;
  assign dataGroup_lo_lo_633 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_634;
  assign dataGroup_lo_lo_634 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_635;
  assign dataGroup_lo_lo_635 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_636;
  assign dataGroup_lo_lo_636 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_637;
  assign dataGroup_lo_lo_637 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_638;
  assign dataGroup_lo_lo_638 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_639;
  assign dataGroup_lo_lo_639 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_640;
  assign dataGroup_lo_lo_640 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_641;
  assign dataGroup_lo_lo_641 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_642;
  assign dataGroup_lo_lo_642 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_643;
  assign dataGroup_lo_lo_643 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_644;
  assign dataGroup_lo_lo_644 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_645;
  assign dataGroup_lo_lo_645 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_646;
  assign dataGroup_lo_lo_646 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_647;
  assign dataGroup_lo_lo_647 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_648;
  assign dataGroup_lo_lo_648 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_649;
  assign dataGroup_lo_lo_649 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_650;
  assign dataGroup_lo_lo_650 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_651;
  assign dataGroup_lo_lo_651 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_652;
  assign dataGroup_lo_lo_652 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_653;
  assign dataGroup_lo_lo_653 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_654;
  assign dataGroup_lo_lo_654 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_655;
  assign dataGroup_lo_lo_655 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_656;
  assign dataGroup_lo_lo_656 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_657;
  assign dataGroup_lo_lo_657 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_658;
  assign dataGroup_lo_lo_658 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_659;
  assign dataGroup_lo_lo_659 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_660;
  assign dataGroup_lo_lo_660 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_661;
  assign dataGroup_lo_lo_661 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_662;
  assign dataGroup_lo_lo_662 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_663;
  assign dataGroup_lo_lo_663 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_664;
  assign dataGroup_lo_lo_664 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_665;
  assign dataGroup_lo_lo_665 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_666;
  assign dataGroup_lo_lo_666 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_667;
  assign dataGroup_lo_lo_667 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_668;
  assign dataGroup_lo_lo_668 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_669;
  assign dataGroup_lo_lo_669 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_670;
  assign dataGroup_lo_lo_670 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_671;
  assign dataGroup_lo_lo_671 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_672;
  assign dataGroup_lo_lo_672 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_673;
  assign dataGroup_lo_lo_673 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_674;
  assign dataGroup_lo_lo_674 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_675;
  assign dataGroup_lo_lo_675 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_676;
  assign dataGroup_lo_lo_676 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_677;
  assign dataGroup_lo_lo_677 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_678;
  assign dataGroup_lo_lo_678 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_679;
  assign dataGroup_lo_lo_679 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_680;
  assign dataGroup_lo_lo_680 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_681;
  assign dataGroup_lo_lo_681 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_682;
  assign dataGroup_lo_lo_682 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_683;
  assign dataGroup_lo_lo_683 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_684;
  assign dataGroup_lo_lo_684 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_685;
  assign dataGroup_lo_lo_685 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_686;
  assign dataGroup_lo_lo_686 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_687;
  assign dataGroup_lo_lo_687 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_688;
  assign dataGroup_lo_lo_688 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_689;
  assign dataGroup_lo_lo_689 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_690;
  assign dataGroup_lo_lo_690 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_691;
  assign dataGroup_lo_lo_691 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_692;
  assign dataGroup_lo_lo_692 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_693;
  assign dataGroup_lo_lo_693 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_694;
  assign dataGroup_lo_lo_694 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_695;
  assign dataGroup_lo_lo_695 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_696;
  assign dataGroup_lo_lo_696 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_697;
  assign dataGroup_lo_lo_697 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_698;
  assign dataGroup_lo_lo_698 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_699;
  assign dataGroup_lo_lo_699 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_700;
  assign dataGroup_lo_lo_700 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_701;
  assign dataGroup_lo_lo_701 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_702;
  assign dataGroup_lo_lo_702 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_703;
  assign dataGroup_lo_lo_703 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_704;
  assign dataGroup_lo_lo_704 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_705;
  assign dataGroup_lo_lo_705 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_706;
  assign dataGroup_lo_lo_706 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_707;
  assign dataGroup_lo_lo_707 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_708;
  assign dataGroup_lo_lo_708 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_709;
  assign dataGroup_lo_lo_709 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_710;
  assign dataGroup_lo_lo_710 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_711;
  assign dataGroup_lo_lo_711 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_712;
  assign dataGroup_lo_lo_712 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_713;
  assign dataGroup_lo_lo_713 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_714;
  assign dataGroup_lo_lo_714 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_715;
  assign dataGroup_lo_lo_715 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_716;
  assign dataGroup_lo_lo_716 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_717;
  assign dataGroup_lo_lo_717 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_718;
  assign dataGroup_lo_lo_718 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_719;
  assign dataGroup_lo_lo_719 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_720;
  assign dataGroup_lo_lo_720 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_721;
  assign dataGroup_lo_lo_721 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_722;
  assign dataGroup_lo_lo_722 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_723;
  assign dataGroup_lo_lo_723 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_724;
  assign dataGroup_lo_lo_724 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_725;
  assign dataGroup_lo_lo_725 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_726;
  assign dataGroup_lo_lo_726 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_727;
  assign dataGroup_lo_lo_727 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_728;
  assign dataGroup_lo_lo_728 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_729;
  assign dataGroup_lo_lo_729 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_730;
  assign dataGroup_lo_lo_730 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_731;
  assign dataGroup_lo_lo_731 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_732;
  assign dataGroup_lo_lo_732 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_733;
  assign dataGroup_lo_lo_733 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_734;
  assign dataGroup_lo_lo_734 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_735;
  assign dataGroup_lo_lo_735 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_736;
  assign dataGroup_lo_lo_736 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_737;
  assign dataGroup_lo_lo_737 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_738;
  assign dataGroup_lo_lo_738 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_739;
  assign dataGroup_lo_lo_739 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_740;
  assign dataGroup_lo_lo_740 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_741;
  assign dataGroup_lo_lo_741 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_742;
  assign dataGroup_lo_lo_742 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_743;
  assign dataGroup_lo_lo_743 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_744;
  assign dataGroup_lo_lo_744 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_745;
  assign dataGroup_lo_lo_745 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_746;
  assign dataGroup_lo_lo_746 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_747;
  assign dataGroup_lo_lo_747 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_748;
  assign dataGroup_lo_lo_748 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_749;
  assign dataGroup_lo_lo_749 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_750;
  assign dataGroup_lo_lo_750 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_751;
  assign dataGroup_lo_lo_751 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_752;
  assign dataGroup_lo_lo_752 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_753;
  assign dataGroup_lo_lo_753 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_754;
  assign dataGroup_lo_lo_754 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_755;
  assign dataGroup_lo_lo_755 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_756;
  assign dataGroup_lo_lo_756 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_757;
  assign dataGroup_lo_lo_757 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_758;
  assign dataGroup_lo_lo_758 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_759;
  assign dataGroup_lo_lo_759 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_760;
  assign dataGroup_lo_lo_760 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_761;
  assign dataGroup_lo_lo_761 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_762;
  assign dataGroup_lo_lo_762 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_763;
  assign dataGroup_lo_lo_763 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_764;
  assign dataGroup_lo_lo_764 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_765;
  assign dataGroup_lo_lo_765 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_766;
  assign dataGroup_lo_lo_766 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_767;
  assign dataGroup_lo_lo_767 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_768;
  assign dataGroup_lo_lo_768 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_769;
  assign dataGroup_lo_lo_769 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_770;
  assign dataGroup_lo_lo_770 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_771;
  assign dataGroup_lo_lo_771 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_772;
  assign dataGroup_lo_lo_772 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_773;
  assign dataGroup_lo_lo_773 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_774;
  assign dataGroup_lo_lo_774 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_775;
  assign dataGroup_lo_lo_775 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_776;
  assign dataGroup_lo_lo_776 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_777;
  assign dataGroup_lo_lo_777 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_778;
  assign dataGroup_lo_lo_778 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_779;
  assign dataGroup_lo_lo_779 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_780;
  assign dataGroup_lo_lo_780 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_781;
  assign dataGroup_lo_lo_781 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_782;
  assign dataGroup_lo_lo_782 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_783;
  assign dataGroup_lo_lo_783 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_784;
  assign dataGroup_lo_lo_784 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_785;
  assign dataGroup_lo_lo_785 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_786;
  assign dataGroup_lo_lo_786 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_787;
  assign dataGroup_lo_lo_787 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_788;
  assign dataGroup_lo_lo_788 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_789;
  assign dataGroup_lo_lo_789 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_790;
  assign dataGroup_lo_lo_790 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_791;
  assign dataGroup_lo_lo_791 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_792;
  assign dataGroup_lo_lo_792 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_793;
  assign dataGroup_lo_lo_793 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_794;
  assign dataGroup_lo_lo_794 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_795;
  assign dataGroup_lo_lo_795 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_796;
  assign dataGroup_lo_lo_796 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_797;
  assign dataGroup_lo_lo_797 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_798;
  assign dataGroup_lo_lo_798 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_799;
  assign dataGroup_lo_lo_799 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_800;
  assign dataGroup_lo_lo_800 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_801;
  assign dataGroup_lo_lo_801 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_802;
  assign dataGroup_lo_lo_802 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_803;
  assign dataGroup_lo_lo_803 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_804;
  assign dataGroup_lo_lo_804 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_805;
  assign dataGroup_lo_lo_805 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_806;
  assign dataGroup_lo_lo_806 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_807;
  assign dataGroup_lo_lo_807 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_808;
  assign dataGroup_lo_lo_808 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_809;
  assign dataGroup_lo_lo_809 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_810;
  assign dataGroup_lo_lo_810 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_811;
  assign dataGroup_lo_lo_811 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_812;
  assign dataGroup_lo_lo_812 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_813;
  assign dataGroup_lo_lo_813 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_814;
  assign dataGroup_lo_lo_814 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_815;
  assign dataGroup_lo_lo_815 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_816;
  assign dataGroup_lo_lo_816 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_817;
  assign dataGroup_lo_lo_817 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_818;
  assign dataGroup_lo_lo_818 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_819;
  assign dataGroup_lo_lo_819 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_820;
  assign dataGroup_lo_lo_820 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_821;
  assign dataGroup_lo_lo_821 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_822;
  assign dataGroup_lo_lo_822 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_823;
  assign dataGroup_lo_lo_823 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_824;
  assign dataGroup_lo_lo_824 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_825;
  assign dataGroup_lo_lo_825 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_826;
  assign dataGroup_lo_lo_826 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_827;
  assign dataGroup_lo_lo_827 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_828;
  assign dataGroup_lo_lo_828 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_829;
  assign dataGroup_lo_lo_829 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_830;
  assign dataGroup_lo_lo_830 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_831;
  assign dataGroup_lo_lo_831 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_832;
  assign dataGroup_lo_lo_832 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_833;
  assign dataGroup_lo_lo_833 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_834;
  assign dataGroup_lo_lo_834 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_835;
  assign dataGroup_lo_lo_835 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_836;
  assign dataGroup_lo_lo_836 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_837;
  assign dataGroup_lo_lo_837 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_838;
  assign dataGroup_lo_lo_838 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_839;
  assign dataGroup_lo_lo_839 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_840;
  assign dataGroup_lo_lo_840 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_841;
  assign dataGroup_lo_lo_841 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_842;
  assign dataGroup_lo_lo_842 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_843;
  assign dataGroup_lo_lo_843 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_844;
  assign dataGroup_lo_lo_844 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_845;
  assign dataGroup_lo_lo_845 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_846;
  assign dataGroup_lo_lo_846 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_847;
  assign dataGroup_lo_lo_847 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_848;
  assign dataGroup_lo_lo_848 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_849;
  assign dataGroup_lo_lo_849 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_850;
  assign dataGroup_lo_lo_850 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_851;
  assign dataGroup_lo_lo_851 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_852;
  assign dataGroup_lo_lo_852 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_853;
  assign dataGroup_lo_lo_853 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_854;
  assign dataGroup_lo_lo_854 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_855;
  assign dataGroup_lo_lo_855 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_856;
  assign dataGroup_lo_lo_856 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_857;
  assign dataGroup_lo_lo_857 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_858;
  assign dataGroup_lo_lo_858 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_859;
  assign dataGroup_lo_lo_859 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_860;
  assign dataGroup_lo_lo_860 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_861;
  assign dataGroup_lo_lo_861 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_862;
  assign dataGroup_lo_lo_862 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_863;
  assign dataGroup_lo_lo_863 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_864;
  assign dataGroup_lo_lo_864 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_865;
  assign dataGroup_lo_lo_865 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_866;
  assign dataGroup_lo_lo_866 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_867;
  assign dataGroup_lo_lo_867 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_868;
  assign dataGroup_lo_lo_868 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_869;
  assign dataGroup_lo_lo_869 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_870;
  assign dataGroup_lo_lo_870 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_871;
  assign dataGroup_lo_lo_871 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_872;
  assign dataGroup_lo_lo_872 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_873;
  assign dataGroup_lo_lo_873 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_874;
  assign dataGroup_lo_lo_874 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_875;
  assign dataGroup_lo_lo_875 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_876;
  assign dataGroup_lo_lo_876 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_877;
  assign dataGroup_lo_lo_877 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_878;
  assign dataGroup_lo_lo_878 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_879;
  assign dataGroup_lo_lo_879 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_880;
  assign dataGroup_lo_lo_880 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_881;
  assign dataGroup_lo_lo_881 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_882;
  assign dataGroup_lo_lo_882 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_883;
  assign dataGroup_lo_lo_883 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_884;
  assign dataGroup_lo_lo_884 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_885;
  assign dataGroup_lo_lo_885 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_886;
  assign dataGroup_lo_lo_886 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_887;
  assign dataGroup_lo_lo_887 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_888;
  assign dataGroup_lo_lo_888 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_889;
  assign dataGroup_lo_lo_889 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_890;
  assign dataGroup_lo_lo_890 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_891;
  assign dataGroup_lo_lo_891 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_892;
  assign dataGroup_lo_lo_892 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_893;
  assign dataGroup_lo_lo_893 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_894;
  assign dataGroup_lo_lo_894 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_895;
  assign dataGroup_lo_lo_895 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_896;
  assign dataGroup_lo_lo_896 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_897;
  assign dataGroup_lo_lo_897 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_898;
  assign dataGroup_lo_lo_898 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_899;
  assign dataGroup_lo_lo_899 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_900;
  assign dataGroup_lo_lo_900 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_901;
  assign dataGroup_lo_lo_901 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_902;
  assign dataGroup_lo_lo_902 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_903;
  assign dataGroup_lo_lo_903 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_904;
  assign dataGroup_lo_lo_904 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_905;
  assign dataGroup_lo_lo_905 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_906;
  assign dataGroup_lo_lo_906 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_907;
  assign dataGroup_lo_lo_907 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_908;
  assign dataGroup_lo_lo_908 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_909;
  assign dataGroup_lo_lo_909 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_910;
  assign dataGroup_lo_lo_910 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_911;
  assign dataGroup_lo_lo_911 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_912;
  assign dataGroup_lo_lo_912 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_913;
  assign dataGroup_lo_lo_913 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_914;
  assign dataGroup_lo_lo_914 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_915;
  assign dataGroup_lo_lo_915 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_916;
  assign dataGroup_lo_lo_916 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_917;
  assign dataGroup_lo_lo_917 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_918;
  assign dataGroup_lo_lo_918 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_919;
  assign dataGroup_lo_lo_919 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_920;
  assign dataGroup_lo_lo_920 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_921;
  assign dataGroup_lo_lo_921 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_922;
  assign dataGroup_lo_lo_922 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_923;
  assign dataGroup_lo_lo_923 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_924;
  assign dataGroup_lo_lo_924 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_925;
  assign dataGroup_lo_lo_925 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_926;
  assign dataGroup_lo_lo_926 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_927;
  assign dataGroup_lo_lo_927 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_928;
  assign dataGroup_lo_lo_928 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_929;
  assign dataGroup_lo_lo_929 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_930;
  assign dataGroup_lo_lo_930 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_931;
  assign dataGroup_lo_lo_931 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_932;
  assign dataGroup_lo_lo_932 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_933;
  assign dataGroup_lo_lo_933 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_934;
  assign dataGroup_lo_lo_934 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_935;
  assign dataGroup_lo_lo_935 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_936;
  assign dataGroup_lo_lo_936 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_937;
  assign dataGroup_lo_lo_937 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_938;
  assign dataGroup_lo_lo_938 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_939;
  assign dataGroup_lo_lo_939 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_940;
  assign dataGroup_lo_lo_940 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_941;
  assign dataGroup_lo_lo_941 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_942;
  assign dataGroup_lo_lo_942 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_943;
  assign dataGroup_lo_lo_943 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_944;
  assign dataGroup_lo_lo_944 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_945;
  assign dataGroup_lo_lo_945 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_946;
  assign dataGroup_lo_lo_946 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_947;
  assign dataGroup_lo_lo_947 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_948;
  assign dataGroup_lo_lo_948 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_949;
  assign dataGroup_lo_lo_949 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_950;
  assign dataGroup_lo_lo_950 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_951;
  assign dataGroup_lo_lo_951 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_952;
  assign dataGroup_lo_lo_952 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_953;
  assign dataGroup_lo_lo_953 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_954;
  assign dataGroup_lo_lo_954 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_955;
  assign dataGroup_lo_lo_955 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_956;
  assign dataGroup_lo_lo_956 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_957;
  assign dataGroup_lo_lo_957 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_958;
  assign dataGroup_lo_lo_958 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_959;
  assign dataGroup_lo_lo_959 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_960;
  assign dataGroup_lo_lo_960 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_961;
  assign dataGroup_lo_lo_961 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_962;
  assign dataGroup_lo_lo_962 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_963;
  assign dataGroup_lo_lo_963 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_964;
  assign dataGroup_lo_lo_964 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_965;
  assign dataGroup_lo_lo_965 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_966;
  assign dataGroup_lo_lo_966 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_967;
  assign dataGroup_lo_lo_967 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_968;
  assign dataGroup_lo_lo_968 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_969;
  assign dataGroup_lo_lo_969 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_970;
  assign dataGroup_lo_lo_970 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_971;
  assign dataGroup_lo_lo_971 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_972;
  assign dataGroup_lo_lo_972 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_973;
  assign dataGroup_lo_lo_973 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_974;
  assign dataGroup_lo_lo_974 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_975;
  assign dataGroup_lo_lo_975 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_976;
  assign dataGroup_lo_lo_976 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_977;
  assign dataGroup_lo_lo_977 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_978;
  assign dataGroup_lo_lo_978 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_979;
  assign dataGroup_lo_lo_979 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_980;
  assign dataGroup_lo_lo_980 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_981;
  assign dataGroup_lo_lo_981 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_982;
  assign dataGroup_lo_lo_982 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_983;
  assign dataGroup_lo_lo_983 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_984;
  assign dataGroup_lo_lo_984 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_985;
  assign dataGroup_lo_lo_985 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_986;
  assign dataGroup_lo_lo_986 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_987;
  assign dataGroup_lo_lo_987 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_988;
  assign dataGroup_lo_lo_988 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_989;
  assign dataGroup_lo_lo_989 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_990;
  assign dataGroup_lo_lo_990 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_991;
  assign dataGroup_lo_lo_991 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_992;
  assign dataGroup_lo_lo_992 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_993;
  assign dataGroup_lo_lo_993 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_994;
  assign dataGroup_lo_lo_994 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_995;
  assign dataGroup_lo_lo_995 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_996;
  assign dataGroup_lo_lo_996 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_997;
  assign dataGroup_lo_lo_997 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_998;
  assign dataGroup_lo_lo_998 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_999;
  assign dataGroup_lo_lo_999 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1000;
  assign dataGroup_lo_lo_1000 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1001;
  assign dataGroup_lo_lo_1001 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1002;
  assign dataGroup_lo_lo_1002 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1003;
  assign dataGroup_lo_lo_1003 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1004;
  assign dataGroup_lo_lo_1004 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1005;
  assign dataGroup_lo_lo_1005 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1006;
  assign dataGroup_lo_lo_1006 = _GEN_3;
  wire [255:0]  dataGroup_lo_lo_1007;
  assign dataGroup_lo_lo_1007 = _GEN_3;
  wire [255:0]  _GEN_4 = {dataSelect_3, dataSelect_2};
  wire [255:0]  dataGroup_lo_hi;
  assign dataGroup_lo_hi = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1;
  assign dataGroup_lo_hi_1 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_2;
  assign dataGroup_lo_hi_2 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_3;
  assign dataGroup_lo_hi_3 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_4;
  assign dataGroup_lo_hi_4 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_5;
  assign dataGroup_lo_hi_5 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_6;
  assign dataGroup_lo_hi_6 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_7;
  assign dataGroup_lo_hi_7 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_8;
  assign dataGroup_lo_hi_8 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_9;
  assign dataGroup_lo_hi_9 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_10;
  assign dataGroup_lo_hi_10 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_11;
  assign dataGroup_lo_hi_11 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_12;
  assign dataGroup_lo_hi_12 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_13;
  assign dataGroup_lo_hi_13 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_14;
  assign dataGroup_lo_hi_14 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_15;
  assign dataGroup_lo_hi_15 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_16;
  assign dataGroup_lo_hi_16 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_17;
  assign dataGroup_lo_hi_17 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_18;
  assign dataGroup_lo_hi_18 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_19;
  assign dataGroup_lo_hi_19 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_20;
  assign dataGroup_lo_hi_20 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_21;
  assign dataGroup_lo_hi_21 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_22;
  assign dataGroup_lo_hi_22 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_23;
  assign dataGroup_lo_hi_23 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_24;
  assign dataGroup_lo_hi_24 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_25;
  assign dataGroup_lo_hi_25 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_26;
  assign dataGroup_lo_hi_26 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_27;
  assign dataGroup_lo_hi_27 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_28;
  assign dataGroup_lo_hi_28 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_29;
  assign dataGroup_lo_hi_29 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_30;
  assign dataGroup_lo_hi_30 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_31;
  assign dataGroup_lo_hi_31 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_32;
  assign dataGroup_lo_hi_32 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_33;
  assign dataGroup_lo_hi_33 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_34;
  assign dataGroup_lo_hi_34 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_35;
  assign dataGroup_lo_hi_35 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_36;
  assign dataGroup_lo_hi_36 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_37;
  assign dataGroup_lo_hi_37 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_38;
  assign dataGroup_lo_hi_38 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_39;
  assign dataGroup_lo_hi_39 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_40;
  assign dataGroup_lo_hi_40 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_41;
  assign dataGroup_lo_hi_41 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_42;
  assign dataGroup_lo_hi_42 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_43;
  assign dataGroup_lo_hi_43 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_44;
  assign dataGroup_lo_hi_44 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_45;
  assign dataGroup_lo_hi_45 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_46;
  assign dataGroup_lo_hi_46 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_47;
  assign dataGroup_lo_hi_47 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_48;
  assign dataGroup_lo_hi_48 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_49;
  assign dataGroup_lo_hi_49 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_50;
  assign dataGroup_lo_hi_50 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_51;
  assign dataGroup_lo_hi_51 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_52;
  assign dataGroup_lo_hi_52 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_53;
  assign dataGroup_lo_hi_53 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_54;
  assign dataGroup_lo_hi_54 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_55;
  assign dataGroup_lo_hi_55 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_56;
  assign dataGroup_lo_hi_56 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_57;
  assign dataGroup_lo_hi_57 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_58;
  assign dataGroup_lo_hi_58 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_59;
  assign dataGroup_lo_hi_59 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_60;
  assign dataGroup_lo_hi_60 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_61;
  assign dataGroup_lo_hi_61 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_62;
  assign dataGroup_lo_hi_62 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_63;
  assign dataGroup_lo_hi_63 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_64;
  assign dataGroup_lo_hi_64 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_65;
  assign dataGroup_lo_hi_65 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_66;
  assign dataGroup_lo_hi_66 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_67;
  assign dataGroup_lo_hi_67 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_68;
  assign dataGroup_lo_hi_68 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_69;
  assign dataGroup_lo_hi_69 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_70;
  assign dataGroup_lo_hi_70 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_71;
  assign dataGroup_lo_hi_71 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_72;
  assign dataGroup_lo_hi_72 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_73;
  assign dataGroup_lo_hi_73 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_74;
  assign dataGroup_lo_hi_74 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_75;
  assign dataGroup_lo_hi_75 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_76;
  assign dataGroup_lo_hi_76 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_77;
  assign dataGroup_lo_hi_77 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_78;
  assign dataGroup_lo_hi_78 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_79;
  assign dataGroup_lo_hi_79 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_80;
  assign dataGroup_lo_hi_80 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_81;
  assign dataGroup_lo_hi_81 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_82;
  assign dataGroup_lo_hi_82 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_83;
  assign dataGroup_lo_hi_83 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_84;
  assign dataGroup_lo_hi_84 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_85;
  assign dataGroup_lo_hi_85 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_86;
  assign dataGroup_lo_hi_86 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_87;
  assign dataGroup_lo_hi_87 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_88;
  assign dataGroup_lo_hi_88 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_89;
  assign dataGroup_lo_hi_89 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_90;
  assign dataGroup_lo_hi_90 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_91;
  assign dataGroup_lo_hi_91 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_92;
  assign dataGroup_lo_hi_92 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_93;
  assign dataGroup_lo_hi_93 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_94;
  assign dataGroup_lo_hi_94 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_95;
  assign dataGroup_lo_hi_95 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_96;
  assign dataGroup_lo_hi_96 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_97;
  assign dataGroup_lo_hi_97 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_98;
  assign dataGroup_lo_hi_98 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_99;
  assign dataGroup_lo_hi_99 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_100;
  assign dataGroup_lo_hi_100 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_101;
  assign dataGroup_lo_hi_101 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_102;
  assign dataGroup_lo_hi_102 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_103;
  assign dataGroup_lo_hi_103 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_104;
  assign dataGroup_lo_hi_104 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_105;
  assign dataGroup_lo_hi_105 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_106;
  assign dataGroup_lo_hi_106 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_107;
  assign dataGroup_lo_hi_107 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_108;
  assign dataGroup_lo_hi_108 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_109;
  assign dataGroup_lo_hi_109 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_110;
  assign dataGroup_lo_hi_110 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_111;
  assign dataGroup_lo_hi_111 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_112;
  assign dataGroup_lo_hi_112 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_113;
  assign dataGroup_lo_hi_113 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_114;
  assign dataGroup_lo_hi_114 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_115;
  assign dataGroup_lo_hi_115 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_116;
  assign dataGroup_lo_hi_116 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_117;
  assign dataGroup_lo_hi_117 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_118;
  assign dataGroup_lo_hi_118 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_119;
  assign dataGroup_lo_hi_119 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_120;
  assign dataGroup_lo_hi_120 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_121;
  assign dataGroup_lo_hi_121 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_122;
  assign dataGroup_lo_hi_122 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_123;
  assign dataGroup_lo_hi_123 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_124;
  assign dataGroup_lo_hi_124 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_125;
  assign dataGroup_lo_hi_125 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_126;
  assign dataGroup_lo_hi_126 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_127;
  assign dataGroup_lo_hi_127 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_128;
  assign dataGroup_lo_hi_128 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_129;
  assign dataGroup_lo_hi_129 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_130;
  assign dataGroup_lo_hi_130 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_131;
  assign dataGroup_lo_hi_131 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_132;
  assign dataGroup_lo_hi_132 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_133;
  assign dataGroup_lo_hi_133 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_134;
  assign dataGroup_lo_hi_134 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_135;
  assign dataGroup_lo_hi_135 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_136;
  assign dataGroup_lo_hi_136 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_137;
  assign dataGroup_lo_hi_137 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_138;
  assign dataGroup_lo_hi_138 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_139;
  assign dataGroup_lo_hi_139 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_140;
  assign dataGroup_lo_hi_140 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_141;
  assign dataGroup_lo_hi_141 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_142;
  assign dataGroup_lo_hi_142 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_143;
  assign dataGroup_lo_hi_143 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_144;
  assign dataGroup_lo_hi_144 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_145;
  assign dataGroup_lo_hi_145 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_146;
  assign dataGroup_lo_hi_146 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_147;
  assign dataGroup_lo_hi_147 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_148;
  assign dataGroup_lo_hi_148 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_149;
  assign dataGroup_lo_hi_149 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_150;
  assign dataGroup_lo_hi_150 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_151;
  assign dataGroup_lo_hi_151 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_152;
  assign dataGroup_lo_hi_152 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_153;
  assign dataGroup_lo_hi_153 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_154;
  assign dataGroup_lo_hi_154 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_155;
  assign dataGroup_lo_hi_155 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_156;
  assign dataGroup_lo_hi_156 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_157;
  assign dataGroup_lo_hi_157 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_158;
  assign dataGroup_lo_hi_158 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_159;
  assign dataGroup_lo_hi_159 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_160;
  assign dataGroup_lo_hi_160 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_161;
  assign dataGroup_lo_hi_161 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_162;
  assign dataGroup_lo_hi_162 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_163;
  assign dataGroup_lo_hi_163 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_164;
  assign dataGroup_lo_hi_164 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_165;
  assign dataGroup_lo_hi_165 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_166;
  assign dataGroup_lo_hi_166 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_167;
  assign dataGroup_lo_hi_167 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_168;
  assign dataGroup_lo_hi_168 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_169;
  assign dataGroup_lo_hi_169 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_170;
  assign dataGroup_lo_hi_170 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_171;
  assign dataGroup_lo_hi_171 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_172;
  assign dataGroup_lo_hi_172 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_173;
  assign dataGroup_lo_hi_173 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_174;
  assign dataGroup_lo_hi_174 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_175;
  assign dataGroup_lo_hi_175 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_176;
  assign dataGroup_lo_hi_176 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_177;
  assign dataGroup_lo_hi_177 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_178;
  assign dataGroup_lo_hi_178 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_179;
  assign dataGroup_lo_hi_179 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_180;
  assign dataGroup_lo_hi_180 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_181;
  assign dataGroup_lo_hi_181 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_182;
  assign dataGroup_lo_hi_182 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_183;
  assign dataGroup_lo_hi_183 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_184;
  assign dataGroup_lo_hi_184 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_185;
  assign dataGroup_lo_hi_185 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_186;
  assign dataGroup_lo_hi_186 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_187;
  assign dataGroup_lo_hi_187 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_188;
  assign dataGroup_lo_hi_188 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_189;
  assign dataGroup_lo_hi_189 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_190;
  assign dataGroup_lo_hi_190 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_191;
  assign dataGroup_lo_hi_191 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_192;
  assign dataGroup_lo_hi_192 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_193;
  assign dataGroup_lo_hi_193 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_194;
  assign dataGroup_lo_hi_194 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_195;
  assign dataGroup_lo_hi_195 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_196;
  assign dataGroup_lo_hi_196 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_197;
  assign dataGroup_lo_hi_197 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_198;
  assign dataGroup_lo_hi_198 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_199;
  assign dataGroup_lo_hi_199 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_200;
  assign dataGroup_lo_hi_200 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_201;
  assign dataGroup_lo_hi_201 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_202;
  assign dataGroup_lo_hi_202 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_203;
  assign dataGroup_lo_hi_203 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_204;
  assign dataGroup_lo_hi_204 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_205;
  assign dataGroup_lo_hi_205 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_206;
  assign dataGroup_lo_hi_206 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_207;
  assign dataGroup_lo_hi_207 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_208;
  assign dataGroup_lo_hi_208 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_209;
  assign dataGroup_lo_hi_209 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_210;
  assign dataGroup_lo_hi_210 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_211;
  assign dataGroup_lo_hi_211 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_212;
  assign dataGroup_lo_hi_212 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_213;
  assign dataGroup_lo_hi_213 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_214;
  assign dataGroup_lo_hi_214 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_215;
  assign dataGroup_lo_hi_215 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_216;
  assign dataGroup_lo_hi_216 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_217;
  assign dataGroup_lo_hi_217 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_218;
  assign dataGroup_lo_hi_218 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_219;
  assign dataGroup_lo_hi_219 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_220;
  assign dataGroup_lo_hi_220 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_221;
  assign dataGroup_lo_hi_221 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_222;
  assign dataGroup_lo_hi_222 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_223;
  assign dataGroup_lo_hi_223 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_224;
  assign dataGroup_lo_hi_224 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_225;
  assign dataGroup_lo_hi_225 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_226;
  assign dataGroup_lo_hi_226 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_227;
  assign dataGroup_lo_hi_227 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_228;
  assign dataGroup_lo_hi_228 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_229;
  assign dataGroup_lo_hi_229 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_230;
  assign dataGroup_lo_hi_230 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_231;
  assign dataGroup_lo_hi_231 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_232;
  assign dataGroup_lo_hi_232 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_233;
  assign dataGroup_lo_hi_233 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_234;
  assign dataGroup_lo_hi_234 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_235;
  assign dataGroup_lo_hi_235 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_236;
  assign dataGroup_lo_hi_236 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_237;
  assign dataGroup_lo_hi_237 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_238;
  assign dataGroup_lo_hi_238 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_239;
  assign dataGroup_lo_hi_239 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_240;
  assign dataGroup_lo_hi_240 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_241;
  assign dataGroup_lo_hi_241 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_242;
  assign dataGroup_lo_hi_242 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_243;
  assign dataGroup_lo_hi_243 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_244;
  assign dataGroup_lo_hi_244 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_245;
  assign dataGroup_lo_hi_245 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_246;
  assign dataGroup_lo_hi_246 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_247;
  assign dataGroup_lo_hi_247 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_248;
  assign dataGroup_lo_hi_248 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_249;
  assign dataGroup_lo_hi_249 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_250;
  assign dataGroup_lo_hi_250 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_251;
  assign dataGroup_lo_hi_251 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_252;
  assign dataGroup_lo_hi_252 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_253;
  assign dataGroup_lo_hi_253 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_254;
  assign dataGroup_lo_hi_254 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_255;
  assign dataGroup_lo_hi_255 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_256;
  assign dataGroup_lo_hi_256 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_257;
  assign dataGroup_lo_hi_257 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_258;
  assign dataGroup_lo_hi_258 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_259;
  assign dataGroup_lo_hi_259 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_260;
  assign dataGroup_lo_hi_260 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_261;
  assign dataGroup_lo_hi_261 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_262;
  assign dataGroup_lo_hi_262 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_263;
  assign dataGroup_lo_hi_263 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_264;
  assign dataGroup_lo_hi_264 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_265;
  assign dataGroup_lo_hi_265 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_266;
  assign dataGroup_lo_hi_266 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_267;
  assign dataGroup_lo_hi_267 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_268;
  assign dataGroup_lo_hi_268 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_269;
  assign dataGroup_lo_hi_269 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_270;
  assign dataGroup_lo_hi_270 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_271;
  assign dataGroup_lo_hi_271 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_272;
  assign dataGroup_lo_hi_272 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_273;
  assign dataGroup_lo_hi_273 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_274;
  assign dataGroup_lo_hi_274 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_275;
  assign dataGroup_lo_hi_275 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_276;
  assign dataGroup_lo_hi_276 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_277;
  assign dataGroup_lo_hi_277 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_278;
  assign dataGroup_lo_hi_278 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_279;
  assign dataGroup_lo_hi_279 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_280;
  assign dataGroup_lo_hi_280 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_281;
  assign dataGroup_lo_hi_281 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_282;
  assign dataGroup_lo_hi_282 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_283;
  assign dataGroup_lo_hi_283 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_284;
  assign dataGroup_lo_hi_284 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_285;
  assign dataGroup_lo_hi_285 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_286;
  assign dataGroup_lo_hi_286 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_287;
  assign dataGroup_lo_hi_287 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_288;
  assign dataGroup_lo_hi_288 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_289;
  assign dataGroup_lo_hi_289 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_290;
  assign dataGroup_lo_hi_290 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_291;
  assign dataGroup_lo_hi_291 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_292;
  assign dataGroup_lo_hi_292 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_293;
  assign dataGroup_lo_hi_293 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_294;
  assign dataGroup_lo_hi_294 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_295;
  assign dataGroup_lo_hi_295 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_296;
  assign dataGroup_lo_hi_296 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_297;
  assign dataGroup_lo_hi_297 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_298;
  assign dataGroup_lo_hi_298 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_299;
  assign dataGroup_lo_hi_299 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_300;
  assign dataGroup_lo_hi_300 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_301;
  assign dataGroup_lo_hi_301 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_302;
  assign dataGroup_lo_hi_302 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_303;
  assign dataGroup_lo_hi_303 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_304;
  assign dataGroup_lo_hi_304 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_305;
  assign dataGroup_lo_hi_305 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_306;
  assign dataGroup_lo_hi_306 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_307;
  assign dataGroup_lo_hi_307 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_308;
  assign dataGroup_lo_hi_308 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_309;
  assign dataGroup_lo_hi_309 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_310;
  assign dataGroup_lo_hi_310 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_311;
  assign dataGroup_lo_hi_311 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_312;
  assign dataGroup_lo_hi_312 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_313;
  assign dataGroup_lo_hi_313 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_314;
  assign dataGroup_lo_hi_314 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_315;
  assign dataGroup_lo_hi_315 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_316;
  assign dataGroup_lo_hi_316 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_317;
  assign dataGroup_lo_hi_317 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_318;
  assign dataGroup_lo_hi_318 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_319;
  assign dataGroup_lo_hi_319 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_320;
  assign dataGroup_lo_hi_320 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_321;
  assign dataGroup_lo_hi_321 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_322;
  assign dataGroup_lo_hi_322 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_323;
  assign dataGroup_lo_hi_323 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_324;
  assign dataGroup_lo_hi_324 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_325;
  assign dataGroup_lo_hi_325 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_326;
  assign dataGroup_lo_hi_326 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_327;
  assign dataGroup_lo_hi_327 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_328;
  assign dataGroup_lo_hi_328 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_329;
  assign dataGroup_lo_hi_329 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_330;
  assign dataGroup_lo_hi_330 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_331;
  assign dataGroup_lo_hi_331 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_332;
  assign dataGroup_lo_hi_332 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_333;
  assign dataGroup_lo_hi_333 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_334;
  assign dataGroup_lo_hi_334 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_335;
  assign dataGroup_lo_hi_335 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_336;
  assign dataGroup_lo_hi_336 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_337;
  assign dataGroup_lo_hi_337 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_338;
  assign dataGroup_lo_hi_338 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_339;
  assign dataGroup_lo_hi_339 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_340;
  assign dataGroup_lo_hi_340 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_341;
  assign dataGroup_lo_hi_341 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_342;
  assign dataGroup_lo_hi_342 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_343;
  assign dataGroup_lo_hi_343 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_344;
  assign dataGroup_lo_hi_344 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_345;
  assign dataGroup_lo_hi_345 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_346;
  assign dataGroup_lo_hi_346 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_347;
  assign dataGroup_lo_hi_347 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_348;
  assign dataGroup_lo_hi_348 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_349;
  assign dataGroup_lo_hi_349 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_350;
  assign dataGroup_lo_hi_350 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_351;
  assign dataGroup_lo_hi_351 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_352;
  assign dataGroup_lo_hi_352 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_353;
  assign dataGroup_lo_hi_353 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_354;
  assign dataGroup_lo_hi_354 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_355;
  assign dataGroup_lo_hi_355 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_356;
  assign dataGroup_lo_hi_356 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_357;
  assign dataGroup_lo_hi_357 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_358;
  assign dataGroup_lo_hi_358 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_359;
  assign dataGroup_lo_hi_359 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_360;
  assign dataGroup_lo_hi_360 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_361;
  assign dataGroup_lo_hi_361 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_362;
  assign dataGroup_lo_hi_362 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_363;
  assign dataGroup_lo_hi_363 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_364;
  assign dataGroup_lo_hi_364 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_365;
  assign dataGroup_lo_hi_365 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_366;
  assign dataGroup_lo_hi_366 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_367;
  assign dataGroup_lo_hi_367 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_368;
  assign dataGroup_lo_hi_368 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_369;
  assign dataGroup_lo_hi_369 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_370;
  assign dataGroup_lo_hi_370 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_371;
  assign dataGroup_lo_hi_371 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_372;
  assign dataGroup_lo_hi_372 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_373;
  assign dataGroup_lo_hi_373 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_374;
  assign dataGroup_lo_hi_374 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_375;
  assign dataGroup_lo_hi_375 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_376;
  assign dataGroup_lo_hi_376 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_377;
  assign dataGroup_lo_hi_377 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_378;
  assign dataGroup_lo_hi_378 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_379;
  assign dataGroup_lo_hi_379 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_380;
  assign dataGroup_lo_hi_380 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_381;
  assign dataGroup_lo_hi_381 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_382;
  assign dataGroup_lo_hi_382 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_383;
  assign dataGroup_lo_hi_383 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_384;
  assign dataGroup_lo_hi_384 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_385;
  assign dataGroup_lo_hi_385 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_386;
  assign dataGroup_lo_hi_386 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_387;
  assign dataGroup_lo_hi_387 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_388;
  assign dataGroup_lo_hi_388 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_389;
  assign dataGroup_lo_hi_389 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_390;
  assign dataGroup_lo_hi_390 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_391;
  assign dataGroup_lo_hi_391 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_392;
  assign dataGroup_lo_hi_392 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_393;
  assign dataGroup_lo_hi_393 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_394;
  assign dataGroup_lo_hi_394 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_395;
  assign dataGroup_lo_hi_395 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_396;
  assign dataGroup_lo_hi_396 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_397;
  assign dataGroup_lo_hi_397 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_398;
  assign dataGroup_lo_hi_398 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_399;
  assign dataGroup_lo_hi_399 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_400;
  assign dataGroup_lo_hi_400 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_401;
  assign dataGroup_lo_hi_401 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_402;
  assign dataGroup_lo_hi_402 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_403;
  assign dataGroup_lo_hi_403 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_404;
  assign dataGroup_lo_hi_404 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_405;
  assign dataGroup_lo_hi_405 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_406;
  assign dataGroup_lo_hi_406 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_407;
  assign dataGroup_lo_hi_407 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_408;
  assign dataGroup_lo_hi_408 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_409;
  assign dataGroup_lo_hi_409 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_410;
  assign dataGroup_lo_hi_410 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_411;
  assign dataGroup_lo_hi_411 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_412;
  assign dataGroup_lo_hi_412 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_413;
  assign dataGroup_lo_hi_413 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_414;
  assign dataGroup_lo_hi_414 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_415;
  assign dataGroup_lo_hi_415 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_416;
  assign dataGroup_lo_hi_416 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_417;
  assign dataGroup_lo_hi_417 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_418;
  assign dataGroup_lo_hi_418 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_419;
  assign dataGroup_lo_hi_419 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_420;
  assign dataGroup_lo_hi_420 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_421;
  assign dataGroup_lo_hi_421 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_422;
  assign dataGroup_lo_hi_422 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_423;
  assign dataGroup_lo_hi_423 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_424;
  assign dataGroup_lo_hi_424 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_425;
  assign dataGroup_lo_hi_425 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_426;
  assign dataGroup_lo_hi_426 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_427;
  assign dataGroup_lo_hi_427 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_428;
  assign dataGroup_lo_hi_428 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_429;
  assign dataGroup_lo_hi_429 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_430;
  assign dataGroup_lo_hi_430 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_431;
  assign dataGroup_lo_hi_431 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_432;
  assign dataGroup_lo_hi_432 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_433;
  assign dataGroup_lo_hi_433 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_434;
  assign dataGroup_lo_hi_434 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_435;
  assign dataGroup_lo_hi_435 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_436;
  assign dataGroup_lo_hi_436 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_437;
  assign dataGroup_lo_hi_437 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_438;
  assign dataGroup_lo_hi_438 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_439;
  assign dataGroup_lo_hi_439 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_440;
  assign dataGroup_lo_hi_440 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_441;
  assign dataGroup_lo_hi_441 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_442;
  assign dataGroup_lo_hi_442 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_443;
  assign dataGroup_lo_hi_443 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_444;
  assign dataGroup_lo_hi_444 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_445;
  assign dataGroup_lo_hi_445 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_446;
  assign dataGroup_lo_hi_446 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_447;
  assign dataGroup_lo_hi_447 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_448;
  assign dataGroup_lo_hi_448 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_449;
  assign dataGroup_lo_hi_449 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_450;
  assign dataGroup_lo_hi_450 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_451;
  assign dataGroup_lo_hi_451 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_452;
  assign dataGroup_lo_hi_452 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_453;
  assign dataGroup_lo_hi_453 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_454;
  assign dataGroup_lo_hi_454 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_455;
  assign dataGroup_lo_hi_455 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_456;
  assign dataGroup_lo_hi_456 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_457;
  assign dataGroup_lo_hi_457 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_458;
  assign dataGroup_lo_hi_458 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_459;
  assign dataGroup_lo_hi_459 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_460;
  assign dataGroup_lo_hi_460 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_461;
  assign dataGroup_lo_hi_461 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_462;
  assign dataGroup_lo_hi_462 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_463;
  assign dataGroup_lo_hi_463 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_464;
  assign dataGroup_lo_hi_464 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_465;
  assign dataGroup_lo_hi_465 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_466;
  assign dataGroup_lo_hi_466 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_467;
  assign dataGroup_lo_hi_467 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_468;
  assign dataGroup_lo_hi_468 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_469;
  assign dataGroup_lo_hi_469 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_470;
  assign dataGroup_lo_hi_470 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_471;
  assign dataGroup_lo_hi_471 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_472;
  assign dataGroup_lo_hi_472 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_473;
  assign dataGroup_lo_hi_473 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_474;
  assign dataGroup_lo_hi_474 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_475;
  assign dataGroup_lo_hi_475 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_476;
  assign dataGroup_lo_hi_476 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_477;
  assign dataGroup_lo_hi_477 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_478;
  assign dataGroup_lo_hi_478 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_479;
  assign dataGroup_lo_hi_479 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_480;
  assign dataGroup_lo_hi_480 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_481;
  assign dataGroup_lo_hi_481 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_482;
  assign dataGroup_lo_hi_482 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_483;
  assign dataGroup_lo_hi_483 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_484;
  assign dataGroup_lo_hi_484 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_485;
  assign dataGroup_lo_hi_485 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_486;
  assign dataGroup_lo_hi_486 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_487;
  assign dataGroup_lo_hi_487 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_488;
  assign dataGroup_lo_hi_488 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_489;
  assign dataGroup_lo_hi_489 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_490;
  assign dataGroup_lo_hi_490 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_491;
  assign dataGroup_lo_hi_491 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_492;
  assign dataGroup_lo_hi_492 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_493;
  assign dataGroup_lo_hi_493 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_494;
  assign dataGroup_lo_hi_494 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_495;
  assign dataGroup_lo_hi_495 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_496;
  assign dataGroup_lo_hi_496 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_497;
  assign dataGroup_lo_hi_497 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_498;
  assign dataGroup_lo_hi_498 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_499;
  assign dataGroup_lo_hi_499 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_500;
  assign dataGroup_lo_hi_500 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_501;
  assign dataGroup_lo_hi_501 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_502;
  assign dataGroup_lo_hi_502 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_503;
  assign dataGroup_lo_hi_503 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_504;
  assign dataGroup_lo_hi_504 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_505;
  assign dataGroup_lo_hi_505 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_506;
  assign dataGroup_lo_hi_506 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_507;
  assign dataGroup_lo_hi_507 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_508;
  assign dataGroup_lo_hi_508 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_509;
  assign dataGroup_lo_hi_509 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_510;
  assign dataGroup_lo_hi_510 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_511;
  assign dataGroup_lo_hi_511 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_512;
  assign dataGroup_lo_hi_512 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_513;
  assign dataGroup_lo_hi_513 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_514;
  assign dataGroup_lo_hi_514 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_515;
  assign dataGroup_lo_hi_515 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_516;
  assign dataGroup_lo_hi_516 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_517;
  assign dataGroup_lo_hi_517 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_518;
  assign dataGroup_lo_hi_518 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_519;
  assign dataGroup_lo_hi_519 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_520;
  assign dataGroup_lo_hi_520 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_521;
  assign dataGroup_lo_hi_521 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_522;
  assign dataGroup_lo_hi_522 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_523;
  assign dataGroup_lo_hi_523 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_524;
  assign dataGroup_lo_hi_524 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_525;
  assign dataGroup_lo_hi_525 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_526;
  assign dataGroup_lo_hi_526 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_527;
  assign dataGroup_lo_hi_527 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_528;
  assign dataGroup_lo_hi_528 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_529;
  assign dataGroup_lo_hi_529 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_530;
  assign dataGroup_lo_hi_530 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_531;
  assign dataGroup_lo_hi_531 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_532;
  assign dataGroup_lo_hi_532 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_533;
  assign dataGroup_lo_hi_533 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_534;
  assign dataGroup_lo_hi_534 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_535;
  assign dataGroup_lo_hi_535 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_536;
  assign dataGroup_lo_hi_536 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_537;
  assign dataGroup_lo_hi_537 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_538;
  assign dataGroup_lo_hi_538 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_539;
  assign dataGroup_lo_hi_539 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_540;
  assign dataGroup_lo_hi_540 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_541;
  assign dataGroup_lo_hi_541 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_542;
  assign dataGroup_lo_hi_542 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_543;
  assign dataGroup_lo_hi_543 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_544;
  assign dataGroup_lo_hi_544 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_545;
  assign dataGroup_lo_hi_545 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_546;
  assign dataGroup_lo_hi_546 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_547;
  assign dataGroup_lo_hi_547 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_548;
  assign dataGroup_lo_hi_548 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_549;
  assign dataGroup_lo_hi_549 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_550;
  assign dataGroup_lo_hi_550 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_551;
  assign dataGroup_lo_hi_551 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_552;
  assign dataGroup_lo_hi_552 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_553;
  assign dataGroup_lo_hi_553 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_554;
  assign dataGroup_lo_hi_554 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_555;
  assign dataGroup_lo_hi_555 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_556;
  assign dataGroup_lo_hi_556 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_557;
  assign dataGroup_lo_hi_557 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_558;
  assign dataGroup_lo_hi_558 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_559;
  assign dataGroup_lo_hi_559 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_560;
  assign dataGroup_lo_hi_560 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_561;
  assign dataGroup_lo_hi_561 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_562;
  assign dataGroup_lo_hi_562 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_563;
  assign dataGroup_lo_hi_563 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_564;
  assign dataGroup_lo_hi_564 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_565;
  assign dataGroup_lo_hi_565 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_566;
  assign dataGroup_lo_hi_566 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_567;
  assign dataGroup_lo_hi_567 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_568;
  assign dataGroup_lo_hi_568 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_569;
  assign dataGroup_lo_hi_569 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_570;
  assign dataGroup_lo_hi_570 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_571;
  assign dataGroup_lo_hi_571 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_572;
  assign dataGroup_lo_hi_572 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_573;
  assign dataGroup_lo_hi_573 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_574;
  assign dataGroup_lo_hi_574 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_575;
  assign dataGroup_lo_hi_575 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_576;
  assign dataGroup_lo_hi_576 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_577;
  assign dataGroup_lo_hi_577 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_578;
  assign dataGroup_lo_hi_578 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_579;
  assign dataGroup_lo_hi_579 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_580;
  assign dataGroup_lo_hi_580 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_581;
  assign dataGroup_lo_hi_581 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_582;
  assign dataGroup_lo_hi_582 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_583;
  assign dataGroup_lo_hi_583 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_584;
  assign dataGroup_lo_hi_584 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_585;
  assign dataGroup_lo_hi_585 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_586;
  assign dataGroup_lo_hi_586 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_587;
  assign dataGroup_lo_hi_587 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_588;
  assign dataGroup_lo_hi_588 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_589;
  assign dataGroup_lo_hi_589 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_590;
  assign dataGroup_lo_hi_590 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_591;
  assign dataGroup_lo_hi_591 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_592;
  assign dataGroup_lo_hi_592 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_593;
  assign dataGroup_lo_hi_593 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_594;
  assign dataGroup_lo_hi_594 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_595;
  assign dataGroup_lo_hi_595 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_596;
  assign dataGroup_lo_hi_596 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_597;
  assign dataGroup_lo_hi_597 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_598;
  assign dataGroup_lo_hi_598 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_599;
  assign dataGroup_lo_hi_599 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_600;
  assign dataGroup_lo_hi_600 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_601;
  assign dataGroup_lo_hi_601 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_602;
  assign dataGroup_lo_hi_602 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_603;
  assign dataGroup_lo_hi_603 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_604;
  assign dataGroup_lo_hi_604 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_605;
  assign dataGroup_lo_hi_605 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_606;
  assign dataGroup_lo_hi_606 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_607;
  assign dataGroup_lo_hi_607 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_608;
  assign dataGroup_lo_hi_608 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_609;
  assign dataGroup_lo_hi_609 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_610;
  assign dataGroup_lo_hi_610 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_611;
  assign dataGroup_lo_hi_611 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_612;
  assign dataGroup_lo_hi_612 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_613;
  assign dataGroup_lo_hi_613 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_614;
  assign dataGroup_lo_hi_614 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_615;
  assign dataGroup_lo_hi_615 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_616;
  assign dataGroup_lo_hi_616 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_617;
  assign dataGroup_lo_hi_617 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_618;
  assign dataGroup_lo_hi_618 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_619;
  assign dataGroup_lo_hi_619 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_620;
  assign dataGroup_lo_hi_620 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_621;
  assign dataGroup_lo_hi_621 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_622;
  assign dataGroup_lo_hi_622 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_623;
  assign dataGroup_lo_hi_623 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_624;
  assign dataGroup_lo_hi_624 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_625;
  assign dataGroup_lo_hi_625 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_626;
  assign dataGroup_lo_hi_626 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_627;
  assign dataGroup_lo_hi_627 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_628;
  assign dataGroup_lo_hi_628 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_629;
  assign dataGroup_lo_hi_629 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_630;
  assign dataGroup_lo_hi_630 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_631;
  assign dataGroup_lo_hi_631 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_632;
  assign dataGroup_lo_hi_632 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_633;
  assign dataGroup_lo_hi_633 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_634;
  assign dataGroup_lo_hi_634 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_635;
  assign dataGroup_lo_hi_635 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_636;
  assign dataGroup_lo_hi_636 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_637;
  assign dataGroup_lo_hi_637 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_638;
  assign dataGroup_lo_hi_638 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_639;
  assign dataGroup_lo_hi_639 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_640;
  assign dataGroup_lo_hi_640 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_641;
  assign dataGroup_lo_hi_641 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_642;
  assign dataGroup_lo_hi_642 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_643;
  assign dataGroup_lo_hi_643 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_644;
  assign dataGroup_lo_hi_644 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_645;
  assign dataGroup_lo_hi_645 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_646;
  assign dataGroup_lo_hi_646 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_647;
  assign dataGroup_lo_hi_647 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_648;
  assign dataGroup_lo_hi_648 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_649;
  assign dataGroup_lo_hi_649 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_650;
  assign dataGroup_lo_hi_650 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_651;
  assign dataGroup_lo_hi_651 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_652;
  assign dataGroup_lo_hi_652 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_653;
  assign dataGroup_lo_hi_653 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_654;
  assign dataGroup_lo_hi_654 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_655;
  assign dataGroup_lo_hi_655 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_656;
  assign dataGroup_lo_hi_656 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_657;
  assign dataGroup_lo_hi_657 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_658;
  assign dataGroup_lo_hi_658 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_659;
  assign dataGroup_lo_hi_659 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_660;
  assign dataGroup_lo_hi_660 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_661;
  assign dataGroup_lo_hi_661 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_662;
  assign dataGroup_lo_hi_662 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_663;
  assign dataGroup_lo_hi_663 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_664;
  assign dataGroup_lo_hi_664 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_665;
  assign dataGroup_lo_hi_665 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_666;
  assign dataGroup_lo_hi_666 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_667;
  assign dataGroup_lo_hi_667 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_668;
  assign dataGroup_lo_hi_668 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_669;
  assign dataGroup_lo_hi_669 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_670;
  assign dataGroup_lo_hi_670 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_671;
  assign dataGroup_lo_hi_671 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_672;
  assign dataGroup_lo_hi_672 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_673;
  assign dataGroup_lo_hi_673 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_674;
  assign dataGroup_lo_hi_674 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_675;
  assign dataGroup_lo_hi_675 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_676;
  assign dataGroup_lo_hi_676 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_677;
  assign dataGroup_lo_hi_677 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_678;
  assign dataGroup_lo_hi_678 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_679;
  assign dataGroup_lo_hi_679 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_680;
  assign dataGroup_lo_hi_680 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_681;
  assign dataGroup_lo_hi_681 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_682;
  assign dataGroup_lo_hi_682 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_683;
  assign dataGroup_lo_hi_683 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_684;
  assign dataGroup_lo_hi_684 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_685;
  assign dataGroup_lo_hi_685 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_686;
  assign dataGroup_lo_hi_686 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_687;
  assign dataGroup_lo_hi_687 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_688;
  assign dataGroup_lo_hi_688 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_689;
  assign dataGroup_lo_hi_689 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_690;
  assign dataGroup_lo_hi_690 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_691;
  assign dataGroup_lo_hi_691 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_692;
  assign dataGroup_lo_hi_692 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_693;
  assign dataGroup_lo_hi_693 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_694;
  assign dataGroup_lo_hi_694 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_695;
  assign dataGroup_lo_hi_695 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_696;
  assign dataGroup_lo_hi_696 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_697;
  assign dataGroup_lo_hi_697 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_698;
  assign dataGroup_lo_hi_698 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_699;
  assign dataGroup_lo_hi_699 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_700;
  assign dataGroup_lo_hi_700 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_701;
  assign dataGroup_lo_hi_701 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_702;
  assign dataGroup_lo_hi_702 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_703;
  assign dataGroup_lo_hi_703 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_704;
  assign dataGroup_lo_hi_704 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_705;
  assign dataGroup_lo_hi_705 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_706;
  assign dataGroup_lo_hi_706 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_707;
  assign dataGroup_lo_hi_707 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_708;
  assign dataGroup_lo_hi_708 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_709;
  assign dataGroup_lo_hi_709 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_710;
  assign dataGroup_lo_hi_710 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_711;
  assign dataGroup_lo_hi_711 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_712;
  assign dataGroup_lo_hi_712 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_713;
  assign dataGroup_lo_hi_713 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_714;
  assign dataGroup_lo_hi_714 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_715;
  assign dataGroup_lo_hi_715 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_716;
  assign dataGroup_lo_hi_716 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_717;
  assign dataGroup_lo_hi_717 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_718;
  assign dataGroup_lo_hi_718 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_719;
  assign dataGroup_lo_hi_719 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_720;
  assign dataGroup_lo_hi_720 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_721;
  assign dataGroup_lo_hi_721 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_722;
  assign dataGroup_lo_hi_722 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_723;
  assign dataGroup_lo_hi_723 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_724;
  assign dataGroup_lo_hi_724 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_725;
  assign dataGroup_lo_hi_725 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_726;
  assign dataGroup_lo_hi_726 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_727;
  assign dataGroup_lo_hi_727 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_728;
  assign dataGroup_lo_hi_728 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_729;
  assign dataGroup_lo_hi_729 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_730;
  assign dataGroup_lo_hi_730 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_731;
  assign dataGroup_lo_hi_731 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_732;
  assign dataGroup_lo_hi_732 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_733;
  assign dataGroup_lo_hi_733 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_734;
  assign dataGroup_lo_hi_734 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_735;
  assign dataGroup_lo_hi_735 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_736;
  assign dataGroup_lo_hi_736 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_737;
  assign dataGroup_lo_hi_737 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_738;
  assign dataGroup_lo_hi_738 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_739;
  assign dataGroup_lo_hi_739 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_740;
  assign dataGroup_lo_hi_740 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_741;
  assign dataGroup_lo_hi_741 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_742;
  assign dataGroup_lo_hi_742 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_743;
  assign dataGroup_lo_hi_743 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_744;
  assign dataGroup_lo_hi_744 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_745;
  assign dataGroup_lo_hi_745 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_746;
  assign dataGroup_lo_hi_746 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_747;
  assign dataGroup_lo_hi_747 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_748;
  assign dataGroup_lo_hi_748 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_749;
  assign dataGroup_lo_hi_749 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_750;
  assign dataGroup_lo_hi_750 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_751;
  assign dataGroup_lo_hi_751 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_752;
  assign dataGroup_lo_hi_752 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_753;
  assign dataGroup_lo_hi_753 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_754;
  assign dataGroup_lo_hi_754 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_755;
  assign dataGroup_lo_hi_755 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_756;
  assign dataGroup_lo_hi_756 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_757;
  assign dataGroup_lo_hi_757 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_758;
  assign dataGroup_lo_hi_758 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_759;
  assign dataGroup_lo_hi_759 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_760;
  assign dataGroup_lo_hi_760 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_761;
  assign dataGroup_lo_hi_761 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_762;
  assign dataGroup_lo_hi_762 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_763;
  assign dataGroup_lo_hi_763 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_764;
  assign dataGroup_lo_hi_764 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_765;
  assign dataGroup_lo_hi_765 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_766;
  assign dataGroup_lo_hi_766 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_767;
  assign dataGroup_lo_hi_767 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_768;
  assign dataGroup_lo_hi_768 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_769;
  assign dataGroup_lo_hi_769 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_770;
  assign dataGroup_lo_hi_770 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_771;
  assign dataGroup_lo_hi_771 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_772;
  assign dataGroup_lo_hi_772 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_773;
  assign dataGroup_lo_hi_773 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_774;
  assign dataGroup_lo_hi_774 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_775;
  assign dataGroup_lo_hi_775 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_776;
  assign dataGroup_lo_hi_776 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_777;
  assign dataGroup_lo_hi_777 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_778;
  assign dataGroup_lo_hi_778 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_779;
  assign dataGroup_lo_hi_779 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_780;
  assign dataGroup_lo_hi_780 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_781;
  assign dataGroup_lo_hi_781 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_782;
  assign dataGroup_lo_hi_782 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_783;
  assign dataGroup_lo_hi_783 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_784;
  assign dataGroup_lo_hi_784 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_785;
  assign dataGroup_lo_hi_785 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_786;
  assign dataGroup_lo_hi_786 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_787;
  assign dataGroup_lo_hi_787 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_788;
  assign dataGroup_lo_hi_788 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_789;
  assign dataGroup_lo_hi_789 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_790;
  assign dataGroup_lo_hi_790 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_791;
  assign dataGroup_lo_hi_791 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_792;
  assign dataGroup_lo_hi_792 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_793;
  assign dataGroup_lo_hi_793 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_794;
  assign dataGroup_lo_hi_794 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_795;
  assign dataGroup_lo_hi_795 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_796;
  assign dataGroup_lo_hi_796 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_797;
  assign dataGroup_lo_hi_797 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_798;
  assign dataGroup_lo_hi_798 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_799;
  assign dataGroup_lo_hi_799 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_800;
  assign dataGroup_lo_hi_800 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_801;
  assign dataGroup_lo_hi_801 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_802;
  assign dataGroup_lo_hi_802 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_803;
  assign dataGroup_lo_hi_803 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_804;
  assign dataGroup_lo_hi_804 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_805;
  assign dataGroup_lo_hi_805 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_806;
  assign dataGroup_lo_hi_806 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_807;
  assign dataGroup_lo_hi_807 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_808;
  assign dataGroup_lo_hi_808 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_809;
  assign dataGroup_lo_hi_809 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_810;
  assign dataGroup_lo_hi_810 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_811;
  assign dataGroup_lo_hi_811 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_812;
  assign dataGroup_lo_hi_812 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_813;
  assign dataGroup_lo_hi_813 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_814;
  assign dataGroup_lo_hi_814 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_815;
  assign dataGroup_lo_hi_815 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_816;
  assign dataGroup_lo_hi_816 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_817;
  assign dataGroup_lo_hi_817 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_818;
  assign dataGroup_lo_hi_818 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_819;
  assign dataGroup_lo_hi_819 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_820;
  assign dataGroup_lo_hi_820 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_821;
  assign dataGroup_lo_hi_821 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_822;
  assign dataGroup_lo_hi_822 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_823;
  assign dataGroup_lo_hi_823 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_824;
  assign dataGroup_lo_hi_824 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_825;
  assign dataGroup_lo_hi_825 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_826;
  assign dataGroup_lo_hi_826 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_827;
  assign dataGroup_lo_hi_827 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_828;
  assign dataGroup_lo_hi_828 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_829;
  assign dataGroup_lo_hi_829 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_830;
  assign dataGroup_lo_hi_830 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_831;
  assign dataGroup_lo_hi_831 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_832;
  assign dataGroup_lo_hi_832 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_833;
  assign dataGroup_lo_hi_833 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_834;
  assign dataGroup_lo_hi_834 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_835;
  assign dataGroup_lo_hi_835 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_836;
  assign dataGroup_lo_hi_836 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_837;
  assign dataGroup_lo_hi_837 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_838;
  assign dataGroup_lo_hi_838 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_839;
  assign dataGroup_lo_hi_839 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_840;
  assign dataGroup_lo_hi_840 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_841;
  assign dataGroup_lo_hi_841 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_842;
  assign dataGroup_lo_hi_842 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_843;
  assign dataGroup_lo_hi_843 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_844;
  assign dataGroup_lo_hi_844 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_845;
  assign dataGroup_lo_hi_845 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_846;
  assign dataGroup_lo_hi_846 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_847;
  assign dataGroup_lo_hi_847 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_848;
  assign dataGroup_lo_hi_848 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_849;
  assign dataGroup_lo_hi_849 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_850;
  assign dataGroup_lo_hi_850 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_851;
  assign dataGroup_lo_hi_851 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_852;
  assign dataGroup_lo_hi_852 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_853;
  assign dataGroup_lo_hi_853 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_854;
  assign dataGroup_lo_hi_854 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_855;
  assign dataGroup_lo_hi_855 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_856;
  assign dataGroup_lo_hi_856 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_857;
  assign dataGroup_lo_hi_857 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_858;
  assign dataGroup_lo_hi_858 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_859;
  assign dataGroup_lo_hi_859 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_860;
  assign dataGroup_lo_hi_860 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_861;
  assign dataGroup_lo_hi_861 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_862;
  assign dataGroup_lo_hi_862 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_863;
  assign dataGroup_lo_hi_863 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_864;
  assign dataGroup_lo_hi_864 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_865;
  assign dataGroup_lo_hi_865 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_866;
  assign dataGroup_lo_hi_866 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_867;
  assign dataGroup_lo_hi_867 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_868;
  assign dataGroup_lo_hi_868 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_869;
  assign dataGroup_lo_hi_869 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_870;
  assign dataGroup_lo_hi_870 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_871;
  assign dataGroup_lo_hi_871 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_872;
  assign dataGroup_lo_hi_872 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_873;
  assign dataGroup_lo_hi_873 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_874;
  assign dataGroup_lo_hi_874 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_875;
  assign dataGroup_lo_hi_875 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_876;
  assign dataGroup_lo_hi_876 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_877;
  assign dataGroup_lo_hi_877 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_878;
  assign dataGroup_lo_hi_878 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_879;
  assign dataGroup_lo_hi_879 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_880;
  assign dataGroup_lo_hi_880 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_881;
  assign dataGroup_lo_hi_881 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_882;
  assign dataGroup_lo_hi_882 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_883;
  assign dataGroup_lo_hi_883 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_884;
  assign dataGroup_lo_hi_884 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_885;
  assign dataGroup_lo_hi_885 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_886;
  assign dataGroup_lo_hi_886 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_887;
  assign dataGroup_lo_hi_887 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_888;
  assign dataGroup_lo_hi_888 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_889;
  assign dataGroup_lo_hi_889 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_890;
  assign dataGroup_lo_hi_890 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_891;
  assign dataGroup_lo_hi_891 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_892;
  assign dataGroup_lo_hi_892 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_893;
  assign dataGroup_lo_hi_893 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_894;
  assign dataGroup_lo_hi_894 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_895;
  assign dataGroup_lo_hi_895 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_896;
  assign dataGroup_lo_hi_896 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_897;
  assign dataGroup_lo_hi_897 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_898;
  assign dataGroup_lo_hi_898 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_899;
  assign dataGroup_lo_hi_899 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_900;
  assign dataGroup_lo_hi_900 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_901;
  assign dataGroup_lo_hi_901 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_902;
  assign dataGroup_lo_hi_902 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_903;
  assign dataGroup_lo_hi_903 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_904;
  assign dataGroup_lo_hi_904 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_905;
  assign dataGroup_lo_hi_905 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_906;
  assign dataGroup_lo_hi_906 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_907;
  assign dataGroup_lo_hi_907 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_908;
  assign dataGroup_lo_hi_908 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_909;
  assign dataGroup_lo_hi_909 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_910;
  assign dataGroup_lo_hi_910 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_911;
  assign dataGroup_lo_hi_911 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_912;
  assign dataGroup_lo_hi_912 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_913;
  assign dataGroup_lo_hi_913 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_914;
  assign dataGroup_lo_hi_914 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_915;
  assign dataGroup_lo_hi_915 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_916;
  assign dataGroup_lo_hi_916 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_917;
  assign dataGroup_lo_hi_917 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_918;
  assign dataGroup_lo_hi_918 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_919;
  assign dataGroup_lo_hi_919 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_920;
  assign dataGroup_lo_hi_920 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_921;
  assign dataGroup_lo_hi_921 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_922;
  assign dataGroup_lo_hi_922 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_923;
  assign dataGroup_lo_hi_923 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_924;
  assign dataGroup_lo_hi_924 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_925;
  assign dataGroup_lo_hi_925 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_926;
  assign dataGroup_lo_hi_926 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_927;
  assign dataGroup_lo_hi_927 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_928;
  assign dataGroup_lo_hi_928 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_929;
  assign dataGroup_lo_hi_929 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_930;
  assign dataGroup_lo_hi_930 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_931;
  assign dataGroup_lo_hi_931 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_932;
  assign dataGroup_lo_hi_932 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_933;
  assign dataGroup_lo_hi_933 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_934;
  assign dataGroup_lo_hi_934 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_935;
  assign dataGroup_lo_hi_935 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_936;
  assign dataGroup_lo_hi_936 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_937;
  assign dataGroup_lo_hi_937 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_938;
  assign dataGroup_lo_hi_938 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_939;
  assign dataGroup_lo_hi_939 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_940;
  assign dataGroup_lo_hi_940 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_941;
  assign dataGroup_lo_hi_941 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_942;
  assign dataGroup_lo_hi_942 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_943;
  assign dataGroup_lo_hi_943 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_944;
  assign dataGroup_lo_hi_944 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_945;
  assign dataGroup_lo_hi_945 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_946;
  assign dataGroup_lo_hi_946 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_947;
  assign dataGroup_lo_hi_947 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_948;
  assign dataGroup_lo_hi_948 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_949;
  assign dataGroup_lo_hi_949 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_950;
  assign dataGroup_lo_hi_950 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_951;
  assign dataGroup_lo_hi_951 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_952;
  assign dataGroup_lo_hi_952 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_953;
  assign dataGroup_lo_hi_953 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_954;
  assign dataGroup_lo_hi_954 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_955;
  assign dataGroup_lo_hi_955 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_956;
  assign dataGroup_lo_hi_956 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_957;
  assign dataGroup_lo_hi_957 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_958;
  assign dataGroup_lo_hi_958 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_959;
  assign dataGroup_lo_hi_959 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_960;
  assign dataGroup_lo_hi_960 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_961;
  assign dataGroup_lo_hi_961 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_962;
  assign dataGroup_lo_hi_962 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_963;
  assign dataGroup_lo_hi_963 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_964;
  assign dataGroup_lo_hi_964 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_965;
  assign dataGroup_lo_hi_965 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_966;
  assign dataGroup_lo_hi_966 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_967;
  assign dataGroup_lo_hi_967 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_968;
  assign dataGroup_lo_hi_968 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_969;
  assign dataGroup_lo_hi_969 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_970;
  assign dataGroup_lo_hi_970 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_971;
  assign dataGroup_lo_hi_971 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_972;
  assign dataGroup_lo_hi_972 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_973;
  assign dataGroup_lo_hi_973 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_974;
  assign dataGroup_lo_hi_974 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_975;
  assign dataGroup_lo_hi_975 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_976;
  assign dataGroup_lo_hi_976 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_977;
  assign dataGroup_lo_hi_977 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_978;
  assign dataGroup_lo_hi_978 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_979;
  assign dataGroup_lo_hi_979 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_980;
  assign dataGroup_lo_hi_980 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_981;
  assign dataGroup_lo_hi_981 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_982;
  assign dataGroup_lo_hi_982 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_983;
  assign dataGroup_lo_hi_983 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_984;
  assign dataGroup_lo_hi_984 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_985;
  assign dataGroup_lo_hi_985 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_986;
  assign dataGroup_lo_hi_986 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_987;
  assign dataGroup_lo_hi_987 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_988;
  assign dataGroup_lo_hi_988 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_989;
  assign dataGroup_lo_hi_989 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_990;
  assign dataGroup_lo_hi_990 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_991;
  assign dataGroup_lo_hi_991 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_992;
  assign dataGroup_lo_hi_992 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_993;
  assign dataGroup_lo_hi_993 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_994;
  assign dataGroup_lo_hi_994 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_995;
  assign dataGroup_lo_hi_995 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_996;
  assign dataGroup_lo_hi_996 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_997;
  assign dataGroup_lo_hi_997 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_998;
  assign dataGroup_lo_hi_998 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_999;
  assign dataGroup_lo_hi_999 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1000;
  assign dataGroup_lo_hi_1000 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1001;
  assign dataGroup_lo_hi_1001 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1002;
  assign dataGroup_lo_hi_1002 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1003;
  assign dataGroup_lo_hi_1003 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1004;
  assign dataGroup_lo_hi_1004 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1005;
  assign dataGroup_lo_hi_1005 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1006;
  assign dataGroup_lo_hi_1006 = _GEN_4;
  wire [255:0]  dataGroup_lo_hi_1007;
  assign dataGroup_lo_hi_1007 = _GEN_4;
  wire [511:0]  dataGroup_lo = {dataGroup_lo_hi, dataGroup_lo_lo};
  wire [255:0]  _GEN_5 = {dataSelect_5, dataSelect_4};
  wire [255:0]  dataGroup_hi_lo;
  assign dataGroup_hi_lo = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1;
  assign dataGroup_hi_lo_1 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_2;
  assign dataGroup_hi_lo_2 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_3;
  assign dataGroup_hi_lo_3 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_4;
  assign dataGroup_hi_lo_4 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_5;
  assign dataGroup_hi_lo_5 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_6;
  assign dataGroup_hi_lo_6 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_7;
  assign dataGroup_hi_lo_7 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_8;
  assign dataGroup_hi_lo_8 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_9;
  assign dataGroup_hi_lo_9 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_10;
  assign dataGroup_hi_lo_10 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_11;
  assign dataGroup_hi_lo_11 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_12;
  assign dataGroup_hi_lo_12 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_13;
  assign dataGroup_hi_lo_13 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_14;
  assign dataGroup_hi_lo_14 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_15;
  assign dataGroup_hi_lo_15 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_16;
  assign dataGroup_hi_lo_16 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_17;
  assign dataGroup_hi_lo_17 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_18;
  assign dataGroup_hi_lo_18 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_19;
  assign dataGroup_hi_lo_19 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_20;
  assign dataGroup_hi_lo_20 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_21;
  assign dataGroup_hi_lo_21 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_22;
  assign dataGroup_hi_lo_22 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_23;
  assign dataGroup_hi_lo_23 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_24;
  assign dataGroup_hi_lo_24 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_25;
  assign dataGroup_hi_lo_25 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_26;
  assign dataGroup_hi_lo_26 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_27;
  assign dataGroup_hi_lo_27 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_28;
  assign dataGroup_hi_lo_28 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_29;
  assign dataGroup_hi_lo_29 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_30;
  assign dataGroup_hi_lo_30 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_31;
  assign dataGroup_hi_lo_31 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_32;
  assign dataGroup_hi_lo_32 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_33;
  assign dataGroup_hi_lo_33 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_34;
  assign dataGroup_hi_lo_34 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_35;
  assign dataGroup_hi_lo_35 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_36;
  assign dataGroup_hi_lo_36 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_37;
  assign dataGroup_hi_lo_37 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_38;
  assign dataGroup_hi_lo_38 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_39;
  assign dataGroup_hi_lo_39 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_40;
  assign dataGroup_hi_lo_40 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_41;
  assign dataGroup_hi_lo_41 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_42;
  assign dataGroup_hi_lo_42 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_43;
  assign dataGroup_hi_lo_43 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_44;
  assign dataGroup_hi_lo_44 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_45;
  assign dataGroup_hi_lo_45 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_46;
  assign dataGroup_hi_lo_46 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_47;
  assign dataGroup_hi_lo_47 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_48;
  assign dataGroup_hi_lo_48 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_49;
  assign dataGroup_hi_lo_49 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_50;
  assign dataGroup_hi_lo_50 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_51;
  assign dataGroup_hi_lo_51 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_52;
  assign dataGroup_hi_lo_52 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_53;
  assign dataGroup_hi_lo_53 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_54;
  assign dataGroup_hi_lo_54 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_55;
  assign dataGroup_hi_lo_55 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_56;
  assign dataGroup_hi_lo_56 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_57;
  assign dataGroup_hi_lo_57 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_58;
  assign dataGroup_hi_lo_58 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_59;
  assign dataGroup_hi_lo_59 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_60;
  assign dataGroup_hi_lo_60 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_61;
  assign dataGroup_hi_lo_61 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_62;
  assign dataGroup_hi_lo_62 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_63;
  assign dataGroup_hi_lo_63 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_64;
  assign dataGroup_hi_lo_64 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_65;
  assign dataGroup_hi_lo_65 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_66;
  assign dataGroup_hi_lo_66 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_67;
  assign dataGroup_hi_lo_67 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_68;
  assign dataGroup_hi_lo_68 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_69;
  assign dataGroup_hi_lo_69 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_70;
  assign dataGroup_hi_lo_70 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_71;
  assign dataGroup_hi_lo_71 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_72;
  assign dataGroup_hi_lo_72 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_73;
  assign dataGroup_hi_lo_73 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_74;
  assign dataGroup_hi_lo_74 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_75;
  assign dataGroup_hi_lo_75 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_76;
  assign dataGroup_hi_lo_76 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_77;
  assign dataGroup_hi_lo_77 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_78;
  assign dataGroup_hi_lo_78 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_79;
  assign dataGroup_hi_lo_79 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_80;
  assign dataGroup_hi_lo_80 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_81;
  assign dataGroup_hi_lo_81 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_82;
  assign dataGroup_hi_lo_82 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_83;
  assign dataGroup_hi_lo_83 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_84;
  assign dataGroup_hi_lo_84 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_85;
  assign dataGroup_hi_lo_85 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_86;
  assign dataGroup_hi_lo_86 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_87;
  assign dataGroup_hi_lo_87 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_88;
  assign dataGroup_hi_lo_88 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_89;
  assign dataGroup_hi_lo_89 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_90;
  assign dataGroup_hi_lo_90 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_91;
  assign dataGroup_hi_lo_91 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_92;
  assign dataGroup_hi_lo_92 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_93;
  assign dataGroup_hi_lo_93 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_94;
  assign dataGroup_hi_lo_94 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_95;
  assign dataGroup_hi_lo_95 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_96;
  assign dataGroup_hi_lo_96 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_97;
  assign dataGroup_hi_lo_97 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_98;
  assign dataGroup_hi_lo_98 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_99;
  assign dataGroup_hi_lo_99 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_100;
  assign dataGroup_hi_lo_100 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_101;
  assign dataGroup_hi_lo_101 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_102;
  assign dataGroup_hi_lo_102 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_103;
  assign dataGroup_hi_lo_103 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_104;
  assign dataGroup_hi_lo_104 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_105;
  assign dataGroup_hi_lo_105 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_106;
  assign dataGroup_hi_lo_106 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_107;
  assign dataGroup_hi_lo_107 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_108;
  assign dataGroup_hi_lo_108 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_109;
  assign dataGroup_hi_lo_109 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_110;
  assign dataGroup_hi_lo_110 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_111;
  assign dataGroup_hi_lo_111 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_112;
  assign dataGroup_hi_lo_112 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_113;
  assign dataGroup_hi_lo_113 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_114;
  assign dataGroup_hi_lo_114 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_115;
  assign dataGroup_hi_lo_115 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_116;
  assign dataGroup_hi_lo_116 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_117;
  assign dataGroup_hi_lo_117 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_118;
  assign dataGroup_hi_lo_118 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_119;
  assign dataGroup_hi_lo_119 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_120;
  assign dataGroup_hi_lo_120 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_121;
  assign dataGroup_hi_lo_121 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_122;
  assign dataGroup_hi_lo_122 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_123;
  assign dataGroup_hi_lo_123 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_124;
  assign dataGroup_hi_lo_124 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_125;
  assign dataGroup_hi_lo_125 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_126;
  assign dataGroup_hi_lo_126 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_127;
  assign dataGroup_hi_lo_127 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_128;
  assign dataGroup_hi_lo_128 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_129;
  assign dataGroup_hi_lo_129 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_130;
  assign dataGroup_hi_lo_130 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_131;
  assign dataGroup_hi_lo_131 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_132;
  assign dataGroup_hi_lo_132 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_133;
  assign dataGroup_hi_lo_133 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_134;
  assign dataGroup_hi_lo_134 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_135;
  assign dataGroup_hi_lo_135 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_136;
  assign dataGroup_hi_lo_136 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_137;
  assign dataGroup_hi_lo_137 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_138;
  assign dataGroup_hi_lo_138 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_139;
  assign dataGroup_hi_lo_139 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_140;
  assign dataGroup_hi_lo_140 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_141;
  assign dataGroup_hi_lo_141 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_142;
  assign dataGroup_hi_lo_142 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_143;
  assign dataGroup_hi_lo_143 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_144;
  assign dataGroup_hi_lo_144 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_145;
  assign dataGroup_hi_lo_145 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_146;
  assign dataGroup_hi_lo_146 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_147;
  assign dataGroup_hi_lo_147 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_148;
  assign dataGroup_hi_lo_148 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_149;
  assign dataGroup_hi_lo_149 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_150;
  assign dataGroup_hi_lo_150 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_151;
  assign dataGroup_hi_lo_151 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_152;
  assign dataGroup_hi_lo_152 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_153;
  assign dataGroup_hi_lo_153 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_154;
  assign dataGroup_hi_lo_154 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_155;
  assign dataGroup_hi_lo_155 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_156;
  assign dataGroup_hi_lo_156 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_157;
  assign dataGroup_hi_lo_157 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_158;
  assign dataGroup_hi_lo_158 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_159;
  assign dataGroup_hi_lo_159 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_160;
  assign dataGroup_hi_lo_160 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_161;
  assign dataGroup_hi_lo_161 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_162;
  assign dataGroup_hi_lo_162 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_163;
  assign dataGroup_hi_lo_163 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_164;
  assign dataGroup_hi_lo_164 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_165;
  assign dataGroup_hi_lo_165 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_166;
  assign dataGroup_hi_lo_166 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_167;
  assign dataGroup_hi_lo_167 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_168;
  assign dataGroup_hi_lo_168 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_169;
  assign dataGroup_hi_lo_169 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_170;
  assign dataGroup_hi_lo_170 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_171;
  assign dataGroup_hi_lo_171 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_172;
  assign dataGroup_hi_lo_172 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_173;
  assign dataGroup_hi_lo_173 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_174;
  assign dataGroup_hi_lo_174 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_175;
  assign dataGroup_hi_lo_175 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_176;
  assign dataGroup_hi_lo_176 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_177;
  assign dataGroup_hi_lo_177 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_178;
  assign dataGroup_hi_lo_178 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_179;
  assign dataGroup_hi_lo_179 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_180;
  assign dataGroup_hi_lo_180 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_181;
  assign dataGroup_hi_lo_181 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_182;
  assign dataGroup_hi_lo_182 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_183;
  assign dataGroup_hi_lo_183 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_184;
  assign dataGroup_hi_lo_184 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_185;
  assign dataGroup_hi_lo_185 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_186;
  assign dataGroup_hi_lo_186 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_187;
  assign dataGroup_hi_lo_187 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_188;
  assign dataGroup_hi_lo_188 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_189;
  assign dataGroup_hi_lo_189 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_190;
  assign dataGroup_hi_lo_190 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_191;
  assign dataGroup_hi_lo_191 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_192;
  assign dataGroup_hi_lo_192 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_193;
  assign dataGroup_hi_lo_193 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_194;
  assign dataGroup_hi_lo_194 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_195;
  assign dataGroup_hi_lo_195 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_196;
  assign dataGroup_hi_lo_196 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_197;
  assign dataGroup_hi_lo_197 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_198;
  assign dataGroup_hi_lo_198 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_199;
  assign dataGroup_hi_lo_199 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_200;
  assign dataGroup_hi_lo_200 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_201;
  assign dataGroup_hi_lo_201 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_202;
  assign dataGroup_hi_lo_202 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_203;
  assign dataGroup_hi_lo_203 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_204;
  assign dataGroup_hi_lo_204 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_205;
  assign dataGroup_hi_lo_205 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_206;
  assign dataGroup_hi_lo_206 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_207;
  assign dataGroup_hi_lo_207 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_208;
  assign dataGroup_hi_lo_208 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_209;
  assign dataGroup_hi_lo_209 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_210;
  assign dataGroup_hi_lo_210 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_211;
  assign dataGroup_hi_lo_211 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_212;
  assign dataGroup_hi_lo_212 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_213;
  assign dataGroup_hi_lo_213 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_214;
  assign dataGroup_hi_lo_214 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_215;
  assign dataGroup_hi_lo_215 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_216;
  assign dataGroup_hi_lo_216 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_217;
  assign dataGroup_hi_lo_217 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_218;
  assign dataGroup_hi_lo_218 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_219;
  assign dataGroup_hi_lo_219 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_220;
  assign dataGroup_hi_lo_220 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_221;
  assign dataGroup_hi_lo_221 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_222;
  assign dataGroup_hi_lo_222 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_223;
  assign dataGroup_hi_lo_223 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_224;
  assign dataGroup_hi_lo_224 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_225;
  assign dataGroup_hi_lo_225 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_226;
  assign dataGroup_hi_lo_226 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_227;
  assign dataGroup_hi_lo_227 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_228;
  assign dataGroup_hi_lo_228 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_229;
  assign dataGroup_hi_lo_229 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_230;
  assign dataGroup_hi_lo_230 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_231;
  assign dataGroup_hi_lo_231 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_232;
  assign dataGroup_hi_lo_232 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_233;
  assign dataGroup_hi_lo_233 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_234;
  assign dataGroup_hi_lo_234 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_235;
  assign dataGroup_hi_lo_235 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_236;
  assign dataGroup_hi_lo_236 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_237;
  assign dataGroup_hi_lo_237 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_238;
  assign dataGroup_hi_lo_238 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_239;
  assign dataGroup_hi_lo_239 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_240;
  assign dataGroup_hi_lo_240 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_241;
  assign dataGroup_hi_lo_241 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_242;
  assign dataGroup_hi_lo_242 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_243;
  assign dataGroup_hi_lo_243 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_244;
  assign dataGroup_hi_lo_244 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_245;
  assign dataGroup_hi_lo_245 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_246;
  assign dataGroup_hi_lo_246 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_247;
  assign dataGroup_hi_lo_247 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_248;
  assign dataGroup_hi_lo_248 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_249;
  assign dataGroup_hi_lo_249 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_250;
  assign dataGroup_hi_lo_250 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_251;
  assign dataGroup_hi_lo_251 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_252;
  assign dataGroup_hi_lo_252 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_253;
  assign dataGroup_hi_lo_253 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_254;
  assign dataGroup_hi_lo_254 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_255;
  assign dataGroup_hi_lo_255 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_256;
  assign dataGroup_hi_lo_256 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_257;
  assign dataGroup_hi_lo_257 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_258;
  assign dataGroup_hi_lo_258 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_259;
  assign dataGroup_hi_lo_259 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_260;
  assign dataGroup_hi_lo_260 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_261;
  assign dataGroup_hi_lo_261 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_262;
  assign dataGroup_hi_lo_262 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_263;
  assign dataGroup_hi_lo_263 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_264;
  assign dataGroup_hi_lo_264 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_265;
  assign dataGroup_hi_lo_265 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_266;
  assign dataGroup_hi_lo_266 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_267;
  assign dataGroup_hi_lo_267 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_268;
  assign dataGroup_hi_lo_268 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_269;
  assign dataGroup_hi_lo_269 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_270;
  assign dataGroup_hi_lo_270 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_271;
  assign dataGroup_hi_lo_271 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_272;
  assign dataGroup_hi_lo_272 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_273;
  assign dataGroup_hi_lo_273 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_274;
  assign dataGroup_hi_lo_274 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_275;
  assign dataGroup_hi_lo_275 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_276;
  assign dataGroup_hi_lo_276 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_277;
  assign dataGroup_hi_lo_277 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_278;
  assign dataGroup_hi_lo_278 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_279;
  assign dataGroup_hi_lo_279 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_280;
  assign dataGroup_hi_lo_280 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_281;
  assign dataGroup_hi_lo_281 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_282;
  assign dataGroup_hi_lo_282 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_283;
  assign dataGroup_hi_lo_283 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_284;
  assign dataGroup_hi_lo_284 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_285;
  assign dataGroup_hi_lo_285 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_286;
  assign dataGroup_hi_lo_286 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_287;
  assign dataGroup_hi_lo_287 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_288;
  assign dataGroup_hi_lo_288 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_289;
  assign dataGroup_hi_lo_289 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_290;
  assign dataGroup_hi_lo_290 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_291;
  assign dataGroup_hi_lo_291 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_292;
  assign dataGroup_hi_lo_292 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_293;
  assign dataGroup_hi_lo_293 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_294;
  assign dataGroup_hi_lo_294 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_295;
  assign dataGroup_hi_lo_295 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_296;
  assign dataGroup_hi_lo_296 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_297;
  assign dataGroup_hi_lo_297 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_298;
  assign dataGroup_hi_lo_298 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_299;
  assign dataGroup_hi_lo_299 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_300;
  assign dataGroup_hi_lo_300 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_301;
  assign dataGroup_hi_lo_301 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_302;
  assign dataGroup_hi_lo_302 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_303;
  assign dataGroup_hi_lo_303 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_304;
  assign dataGroup_hi_lo_304 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_305;
  assign dataGroup_hi_lo_305 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_306;
  assign dataGroup_hi_lo_306 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_307;
  assign dataGroup_hi_lo_307 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_308;
  assign dataGroup_hi_lo_308 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_309;
  assign dataGroup_hi_lo_309 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_310;
  assign dataGroup_hi_lo_310 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_311;
  assign dataGroup_hi_lo_311 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_312;
  assign dataGroup_hi_lo_312 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_313;
  assign dataGroup_hi_lo_313 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_314;
  assign dataGroup_hi_lo_314 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_315;
  assign dataGroup_hi_lo_315 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_316;
  assign dataGroup_hi_lo_316 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_317;
  assign dataGroup_hi_lo_317 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_318;
  assign dataGroup_hi_lo_318 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_319;
  assign dataGroup_hi_lo_319 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_320;
  assign dataGroup_hi_lo_320 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_321;
  assign dataGroup_hi_lo_321 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_322;
  assign dataGroup_hi_lo_322 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_323;
  assign dataGroup_hi_lo_323 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_324;
  assign dataGroup_hi_lo_324 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_325;
  assign dataGroup_hi_lo_325 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_326;
  assign dataGroup_hi_lo_326 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_327;
  assign dataGroup_hi_lo_327 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_328;
  assign dataGroup_hi_lo_328 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_329;
  assign dataGroup_hi_lo_329 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_330;
  assign dataGroup_hi_lo_330 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_331;
  assign dataGroup_hi_lo_331 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_332;
  assign dataGroup_hi_lo_332 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_333;
  assign dataGroup_hi_lo_333 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_334;
  assign dataGroup_hi_lo_334 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_335;
  assign dataGroup_hi_lo_335 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_336;
  assign dataGroup_hi_lo_336 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_337;
  assign dataGroup_hi_lo_337 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_338;
  assign dataGroup_hi_lo_338 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_339;
  assign dataGroup_hi_lo_339 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_340;
  assign dataGroup_hi_lo_340 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_341;
  assign dataGroup_hi_lo_341 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_342;
  assign dataGroup_hi_lo_342 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_343;
  assign dataGroup_hi_lo_343 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_344;
  assign dataGroup_hi_lo_344 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_345;
  assign dataGroup_hi_lo_345 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_346;
  assign dataGroup_hi_lo_346 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_347;
  assign dataGroup_hi_lo_347 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_348;
  assign dataGroup_hi_lo_348 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_349;
  assign dataGroup_hi_lo_349 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_350;
  assign dataGroup_hi_lo_350 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_351;
  assign dataGroup_hi_lo_351 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_352;
  assign dataGroup_hi_lo_352 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_353;
  assign dataGroup_hi_lo_353 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_354;
  assign dataGroup_hi_lo_354 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_355;
  assign dataGroup_hi_lo_355 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_356;
  assign dataGroup_hi_lo_356 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_357;
  assign dataGroup_hi_lo_357 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_358;
  assign dataGroup_hi_lo_358 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_359;
  assign dataGroup_hi_lo_359 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_360;
  assign dataGroup_hi_lo_360 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_361;
  assign dataGroup_hi_lo_361 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_362;
  assign dataGroup_hi_lo_362 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_363;
  assign dataGroup_hi_lo_363 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_364;
  assign dataGroup_hi_lo_364 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_365;
  assign dataGroup_hi_lo_365 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_366;
  assign dataGroup_hi_lo_366 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_367;
  assign dataGroup_hi_lo_367 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_368;
  assign dataGroup_hi_lo_368 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_369;
  assign dataGroup_hi_lo_369 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_370;
  assign dataGroup_hi_lo_370 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_371;
  assign dataGroup_hi_lo_371 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_372;
  assign dataGroup_hi_lo_372 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_373;
  assign dataGroup_hi_lo_373 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_374;
  assign dataGroup_hi_lo_374 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_375;
  assign dataGroup_hi_lo_375 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_376;
  assign dataGroup_hi_lo_376 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_377;
  assign dataGroup_hi_lo_377 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_378;
  assign dataGroup_hi_lo_378 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_379;
  assign dataGroup_hi_lo_379 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_380;
  assign dataGroup_hi_lo_380 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_381;
  assign dataGroup_hi_lo_381 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_382;
  assign dataGroup_hi_lo_382 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_383;
  assign dataGroup_hi_lo_383 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_384;
  assign dataGroup_hi_lo_384 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_385;
  assign dataGroup_hi_lo_385 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_386;
  assign dataGroup_hi_lo_386 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_387;
  assign dataGroup_hi_lo_387 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_388;
  assign dataGroup_hi_lo_388 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_389;
  assign dataGroup_hi_lo_389 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_390;
  assign dataGroup_hi_lo_390 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_391;
  assign dataGroup_hi_lo_391 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_392;
  assign dataGroup_hi_lo_392 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_393;
  assign dataGroup_hi_lo_393 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_394;
  assign dataGroup_hi_lo_394 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_395;
  assign dataGroup_hi_lo_395 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_396;
  assign dataGroup_hi_lo_396 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_397;
  assign dataGroup_hi_lo_397 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_398;
  assign dataGroup_hi_lo_398 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_399;
  assign dataGroup_hi_lo_399 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_400;
  assign dataGroup_hi_lo_400 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_401;
  assign dataGroup_hi_lo_401 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_402;
  assign dataGroup_hi_lo_402 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_403;
  assign dataGroup_hi_lo_403 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_404;
  assign dataGroup_hi_lo_404 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_405;
  assign dataGroup_hi_lo_405 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_406;
  assign dataGroup_hi_lo_406 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_407;
  assign dataGroup_hi_lo_407 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_408;
  assign dataGroup_hi_lo_408 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_409;
  assign dataGroup_hi_lo_409 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_410;
  assign dataGroup_hi_lo_410 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_411;
  assign dataGroup_hi_lo_411 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_412;
  assign dataGroup_hi_lo_412 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_413;
  assign dataGroup_hi_lo_413 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_414;
  assign dataGroup_hi_lo_414 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_415;
  assign dataGroup_hi_lo_415 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_416;
  assign dataGroup_hi_lo_416 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_417;
  assign dataGroup_hi_lo_417 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_418;
  assign dataGroup_hi_lo_418 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_419;
  assign dataGroup_hi_lo_419 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_420;
  assign dataGroup_hi_lo_420 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_421;
  assign dataGroup_hi_lo_421 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_422;
  assign dataGroup_hi_lo_422 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_423;
  assign dataGroup_hi_lo_423 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_424;
  assign dataGroup_hi_lo_424 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_425;
  assign dataGroup_hi_lo_425 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_426;
  assign dataGroup_hi_lo_426 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_427;
  assign dataGroup_hi_lo_427 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_428;
  assign dataGroup_hi_lo_428 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_429;
  assign dataGroup_hi_lo_429 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_430;
  assign dataGroup_hi_lo_430 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_431;
  assign dataGroup_hi_lo_431 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_432;
  assign dataGroup_hi_lo_432 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_433;
  assign dataGroup_hi_lo_433 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_434;
  assign dataGroup_hi_lo_434 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_435;
  assign dataGroup_hi_lo_435 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_436;
  assign dataGroup_hi_lo_436 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_437;
  assign dataGroup_hi_lo_437 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_438;
  assign dataGroup_hi_lo_438 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_439;
  assign dataGroup_hi_lo_439 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_440;
  assign dataGroup_hi_lo_440 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_441;
  assign dataGroup_hi_lo_441 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_442;
  assign dataGroup_hi_lo_442 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_443;
  assign dataGroup_hi_lo_443 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_444;
  assign dataGroup_hi_lo_444 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_445;
  assign dataGroup_hi_lo_445 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_446;
  assign dataGroup_hi_lo_446 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_447;
  assign dataGroup_hi_lo_447 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_448;
  assign dataGroup_hi_lo_448 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_449;
  assign dataGroup_hi_lo_449 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_450;
  assign dataGroup_hi_lo_450 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_451;
  assign dataGroup_hi_lo_451 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_452;
  assign dataGroup_hi_lo_452 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_453;
  assign dataGroup_hi_lo_453 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_454;
  assign dataGroup_hi_lo_454 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_455;
  assign dataGroup_hi_lo_455 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_456;
  assign dataGroup_hi_lo_456 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_457;
  assign dataGroup_hi_lo_457 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_458;
  assign dataGroup_hi_lo_458 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_459;
  assign dataGroup_hi_lo_459 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_460;
  assign dataGroup_hi_lo_460 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_461;
  assign dataGroup_hi_lo_461 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_462;
  assign dataGroup_hi_lo_462 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_463;
  assign dataGroup_hi_lo_463 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_464;
  assign dataGroup_hi_lo_464 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_465;
  assign dataGroup_hi_lo_465 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_466;
  assign dataGroup_hi_lo_466 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_467;
  assign dataGroup_hi_lo_467 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_468;
  assign dataGroup_hi_lo_468 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_469;
  assign dataGroup_hi_lo_469 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_470;
  assign dataGroup_hi_lo_470 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_471;
  assign dataGroup_hi_lo_471 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_472;
  assign dataGroup_hi_lo_472 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_473;
  assign dataGroup_hi_lo_473 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_474;
  assign dataGroup_hi_lo_474 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_475;
  assign dataGroup_hi_lo_475 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_476;
  assign dataGroup_hi_lo_476 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_477;
  assign dataGroup_hi_lo_477 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_478;
  assign dataGroup_hi_lo_478 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_479;
  assign dataGroup_hi_lo_479 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_480;
  assign dataGroup_hi_lo_480 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_481;
  assign dataGroup_hi_lo_481 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_482;
  assign dataGroup_hi_lo_482 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_483;
  assign dataGroup_hi_lo_483 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_484;
  assign dataGroup_hi_lo_484 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_485;
  assign dataGroup_hi_lo_485 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_486;
  assign dataGroup_hi_lo_486 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_487;
  assign dataGroup_hi_lo_487 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_488;
  assign dataGroup_hi_lo_488 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_489;
  assign dataGroup_hi_lo_489 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_490;
  assign dataGroup_hi_lo_490 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_491;
  assign dataGroup_hi_lo_491 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_492;
  assign dataGroup_hi_lo_492 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_493;
  assign dataGroup_hi_lo_493 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_494;
  assign dataGroup_hi_lo_494 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_495;
  assign dataGroup_hi_lo_495 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_496;
  assign dataGroup_hi_lo_496 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_497;
  assign dataGroup_hi_lo_497 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_498;
  assign dataGroup_hi_lo_498 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_499;
  assign dataGroup_hi_lo_499 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_500;
  assign dataGroup_hi_lo_500 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_501;
  assign dataGroup_hi_lo_501 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_502;
  assign dataGroup_hi_lo_502 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_503;
  assign dataGroup_hi_lo_503 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_504;
  assign dataGroup_hi_lo_504 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_505;
  assign dataGroup_hi_lo_505 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_506;
  assign dataGroup_hi_lo_506 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_507;
  assign dataGroup_hi_lo_507 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_508;
  assign dataGroup_hi_lo_508 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_509;
  assign dataGroup_hi_lo_509 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_510;
  assign dataGroup_hi_lo_510 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_511;
  assign dataGroup_hi_lo_511 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_512;
  assign dataGroup_hi_lo_512 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_513;
  assign dataGroup_hi_lo_513 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_514;
  assign dataGroup_hi_lo_514 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_515;
  assign dataGroup_hi_lo_515 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_516;
  assign dataGroup_hi_lo_516 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_517;
  assign dataGroup_hi_lo_517 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_518;
  assign dataGroup_hi_lo_518 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_519;
  assign dataGroup_hi_lo_519 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_520;
  assign dataGroup_hi_lo_520 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_521;
  assign dataGroup_hi_lo_521 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_522;
  assign dataGroup_hi_lo_522 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_523;
  assign dataGroup_hi_lo_523 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_524;
  assign dataGroup_hi_lo_524 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_525;
  assign dataGroup_hi_lo_525 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_526;
  assign dataGroup_hi_lo_526 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_527;
  assign dataGroup_hi_lo_527 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_528;
  assign dataGroup_hi_lo_528 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_529;
  assign dataGroup_hi_lo_529 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_530;
  assign dataGroup_hi_lo_530 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_531;
  assign dataGroup_hi_lo_531 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_532;
  assign dataGroup_hi_lo_532 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_533;
  assign dataGroup_hi_lo_533 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_534;
  assign dataGroup_hi_lo_534 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_535;
  assign dataGroup_hi_lo_535 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_536;
  assign dataGroup_hi_lo_536 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_537;
  assign dataGroup_hi_lo_537 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_538;
  assign dataGroup_hi_lo_538 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_539;
  assign dataGroup_hi_lo_539 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_540;
  assign dataGroup_hi_lo_540 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_541;
  assign dataGroup_hi_lo_541 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_542;
  assign dataGroup_hi_lo_542 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_543;
  assign dataGroup_hi_lo_543 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_544;
  assign dataGroup_hi_lo_544 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_545;
  assign dataGroup_hi_lo_545 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_546;
  assign dataGroup_hi_lo_546 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_547;
  assign dataGroup_hi_lo_547 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_548;
  assign dataGroup_hi_lo_548 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_549;
  assign dataGroup_hi_lo_549 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_550;
  assign dataGroup_hi_lo_550 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_551;
  assign dataGroup_hi_lo_551 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_552;
  assign dataGroup_hi_lo_552 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_553;
  assign dataGroup_hi_lo_553 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_554;
  assign dataGroup_hi_lo_554 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_555;
  assign dataGroup_hi_lo_555 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_556;
  assign dataGroup_hi_lo_556 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_557;
  assign dataGroup_hi_lo_557 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_558;
  assign dataGroup_hi_lo_558 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_559;
  assign dataGroup_hi_lo_559 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_560;
  assign dataGroup_hi_lo_560 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_561;
  assign dataGroup_hi_lo_561 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_562;
  assign dataGroup_hi_lo_562 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_563;
  assign dataGroup_hi_lo_563 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_564;
  assign dataGroup_hi_lo_564 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_565;
  assign dataGroup_hi_lo_565 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_566;
  assign dataGroup_hi_lo_566 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_567;
  assign dataGroup_hi_lo_567 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_568;
  assign dataGroup_hi_lo_568 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_569;
  assign dataGroup_hi_lo_569 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_570;
  assign dataGroup_hi_lo_570 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_571;
  assign dataGroup_hi_lo_571 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_572;
  assign dataGroup_hi_lo_572 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_573;
  assign dataGroup_hi_lo_573 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_574;
  assign dataGroup_hi_lo_574 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_575;
  assign dataGroup_hi_lo_575 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_576;
  assign dataGroup_hi_lo_576 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_577;
  assign dataGroup_hi_lo_577 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_578;
  assign dataGroup_hi_lo_578 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_579;
  assign dataGroup_hi_lo_579 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_580;
  assign dataGroup_hi_lo_580 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_581;
  assign dataGroup_hi_lo_581 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_582;
  assign dataGroup_hi_lo_582 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_583;
  assign dataGroup_hi_lo_583 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_584;
  assign dataGroup_hi_lo_584 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_585;
  assign dataGroup_hi_lo_585 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_586;
  assign dataGroup_hi_lo_586 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_587;
  assign dataGroup_hi_lo_587 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_588;
  assign dataGroup_hi_lo_588 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_589;
  assign dataGroup_hi_lo_589 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_590;
  assign dataGroup_hi_lo_590 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_591;
  assign dataGroup_hi_lo_591 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_592;
  assign dataGroup_hi_lo_592 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_593;
  assign dataGroup_hi_lo_593 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_594;
  assign dataGroup_hi_lo_594 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_595;
  assign dataGroup_hi_lo_595 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_596;
  assign dataGroup_hi_lo_596 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_597;
  assign dataGroup_hi_lo_597 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_598;
  assign dataGroup_hi_lo_598 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_599;
  assign dataGroup_hi_lo_599 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_600;
  assign dataGroup_hi_lo_600 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_601;
  assign dataGroup_hi_lo_601 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_602;
  assign dataGroup_hi_lo_602 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_603;
  assign dataGroup_hi_lo_603 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_604;
  assign dataGroup_hi_lo_604 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_605;
  assign dataGroup_hi_lo_605 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_606;
  assign dataGroup_hi_lo_606 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_607;
  assign dataGroup_hi_lo_607 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_608;
  assign dataGroup_hi_lo_608 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_609;
  assign dataGroup_hi_lo_609 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_610;
  assign dataGroup_hi_lo_610 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_611;
  assign dataGroup_hi_lo_611 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_612;
  assign dataGroup_hi_lo_612 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_613;
  assign dataGroup_hi_lo_613 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_614;
  assign dataGroup_hi_lo_614 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_615;
  assign dataGroup_hi_lo_615 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_616;
  assign dataGroup_hi_lo_616 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_617;
  assign dataGroup_hi_lo_617 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_618;
  assign dataGroup_hi_lo_618 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_619;
  assign dataGroup_hi_lo_619 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_620;
  assign dataGroup_hi_lo_620 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_621;
  assign dataGroup_hi_lo_621 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_622;
  assign dataGroup_hi_lo_622 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_623;
  assign dataGroup_hi_lo_623 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_624;
  assign dataGroup_hi_lo_624 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_625;
  assign dataGroup_hi_lo_625 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_626;
  assign dataGroup_hi_lo_626 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_627;
  assign dataGroup_hi_lo_627 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_628;
  assign dataGroup_hi_lo_628 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_629;
  assign dataGroup_hi_lo_629 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_630;
  assign dataGroup_hi_lo_630 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_631;
  assign dataGroup_hi_lo_631 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_632;
  assign dataGroup_hi_lo_632 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_633;
  assign dataGroup_hi_lo_633 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_634;
  assign dataGroup_hi_lo_634 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_635;
  assign dataGroup_hi_lo_635 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_636;
  assign dataGroup_hi_lo_636 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_637;
  assign dataGroup_hi_lo_637 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_638;
  assign dataGroup_hi_lo_638 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_639;
  assign dataGroup_hi_lo_639 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_640;
  assign dataGroup_hi_lo_640 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_641;
  assign dataGroup_hi_lo_641 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_642;
  assign dataGroup_hi_lo_642 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_643;
  assign dataGroup_hi_lo_643 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_644;
  assign dataGroup_hi_lo_644 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_645;
  assign dataGroup_hi_lo_645 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_646;
  assign dataGroup_hi_lo_646 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_647;
  assign dataGroup_hi_lo_647 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_648;
  assign dataGroup_hi_lo_648 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_649;
  assign dataGroup_hi_lo_649 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_650;
  assign dataGroup_hi_lo_650 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_651;
  assign dataGroup_hi_lo_651 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_652;
  assign dataGroup_hi_lo_652 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_653;
  assign dataGroup_hi_lo_653 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_654;
  assign dataGroup_hi_lo_654 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_655;
  assign dataGroup_hi_lo_655 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_656;
  assign dataGroup_hi_lo_656 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_657;
  assign dataGroup_hi_lo_657 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_658;
  assign dataGroup_hi_lo_658 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_659;
  assign dataGroup_hi_lo_659 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_660;
  assign dataGroup_hi_lo_660 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_661;
  assign dataGroup_hi_lo_661 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_662;
  assign dataGroup_hi_lo_662 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_663;
  assign dataGroup_hi_lo_663 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_664;
  assign dataGroup_hi_lo_664 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_665;
  assign dataGroup_hi_lo_665 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_666;
  assign dataGroup_hi_lo_666 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_667;
  assign dataGroup_hi_lo_667 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_668;
  assign dataGroup_hi_lo_668 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_669;
  assign dataGroup_hi_lo_669 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_670;
  assign dataGroup_hi_lo_670 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_671;
  assign dataGroup_hi_lo_671 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_672;
  assign dataGroup_hi_lo_672 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_673;
  assign dataGroup_hi_lo_673 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_674;
  assign dataGroup_hi_lo_674 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_675;
  assign dataGroup_hi_lo_675 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_676;
  assign dataGroup_hi_lo_676 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_677;
  assign dataGroup_hi_lo_677 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_678;
  assign dataGroup_hi_lo_678 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_679;
  assign dataGroup_hi_lo_679 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_680;
  assign dataGroup_hi_lo_680 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_681;
  assign dataGroup_hi_lo_681 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_682;
  assign dataGroup_hi_lo_682 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_683;
  assign dataGroup_hi_lo_683 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_684;
  assign dataGroup_hi_lo_684 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_685;
  assign dataGroup_hi_lo_685 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_686;
  assign dataGroup_hi_lo_686 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_687;
  assign dataGroup_hi_lo_687 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_688;
  assign dataGroup_hi_lo_688 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_689;
  assign dataGroup_hi_lo_689 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_690;
  assign dataGroup_hi_lo_690 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_691;
  assign dataGroup_hi_lo_691 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_692;
  assign dataGroup_hi_lo_692 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_693;
  assign dataGroup_hi_lo_693 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_694;
  assign dataGroup_hi_lo_694 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_695;
  assign dataGroup_hi_lo_695 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_696;
  assign dataGroup_hi_lo_696 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_697;
  assign dataGroup_hi_lo_697 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_698;
  assign dataGroup_hi_lo_698 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_699;
  assign dataGroup_hi_lo_699 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_700;
  assign dataGroup_hi_lo_700 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_701;
  assign dataGroup_hi_lo_701 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_702;
  assign dataGroup_hi_lo_702 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_703;
  assign dataGroup_hi_lo_703 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_704;
  assign dataGroup_hi_lo_704 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_705;
  assign dataGroup_hi_lo_705 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_706;
  assign dataGroup_hi_lo_706 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_707;
  assign dataGroup_hi_lo_707 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_708;
  assign dataGroup_hi_lo_708 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_709;
  assign dataGroup_hi_lo_709 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_710;
  assign dataGroup_hi_lo_710 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_711;
  assign dataGroup_hi_lo_711 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_712;
  assign dataGroup_hi_lo_712 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_713;
  assign dataGroup_hi_lo_713 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_714;
  assign dataGroup_hi_lo_714 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_715;
  assign dataGroup_hi_lo_715 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_716;
  assign dataGroup_hi_lo_716 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_717;
  assign dataGroup_hi_lo_717 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_718;
  assign dataGroup_hi_lo_718 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_719;
  assign dataGroup_hi_lo_719 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_720;
  assign dataGroup_hi_lo_720 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_721;
  assign dataGroup_hi_lo_721 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_722;
  assign dataGroup_hi_lo_722 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_723;
  assign dataGroup_hi_lo_723 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_724;
  assign dataGroup_hi_lo_724 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_725;
  assign dataGroup_hi_lo_725 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_726;
  assign dataGroup_hi_lo_726 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_727;
  assign dataGroup_hi_lo_727 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_728;
  assign dataGroup_hi_lo_728 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_729;
  assign dataGroup_hi_lo_729 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_730;
  assign dataGroup_hi_lo_730 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_731;
  assign dataGroup_hi_lo_731 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_732;
  assign dataGroup_hi_lo_732 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_733;
  assign dataGroup_hi_lo_733 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_734;
  assign dataGroup_hi_lo_734 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_735;
  assign dataGroup_hi_lo_735 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_736;
  assign dataGroup_hi_lo_736 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_737;
  assign dataGroup_hi_lo_737 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_738;
  assign dataGroup_hi_lo_738 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_739;
  assign dataGroup_hi_lo_739 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_740;
  assign dataGroup_hi_lo_740 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_741;
  assign dataGroup_hi_lo_741 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_742;
  assign dataGroup_hi_lo_742 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_743;
  assign dataGroup_hi_lo_743 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_744;
  assign dataGroup_hi_lo_744 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_745;
  assign dataGroup_hi_lo_745 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_746;
  assign dataGroup_hi_lo_746 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_747;
  assign dataGroup_hi_lo_747 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_748;
  assign dataGroup_hi_lo_748 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_749;
  assign dataGroup_hi_lo_749 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_750;
  assign dataGroup_hi_lo_750 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_751;
  assign dataGroup_hi_lo_751 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_752;
  assign dataGroup_hi_lo_752 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_753;
  assign dataGroup_hi_lo_753 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_754;
  assign dataGroup_hi_lo_754 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_755;
  assign dataGroup_hi_lo_755 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_756;
  assign dataGroup_hi_lo_756 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_757;
  assign dataGroup_hi_lo_757 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_758;
  assign dataGroup_hi_lo_758 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_759;
  assign dataGroup_hi_lo_759 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_760;
  assign dataGroup_hi_lo_760 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_761;
  assign dataGroup_hi_lo_761 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_762;
  assign dataGroup_hi_lo_762 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_763;
  assign dataGroup_hi_lo_763 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_764;
  assign dataGroup_hi_lo_764 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_765;
  assign dataGroup_hi_lo_765 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_766;
  assign dataGroup_hi_lo_766 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_767;
  assign dataGroup_hi_lo_767 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_768;
  assign dataGroup_hi_lo_768 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_769;
  assign dataGroup_hi_lo_769 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_770;
  assign dataGroup_hi_lo_770 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_771;
  assign dataGroup_hi_lo_771 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_772;
  assign dataGroup_hi_lo_772 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_773;
  assign dataGroup_hi_lo_773 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_774;
  assign dataGroup_hi_lo_774 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_775;
  assign dataGroup_hi_lo_775 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_776;
  assign dataGroup_hi_lo_776 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_777;
  assign dataGroup_hi_lo_777 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_778;
  assign dataGroup_hi_lo_778 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_779;
  assign dataGroup_hi_lo_779 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_780;
  assign dataGroup_hi_lo_780 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_781;
  assign dataGroup_hi_lo_781 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_782;
  assign dataGroup_hi_lo_782 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_783;
  assign dataGroup_hi_lo_783 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_784;
  assign dataGroup_hi_lo_784 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_785;
  assign dataGroup_hi_lo_785 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_786;
  assign dataGroup_hi_lo_786 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_787;
  assign dataGroup_hi_lo_787 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_788;
  assign dataGroup_hi_lo_788 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_789;
  assign dataGroup_hi_lo_789 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_790;
  assign dataGroup_hi_lo_790 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_791;
  assign dataGroup_hi_lo_791 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_792;
  assign dataGroup_hi_lo_792 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_793;
  assign dataGroup_hi_lo_793 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_794;
  assign dataGroup_hi_lo_794 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_795;
  assign dataGroup_hi_lo_795 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_796;
  assign dataGroup_hi_lo_796 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_797;
  assign dataGroup_hi_lo_797 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_798;
  assign dataGroup_hi_lo_798 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_799;
  assign dataGroup_hi_lo_799 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_800;
  assign dataGroup_hi_lo_800 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_801;
  assign dataGroup_hi_lo_801 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_802;
  assign dataGroup_hi_lo_802 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_803;
  assign dataGroup_hi_lo_803 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_804;
  assign dataGroup_hi_lo_804 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_805;
  assign dataGroup_hi_lo_805 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_806;
  assign dataGroup_hi_lo_806 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_807;
  assign dataGroup_hi_lo_807 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_808;
  assign dataGroup_hi_lo_808 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_809;
  assign dataGroup_hi_lo_809 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_810;
  assign dataGroup_hi_lo_810 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_811;
  assign dataGroup_hi_lo_811 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_812;
  assign dataGroup_hi_lo_812 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_813;
  assign dataGroup_hi_lo_813 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_814;
  assign dataGroup_hi_lo_814 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_815;
  assign dataGroup_hi_lo_815 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_816;
  assign dataGroup_hi_lo_816 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_817;
  assign dataGroup_hi_lo_817 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_818;
  assign dataGroup_hi_lo_818 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_819;
  assign dataGroup_hi_lo_819 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_820;
  assign dataGroup_hi_lo_820 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_821;
  assign dataGroup_hi_lo_821 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_822;
  assign dataGroup_hi_lo_822 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_823;
  assign dataGroup_hi_lo_823 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_824;
  assign dataGroup_hi_lo_824 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_825;
  assign dataGroup_hi_lo_825 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_826;
  assign dataGroup_hi_lo_826 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_827;
  assign dataGroup_hi_lo_827 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_828;
  assign dataGroup_hi_lo_828 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_829;
  assign dataGroup_hi_lo_829 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_830;
  assign dataGroup_hi_lo_830 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_831;
  assign dataGroup_hi_lo_831 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_832;
  assign dataGroup_hi_lo_832 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_833;
  assign dataGroup_hi_lo_833 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_834;
  assign dataGroup_hi_lo_834 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_835;
  assign dataGroup_hi_lo_835 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_836;
  assign dataGroup_hi_lo_836 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_837;
  assign dataGroup_hi_lo_837 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_838;
  assign dataGroup_hi_lo_838 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_839;
  assign dataGroup_hi_lo_839 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_840;
  assign dataGroup_hi_lo_840 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_841;
  assign dataGroup_hi_lo_841 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_842;
  assign dataGroup_hi_lo_842 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_843;
  assign dataGroup_hi_lo_843 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_844;
  assign dataGroup_hi_lo_844 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_845;
  assign dataGroup_hi_lo_845 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_846;
  assign dataGroup_hi_lo_846 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_847;
  assign dataGroup_hi_lo_847 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_848;
  assign dataGroup_hi_lo_848 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_849;
  assign dataGroup_hi_lo_849 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_850;
  assign dataGroup_hi_lo_850 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_851;
  assign dataGroup_hi_lo_851 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_852;
  assign dataGroup_hi_lo_852 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_853;
  assign dataGroup_hi_lo_853 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_854;
  assign dataGroup_hi_lo_854 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_855;
  assign dataGroup_hi_lo_855 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_856;
  assign dataGroup_hi_lo_856 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_857;
  assign dataGroup_hi_lo_857 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_858;
  assign dataGroup_hi_lo_858 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_859;
  assign dataGroup_hi_lo_859 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_860;
  assign dataGroup_hi_lo_860 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_861;
  assign dataGroup_hi_lo_861 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_862;
  assign dataGroup_hi_lo_862 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_863;
  assign dataGroup_hi_lo_863 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_864;
  assign dataGroup_hi_lo_864 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_865;
  assign dataGroup_hi_lo_865 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_866;
  assign dataGroup_hi_lo_866 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_867;
  assign dataGroup_hi_lo_867 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_868;
  assign dataGroup_hi_lo_868 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_869;
  assign dataGroup_hi_lo_869 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_870;
  assign dataGroup_hi_lo_870 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_871;
  assign dataGroup_hi_lo_871 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_872;
  assign dataGroup_hi_lo_872 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_873;
  assign dataGroup_hi_lo_873 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_874;
  assign dataGroup_hi_lo_874 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_875;
  assign dataGroup_hi_lo_875 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_876;
  assign dataGroup_hi_lo_876 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_877;
  assign dataGroup_hi_lo_877 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_878;
  assign dataGroup_hi_lo_878 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_879;
  assign dataGroup_hi_lo_879 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_880;
  assign dataGroup_hi_lo_880 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_881;
  assign dataGroup_hi_lo_881 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_882;
  assign dataGroup_hi_lo_882 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_883;
  assign dataGroup_hi_lo_883 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_884;
  assign dataGroup_hi_lo_884 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_885;
  assign dataGroup_hi_lo_885 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_886;
  assign dataGroup_hi_lo_886 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_887;
  assign dataGroup_hi_lo_887 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_888;
  assign dataGroup_hi_lo_888 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_889;
  assign dataGroup_hi_lo_889 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_890;
  assign dataGroup_hi_lo_890 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_891;
  assign dataGroup_hi_lo_891 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_892;
  assign dataGroup_hi_lo_892 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_893;
  assign dataGroup_hi_lo_893 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_894;
  assign dataGroup_hi_lo_894 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_895;
  assign dataGroup_hi_lo_895 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_896;
  assign dataGroup_hi_lo_896 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_897;
  assign dataGroup_hi_lo_897 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_898;
  assign dataGroup_hi_lo_898 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_899;
  assign dataGroup_hi_lo_899 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_900;
  assign dataGroup_hi_lo_900 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_901;
  assign dataGroup_hi_lo_901 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_902;
  assign dataGroup_hi_lo_902 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_903;
  assign dataGroup_hi_lo_903 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_904;
  assign dataGroup_hi_lo_904 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_905;
  assign dataGroup_hi_lo_905 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_906;
  assign dataGroup_hi_lo_906 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_907;
  assign dataGroup_hi_lo_907 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_908;
  assign dataGroup_hi_lo_908 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_909;
  assign dataGroup_hi_lo_909 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_910;
  assign dataGroup_hi_lo_910 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_911;
  assign dataGroup_hi_lo_911 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_912;
  assign dataGroup_hi_lo_912 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_913;
  assign dataGroup_hi_lo_913 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_914;
  assign dataGroup_hi_lo_914 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_915;
  assign dataGroup_hi_lo_915 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_916;
  assign dataGroup_hi_lo_916 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_917;
  assign dataGroup_hi_lo_917 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_918;
  assign dataGroup_hi_lo_918 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_919;
  assign dataGroup_hi_lo_919 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_920;
  assign dataGroup_hi_lo_920 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_921;
  assign dataGroup_hi_lo_921 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_922;
  assign dataGroup_hi_lo_922 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_923;
  assign dataGroup_hi_lo_923 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_924;
  assign dataGroup_hi_lo_924 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_925;
  assign dataGroup_hi_lo_925 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_926;
  assign dataGroup_hi_lo_926 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_927;
  assign dataGroup_hi_lo_927 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_928;
  assign dataGroup_hi_lo_928 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_929;
  assign dataGroup_hi_lo_929 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_930;
  assign dataGroup_hi_lo_930 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_931;
  assign dataGroup_hi_lo_931 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_932;
  assign dataGroup_hi_lo_932 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_933;
  assign dataGroup_hi_lo_933 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_934;
  assign dataGroup_hi_lo_934 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_935;
  assign dataGroup_hi_lo_935 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_936;
  assign dataGroup_hi_lo_936 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_937;
  assign dataGroup_hi_lo_937 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_938;
  assign dataGroup_hi_lo_938 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_939;
  assign dataGroup_hi_lo_939 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_940;
  assign dataGroup_hi_lo_940 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_941;
  assign dataGroup_hi_lo_941 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_942;
  assign dataGroup_hi_lo_942 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_943;
  assign dataGroup_hi_lo_943 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_944;
  assign dataGroup_hi_lo_944 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_945;
  assign dataGroup_hi_lo_945 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_946;
  assign dataGroup_hi_lo_946 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_947;
  assign dataGroup_hi_lo_947 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_948;
  assign dataGroup_hi_lo_948 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_949;
  assign dataGroup_hi_lo_949 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_950;
  assign dataGroup_hi_lo_950 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_951;
  assign dataGroup_hi_lo_951 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_952;
  assign dataGroup_hi_lo_952 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_953;
  assign dataGroup_hi_lo_953 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_954;
  assign dataGroup_hi_lo_954 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_955;
  assign dataGroup_hi_lo_955 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_956;
  assign dataGroup_hi_lo_956 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_957;
  assign dataGroup_hi_lo_957 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_958;
  assign dataGroup_hi_lo_958 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_959;
  assign dataGroup_hi_lo_959 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_960;
  assign dataGroup_hi_lo_960 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_961;
  assign dataGroup_hi_lo_961 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_962;
  assign dataGroup_hi_lo_962 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_963;
  assign dataGroup_hi_lo_963 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_964;
  assign dataGroup_hi_lo_964 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_965;
  assign dataGroup_hi_lo_965 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_966;
  assign dataGroup_hi_lo_966 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_967;
  assign dataGroup_hi_lo_967 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_968;
  assign dataGroup_hi_lo_968 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_969;
  assign dataGroup_hi_lo_969 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_970;
  assign dataGroup_hi_lo_970 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_971;
  assign dataGroup_hi_lo_971 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_972;
  assign dataGroup_hi_lo_972 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_973;
  assign dataGroup_hi_lo_973 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_974;
  assign dataGroup_hi_lo_974 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_975;
  assign dataGroup_hi_lo_975 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_976;
  assign dataGroup_hi_lo_976 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_977;
  assign dataGroup_hi_lo_977 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_978;
  assign dataGroup_hi_lo_978 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_979;
  assign dataGroup_hi_lo_979 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_980;
  assign dataGroup_hi_lo_980 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_981;
  assign dataGroup_hi_lo_981 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_982;
  assign dataGroup_hi_lo_982 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_983;
  assign dataGroup_hi_lo_983 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_984;
  assign dataGroup_hi_lo_984 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_985;
  assign dataGroup_hi_lo_985 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_986;
  assign dataGroup_hi_lo_986 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_987;
  assign dataGroup_hi_lo_987 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_988;
  assign dataGroup_hi_lo_988 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_989;
  assign dataGroup_hi_lo_989 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_990;
  assign dataGroup_hi_lo_990 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_991;
  assign dataGroup_hi_lo_991 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_992;
  assign dataGroup_hi_lo_992 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_993;
  assign dataGroup_hi_lo_993 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_994;
  assign dataGroup_hi_lo_994 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_995;
  assign dataGroup_hi_lo_995 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_996;
  assign dataGroup_hi_lo_996 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_997;
  assign dataGroup_hi_lo_997 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_998;
  assign dataGroup_hi_lo_998 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_999;
  assign dataGroup_hi_lo_999 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1000;
  assign dataGroup_hi_lo_1000 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1001;
  assign dataGroup_hi_lo_1001 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1002;
  assign dataGroup_hi_lo_1002 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1003;
  assign dataGroup_hi_lo_1003 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1004;
  assign dataGroup_hi_lo_1004 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1005;
  assign dataGroup_hi_lo_1005 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1006;
  assign dataGroup_hi_lo_1006 = _GEN_5;
  wire [255:0]  dataGroup_hi_lo_1007;
  assign dataGroup_hi_lo_1007 = _GEN_5;
  wire [255:0]  _GEN_6 = {dataSelect_7, dataSelect_6};
  wire [255:0]  dataGroup_hi_hi;
  assign dataGroup_hi_hi = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1;
  assign dataGroup_hi_hi_1 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_2;
  assign dataGroup_hi_hi_2 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_3;
  assign dataGroup_hi_hi_3 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_4;
  assign dataGroup_hi_hi_4 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_5;
  assign dataGroup_hi_hi_5 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_6;
  assign dataGroup_hi_hi_6 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_7;
  assign dataGroup_hi_hi_7 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_8;
  assign dataGroup_hi_hi_8 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_9;
  assign dataGroup_hi_hi_9 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_10;
  assign dataGroup_hi_hi_10 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_11;
  assign dataGroup_hi_hi_11 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_12;
  assign dataGroup_hi_hi_12 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_13;
  assign dataGroup_hi_hi_13 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_14;
  assign dataGroup_hi_hi_14 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_15;
  assign dataGroup_hi_hi_15 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_16;
  assign dataGroup_hi_hi_16 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_17;
  assign dataGroup_hi_hi_17 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_18;
  assign dataGroup_hi_hi_18 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_19;
  assign dataGroup_hi_hi_19 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_20;
  assign dataGroup_hi_hi_20 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_21;
  assign dataGroup_hi_hi_21 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_22;
  assign dataGroup_hi_hi_22 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_23;
  assign dataGroup_hi_hi_23 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_24;
  assign dataGroup_hi_hi_24 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_25;
  assign dataGroup_hi_hi_25 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_26;
  assign dataGroup_hi_hi_26 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_27;
  assign dataGroup_hi_hi_27 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_28;
  assign dataGroup_hi_hi_28 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_29;
  assign dataGroup_hi_hi_29 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_30;
  assign dataGroup_hi_hi_30 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_31;
  assign dataGroup_hi_hi_31 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_32;
  assign dataGroup_hi_hi_32 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_33;
  assign dataGroup_hi_hi_33 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_34;
  assign dataGroup_hi_hi_34 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_35;
  assign dataGroup_hi_hi_35 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_36;
  assign dataGroup_hi_hi_36 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_37;
  assign dataGroup_hi_hi_37 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_38;
  assign dataGroup_hi_hi_38 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_39;
  assign dataGroup_hi_hi_39 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_40;
  assign dataGroup_hi_hi_40 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_41;
  assign dataGroup_hi_hi_41 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_42;
  assign dataGroup_hi_hi_42 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_43;
  assign dataGroup_hi_hi_43 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_44;
  assign dataGroup_hi_hi_44 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_45;
  assign dataGroup_hi_hi_45 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_46;
  assign dataGroup_hi_hi_46 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_47;
  assign dataGroup_hi_hi_47 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_48;
  assign dataGroup_hi_hi_48 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_49;
  assign dataGroup_hi_hi_49 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_50;
  assign dataGroup_hi_hi_50 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_51;
  assign dataGroup_hi_hi_51 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_52;
  assign dataGroup_hi_hi_52 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_53;
  assign dataGroup_hi_hi_53 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_54;
  assign dataGroup_hi_hi_54 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_55;
  assign dataGroup_hi_hi_55 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_56;
  assign dataGroup_hi_hi_56 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_57;
  assign dataGroup_hi_hi_57 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_58;
  assign dataGroup_hi_hi_58 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_59;
  assign dataGroup_hi_hi_59 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_60;
  assign dataGroup_hi_hi_60 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_61;
  assign dataGroup_hi_hi_61 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_62;
  assign dataGroup_hi_hi_62 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_63;
  assign dataGroup_hi_hi_63 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_64;
  assign dataGroup_hi_hi_64 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_65;
  assign dataGroup_hi_hi_65 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_66;
  assign dataGroup_hi_hi_66 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_67;
  assign dataGroup_hi_hi_67 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_68;
  assign dataGroup_hi_hi_68 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_69;
  assign dataGroup_hi_hi_69 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_70;
  assign dataGroup_hi_hi_70 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_71;
  assign dataGroup_hi_hi_71 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_72;
  assign dataGroup_hi_hi_72 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_73;
  assign dataGroup_hi_hi_73 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_74;
  assign dataGroup_hi_hi_74 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_75;
  assign dataGroup_hi_hi_75 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_76;
  assign dataGroup_hi_hi_76 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_77;
  assign dataGroup_hi_hi_77 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_78;
  assign dataGroup_hi_hi_78 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_79;
  assign dataGroup_hi_hi_79 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_80;
  assign dataGroup_hi_hi_80 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_81;
  assign dataGroup_hi_hi_81 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_82;
  assign dataGroup_hi_hi_82 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_83;
  assign dataGroup_hi_hi_83 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_84;
  assign dataGroup_hi_hi_84 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_85;
  assign dataGroup_hi_hi_85 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_86;
  assign dataGroup_hi_hi_86 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_87;
  assign dataGroup_hi_hi_87 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_88;
  assign dataGroup_hi_hi_88 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_89;
  assign dataGroup_hi_hi_89 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_90;
  assign dataGroup_hi_hi_90 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_91;
  assign dataGroup_hi_hi_91 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_92;
  assign dataGroup_hi_hi_92 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_93;
  assign dataGroup_hi_hi_93 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_94;
  assign dataGroup_hi_hi_94 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_95;
  assign dataGroup_hi_hi_95 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_96;
  assign dataGroup_hi_hi_96 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_97;
  assign dataGroup_hi_hi_97 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_98;
  assign dataGroup_hi_hi_98 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_99;
  assign dataGroup_hi_hi_99 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_100;
  assign dataGroup_hi_hi_100 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_101;
  assign dataGroup_hi_hi_101 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_102;
  assign dataGroup_hi_hi_102 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_103;
  assign dataGroup_hi_hi_103 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_104;
  assign dataGroup_hi_hi_104 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_105;
  assign dataGroup_hi_hi_105 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_106;
  assign dataGroup_hi_hi_106 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_107;
  assign dataGroup_hi_hi_107 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_108;
  assign dataGroup_hi_hi_108 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_109;
  assign dataGroup_hi_hi_109 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_110;
  assign dataGroup_hi_hi_110 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_111;
  assign dataGroup_hi_hi_111 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_112;
  assign dataGroup_hi_hi_112 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_113;
  assign dataGroup_hi_hi_113 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_114;
  assign dataGroup_hi_hi_114 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_115;
  assign dataGroup_hi_hi_115 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_116;
  assign dataGroup_hi_hi_116 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_117;
  assign dataGroup_hi_hi_117 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_118;
  assign dataGroup_hi_hi_118 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_119;
  assign dataGroup_hi_hi_119 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_120;
  assign dataGroup_hi_hi_120 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_121;
  assign dataGroup_hi_hi_121 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_122;
  assign dataGroup_hi_hi_122 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_123;
  assign dataGroup_hi_hi_123 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_124;
  assign dataGroup_hi_hi_124 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_125;
  assign dataGroup_hi_hi_125 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_126;
  assign dataGroup_hi_hi_126 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_127;
  assign dataGroup_hi_hi_127 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_128;
  assign dataGroup_hi_hi_128 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_129;
  assign dataGroup_hi_hi_129 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_130;
  assign dataGroup_hi_hi_130 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_131;
  assign dataGroup_hi_hi_131 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_132;
  assign dataGroup_hi_hi_132 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_133;
  assign dataGroup_hi_hi_133 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_134;
  assign dataGroup_hi_hi_134 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_135;
  assign dataGroup_hi_hi_135 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_136;
  assign dataGroup_hi_hi_136 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_137;
  assign dataGroup_hi_hi_137 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_138;
  assign dataGroup_hi_hi_138 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_139;
  assign dataGroup_hi_hi_139 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_140;
  assign dataGroup_hi_hi_140 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_141;
  assign dataGroup_hi_hi_141 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_142;
  assign dataGroup_hi_hi_142 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_143;
  assign dataGroup_hi_hi_143 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_144;
  assign dataGroup_hi_hi_144 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_145;
  assign dataGroup_hi_hi_145 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_146;
  assign dataGroup_hi_hi_146 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_147;
  assign dataGroup_hi_hi_147 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_148;
  assign dataGroup_hi_hi_148 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_149;
  assign dataGroup_hi_hi_149 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_150;
  assign dataGroup_hi_hi_150 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_151;
  assign dataGroup_hi_hi_151 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_152;
  assign dataGroup_hi_hi_152 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_153;
  assign dataGroup_hi_hi_153 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_154;
  assign dataGroup_hi_hi_154 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_155;
  assign dataGroup_hi_hi_155 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_156;
  assign dataGroup_hi_hi_156 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_157;
  assign dataGroup_hi_hi_157 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_158;
  assign dataGroup_hi_hi_158 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_159;
  assign dataGroup_hi_hi_159 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_160;
  assign dataGroup_hi_hi_160 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_161;
  assign dataGroup_hi_hi_161 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_162;
  assign dataGroup_hi_hi_162 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_163;
  assign dataGroup_hi_hi_163 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_164;
  assign dataGroup_hi_hi_164 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_165;
  assign dataGroup_hi_hi_165 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_166;
  assign dataGroup_hi_hi_166 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_167;
  assign dataGroup_hi_hi_167 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_168;
  assign dataGroup_hi_hi_168 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_169;
  assign dataGroup_hi_hi_169 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_170;
  assign dataGroup_hi_hi_170 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_171;
  assign dataGroup_hi_hi_171 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_172;
  assign dataGroup_hi_hi_172 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_173;
  assign dataGroup_hi_hi_173 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_174;
  assign dataGroup_hi_hi_174 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_175;
  assign dataGroup_hi_hi_175 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_176;
  assign dataGroup_hi_hi_176 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_177;
  assign dataGroup_hi_hi_177 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_178;
  assign dataGroup_hi_hi_178 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_179;
  assign dataGroup_hi_hi_179 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_180;
  assign dataGroup_hi_hi_180 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_181;
  assign dataGroup_hi_hi_181 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_182;
  assign dataGroup_hi_hi_182 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_183;
  assign dataGroup_hi_hi_183 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_184;
  assign dataGroup_hi_hi_184 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_185;
  assign dataGroup_hi_hi_185 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_186;
  assign dataGroup_hi_hi_186 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_187;
  assign dataGroup_hi_hi_187 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_188;
  assign dataGroup_hi_hi_188 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_189;
  assign dataGroup_hi_hi_189 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_190;
  assign dataGroup_hi_hi_190 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_191;
  assign dataGroup_hi_hi_191 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_192;
  assign dataGroup_hi_hi_192 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_193;
  assign dataGroup_hi_hi_193 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_194;
  assign dataGroup_hi_hi_194 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_195;
  assign dataGroup_hi_hi_195 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_196;
  assign dataGroup_hi_hi_196 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_197;
  assign dataGroup_hi_hi_197 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_198;
  assign dataGroup_hi_hi_198 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_199;
  assign dataGroup_hi_hi_199 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_200;
  assign dataGroup_hi_hi_200 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_201;
  assign dataGroup_hi_hi_201 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_202;
  assign dataGroup_hi_hi_202 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_203;
  assign dataGroup_hi_hi_203 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_204;
  assign dataGroup_hi_hi_204 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_205;
  assign dataGroup_hi_hi_205 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_206;
  assign dataGroup_hi_hi_206 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_207;
  assign dataGroup_hi_hi_207 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_208;
  assign dataGroup_hi_hi_208 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_209;
  assign dataGroup_hi_hi_209 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_210;
  assign dataGroup_hi_hi_210 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_211;
  assign dataGroup_hi_hi_211 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_212;
  assign dataGroup_hi_hi_212 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_213;
  assign dataGroup_hi_hi_213 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_214;
  assign dataGroup_hi_hi_214 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_215;
  assign dataGroup_hi_hi_215 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_216;
  assign dataGroup_hi_hi_216 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_217;
  assign dataGroup_hi_hi_217 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_218;
  assign dataGroup_hi_hi_218 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_219;
  assign dataGroup_hi_hi_219 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_220;
  assign dataGroup_hi_hi_220 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_221;
  assign dataGroup_hi_hi_221 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_222;
  assign dataGroup_hi_hi_222 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_223;
  assign dataGroup_hi_hi_223 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_224;
  assign dataGroup_hi_hi_224 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_225;
  assign dataGroup_hi_hi_225 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_226;
  assign dataGroup_hi_hi_226 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_227;
  assign dataGroup_hi_hi_227 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_228;
  assign dataGroup_hi_hi_228 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_229;
  assign dataGroup_hi_hi_229 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_230;
  assign dataGroup_hi_hi_230 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_231;
  assign dataGroup_hi_hi_231 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_232;
  assign dataGroup_hi_hi_232 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_233;
  assign dataGroup_hi_hi_233 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_234;
  assign dataGroup_hi_hi_234 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_235;
  assign dataGroup_hi_hi_235 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_236;
  assign dataGroup_hi_hi_236 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_237;
  assign dataGroup_hi_hi_237 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_238;
  assign dataGroup_hi_hi_238 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_239;
  assign dataGroup_hi_hi_239 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_240;
  assign dataGroup_hi_hi_240 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_241;
  assign dataGroup_hi_hi_241 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_242;
  assign dataGroup_hi_hi_242 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_243;
  assign dataGroup_hi_hi_243 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_244;
  assign dataGroup_hi_hi_244 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_245;
  assign dataGroup_hi_hi_245 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_246;
  assign dataGroup_hi_hi_246 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_247;
  assign dataGroup_hi_hi_247 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_248;
  assign dataGroup_hi_hi_248 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_249;
  assign dataGroup_hi_hi_249 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_250;
  assign dataGroup_hi_hi_250 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_251;
  assign dataGroup_hi_hi_251 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_252;
  assign dataGroup_hi_hi_252 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_253;
  assign dataGroup_hi_hi_253 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_254;
  assign dataGroup_hi_hi_254 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_255;
  assign dataGroup_hi_hi_255 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_256;
  assign dataGroup_hi_hi_256 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_257;
  assign dataGroup_hi_hi_257 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_258;
  assign dataGroup_hi_hi_258 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_259;
  assign dataGroup_hi_hi_259 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_260;
  assign dataGroup_hi_hi_260 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_261;
  assign dataGroup_hi_hi_261 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_262;
  assign dataGroup_hi_hi_262 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_263;
  assign dataGroup_hi_hi_263 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_264;
  assign dataGroup_hi_hi_264 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_265;
  assign dataGroup_hi_hi_265 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_266;
  assign dataGroup_hi_hi_266 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_267;
  assign dataGroup_hi_hi_267 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_268;
  assign dataGroup_hi_hi_268 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_269;
  assign dataGroup_hi_hi_269 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_270;
  assign dataGroup_hi_hi_270 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_271;
  assign dataGroup_hi_hi_271 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_272;
  assign dataGroup_hi_hi_272 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_273;
  assign dataGroup_hi_hi_273 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_274;
  assign dataGroup_hi_hi_274 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_275;
  assign dataGroup_hi_hi_275 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_276;
  assign dataGroup_hi_hi_276 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_277;
  assign dataGroup_hi_hi_277 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_278;
  assign dataGroup_hi_hi_278 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_279;
  assign dataGroup_hi_hi_279 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_280;
  assign dataGroup_hi_hi_280 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_281;
  assign dataGroup_hi_hi_281 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_282;
  assign dataGroup_hi_hi_282 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_283;
  assign dataGroup_hi_hi_283 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_284;
  assign dataGroup_hi_hi_284 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_285;
  assign dataGroup_hi_hi_285 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_286;
  assign dataGroup_hi_hi_286 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_287;
  assign dataGroup_hi_hi_287 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_288;
  assign dataGroup_hi_hi_288 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_289;
  assign dataGroup_hi_hi_289 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_290;
  assign dataGroup_hi_hi_290 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_291;
  assign dataGroup_hi_hi_291 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_292;
  assign dataGroup_hi_hi_292 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_293;
  assign dataGroup_hi_hi_293 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_294;
  assign dataGroup_hi_hi_294 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_295;
  assign dataGroup_hi_hi_295 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_296;
  assign dataGroup_hi_hi_296 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_297;
  assign dataGroup_hi_hi_297 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_298;
  assign dataGroup_hi_hi_298 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_299;
  assign dataGroup_hi_hi_299 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_300;
  assign dataGroup_hi_hi_300 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_301;
  assign dataGroup_hi_hi_301 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_302;
  assign dataGroup_hi_hi_302 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_303;
  assign dataGroup_hi_hi_303 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_304;
  assign dataGroup_hi_hi_304 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_305;
  assign dataGroup_hi_hi_305 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_306;
  assign dataGroup_hi_hi_306 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_307;
  assign dataGroup_hi_hi_307 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_308;
  assign dataGroup_hi_hi_308 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_309;
  assign dataGroup_hi_hi_309 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_310;
  assign dataGroup_hi_hi_310 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_311;
  assign dataGroup_hi_hi_311 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_312;
  assign dataGroup_hi_hi_312 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_313;
  assign dataGroup_hi_hi_313 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_314;
  assign dataGroup_hi_hi_314 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_315;
  assign dataGroup_hi_hi_315 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_316;
  assign dataGroup_hi_hi_316 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_317;
  assign dataGroup_hi_hi_317 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_318;
  assign dataGroup_hi_hi_318 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_319;
  assign dataGroup_hi_hi_319 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_320;
  assign dataGroup_hi_hi_320 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_321;
  assign dataGroup_hi_hi_321 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_322;
  assign dataGroup_hi_hi_322 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_323;
  assign dataGroup_hi_hi_323 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_324;
  assign dataGroup_hi_hi_324 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_325;
  assign dataGroup_hi_hi_325 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_326;
  assign dataGroup_hi_hi_326 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_327;
  assign dataGroup_hi_hi_327 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_328;
  assign dataGroup_hi_hi_328 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_329;
  assign dataGroup_hi_hi_329 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_330;
  assign dataGroup_hi_hi_330 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_331;
  assign dataGroup_hi_hi_331 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_332;
  assign dataGroup_hi_hi_332 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_333;
  assign dataGroup_hi_hi_333 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_334;
  assign dataGroup_hi_hi_334 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_335;
  assign dataGroup_hi_hi_335 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_336;
  assign dataGroup_hi_hi_336 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_337;
  assign dataGroup_hi_hi_337 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_338;
  assign dataGroup_hi_hi_338 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_339;
  assign dataGroup_hi_hi_339 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_340;
  assign dataGroup_hi_hi_340 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_341;
  assign dataGroup_hi_hi_341 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_342;
  assign dataGroup_hi_hi_342 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_343;
  assign dataGroup_hi_hi_343 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_344;
  assign dataGroup_hi_hi_344 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_345;
  assign dataGroup_hi_hi_345 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_346;
  assign dataGroup_hi_hi_346 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_347;
  assign dataGroup_hi_hi_347 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_348;
  assign dataGroup_hi_hi_348 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_349;
  assign dataGroup_hi_hi_349 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_350;
  assign dataGroup_hi_hi_350 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_351;
  assign dataGroup_hi_hi_351 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_352;
  assign dataGroup_hi_hi_352 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_353;
  assign dataGroup_hi_hi_353 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_354;
  assign dataGroup_hi_hi_354 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_355;
  assign dataGroup_hi_hi_355 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_356;
  assign dataGroup_hi_hi_356 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_357;
  assign dataGroup_hi_hi_357 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_358;
  assign dataGroup_hi_hi_358 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_359;
  assign dataGroup_hi_hi_359 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_360;
  assign dataGroup_hi_hi_360 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_361;
  assign dataGroup_hi_hi_361 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_362;
  assign dataGroup_hi_hi_362 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_363;
  assign dataGroup_hi_hi_363 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_364;
  assign dataGroup_hi_hi_364 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_365;
  assign dataGroup_hi_hi_365 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_366;
  assign dataGroup_hi_hi_366 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_367;
  assign dataGroup_hi_hi_367 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_368;
  assign dataGroup_hi_hi_368 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_369;
  assign dataGroup_hi_hi_369 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_370;
  assign dataGroup_hi_hi_370 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_371;
  assign dataGroup_hi_hi_371 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_372;
  assign dataGroup_hi_hi_372 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_373;
  assign dataGroup_hi_hi_373 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_374;
  assign dataGroup_hi_hi_374 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_375;
  assign dataGroup_hi_hi_375 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_376;
  assign dataGroup_hi_hi_376 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_377;
  assign dataGroup_hi_hi_377 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_378;
  assign dataGroup_hi_hi_378 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_379;
  assign dataGroup_hi_hi_379 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_380;
  assign dataGroup_hi_hi_380 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_381;
  assign dataGroup_hi_hi_381 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_382;
  assign dataGroup_hi_hi_382 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_383;
  assign dataGroup_hi_hi_383 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_384;
  assign dataGroup_hi_hi_384 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_385;
  assign dataGroup_hi_hi_385 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_386;
  assign dataGroup_hi_hi_386 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_387;
  assign dataGroup_hi_hi_387 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_388;
  assign dataGroup_hi_hi_388 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_389;
  assign dataGroup_hi_hi_389 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_390;
  assign dataGroup_hi_hi_390 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_391;
  assign dataGroup_hi_hi_391 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_392;
  assign dataGroup_hi_hi_392 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_393;
  assign dataGroup_hi_hi_393 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_394;
  assign dataGroup_hi_hi_394 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_395;
  assign dataGroup_hi_hi_395 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_396;
  assign dataGroup_hi_hi_396 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_397;
  assign dataGroup_hi_hi_397 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_398;
  assign dataGroup_hi_hi_398 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_399;
  assign dataGroup_hi_hi_399 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_400;
  assign dataGroup_hi_hi_400 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_401;
  assign dataGroup_hi_hi_401 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_402;
  assign dataGroup_hi_hi_402 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_403;
  assign dataGroup_hi_hi_403 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_404;
  assign dataGroup_hi_hi_404 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_405;
  assign dataGroup_hi_hi_405 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_406;
  assign dataGroup_hi_hi_406 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_407;
  assign dataGroup_hi_hi_407 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_408;
  assign dataGroup_hi_hi_408 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_409;
  assign dataGroup_hi_hi_409 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_410;
  assign dataGroup_hi_hi_410 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_411;
  assign dataGroup_hi_hi_411 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_412;
  assign dataGroup_hi_hi_412 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_413;
  assign dataGroup_hi_hi_413 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_414;
  assign dataGroup_hi_hi_414 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_415;
  assign dataGroup_hi_hi_415 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_416;
  assign dataGroup_hi_hi_416 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_417;
  assign dataGroup_hi_hi_417 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_418;
  assign dataGroup_hi_hi_418 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_419;
  assign dataGroup_hi_hi_419 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_420;
  assign dataGroup_hi_hi_420 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_421;
  assign dataGroup_hi_hi_421 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_422;
  assign dataGroup_hi_hi_422 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_423;
  assign dataGroup_hi_hi_423 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_424;
  assign dataGroup_hi_hi_424 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_425;
  assign dataGroup_hi_hi_425 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_426;
  assign dataGroup_hi_hi_426 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_427;
  assign dataGroup_hi_hi_427 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_428;
  assign dataGroup_hi_hi_428 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_429;
  assign dataGroup_hi_hi_429 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_430;
  assign dataGroup_hi_hi_430 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_431;
  assign dataGroup_hi_hi_431 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_432;
  assign dataGroup_hi_hi_432 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_433;
  assign dataGroup_hi_hi_433 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_434;
  assign dataGroup_hi_hi_434 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_435;
  assign dataGroup_hi_hi_435 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_436;
  assign dataGroup_hi_hi_436 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_437;
  assign dataGroup_hi_hi_437 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_438;
  assign dataGroup_hi_hi_438 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_439;
  assign dataGroup_hi_hi_439 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_440;
  assign dataGroup_hi_hi_440 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_441;
  assign dataGroup_hi_hi_441 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_442;
  assign dataGroup_hi_hi_442 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_443;
  assign dataGroup_hi_hi_443 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_444;
  assign dataGroup_hi_hi_444 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_445;
  assign dataGroup_hi_hi_445 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_446;
  assign dataGroup_hi_hi_446 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_447;
  assign dataGroup_hi_hi_447 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_448;
  assign dataGroup_hi_hi_448 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_449;
  assign dataGroup_hi_hi_449 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_450;
  assign dataGroup_hi_hi_450 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_451;
  assign dataGroup_hi_hi_451 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_452;
  assign dataGroup_hi_hi_452 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_453;
  assign dataGroup_hi_hi_453 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_454;
  assign dataGroup_hi_hi_454 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_455;
  assign dataGroup_hi_hi_455 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_456;
  assign dataGroup_hi_hi_456 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_457;
  assign dataGroup_hi_hi_457 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_458;
  assign dataGroup_hi_hi_458 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_459;
  assign dataGroup_hi_hi_459 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_460;
  assign dataGroup_hi_hi_460 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_461;
  assign dataGroup_hi_hi_461 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_462;
  assign dataGroup_hi_hi_462 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_463;
  assign dataGroup_hi_hi_463 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_464;
  assign dataGroup_hi_hi_464 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_465;
  assign dataGroup_hi_hi_465 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_466;
  assign dataGroup_hi_hi_466 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_467;
  assign dataGroup_hi_hi_467 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_468;
  assign dataGroup_hi_hi_468 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_469;
  assign dataGroup_hi_hi_469 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_470;
  assign dataGroup_hi_hi_470 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_471;
  assign dataGroup_hi_hi_471 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_472;
  assign dataGroup_hi_hi_472 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_473;
  assign dataGroup_hi_hi_473 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_474;
  assign dataGroup_hi_hi_474 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_475;
  assign dataGroup_hi_hi_475 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_476;
  assign dataGroup_hi_hi_476 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_477;
  assign dataGroup_hi_hi_477 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_478;
  assign dataGroup_hi_hi_478 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_479;
  assign dataGroup_hi_hi_479 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_480;
  assign dataGroup_hi_hi_480 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_481;
  assign dataGroup_hi_hi_481 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_482;
  assign dataGroup_hi_hi_482 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_483;
  assign dataGroup_hi_hi_483 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_484;
  assign dataGroup_hi_hi_484 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_485;
  assign dataGroup_hi_hi_485 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_486;
  assign dataGroup_hi_hi_486 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_487;
  assign dataGroup_hi_hi_487 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_488;
  assign dataGroup_hi_hi_488 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_489;
  assign dataGroup_hi_hi_489 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_490;
  assign dataGroup_hi_hi_490 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_491;
  assign dataGroup_hi_hi_491 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_492;
  assign dataGroup_hi_hi_492 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_493;
  assign dataGroup_hi_hi_493 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_494;
  assign dataGroup_hi_hi_494 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_495;
  assign dataGroup_hi_hi_495 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_496;
  assign dataGroup_hi_hi_496 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_497;
  assign dataGroup_hi_hi_497 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_498;
  assign dataGroup_hi_hi_498 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_499;
  assign dataGroup_hi_hi_499 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_500;
  assign dataGroup_hi_hi_500 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_501;
  assign dataGroup_hi_hi_501 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_502;
  assign dataGroup_hi_hi_502 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_503;
  assign dataGroup_hi_hi_503 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_504;
  assign dataGroup_hi_hi_504 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_505;
  assign dataGroup_hi_hi_505 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_506;
  assign dataGroup_hi_hi_506 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_507;
  assign dataGroup_hi_hi_507 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_508;
  assign dataGroup_hi_hi_508 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_509;
  assign dataGroup_hi_hi_509 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_510;
  assign dataGroup_hi_hi_510 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_511;
  assign dataGroup_hi_hi_511 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_512;
  assign dataGroup_hi_hi_512 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_513;
  assign dataGroup_hi_hi_513 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_514;
  assign dataGroup_hi_hi_514 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_515;
  assign dataGroup_hi_hi_515 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_516;
  assign dataGroup_hi_hi_516 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_517;
  assign dataGroup_hi_hi_517 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_518;
  assign dataGroup_hi_hi_518 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_519;
  assign dataGroup_hi_hi_519 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_520;
  assign dataGroup_hi_hi_520 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_521;
  assign dataGroup_hi_hi_521 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_522;
  assign dataGroup_hi_hi_522 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_523;
  assign dataGroup_hi_hi_523 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_524;
  assign dataGroup_hi_hi_524 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_525;
  assign dataGroup_hi_hi_525 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_526;
  assign dataGroup_hi_hi_526 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_527;
  assign dataGroup_hi_hi_527 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_528;
  assign dataGroup_hi_hi_528 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_529;
  assign dataGroup_hi_hi_529 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_530;
  assign dataGroup_hi_hi_530 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_531;
  assign dataGroup_hi_hi_531 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_532;
  assign dataGroup_hi_hi_532 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_533;
  assign dataGroup_hi_hi_533 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_534;
  assign dataGroup_hi_hi_534 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_535;
  assign dataGroup_hi_hi_535 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_536;
  assign dataGroup_hi_hi_536 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_537;
  assign dataGroup_hi_hi_537 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_538;
  assign dataGroup_hi_hi_538 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_539;
  assign dataGroup_hi_hi_539 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_540;
  assign dataGroup_hi_hi_540 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_541;
  assign dataGroup_hi_hi_541 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_542;
  assign dataGroup_hi_hi_542 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_543;
  assign dataGroup_hi_hi_543 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_544;
  assign dataGroup_hi_hi_544 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_545;
  assign dataGroup_hi_hi_545 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_546;
  assign dataGroup_hi_hi_546 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_547;
  assign dataGroup_hi_hi_547 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_548;
  assign dataGroup_hi_hi_548 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_549;
  assign dataGroup_hi_hi_549 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_550;
  assign dataGroup_hi_hi_550 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_551;
  assign dataGroup_hi_hi_551 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_552;
  assign dataGroup_hi_hi_552 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_553;
  assign dataGroup_hi_hi_553 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_554;
  assign dataGroup_hi_hi_554 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_555;
  assign dataGroup_hi_hi_555 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_556;
  assign dataGroup_hi_hi_556 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_557;
  assign dataGroup_hi_hi_557 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_558;
  assign dataGroup_hi_hi_558 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_559;
  assign dataGroup_hi_hi_559 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_560;
  assign dataGroup_hi_hi_560 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_561;
  assign dataGroup_hi_hi_561 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_562;
  assign dataGroup_hi_hi_562 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_563;
  assign dataGroup_hi_hi_563 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_564;
  assign dataGroup_hi_hi_564 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_565;
  assign dataGroup_hi_hi_565 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_566;
  assign dataGroup_hi_hi_566 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_567;
  assign dataGroup_hi_hi_567 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_568;
  assign dataGroup_hi_hi_568 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_569;
  assign dataGroup_hi_hi_569 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_570;
  assign dataGroup_hi_hi_570 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_571;
  assign dataGroup_hi_hi_571 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_572;
  assign dataGroup_hi_hi_572 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_573;
  assign dataGroup_hi_hi_573 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_574;
  assign dataGroup_hi_hi_574 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_575;
  assign dataGroup_hi_hi_575 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_576;
  assign dataGroup_hi_hi_576 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_577;
  assign dataGroup_hi_hi_577 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_578;
  assign dataGroup_hi_hi_578 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_579;
  assign dataGroup_hi_hi_579 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_580;
  assign dataGroup_hi_hi_580 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_581;
  assign dataGroup_hi_hi_581 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_582;
  assign dataGroup_hi_hi_582 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_583;
  assign dataGroup_hi_hi_583 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_584;
  assign dataGroup_hi_hi_584 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_585;
  assign dataGroup_hi_hi_585 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_586;
  assign dataGroup_hi_hi_586 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_587;
  assign dataGroup_hi_hi_587 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_588;
  assign dataGroup_hi_hi_588 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_589;
  assign dataGroup_hi_hi_589 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_590;
  assign dataGroup_hi_hi_590 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_591;
  assign dataGroup_hi_hi_591 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_592;
  assign dataGroup_hi_hi_592 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_593;
  assign dataGroup_hi_hi_593 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_594;
  assign dataGroup_hi_hi_594 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_595;
  assign dataGroup_hi_hi_595 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_596;
  assign dataGroup_hi_hi_596 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_597;
  assign dataGroup_hi_hi_597 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_598;
  assign dataGroup_hi_hi_598 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_599;
  assign dataGroup_hi_hi_599 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_600;
  assign dataGroup_hi_hi_600 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_601;
  assign dataGroup_hi_hi_601 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_602;
  assign dataGroup_hi_hi_602 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_603;
  assign dataGroup_hi_hi_603 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_604;
  assign dataGroup_hi_hi_604 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_605;
  assign dataGroup_hi_hi_605 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_606;
  assign dataGroup_hi_hi_606 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_607;
  assign dataGroup_hi_hi_607 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_608;
  assign dataGroup_hi_hi_608 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_609;
  assign dataGroup_hi_hi_609 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_610;
  assign dataGroup_hi_hi_610 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_611;
  assign dataGroup_hi_hi_611 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_612;
  assign dataGroup_hi_hi_612 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_613;
  assign dataGroup_hi_hi_613 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_614;
  assign dataGroup_hi_hi_614 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_615;
  assign dataGroup_hi_hi_615 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_616;
  assign dataGroup_hi_hi_616 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_617;
  assign dataGroup_hi_hi_617 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_618;
  assign dataGroup_hi_hi_618 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_619;
  assign dataGroup_hi_hi_619 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_620;
  assign dataGroup_hi_hi_620 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_621;
  assign dataGroup_hi_hi_621 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_622;
  assign dataGroup_hi_hi_622 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_623;
  assign dataGroup_hi_hi_623 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_624;
  assign dataGroup_hi_hi_624 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_625;
  assign dataGroup_hi_hi_625 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_626;
  assign dataGroup_hi_hi_626 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_627;
  assign dataGroup_hi_hi_627 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_628;
  assign dataGroup_hi_hi_628 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_629;
  assign dataGroup_hi_hi_629 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_630;
  assign dataGroup_hi_hi_630 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_631;
  assign dataGroup_hi_hi_631 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_632;
  assign dataGroup_hi_hi_632 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_633;
  assign dataGroup_hi_hi_633 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_634;
  assign dataGroup_hi_hi_634 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_635;
  assign dataGroup_hi_hi_635 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_636;
  assign dataGroup_hi_hi_636 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_637;
  assign dataGroup_hi_hi_637 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_638;
  assign dataGroup_hi_hi_638 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_639;
  assign dataGroup_hi_hi_639 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_640;
  assign dataGroup_hi_hi_640 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_641;
  assign dataGroup_hi_hi_641 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_642;
  assign dataGroup_hi_hi_642 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_643;
  assign dataGroup_hi_hi_643 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_644;
  assign dataGroup_hi_hi_644 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_645;
  assign dataGroup_hi_hi_645 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_646;
  assign dataGroup_hi_hi_646 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_647;
  assign dataGroup_hi_hi_647 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_648;
  assign dataGroup_hi_hi_648 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_649;
  assign dataGroup_hi_hi_649 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_650;
  assign dataGroup_hi_hi_650 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_651;
  assign dataGroup_hi_hi_651 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_652;
  assign dataGroup_hi_hi_652 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_653;
  assign dataGroup_hi_hi_653 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_654;
  assign dataGroup_hi_hi_654 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_655;
  assign dataGroup_hi_hi_655 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_656;
  assign dataGroup_hi_hi_656 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_657;
  assign dataGroup_hi_hi_657 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_658;
  assign dataGroup_hi_hi_658 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_659;
  assign dataGroup_hi_hi_659 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_660;
  assign dataGroup_hi_hi_660 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_661;
  assign dataGroup_hi_hi_661 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_662;
  assign dataGroup_hi_hi_662 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_663;
  assign dataGroup_hi_hi_663 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_664;
  assign dataGroup_hi_hi_664 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_665;
  assign dataGroup_hi_hi_665 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_666;
  assign dataGroup_hi_hi_666 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_667;
  assign dataGroup_hi_hi_667 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_668;
  assign dataGroup_hi_hi_668 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_669;
  assign dataGroup_hi_hi_669 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_670;
  assign dataGroup_hi_hi_670 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_671;
  assign dataGroup_hi_hi_671 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_672;
  assign dataGroup_hi_hi_672 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_673;
  assign dataGroup_hi_hi_673 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_674;
  assign dataGroup_hi_hi_674 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_675;
  assign dataGroup_hi_hi_675 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_676;
  assign dataGroup_hi_hi_676 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_677;
  assign dataGroup_hi_hi_677 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_678;
  assign dataGroup_hi_hi_678 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_679;
  assign dataGroup_hi_hi_679 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_680;
  assign dataGroup_hi_hi_680 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_681;
  assign dataGroup_hi_hi_681 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_682;
  assign dataGroup_hi_hi_682 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_683;
  assign dataGroup_hi_hi_683 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_684;
  assign dataGroup_hi_hi_684 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_685;
  assign dataGroup_hi_hi_685 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_686;
  assign dataGroup_hi_hi_686 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_687;
  assign dataGroup_hi_hi_687 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_688;
  assign dataGroup_hi_hi_688 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_689;
  assign dataGroup_hi_hi_689 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_690;
  assign dataGroup_hi_hi_690 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_691;
  assign dataGroup_hi_hi_691 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_692;
  assign dataGroup_hi_hi_692 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_693;
  assign dataGroup_hi_hi_693 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_694;
  assign dataGroup_hi_hi_694 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_695;
  assign dataGroup_hi_hi_695 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_696;
  assign dataGroup_hi_hi_696 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_697;
  assign dataGroup_hi_hi_697 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_698;
  assign dataGroup_hi_hi_698 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_699;
  assign dataGroup_hi_hi_699 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_700;
  assign dataGroup_hi_hi_700 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_701;
  assign dataGroup_hi_hi_701 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_702;
  assign dataGroup_hi_hi_702 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_703;
  assign dataGroup_hi_hi_703 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_704;
  assign dataGroup_hi_hi_704 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_705;
  assign dataGroup_hi_hi_705 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_706;
  assign dataGroup_hi_hi_706 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_707;
  assign dataGroup_hi_hi_707 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_708;
  assign dataGroup_hi_hi_708 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_709;
  assign dataGroup_hi_hi_709 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_710;
  assign dataGroup_hi_hi_710 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_711;
  assign dataGroup_hi_hi_711 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_712;
  assign dataGroup_hi_hi_712 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_713;
  assign dataGroup_hi_hi_713 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_714;
  assign dataGroup_hi_hi_714 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_715;
  assign dataGroup_hi_hi_715 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_716;
  assign dataGroup_hi_hi_716 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_717;
  assign dataGroup_hi_hi_717 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_718;
  assign dataGroup_hi_hi_718 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_719;
  assign dataGroup_hi_hi_719 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_720;
  assign dataGroup_hi_hi_720 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_721;
  assign dataGroup_hi_hi_721 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_722;
  assign dataGroup_hi_hi_722 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_723;
  assign dataGroup_hi_hi_723 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_724;
  assign dataGroup_hi_hi_724 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_725;
  assign dataGroup_hi_hi_725 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_726;
  assign dataGroup_hi_hi_726 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_727;
  assign dataGroup_hi_hi_727 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_728;
  assign dataGroup_hi_hi_728 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_729;
  assign dataGroup_hi_hi_729 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_730;
  assign dataGroup_hi_hi_730 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_731;
  assign dataGroup_hi_hi_731 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_732;
  assign dataGroup_hi_hi_732 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_733;
  assign dataGroup_hi_hi_733 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_734;
  assign dataGroup_hi_hi_734 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_735;
  assign dataGroup_hi_hi_735 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_736;
  assign dataGroup_hi_hi_736 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_737;
  assign dataGroup_hi_hi_737 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_738;
  assign dataGroup_hi_hi_738 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_739;
  assign dataGroup_hi_hi_739 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_740;
  assign dataGroup_hi_hi_740 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_741;
  assign dataGroup_hi_hi_741 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_742;
  assign dataGroup_hi_hi_742 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_743;
  assign dataGroup_hi_hi_743 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_744;
  assign dataGroup_hi_hi_744 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_745;
  assign dataGroup_hi_hi_745 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_746;
  assign dataGroup_hi_hi_746 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_747;
  assign dataGroup_hi_hi_747 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_748;
  assign dataGroup_hi_hi_748 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_749;
  assign dataGroup_hi_hi_749 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_750;
  assign dataGroup_hi_hi_750 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_751;
  assign dataGroup_hi_hi_751 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_752;
  assign dataGroup_hi_hi_752 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_753;
  assign dataGroup_hi_hi_753 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_754;
  assign dataGroup_hi_hi_754 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_755;
  assign dataGroup_hi_hi_755 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_756;
  assign dataGroup_hi_hi_756 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_757;
  assign dataGroup_hi_hi_757 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_758;
  assign dataGroup_hi_hi_758 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_759;
  assign dataGroup_hi_hi_759 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_760;
  assign dataGroup_hi_hi_760 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_761;
  assign dataGroup_hi_hi_761 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_762;
  assign dataGroup_hi_hi_762 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_763;
  assign dataGroup_hi_hi_763 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_764;
  assign dataGroup_hi_hi_764 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_765;
  assign dataGroup_hi_hi_765 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_766;
  assign dataGroup_hi_hi_766 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_767;
  assign dataGroup_hi_hi_767 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_768;
  assign dataGroup_hi_hi_768 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_769;
  assign dataGroup_hi_hi_769 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_770;
  assign dataGroup_hi_hi_770 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_771;
  assign dataGroup_hi_hi_771 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_772;
  assign dataGroup_hi_hi_772 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_773;
  assign dataGroup_hi_hi_773 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_774;
  assign dataGroup_hi_hi_774 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_775;
  assign dataGroup_hi_hi_775 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_776;
  assign dataGroup_hi_hi_776 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_777;
  assign dataGroup_hi_hi_777 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_778;
  assign dataGroup_hi_hi_778 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_779;
  assign dataGroup_hi_hi_779 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_780;
  assign dataGroup_hi_hi_780 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_781;
  assign dataGroup_hi_hi_781 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_782;
  assign dataGroup_hi_hi_782 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_783;
  assign dataGroup_hi_hi_783 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_784;
  assign dataGroup_hi_hi_784 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_785;
  assign dataGroup_hi_hi_785 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_786;
  assign dataGroup_hi_hi_786 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_787;
  assign dataGroup_hi_hi_787 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_788;
  assign dataGroup_hi_hi_788 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_789;
  assign dataGroup_hi_hi_789 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_790;
  assign dataGroup_hi_hi_790 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_791;
  assign dataGroup_hi_hi_791 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_792;
  assign dataGroup_hi_hi_792 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_793;
  assign dataGroup_hi_hi_793 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_794;
  assign dataGroup_hi_hi_794 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_795;
  assign dataGroup_hi_hi_795 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_796;
  assign dataGroup_hi_hi_796 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_797;
  assign dataGroup_hi_hi_797 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_798;
  assign dataGroup_hi_hi_798 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_799;
  assign dataGroup_hi_hi_799 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_800;
  assign dataGroup_hi_hi_800 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_801;
  assign dataGroup_hi_hi_801 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_802;
  assign dataGroup_hi_hi_802 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_803;
  assign dataGroup_hi_hi_803 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_804;
  assign dataGroup_hi_hi_804 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_805;
  assign dataGroup_hi_hi_805 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_806;
  assign dataGroup_hi_hi_806 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_807;
  assign dataGroup_hi_hi_807 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_808;
  assign dataGroup_hi_hi_808 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_809;
  assign dataGroup_hi_hi_809 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_810;
  assign dataGroup_hi_hi_810 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_811;
  assign dataGroup_hi_hi_811 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_812;
  assign dataGroup_hi_hi_812 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_813;
  assign dataGroup_hi_hi_813 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_814;
  assign dataGroup_hi_hi_814 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_815;
  assign dataGroup_hi_hi_815 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_816;
  assign dataGroup_hi_hi_816 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_817;
  assign dataGroup_hi_hi_817 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_818;
  assign dataGroup_hi_hi_818 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_819;
  assign dataGroup_hi_hi_819 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_820;
  assign dataGroup_hi_hi_820 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_821;
  assign dataGroup_hi_hi_821 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_822;
  assign dataGroup_hi_hi_822 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_823;
  assign dataGroup_hi_hi_823 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_824;
  assign dataGroup_hi_hi_824 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_825;
  assign dataGroup_hi_hi_825 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_826;
  assign dataGroup_hi_hi_826 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_827;
  assign dataGroup_hi_hi_827 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_828;
  assign dataGroup_hi_hi_828 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_829;
  assign dataGroup_hi_hi_829 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_830;
  assign dataGroup_hi_hi_830 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_831;
  assign dataGroup_hi_hi_831 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_832;
  assign dataGroup_hi_hi_832 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_833;
  assign dataGroup_hi_hi_833 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_834;
  assign dataGroup_hi_hi_834 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_835;
  assign dataGroup_hi_hi_835 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_836;
  assign dataGroup_hi_hi_836 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_837;
  assign dataGroup_hi_hi_837 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_838;
  assign dataGroup_hi_hi_838 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_839;
  assign dataGroup_hi_hi_839 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_840;
  assign dataGroup_hi_hi_840 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_841;
  assign dataGroup_hi_hi_841 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_842;
  assign dataGroup_hi_hi_842 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_843;
  assign dataGroup_hi_hi_843 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_844;
  assign dataGroup_hi_hi_844 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_845;
  assign dataGroup_hi_hi_845 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_846;
  assign dataGroup_hi_hi_846 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_847;
  assign dataGroup_hi_hi_847 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_848;
  assign dataGroup_hi_hi_848 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_849;
  assign dataGroup_hi_hi_849 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_850;
  assign dataGroup_hi_hi_850 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_851;
  assign dataGroup_hi_hi_851 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_852;
  assign dataGroup_hi_hi_852 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_853;
  assign dataGroup_hi_hi_853 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_854;
  assign dataGroup_hi_hi_854 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_855;
  assign dataGroup_hi_hi_855 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_856;
  assign dataGroup_hi_hi_856 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_857;
  assign dataGroup_hi_hi_857 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_858;
  assign dataGroup_hi_hi_858 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_859;
  assign dataGroup_hi_hi_859 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_860;
  assign dataGroup_hi_hi_860 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_861;
  assign dataGroup_hi_hi_861 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_862;
  assign dataGroup_hi_hi_862 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_863;
  assign dataGroup_hi_hi_863 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_864;
  assign dataGroup_hi_hi_864 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_865;
  assign dataGroup_hi_hi_865 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_866;
  assign dataGroup_hi_hi_866 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_867;
  assign dataGroup_hi_hi_867 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_868;
  assign dataGroup_hi_hi_868 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_869;
  assign dataGroup_hi_hi_869 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_870;
  assign dataGroup_hi_hi_870 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_871;
  assign dataGroup_hi_hi_871 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_872;
  assign dataGroup_hi_hi_872 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_873;
  assign dataGroup_hi_hi_873 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_874;
  assign dataGroup_hi_hi_874 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_875;
  assign dataGroup_hi_hi_875 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_876;
  assign dataGroup_hi_hi_876 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_877;
  assign dataGroup_hi_hi_877 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_878;
  assign dataGroup_hi_hi_878 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_879;
  assign dataGroup_hi_hi_879 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_880;
  assign dataGroup_hi_hi_880 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_881;
  assign dataGroup_hi_hi_881 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_882;
  assign dataGroup_hi_hi_882 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_883;
  assign dataGroup_hi_hi_883 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_884;
  assign dataGroup_hi_hi_884 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_885;
  assign dataGroup_hi_hi_885 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_886;
  assign dataGroup_hi_hi_886 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_887;
  assign dataGroup_hi_hi_887 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_888;
  assign dataGroup_hi_hi_888 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_889;
  assign dataGroup_hi_hi_889 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_890;
  assign dataGroup_hi_hi_890 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_891;
  assign dataGroup_hi_hi_891 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_892;
  assign dataGroup_hi_hi_892 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_893;
  assign dataGroup_hi_hi_893 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_894;
  assign dataGroup_hi_hi_894 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_895;
  assign dataGroup_hi_hi_895 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_896;
  assign dataGroup_hi_hi_896 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_897;
  assign dataGroup_hi_hi_897 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_898;
  assign dataGroup_hi_hi_898 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_899;
  assign dataGroup_hi_hi_899 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_900;
  assign dataGroup_hi_hi_900 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_901;
  assign dataGroup_hi_hi_901 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_902;
  assign dataGroup_hi_hi_902 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_903;
  assign dataGroup_hi_hi_903 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_904;
  assign dataGroup_hi_hi_904 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_905;
  assign dataGroup_hi_hi_905 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_906;
  assign dataGroup_hi_hi_906 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_907;
  assign dataGroup_hi_hi_907 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_908;
  assign dataGroup_hi_hi_908 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_909;
  assign dataGroup_hi_hi_909 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_910;
  assign dataGroup_hi_hi_910 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_911;
  assign dataGroup_hi_hi_911 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_912;
  assign dataGroup_hi_hi_912 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_913;
  assign dataGroup_hi_hi_913 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_914;
  assign dataGroup_hi_hi_914 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_915;
  assign dataGroup_hi_hi_915 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_916;
  assign dataGroup_hi_hi_916 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_917;
  assign dataGroup_hi_hi_917 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_918;
  assign dataGroup_hi_hi_918 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_919;
  assign dataGroup_hi_hi_919 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_920;
  assign dataGroup_hi_hi_920 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_921;
  assign dataGroup_hi_hi_921 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_922;
  assign dataGroup_hi_hi_922 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_923;
  assign dataGroup_hi_hi_923 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_924;
  assign dataGroup_hi_hi_924 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_925;
  assign dataGroup_hi_hi_925 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_926;
  assign dataGroup_hi_hi_926 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_927;
  assign dataGroup_hi_hi_927 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_928;
  assign dataGroup_hi_hi_928 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_929;
  assign dataGroup_hi_hi_929 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_930;
  assign dataGroup_hi_hi_930 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_931;
  assign dataGroup_hi_hi_931 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_932;
  assign dataGroup_hi_hi_932 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_933;
  assign dataGroup_hi_hi_933 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_934;
  assign dataGroup_hi_hi_934 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_935;
  assign dataGroup_hi_hi_935 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_936;
  assign dataGroup_hi_hi_936 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_937;
  assign dataGroup_hi_hi_937 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_938;
  assign dataGroup_hi_hi_938 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_939;
  assign dataGroup_hi_hi_939 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_940;
  assign dataGroup_hi_hi_940 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_941;
  assign dataGroup_hi_hi_941 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_942;
  assign dataGroup_hi_hi_942 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_943;
  assign dataGroup_hi_hi_943 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_944;
  assign dataGroup_hi_hi_944 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_945;
  assign dataGroup_hi_hi_945 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_946;
  assign dataGroup_hi_hi_946 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_947;
  assign dataGroup_hi_hi_947 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_948;
  assign dataGroup_hi_hi_948 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_949;
  assign dataGroup_hi_hi_949 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_950;
  assign dataGroup_hi_hi_950 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_951;
  assign dataGroup_hi_hi_951 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_952;
  assign dataGroup_hi_hi_952 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_953;
  assign dataGroup_hi_hi_953 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_954;
  assign dataGroup_hi_hi_954 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_955;
  assign dataGroup_hi_hi_955 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_956;
  assign dataGroup_hi_hi_956 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_957;
  assign dataGroup_hi_hi_957 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_958;
  assign dataGroup_hi_hi_958 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_959;
  assign dataGroup_hi_hi_959 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_960;
  assign dataGroup_hi_hi_960 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_961;
  assign dataGroup_hi_hi_961 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_962;
  assign dataGroup_hi_hi_962 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_963;
  assign dataGroup_hi_hi_963 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_964;
  assign dataGroup_hi_hi_964 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_965;
  assign dataGroup_hi_hi_965 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_966;
  assign dataGroup_hi_hi_966 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_967;
  assign dataGroup_hi_hi_967 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_968;
  assign dataGroup_hi_hi_968 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_969;
  assign dataGroup_hi_hi_969 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_970;
  assign dataGroup_hi_hi_970 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_971;
  assign dataGroup_hi_hi_971 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_972;
  assign dataGroup_hi_hi_972 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_973;
  assign dataGroup_hi_hi_973 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_974;
  assign dataGroup_hi_hi_974 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_975;
  assign dataGroup_hi_hi_975 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_976;
  assign dataGroup_hi_hi_976 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_977;
  assign dataGroup_hi_hi_977 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_978;
  assign dataGroup_hi_hi_978 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_979;
  assign dataGroup_hi_hi_979 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_980;
  assign dataGroup_hi_hi_980 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_981;
  assign dataGroup_hi_hi_981 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_982;
  assign dataGroup_hi_hi_982 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_983;
  assign dataGroup_hi_hi_983 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_984;
  assign dataGroup_hi_hi_984 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_985;
  assign dataGroup_hi_hi_985 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_986;
  assign dataGroup_hi_hi_986 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_987;
  assign dataGroup_hi_hi_987 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_988;
  assign dataGroup_hi_hi_988 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_989;
  assign dataGroup_hi_hi_989 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_990;
  assign dataGroup_hi_hi_990 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_991;
  assign dataGroup_hi_hi_991 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_992;
  assign dataGroup_hi_hi_992 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_993;
  assign dataGroup_hi_hi_993 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_994;
  assign dataGroup_hi_hi_994 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_995;
  assign dataGroup_hi_hi_995 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_996;
  assign dataGroup_hi_hi_996 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_997;
  assign dataGroup_hi_hi_997 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_998;
  assign dataGroup_hi_hi_998 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_999;
  assign dataGroup_hi_hi_999 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1000;
  assign dataGroup_hi_hi_1000 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1001;
  assign dataGroup_hi_hi_1001 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1002;
  assign dataGroup_hi_hi_1002 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1003;
  assign dataGroup_hi_hi_1003 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1004;
  assign dataGroup_hi_hi_1004 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1005;
  assign dataGroup_hi_hi_1005 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1006;
  assign dataGroup_hi_hi_1006 = _GEN_6;
  wire [255:0]  dataGroup_hi_hi_1007;
  assign dataGroup_hi_hi_1007 = _GEN_6;
  wire [511:0]  dataGroup_hi = {dataGroup_hi_hi, dataGroup_hi_lo};
  wire [7:0]    dataGroup_0 = dataGroup_lo[7:0];
  wire [511:0]  dataGroup_lo_1 = {dataGroup_lo_hi_1, dataGroup_lo_lo_1};
  wire [511:0]  dataGroup_hi_1 = {dataGroup_hi_hi_1, dataGroup_hi_lo_1};
  wire [7:0]    dataGroup_1 = dataGroup_lo_1[15:8];
  wire [511:0]  dataGroup_lo_2 = {dataGroup_lo_hi_2, dataGroup_lo_lo_2};
  wire [511:0]  dataGroup_hi_2 = {dataGroup_hi_hi_2, dataGroup_hi_lo_2};
  wire [7:0]    dataGroup_2 = dataGroup_lo_2[23:16];
  wire [511:0]  dataGroup_lo_3 = {dataGroup_lo_hi_3, dataGroup_lo_lo_3};
  wire [511:0]  dataGroup_hi_3 = {dataGroup_hi_hi_3, dataGroup_hi_lo_3};
  wire [7:0]    dataGroup_3 = dataGroup_lo_3[31:24];
  wire [511:0]  dataGroup_lo_4 = {dataGroup_lo_hi_4, dataGroup_lo_lo_4};
  wire [511:0]  dataGroup_hi_4 = {dataGroup_hi_hi_4, dataGroup_hi_lo_4};
  wire [7:0]    dataGroup_4 = dataGroup_lo_4[39:32];
  wire [511:0]  dataGroup_lo_5 = {dataGroup_lo_hi_5, dataGroup_lo_lo_5};
  wire [511:0]  dataGroup_hi_5 = {dataGroup_hi_hi_5, dataGroup_hi_lo_5};
  wire [7:0]    dataGroup_5 = dataGroup_lo_5[47:40];
  wire [511:0]  dataGroup_lo_6 = {dataGroup_lo_hi_6, dataGroup_lo_lo_6};
  wire [511:0]  dataGroup_hi_6 = {dataGroup_hi_hi_6, dataGroup_hi_lo_6};
  wire [7:0]    dataGroup_6 = dataGroup_lo_6[55:48];
  wire [511:0]  dataGroup_lo_7 = {dataGroup_lo_hi_7, dataGroup_lo_lo_7};
  wire [511:0]  dataGroup_hi_7 = {dataGroup_hi_hi_7, dataGroup_hi_lo_7};
  wire [7:0]    dataGroup_7 = dataGroup_lo_7[63:56];
  wire [511:0]  dataGroup_lo_8 = {dataGroup_lo_hi_8, dataGroup_lo_lo_8};
  wire [511:0]  dataGroup_hi_8 = {dataGroup_hi_hi_8, dataGroup_hi_lo_8};
  wire [7:0]    dataGroup_8 = dataGroup_lo_8[71:64];
  wire [511:0]  dataGroup_lo_9 = {dataGroup_lo_hi_9, dataGroup_lo_lo_9};
  wire [511:0]  dataGroup_hi_9 = {dataGroup_hi_hi_9, dataGroup_hi_lo_9};
  wire [7:0]    dataGroup_9 = dataGroup_lo_9[79:72];
  wire [511:0]  dataGroup_lo_10 = {dataGroup_lo_hi_10, dataGroup_lo_lo_10};
  wire [511:0]  dataGroup_hi_10 = {dataGroup_hi_hi_10, dataGroup_hi_lo_10};
  wire [7:0]    dataGroup_10 = dataGroup_lo_10[87:80];
  wire [511:0]  dataGroup_lo_11 = {dataGroup_lo_hi_11, dataGroup_lo_lo_11};
  wire [511:0]  dataGroup_hi_11 = {dataGroup_hi_hi_11, dataGroup_hi_lo_11};
  wire [7:0]    dataGroup_11 = dataGroup_lo_11[95:88];
  wire [511:0]  dataGroup_lo_12 = {dataGroup_lo_hi_12, dataGroup_lo_lo_12};
  wire [511:0]  dataGroup_hi_12 = {dataGroup_hi_hi_12, dataGroup_hi_lo_12};
  wire [7:0]    dataGroup_12 = dataGroup_lo_12[103:96];
  wire [511:0]  dataGroup_lo_13 = {dataGroup_lo_hi_13, dataGroup_lo_lo_13};
  wire [511:0]  dataGroup_hi_13 = {dataGroup_hi_hi_13, dataGroup_hi_lo_13};
  wire [7:0]    dataGroup_13 = dataGroup_lo_13[111:104];
  wire [511:0]  dataGroup_lo_14 = {dataGroup_lo_hi_14, dataGroup_lo_lo_14};
  wire [511:0]  dataGroup_hi_14 = {dataGroup_hi_hi_14, dataGroup_hi_lo_14};
  wire [7:0]    dataGroup_14 = dataGroup_lo_14[119:112];
  wire [511:0]  dataGroup_lo_15 = {dataGroup_lo_hi_15, dataGroup_lo_lo_15};
  wire [511:0]  dataGroup_hi_15 = {dataGroup_hi_hi_15, dataGroup_hi_lo_15};
  wire [7:0]    dataGroup_15 = dataGroup_lo_15[127:120];
  wire [15:0]   res_lo_lo_lo = {dataGroup_1, dataGroup_0};
  wire [15:0]   res_lo_lo_hi = {dataGroup_3, dataGroup_2};
  wire [31:0]   res_lo_lo = {res_lo_lo_hi, res_lo_lo_lo};
  wire [15:0]   res_lo_hi_lo = {dataGroup_5, dataGroup_4};
  wire [15:0]   res_lo_hi_hi = {dataGroup_7, dataGroup_6};
  wire [31:0]   res_lo_hi = {res_lo_hi_hi, res_lo_hi_lo};
  wire [63:0]   res_lo = {res_lo_hi, res_lo_lo};
  wire [15:0]   res_hi_lo_lo = {dataGroup_9, dataGroup_8};
  wire [15:0]   res_hi_lo_hi = {dataGroup_11, dataGroup_10};
  wire [31:0]   res_hi_lo = {res_hi_lo_hi, res_hi_lo_lo};
  wire [15:0]   res_hi_hi_lo = {dataGroup_13, dataGroup_12};
  wire [15:0]   res_hi_hi_hi = {dataGroup_15, dataGroup_14};
  wire [31:0]   res_hi_hi = {res_hi_hi_hi, res_hi_hi_lo};
  wire [63:0]   res_hi = {res_hi_hi, res_hi_lo};
  wire [127:0]  res = {res_hi, res_lo};
  wire [255:0]  lo_lo = {128'h0, res};
  wire [511:0]  lo = {256'h0, lo_lo};
  wire [1023:0] regroupLoadData_0_0 = {512'h0, lo};
  wire [511:0]  dataGroup_lo_16 = {dataGroup_lo_hi_16, dataGroup_lo_lo_16};
  wire [511:0]  dataGroup_hi_16 = {dataGroup_hi_hi_16, dataGroup_hi_lo_16};
  wire [7:0]    dataGroup_0_1 = dataGroup_lo_16[7:0];
  wire [511:0]  dataGroup_lo_17 = {dataGroup_lo_hi_17, dataGroup_lo_lo_17};
  wire [511:0]  dataGroup_hi_17 = {dataGroup_hi_hi_17, dataGroup_hi_lo_17};
  wire [7:0]    dataGroup_1_1 = dataGroup_lo_17[23:16];
  wire [511:0]  dataGroup_lo_18 = {dataGroup_lo_hi_18, dataGroup_lo_lo_18};
  wire [511:0]  dataGroup_hi_18 = {dataGroup_hi_hi_18, dataGroup_hi_lo_18};
  wire [7:0]    dataGroup_2_1 = dataGroup_lo_18[39:32];
  wire [511:0]  dataGroup_lo_19 = {dataGroup_lo_hi_19, dataGroup_lo_lo_19};
  wire [511:0]  dataGroup_hi_19 = {dataGroup_hi_hi_19, dataGroup_hi_lo_19};
  wire [7:0]    dataGroup_3_1 = dataGroup_lo_19[55:48];
  wire [511:0]  dataGroup_lo_20 = {dataGroup_lo_hi_20, dataGroup_lo_lo_20};
  wire [511:0]  dataGroup_hi_20 = {dataGroup_hi_hi_20, dataGroup_hi_lo_20};
  wire [7:0]    dataGroup_4_1 = dataGroup_lo_20[71:64];
  wire [511:0]  dataGroup_lo_21 = {dataGroup_lo_hi_21, dataGroup_lo_lo_21};
  wire [511:0]  dataGroup_hi_21 = {dataGroup_hi_hi_21, dataGroup_hi_lo_21};
  wire [7:0]    dataGroup_5_1 = dataGroup_lo_21[87:80];
  wire [511:0]  dataGroup_lo_22 = {dataGroup_lo_hi_22, dataGroup_lo_lo_22};
  wire [511:0]  dataGroup_hi_22 = {dataGroup_hi_hi_22, dataGroup_hi_lo_22};
  wire [7:0]    dataGroup_6_1 = dataGroup_lo_22[103:96];
  wire [511:0]  dataGroup_lo_23 = {dataGroup_lo_hi_23, dataGroup_lo_lo_23};
  wire [511:0]  dataGroup_hi_23 = {dataGroup_hi_hi_23, dataGroup_hi_lo_23};
  wire [7:0]    dataGroup_7_1 = dataGroup_lo_23[119:112];
  wire [511:0]  dataGroup_lo_24 = {dataGroup_lo_hi_24, dataGroup_lo_lo_24};
  wire [511:0]  dataGroup_hi_24 = {dataGroup_hi_hi_24, dataGroup_hi_lo_24};
  wire [7:0]    dataGroup_8_1 = dataGroup_lo_24[135:128];
  wire [511:0]  dataGroup_lo_25 = {dataGroup_lo_hi_25, dataGroup_lo_lo_25};
  wire [511:0]  dataGroup_hi_25 = {dataGroup_hi_hi_25, dataGroup_hi_lo_25};
  wire [7:0]    dataGroup_9_1 = dataGroup_lo_25[151:144];
  wire [511:0]  dataGroup_lo_26 = {dataGroup_lo_hi_26, dataGroup_lo_lo_26};
  wire [511:0]  dataGroup_hi_26 = {dataGroup_hi_hi_26, dataGroup_hi_lo_26};
  wire [7:0]    dataGroup_10_1 = dataGroup_lo_26[167:160];
  wire [511:0]  dataGroup_lo_27 = {dataGroup_lo_hi_27, dataGroup_lo_lo_27};
  wire [511:0]  dataGroup_hi_27 = {dataGroup_hi_hi_27, dataGroup_hi_lo_27};
  wire [7:0]    dataGroup_11_1 = dataGroup_lo_27[183:176];
  wire [511:0]  dataGroup_lo_28 = {dataGroup_lo_hi_28, dataGroup_lo_lo_28};
  wire [511:0]  dataGroup_hi_28 = {dataGroup_hi_hi_28, dataGroup_hi_lo_28};
  wire [7:0]    dataGroup_12_1 = dataGroup_lo_28[199:192];
  wire [511:0]  dataGroup_lo_29 = {dataGroup_lo_hi_29, dataGroup_lo_lo_29};
  wire [511:0]  dataGroup_hi_29 = {dataGroup_hi_hi_29, dataGroup_hi_lo_29};
  wire [7:0]    dataGroup_13_1 = dataGroup_lo_29[215:208];
  wire [511:0]  dataGroup_lo_30 = {dataGroup_lo_hi_30, dataGroup_lo_lo_30};
  wire [511:0]  dataGroup_hi_30 = {dataGroup_hi_hi_30, dataGroup_hi_lo_30};
  wire [7:0]    dataGroup_14_1 = dataGroup_lo_30[231:224];
  wire [511:0]  dataGroup_lo_31 = {dataGroup_lo_hi_31, dataGroup_lo_lo_31};
  wire [511:0]  dataGroup_hi_31 = {dataGroup_hi_hi_31, dataGroup_hi_lo_31};
  wire [7:0]    dataGroup_15_1 = dataGroup_lo_31[247:240];
  wire [15:0]   res_lo_lo_lo_1 = {dataGroup_1_1, dataGroup_0_1};
  wire [15:0]   res_lo_lo_hi_1 = {dataGroup_3_1, dataGroup_2_1};
  wire [31:0]   res_lo_lo_1 = {res_lo_lo_hi_1, res_lo_lo_lo_1};
  wire [15:0]   res_lo_hi_lo_1 = {dataGroup_5_1, dataGroup_4_1};
  wire [15:0]   res_lo_hi_hi_1 = {dataGroup_7_1, dataGroup_6_1};
  wire [31:0]   res_lo_hi_1 = {res_lo_hi_hi_1, res_lo_hi_lo_1};
  wire [63:0]   res_lo_1 = {res_lo_hi_1, res_lo_lo_1};
  wire [15:0]   res_hi_lo_lo_1 = {dataGroup_9_1, dataGroup_8_1};
  wire [15:0]   res_hi_lo_hi_1 = {dataGroup_11_1, dataGroup_10_1};
  wire [31:0]   res_hi_lo_1 = {res_hi_lo_hi_1, res_hi_lo_lo_1};
  wire [15:0]   res_hi_hi_lo_1 = {dataGroup_13_1, dataGroup_12_1};
  wire [15:0]   res_hi_hi_hi_1 = {dataGroup_15_1, dataGroup_14_1};
  wire [31:0]   res_hi_hi_1 = {res_hi_hi_hi_1, res_hi_hi_lo_1};
  wire [63:0]   res_hi_1 = {res_hi_hi_1, res_hi_lo_1};
  wire [127:0]  res_8 = {res_hi_1, res_lo_1};
  wire [511:0]  dataGroup_lo_32 = {dataGroup_lo_hi_32, dataGroup_lo_lo_32};
  wire [511:0]  dataGroup_hi_32 = {dataGroup_hi_hi_32, dataGroup_hi_lo_32};
  wire [7:0]    dataGroup_0_2 = dataGroup_lo_32[15:8];
  wire [511:0]  dataGroup_lo_33 = {dataGroup_lo_hi_33, dataGroup_lo_lo_33};
  wire [511:0]  dataGroup_hi_33 = {dataGroup_hi_hi_33, dataGroup_hi_lo_33};
  wire [7:0]    dataGroup_1_2 = dataGroup_lo_33[31:24];
  wire [511:0]  dataGroup_lo_34 = {dataGroup_lo_hi_34, dataGroup_lo_lo_34};
  wire [511:0]  dataGroup_hi_34 = {dataGroup_hi_hi_34, dataGroup_hi_lo_34};
  wire [7:0]    dataGroup_2_2 = dataGroup_lo_34[47:40];
  wire [511:0]  dataGroup_lo_35 = {dataGroup_lo_hi_35, dataGroup_lo_lo_35};
  wire [511:0]  dataGroup_hi_35 = {dataGroup_hi_hi_35, dataGroup_hi_lo_35};
  wire [7:0]    dataGroup_3_2 = dataGroup_lo_35[63:56];
  wire [511:0]  dataGroup_lo_36 = {dataGroup_lo_hi_36, dataGroup_lo_lo_36};
  wire [511:0]  dataGroup_hi_36 = {dataGroup_hi_hi_36, dataGroup_hi_lo_36};
  wire [7:0]    dataGroup_4_2 = dataGroup_lo_36[79:72];
  wire [511:0]  dataGroup_lo_37 = {dataGroup_lo_hi_37, dataGroup_lo_lo_37};
  wire [511:0]  dataGroup_hi_37 = {dataGroup_hi_hi_37, dataGroup_hi_lo_37};
  wire [7:0]    dataGroup_5_2 = dataGroup_lo_37[95:88];
  wire [511:0]  dataGroup_lo_38 = {dataGroup_lo_hi_38, dataGroup_lo_lo_38};
  wire [511:0]  dataGroup_hi_38 = {dataGroup_hi_hi_38, dataGroup_hi_lo_38};
  wire [7:0]    dataGroup_6_2 = dataGroup_lo_38[111:104];
  wire [511:0]  dataGroup_lo_39 = {dataGroup_lo_hi_39, dataGroup_lo_lo_39};
  wire [511:0]  dataGroup_hi_39 = {dataGroup_hi_hi_39, dataGroup_hi_lo_39};
  wire [7:0]    dataGroup_7_2 = dataGroup_lo_39[127:120];
  wire [511:0]  dataGroup_lo_40 = {dataGroup_lo_hi_40, dataGroup_lo_lo_40};
  wire [511:0]  dataGroup_hi_40 = {dataGroup_hi_hi_40, dataGroup_hi_lo_40};
  wire [7:0]    dataGroup_8_2 = dataGroup_lo_40[143:136];
  wire [511:0]  dataGroup_lo_41 = {dataGroup_lo_hi_41, dataGroup_lo_lo_41};
  wire [511:0]  dataGroup_hi_41 = {dataGroup_hi_hi_41, dataGroup_hi_lo_41};
  wire [7:0]    dataGroup_9_2 = dataGroup_lo_41[159:152];
  wire [511:0]  dataGroup_lo_42 = {dataGroup_lo_hi_42, dataGroup_lo_lo_42};
  wire [511:0]  dataGroup_hi_42 = {dataGroup_hi_hi_42, dataGroup_hi_lo_42};
  wire [7:0]    dataGroup_10_2 = dataGroup_lo_42[175:168];
  wire [511:0]  dataGroup_lo_43 = {dataGroup_lo_hi_43, dataGroup_lo_lo_43};
  wire [511:0]  dataGroup_hi_43 = {dataGroup_hi_hi_43, dataGroup_hi_lo_43};
  wire [7:0]    dataGroup_11_2 = dataGroup_lo_43[191:184];
  wire [511:0]  dataGroup_lo_44 = {dataGroup_lo_hi_44, dataGroup_lo_lo_44};
  wire [511:0]  dataGroup_hi_44 = {dataGroup_hi_hi_44, dataGroup_hi_lo_44};
  wire [7:0]    dataGroup_12_2 = dataGroup_lo_44[207:200];
  wire [511:0]  dataGroup_lo_45 = {dataGroup_lo_hi_45, dataGroup_lo_lo_45};
  wire [511:0]  dataGroup_hi_45 = {dataGroup_hi_hi_45, dataGroup_hi_lo_45};
  wire [7:0]    dataGroup_13_2 = dataGroup_lo_45[223:216];
  wire [511:0]  dataGroup_lo_46 = {dataGroup_lo_hi_46, dataGroup_lo_lo_46};
  wire [511:0]  dataGroup_hi_46 = {dataGroup_hi_hi_46, dataGroup_hi_lo_46};
  wire [7:0]    dataGroup_14_2 = dataGroup_lo_46[239:232];
  wire [511:0]  dataGroup_lo_47 = {dataGroup_lo_hi_47, dataGroup_lo_lo_47};
  wire [511:0]  dataGroup_hi_47 = {dataGroup_hi_hi_47, dataGroup_hi_lo_47};
  wire [7:0]    dataGroup_15_2 = dataGroup_lo_47[255:248];
  wire [15:0]   res_lo_lo_lo_2 = {dataGroup_1_2, dataGroup_0_2};
  wire [15:0]   res_lo_lo_hi_2 = {dataGroup_3_2, dataGroup_2_2};
  wire [31:0]   res_lo_lo_2 = {res_lo_lo_hi_2, res_lo_lo_lo_2};
  wire [15:0]   res_lo_hi_lo_2 = {dataGroup_5_2, dataGroup_4_2};
  wire [15:0]   res_lo_hi_hi_2 = {dataGroup_7_2, dataGroup_6_2};
  wire [31:0]   res_lo_hi_2 = {res_lo_hi_hi_2, res_lo_hi_lo_2};
  wire [63:0]   res_lo_2 = {res_lo_hi_2, res_lo_lo_2};
  wire [15:0]   res_hi_lo_lo_2 = {dataGroup_9_2, dataGroup_8_2};
  wire [15:0]   res_hi_lo_hi_2 = {dataGroup_11_2, dataGroup_10_2};
  wire [31:0]   res_hi_lo_2 = {res_hi_lo_hi_2, res_hi_lo_lo_2};
  wire [15:0]   res_hi_hi_lo_2 = {dataGroup_13_2, dataGroup_12_2};
  wire [15:0]   res_hi_hi_hi_2 = {dataGroup_15_2, dataGroup_14_2};
  wire [31:0]   res_hi_hi_2 = {res_hi_hi_hi_2, res_hi_hi_lo_2};
  wire [63:0]   res_hi_2 = {res_hi_hi_2, res_hi_lo_2};
  wire [127:0]  res_9 = {res_hi_2, res_lo_2};
  wire [255:0]  lo_lo_1 = {res_9, res_8};
  wire [511:0]  lo_1 = {256'h0, lo_lo_1};
  wire [1023:0] regroupLoadData_0_1 = {512'h0, lo_1};
  wire [511:0]  dataGroup_lo_48 = {dataGroup_lo_hi_48, dataGroup_lo_lo_48};
  wire [511:0]  dataGroup_hi_48 = {dataGroup_hi_hi_48, dataGroup_hi_lo_48};
  wire [7:0]    dataGroup_0_3 = dataGroup_lo_48[7:0];
  wire [511:0]  dataGroup_lo_49 = {dataGroup_lo_hi_49, dataGroup_lo_lo_49};
  wire [511:0]  dataGroup_hi_49 = {dataGroup_hi_hi_49, dataGroup_hi_lo_49};
  wire [7:0]    dataGroup_1_3 = dataGroup_lo_49[31:24];
  wire [511:0]  dataGroup_lo_50 = {dataGroup_lo_hi_50, dataGroup_lo_lo_50};
  wire [511:0]  dataGroup_hi_50 = {dataGroup_hi_hi_50, dataGroup_hi_lo_50};
  wire [7:0]    dataGroup_2_3 = dataGroup_lo_50[55:48];
  wire [511:0]  dataGroup_lo_51 = {dataGroup_lo_hi_51, dataGroup_lo_lo_51};
  wire [511:0]  dataGroup_hi_51 = {dataGroup_hi_hi_51, dataGroup_hi_lo_51};
  wire [7:0]    dataGroup_3_3 = dataGroup_lo_51[79:72];
  wire [511:0]  dataGroup_lo_52 = {dataGroup_lo_hi_52, dataGroup_lo_lo_52};
  wire [511:0]  dataGroup_hi_52 = {dataGroup_hi_hi_52, dataGroup_hi_lo_52};
  wire [7:0]    dataGroup_4_3 = dataGroup_lo_52[103:96];
  wire [511:0]  dataGroup_lo_53 = {dataGroup_lo_hi_53, dataGroup_lo_lo_53};
  wire [511:0]  dataGroup_hi_53 = {dataGroup_hi_hi_53, dataGroup_hi_lo_53};
  wire [7:0]    dataGroup_5_3 = dataGroup_lo_53[127:120];
  wire [511:0]  dataGroup_lo_54 = {dataGroup_lo_hi_54, dataGroup_lo_lo_54};
  wire [511:0]  dataGroup_hi_54 = {dataGroup_hi_hi_54, dataGroup_hi_lo_54};
  wire [7:0]    dataGroup_6_3 = dataGroup_lo_54[151:144];
  wire [511:0]  dataGroup_lo_55 = {dataGroup_lo_hi_55, dataGroup_lo_lo_55};
  wire [511:0]  dataGroup_hi_55 = {dataGroup_hi_hi_55, dataGroup_hi_lo_55};
  wire [7:0]    dataGroup_7_3 = dataGroup_lo_55[175:168];
  wire [511:0]  dataGroup_lo_56 = {dataGroup_lo_hi_56, dataGroup_lo_lo_56};
  wire [511:0]  dataGroup_hi_56 = {dataGroup_hi_hi_56, dataGroup_hi_lo_56};
  wire [7:0]    dataGroup_8_3 = dataGroup_lo_56[199:192];
  wire [511:0]  dataGroup_lo_57 = {dataGroup_lo_hi_57, dataGroup_lo_lo_57};
  wire [511:0]  dataGroup_hi_57 = {dataGroup_hi_hi_57, dataGroup_hi_lo_57};
  wire [7:0]    dataGroup_9_3 = dataGroup_lo_57[223:216];
  wire [511:0]  dataGroup_lo_58 = {dataGroup_lo_hi_58, dataGroup_lo_lo_58};
  wire [511:0]  dataGroup_hi_58 = {dataGroup_hi_hi_58, dataGroup_hi_lo_58};
  wire [7:0]    dataGroup_10_3 = dataGroup_lo_58[247:240];
  wire [511:0]  dataGroup_lo_59 = {dataGroup_lo_hi_59, dataGroup_lo_lo_59};
  wire [511:0]  dataGroup_hi_59 = {dataGroup_hi_hi_59, dataGroup_hi_lo_59};
  wire [7:0]    dataGroup_11_3 = dataGroup_lo_59[271:264];
  wire [511:0]  dataGroup_lo_60 = {dataGroup_lo_hi_60, dataGroup_lo_lo_60};
  wire [511:0]  dataGroup_hi_60 = {dataGroup_hi_hi_60, dataGroup_hi_lo_60};
  wire [7:0]    dataGroup_12_3 = dataGroup_lo_60[295:288];
  wire [511:0]  dataGroup_lo_61 = {dataGroup_lo_hi_61, dataGroup_lo_lo_61};
  wire [511:0]  dataGroup_hi_61 = {dataGroup_hi_hi_61, dataGroup_hi_lo_61};
  wire [7:0]    dataGroup_13_3 = dataGroup_lo_61[319:312];
  wire [511:0]  dataGroup_lo_62 = {dataGroup_lo_hi_62, dataGroup_lo_lo_62};
  wire [511:0]  dataGroup_hi_62 = {dataGroup_hi_hi_62, dataGroup_hi_lo_62};
  wire [7:0]    dataGroup_14_3 = dataGroup_lo_62[343:336];
  wire [511:0]  dataGroup_lo_63 = {dataGroup_lo_hi_63, dataGroup_lo_lo_63};
  wire [511:0]  dataGroup_hi_63 = {dataGroup_hi_hi_63, dataGroup_hi_lo_63};
  wire [7:0]    dataGroup_15_3 = dataGroup_lo_63[367:360];
  wire [15:0]   res_lo_lo_lo_3 = {dataGroup_1_3, dataGroup_0_3};
  wire [15:0]   res_lo_lo_hi_3 = {dataGroup_3_3, dataGroup_2_3};
  wire [31:0]   res_lo_lo_3 = {res_lo_lo_hi_3, res_lo_lo_lo_3};
  wire [15:0]   res_lo_hi_lo_3 = {dataGroup_5_3, dataGroup_4_3};
  wire [15:0]   res_lo_hi_hi_3 = {dataGroup_7_3, dataGroup_6_3};
  wire [31:0]   res_lo_hi_3 = {res_lo_hi_hi_3, res_lo_hi_lo_3};
  wire [63:0]   res_lo_3 = {res_lo_hi_3, res_lo_lo_3};
  wire [15:0]   res_hi_lo_lo_3 = {dataGroup_9_3, dataGroup_8_3};
  wire [15:0]   res_hi_lo_hi_3 = {dataGroup_11_3, dataGroup_10_3};
  wire [31:0]   res_hi_lo_3 = {res_hi_lo_hi_3, res_hi_lo_lo_3};
  wire [15:0]   res_hi_hi_lo_3 = {dataGroup_13_3, dataGroup_12_3};
  wire [15:0]   res_hi_hi_hi_3 = {dataGroup_15_3, dataGroup_14_3};
  wire [31:0]   res_hi_hi_3 = {res_hi_hi_hi_3, res_hi_hi_lo_3};
  wire [63:0]   res_hi_3 = {res_hi_hi_3, res_hi_lo_3};
  wire [127:0]  res_16 = {res_hi_3, res_lo_3};
  wire [511:0]  dataGroup_lo_64 = {dataGroup_lo_hi_64, dataGroup_lo_lo_64};
  wire [511:0]  dataGroup_hi_64 = {dataGroup_hi_hi_64, dataGroup_hi_lo_64};
  wire [7:0]    dataGroup_0_4 = dataGroup_lo_64[15:8];
  wire [511:0]  dataGroup_lo_65 = {dataGroup_lo_hi_65, dataGroup_lo_lo_65};
  wire [511:0]  dataGroup_hi_65 = {dataGroup_hi_hi_65, dataGroup_hi_lo_65};
  wire [7:0]    dataGroup_1_4 = dataGroup_lo_65[39:32];
  wire [511:0]  dataGroup_lo_66 = {dataGroup_lo_hi_66, dataGroup_lo_lo_66};
  wire [511:0]  dataGroup_hi_66 = {dataGroup_hi_hi_66, dataGroup_hi_lo_66};
  wire [7:0]    dataGroup_2_4 = dataGroup_lo_66[63:56];
  wire [511:0]  dataGroup_lo_67 = {dataGroup_lo_hi_67, dataGroup_lo_lo_67};
  wire [511:0]  dataGroup_hi_67 = {dataGroup_hi_hi_67, dataGroup_hi_lo_67};
  wire [7:0]    dataGroup_3_4 = dataGroup_lo_67[87:80];
  wire [511:0]  dataGroup_lo_68 = {dataGroup_lo_hi_68, dataGroup_lo_lo_68};
  wire [511:0]  dataGroup_hi_68 = {dataGroup_hi_hi_68, dataGroup_hi_lo_68};
  wire [7:0]    dataGroup_4_4 = dataGroup_lo_68[111:104];
  wire [511:0]  dataGroup_lo_69 = {dataGroup_lo_hi_69, dataGroup_lo_lo_69};
  wire [511:0]  dataGroup_hi_69 = {dataGroup_hi_hi_69, dataGroup_hi_lo_69};
  wire [7:0]    dataGroup_5_4 = dataGroup_lo_69[135:128];
  wire [511:0]  dataGroup_lo_70 = {dataGroup_lo_hi_70, dataGroup_lo_lo_70};
  wire [511:0]  dataGroup_hi_70 = {dataGroup_hi_hi_70, dataGroup_hi_lo_70};
  wire [7:0]    dataGroup_6_4 = dataGroup_lo_70[159:152];
  wire [511:0]  dataGroup_lo_71 = {dataGroup_lo_hi_71, dataGroup_lo_lo_71};
  wire [511:0]  dataGroup_hi_71 = {dataGroup_hi_hi_71, dataGroup_hi_lo_71};
  wire [7:0]    dataGroup_7_4 = dataGroup_lo_71[183:176];
  wire [511:0]  dataGroup_lo_72 = {dataGroup_lo_hi_72, dataGroup_lo_lo_72};
  wire [511:0]  dataGroup_hi_72 = {dataGroup_hi_hi_72, dataGroup_hi_lo_72};
  wire [7:0]    dataGroup_8_4 = dataGroup_lo_72[207:200];
  wire [511:0]  dataGroup_lo_73 = {dataGroup_lo_hi_73, dataGroup_lo_lo_73};
  wire [511:0]  dataGroup_hi_73 = {dataGroup_hi_hi_73, dataGroup_hi_lo_73};
  wire [7:0]    dataGroup_9_4 = dataGroup_lo_73[231:224];
  wire [511:0]  dataGroup_lo_74 = {dataGroup_lo_hi_74, dataGroup_lo_lo_74};
  wire [511:0]  dataGroup_hi_74 = {dataGroup_hi_hi_74, dataGroup_hi_lo_74};
  wire [7:0]    dataGroup_10_4 = dataGroup_lo_74[255:248];
  wire [511:0]  dataGroup_lo_75 = {dataGroup_lo_hi_75, dataGroup_lo_lo_75};
  wire [511:0]  dataGroup_hi_75 = {dataGroup_hi_hi_75, dataGroup_hi_lo_75};
  wire [7:0]    dataGroup_11_4 = dataGroup_lo_75[279:272];
  wire [511:0]  dataGroup_lo_76 = {dataGroup_lo_hi_76, dataGroup_lo_lo_76};
  wire [511:0]  dataGroup_hi_76 = {dataGroup_hi_hi_76, dataGroup_hi_lo_76};
  wire [7:0]    dataGroup_12_4 = dataGroup_lo_76[303:296];
  wire [511:0]  dataGroup_lo_77 = {dataGroup_lo_hi_77, dataGroup_lo_lo_77};
  wire [511:0]  dataGroup_hi_77 = {dataGroup_hi_hi_77, dataGroup_hi_lo_77};
  wire [7:0]    dataGroup_13_4 = dataGroup_lo_77[327:320];
  wire [511:0]  dataGroup_lo_78 = {dataGroup_lo_hi_78, dataGroup_lo_lo_78};
  wire [511:0]  dataGroup_hi_78 = {dataGroup_hi_hi_78, dataGroup_hi_lo_78};
  wire [7:0]    dataGroup_14_4 = dataGroup_lo_78[351:344];
  wire [511:0]  dataGroup_lo_79 = {dataGroup_lo_hi_79, dataGroup_lo_lo_79};
  wire [511:0]  dataGroup_hi_79 = {dataGroup_hi_hi_79, dataGroup_hi_lo_79};
  wire [7:0]    dataGroup_15_4 = dataGroup_lo_79[375:368];
  wire [15:0]   res_lo_lo_lo_4 = {dataGroup_1_4, dataGroup_0_4};
  wire [15:0]   res_lo_lo_hi_4 = {dataGroup_3_4, dataGroup_2_4};
  wire [31:0]   res_lo_lo_4 = {res_lo_lo_hi_4, res_lo_lo_lo_4};
  wire [15:0]   res_lo_hi_lo_4 = {dataGroup_5_4, dataGroup_4_4};
  wire [15:0]   res_lo_hi_hi_4 = {dataGroup_7_4, dataGroup_6_4};
  wire [31:0]   res_lo_hi_4 = {res_lo_hi_hi_4, res_lo_hi_lo_4};
  wire [63:0]   res_lo_4 = {res_lo_hi_4, res_lo_lo_4};
  wire [15:0]   res_hi_lo_lo_4 = {dataGroup_9_4, dataGroup_8_4};
  wire [15:0]   res_hi_lo_hi_4 = {dataGroup_11_4, dataGroup_10_4};
  wire [31:0]   res_hi_lo_4 = {res_hi_lo_hi_4, res_hi_lo_lo_4};
  wire [15:0]   res_hi_hi_lo_4 = {dataGroup_13_4, dataGroup_12_4};
  wire [15:0]   res_hi_hi_hi_4 = {dataGroup_15_4, dataGroup_14_4};
  wire [31:0]   res_hi_hi_4 = {res_hi_hi_hi_4, res_hi_hi_lo_4};
  wire [63:0]   res_hi_4 = {res_hi_hi_4, res_hi_lo_4};
  wire [127:0]  res_17 = {res_hi_4, res_lo_4};
  wire [511:0]  dataGroup_lo_80 = {dataGroup_lo_hi_80, dataGroup_lo_lo_80};
  wire [511:0]  dataGroup_hi_80 = {dataGroup_hi_hi_80, dataGroup_hi_lo_80};
  wire [7:0]    dataGroup_0_5 = dataGroup_lo_80[23:16];
  wire [511:0]  dataGroup_lo_81 = {dataGroup_lo_hi_81, dataGroup_lo_lo_81};
  wire [511:0]  dataGroup_hi_81 = {dataGroup_hi_hi_81, dataGroup_hi_lo_81};
  wire [7:0]    dataGroup_1_5 = dataGroup_lo_81[47:40];
  wire [511:0]  dataGroup_lo_82 = {dataGroup_lo_hi_82, dataGroup_lo_lo_82};
  wire [511:0]  dataGroup_hi_82 = {dataGroup_hi_hi_82, dataGroup_hi_lo_82};
  wire [7:0]    dataGroup_2_5 = dataGroup_lo_82[71:64];
  wire [511:0]  dataGroup_lo_83 = {dataGroup_lo_hi_83, dataGroup_lo_lo_83};
  wire [511:0]  dataGroup_hi_83 = {dataGroup_hi_hi_83, dataGroup_hi_lo_83};
  wire [7:0]    dataGroup_3_5 = dataGroup_lo_83[95:88];
  wire [511:0]  dataGroup_lo_84 = {dataGroup_lo_hi_84, dataGroup_lo_lo_84};
  wire [511:0]  dataGroup_hi_84 = {dataGroup_hi_hi_84, dataGroup_hi_lo_84};
  wire [7:0]    dataGroup_4_5 = dataGroup_lo_84[119:112];
  wire [511:0]  dataGroup_lo_85 = {dataGroup_lo_hi_85, dataGroup_lo_lo_85};
  wire [511:0]  dataGroup_hi_85 = {dataGroup_hi_hi_85, dataGroup_hi_lo_85};
  wire [7:0]    dataGroup_5_5 = dataGroup_lo_85[143:136];
  wire [511:0]  dataGroup_lo_86 = {dataGroup_lo_hi_86, dataGroup_lo_lo_86};
  wire [511:0]  dataGroup_hi_86 = {dataGroup_hi_hi_86, dataGroup_hi_lo_86};
  wire [7:0]    dataGroup_6_5 = dataGroup_lo_86[167:160];
  wire [511:0]  dataGroup_lo_87 = {dataGroup_lo_hi_87, dataGroup_lo_lo_87};
  wire [511:0]  dataGroup_hi_87 = {dataGroup_hi_hi_87, dataGroup_hi_lo_87};
  wire [7:0]    dataGroup_7_5 = dataGroup_lo_87[191:184];
  wire [511:0]  dataGroup_lo_88 = {dataGroup_lo_hi_88, dataGroup_lo_lo_88};
  wire [511:0]  dataGroup_hi_88 = {dataGroup_hi_hi_88, dataGroup_hi_lo_88};
  wire [7:0]    dataGroup_8_5 = dataGroup_lo_88[215:208];
  wire [511:0]  dataGroup_lo_89 = {dataGroup_lo_hi_89, dataGroup_lo_lo_89};
  wire [511:0]  dataGroup_hi_89 = {dataGroup_hi_hi_89, dataGroup_hi_lo_89};
  wire [7:0]    dataGroup_9_5 = dataGroup_lo_89[239:232];
  wire [511:0]  dataGroup_lo_90 = {dataGroup_lo_hi_90, dataGroup_lo_lo_90};
  wire [511:0]  dataGroup_hi_90 = {dataGroup_hi_hi_90, dataGroup_hi_lo_90};
  wire [7:0]    dataGroup_10_5 = dataGroup_lo_90[263:256];
  wire [511:0]  dataGroup_lo_91 = {dataGroup_lo_hi_91, dataGroup_lo_lo_91};
  wire [511:0]  dataGroup_hi_91 = {dataGroup_hi_hi_91, dataGroup_hi_lo_91};
  wire [7:0]    dataGroup_11_5 = dataGroup_lo_91[287:280];
  wire [511:0]  dataGroup_lo_92 = {dataGroup_lo_hi_92, dataGroup_lo_lo_92};
  wire [511:0]  dataGroup_hi_92 = {dataGroup_hi_hi_92, dataGroup_hi_lo_92};
  wire [7:0]    dataGroup_12_5 = dataGroup_lo_92[311:304];
  wire [511:0]  dataGroup_lo_93 = {dataGroup_lo_hi_93, dataGroup_lo_lo_93};
  wire [511:0]  dataGroup_hi_93 = {dataGroup_hi_hi_93, dataGroup_hi_lo_93};
  wire [7:0]    dataGroup_13_5 = dataGroup_lo_93[335:328];
  wire [511:0]  dataGroup_lo_94 = {dataGroup_lo_hi_94, dataGroup_lo_lo_94};
  wire [511:0]  dataGroup_hi_94 = {dataGroup_hi_hi_94, dataGroup_hi_lo_94};
  wire [7:0]    dataGroup_14_5 = dataGroup_lo_94[359:352];
  wire [511:0]  dataGroup_lo_95 = {dataGroup_lo_hi_95, dataGroup_lo_lo_95};
  wire [511:0]  dataGroup_hi_95 = {dataGroup_hi_hi_95, dataGroup_hi_lo_95};
  wire [7:0]    dataGroup_15_5 = dataGroup_lo_95[383:376];
  wire [15:0]   res_lo_lo_lo_5 = {dataGroup_1_5, dataGroup_0_5};
  wire [15:0]   res_lo_lo_hi_5 = {dataGroup_3_5, dataGroup_2_5};
  wire [31:0]   res_lo_lo_5 = {res_lo_lo_hi_5, res_lo_lo_lo_5};
  wire [15:0]   res_lo_hi_lo_5 = {dataGroup_5_5, dataGroup_4_5};
  wire [15:0]   res_lo_hi_hi_5 = {dataGroup_7_5, dataGroup_6_5};
  wire [31:0]   res_lo_hi_5 = {res_lo_hi_hi_5, res_lo_hi_lo_5};
  wire [63:0]   res_lo_5 = {res_lo_hi_5, res_lo_lo_5};
  wire [15:0]   res_hi_lo_lo_5 = {dataGroup_9_5, dataGroup_8_5};
  wire [15:0]   res_hi_lo_hi_5 = {dataGroup_11_5, dataGroup_10_5};
  wire [31:0]   res_hi_lo_5 = {res_hi_lo_hi_5, res_hi_lo_lo_5};
  wire [15:0]   res_hi_hi_lo_5 = {dataGroup_13_5, dataGroup_12_5};
  wire [15:0]   res_hi_hi_hi_5 = {dataGroup_15_5, dataGroup_14_5};
  wire [31:0]   res_hi_hi_5 = {res_hi_hi_hi_5, res_hi_hi_lo_5};
  wire [63:0]   res_hi_5 = {res_hi_hi_5, res_hi_lo_5};
  wire [127:0]  res_18 = {res_hi_5, res_lo_5};
  wire [255:0]  lo_lo_2 = {res_17, res_16};
  wire [255:0]  lo_hi_2 = {128'h0, res_18};
  wire [511:0]  lo_2 = {lo_hi_2, lo_lo_2};
  wire [1023:0] regroupLoadData_0_2 = {512'h0, lo_2};
  wire [511:0]  dataGroup_lo_96 = {dataGroup_lo_hi_96, dataGroup_lo_lo_96};
  wire [511:0]  dataGroup_hi_96 = {dataGroup_hi_hi_96, dataGroup_hi_lo_96};
  wire [7:0]    dataGroup_0_6 = dataGroup_lo_96[7:0];
  wire [511:0]  dataGroup_lo_97 = {dataGroup_lo_hi_97, dataGroup_lo_lo_97};
  wire [511:0]  dataGroup_hi_97 = {dataGroup_hi_hi_97, dataGroup_hi_lo_97};
  wire [7:0]    dataGroup_1_6 = dataGroup_lo_97[39:32];
  wire [511:0]  dataGroup_lo_98 = {dataGroup_lo_hi_98, dataGroup_lo_lo_98};
  wire [511:0]  dataGroup_hi_98 = {dataGroup_hi_hi_98, dataGroup_hi_lo_98};
  wire [7:0]    dataGroup_2_6 = dataGroup_lo_98[71:64];
  wire [511:0]  dataGroup_lo_99 = {dataGroup_lo_hi_99, dataGroup_lo_lo_99};
  wire [511:0]  dataGroup_hi_99 = {dataGroup_hi_hi_99, dataGroup_hi_lo_99};
  wire [7:0]    dataGroup_3_6 = dataGroup_lo_99[103:96];
  wire [511:0]  dataGroup_lo_100 = {dataGroup_lo_hi_100, dataGroup_lo_lo_100};
  wire [511:0]  dataGroup_hi_100 = {dataGroup_hi_hi_100, dataGroup_hi_lo_100};
  wire [7:0]    dataGroup_4_6 = dataGroup_lo_100[135:128];
  wire [511:0]  dataGroup_lo_101 = {dataGroup_lo_hi_101, dataGroup_lo_lo_101};
  wire [511:0]  dataGroup_hi_101 = {dataGroup_hi_hi_101, dataGroup_hi_lo_101};
  wire [7:0]    dataGroup_5_6 = dataGroup_lo_101[167:160];
  wire [511:0]  dataGroup_lo_102 = {dataGroup_lo_hi_102, dataGroup_lo_lo_102};
  wire [511:0]  dataGroup_hi_102 = {dataGroup_hi_hi_102, dataGroup_hi_lo_102};
  wire [7:0]    dataGroup_6_6 = dataGroup_lo_102[199:192];
  wire [511:0]  dataGroup_lo_103 = {dataGroup_lo_hi_103, dataGroup_lo_lo_103};
  wire [511:0]  dataGroup_hi_103 = {dataGroup_hi_hi_103, dataGroup_hi_lo_103};
  wire [7:0]    dataGroup_7_6 = dataGroup_lo_103[231:224];
  wire [511:0]  dataGroup_lo_104 = {dataGroup_lo_hi_104, dataGroup_lo_lo_104};
  wire [511:0]  dataGroup_hi_104 = {dataGroup_hi_hi_104, dataGroup_hi_lo_104};
  wire [7:0]    dataGroup_8_6 = dataGroup_lo_104[263:256];
  wire [511:0]  dataGroup_lo_105 = {dataGroup_lo_hi_105, dataGroup_lo_lo_105};
  wire [511:0]  dataGroup_hi_105 = {dataGroup_hi_hi_105, dataGroup_hi_lo_105};
  wire [7:0]    dataGroup_9_6 = dataGroup_lo_105[295:288];
  wire [511:0]  dataGroup_lo_106 = {dataGroup_lo_hi_106, dataGroup_lo_lo_106};
  wire [511:0]  dataGroup_hi_106 = {dataGroup_hi_hi_106, dataGroup_hi_lo_106};
  wire [7:0]    dataGroup_10_6 = dataGroup_lo_106[327:320];
  wire [511:0]  dataGroup_lo_107 = {dataGroup_lo_hi_107, dataGroup_lo_lo_107};
  wire [511:0]  dataGroup_hi_107 = {dataGroup_hi_hi_107, dataGroup_hi_lo_107};
  wire [7:0]    dataGroup_11_6 = dataGroup_lo_107[359:352];
  wire [511:0]  dataGroup_lo_108 = {dataGroup_lo_hi_108, dataGroup_lo_lo_108};
  wire [511:0]  dataGroup_hi_108 = {dataGroup_hi_hi_108, dataGroup_hi_lo_108};
  wire [7:0]    dataGroup_12_6 = dataGroup_lo_108[391:384];
  wire [511:0]  dataGroup_lo_109 = {dataGroup_lo_hi_109, dataGroup_lo_lo_109};
  wire [511:0]  dataGroup_hi_109 = {dataGroup_hi_hi_109, dataGroup_hi_lo_109};
  wire [7:0]    dataGroup_13_6 = dataGroup_lo_109[423:416];
  wire [511:0]  dataGroup_lo_110 = {dataGroup_lo_hi_110, dataGroup_lo_lo_110};
  wire [511:0]  dataGroup_hi_110 = {dataGroup_hi_hi_110, dataGroup_hi_lo_110};
  wire [7:0]    dataGroup_14_6 = dataGroup_lo_110[455:448];
  wire [511:0]  dataGroup_lo_111 = {dataGroup_lo_hi_111, dataGroup_lo_lo_111};
  wire [511:0]  dataGroup_hi_111 = {dataGroup_hi_hi_111, dataGroup_hi_lo_111};
  wire [7:0]    dataGroup_15_6 = dataGroup_lo_111[487:480];
  wire [15:0]   res_lo_lo_lo_6 = {dataGroup_1_6, dataGroup_0_6};
  wire [15:0]   res_lo_lo_hi_6 = {dataGroup_3_6, dataGroup_2_6};
  wire [31:0]   res_lo_lo_6 = {res_lo_lo_hi_6, res_lo_lo_lo_6};
  wire [15:0]   res_lo_hi_lo_6 = {dataGroup_5_6, dataGroup_4_6};
  wire [15:0]   res_lo_hi_hi_6 = {dataGroup_7_6, dataGroup_6_6};
  wire [31:0]   res_lo_hi_6 = {res_lo_hi_hi_6, res_lo_hi_lo_6};
  wire [63:0]   res_lo_6 = {res_lo_hi_6, res_lo_lo_6};
  wire [15:0]   res_hi_lo_lo_6 = {dataGroup_9_6, dataGroup_8_6};
  wire [15:0]   res_hi_lo_hi_6 = {dataGroup_11_6, dataGroup_10_6};
  wire [31:0]   res_hi_lo_6 = {res_hi_lo_hi_6, res_hi_lo_lo_6};
  wire [15:0]   res_hi_hi_lo_6 = {dataGroup_13_6, dataGroup_12_6};
  wire [15:0]   res_hi_hi_hi_6 = {dataGroup_15_6, dataGroup_14_6};
  wire [31:0]   res_hi_hi_6 = {res_hi_hi_hi_6, res_hi_hi_lo_6};
  wire [63:0]   res_hi_6 = {res_hi_hi_6, res_hi_lo_6};
  wire [127:0]  res_24 = {res_hi_6, res_lo_6};
  wire [511:0]  dataGroup_lo_112 = {dataGroup_lo_hi_112, dataGroup_lo_lo_112};
  wire [511:0]  dataGroup_hi_112 = {dataGroup_hi_hi_112, dataGroup_hi_lo_112};
  wire [7:0]    dataGroup_0_7 = dataGroup_lo_112[15:8];
  wire [511:0]  dataGroup_lo_113 = {dataGroup_lo_hi_113, dataGroup_lo_lo_113};
  wire [511:0]  dataGroup_hi_113 = {dataGroup_hi_hi_113, dataGroup_hi_lo_113};
  wire [7:0]    dataGroup_1_7 = dataGroup_lo_113[47:40];
  wire [511:0]  dataGroup_lo_114 = {dataGroup_lo_hi_114, dataGroup_lo_lo_114};
  wire [511:0]  dataGroup_hi_114 = {dataGroup_hi_hi_114, dataGroup_hi_lo_114};
  wire [7:0]    dataGroup_2_7 = dataGroup_lo_114[79:72];
  wire [511:0]  dataGroup_lo_115 = {dataGroup_lo_hi_115, dataGroup_lo_lo_115};
  wire [511:0]  dataGroup_hi_115 = {dataGroup_hi_hi_115, dataGroup_hi_lo_115};
  wire [7:0]    dataGroup_3_7 = dataGroup_lo_115[111:104];
  wire [511:0]  dataGroup_lo_116 = {dataGroup_lo_hi_116, dataGroup_lo_lo_116};
  wire [511:0]  dataGroup_hi_116 = {dataGroup_hi_hi_116, dataGroup_hi_lo_116};
  wire [7:0]    dataGroup_4_7 = dataGroup_lo_116[143:136];
  wire [511:0]  dataGroup_lo_117 = {dataGroup_lo_hi_117, dataGroup_lo_lo_117};
  wire [511:0]  dataGroup_hi_117 = {dataGroup_hi_hi_117, dataGroup_hi_lo_117};
  wire [7:0]    dataGroup_5_7 = dataGroup_lo_117[175:168];
  wire [511:0]  dataGroup_lo_118 = {dataGroup_lo_hi_118, dataGroup_lo_lo_118};
  wire [511:0]  dataGroup_hi_118 = {dataGroup_hi_hi_118, dataGroup_hi_lo_118};
  wire [7:0]    dataGroup_6_7 = dataGroup_lo_118[207:200];
  wire [511:0]  dataGroup_lo_119 = {dataGroup_lo_hi_119, dataGroup_lo_lo_119};
  wire [511:0]  dataGroup_hi_119 = {dataGroup_hi_hi_119, dataGroup_hi_lo_119};
  wire [7:0]    dataGroup_7_7 = dataGroup_lo_119[239:232];
  wire [511:0]  dataGroup_lo_120 = {dataGroup_lo_hi_120, dataGroup_lo_lo_120};
  wire [511:0]  dataGroup_hi_120 = {dataGroup_hi_hi_120, dataGroup_hi_lo_120};
  wire [7:0]    dataGroup_8_7 = dataGroup_lo_120[271:264];
  wire [511:0]  dataGroup_lo_121 = {dataGroup_lo_hi_121, dataGroup_lo_lo_121};
  wire [511:0]  dataGroup_hi_121 = {dataGroup_hi_hi_121, dataGroup_hi_lo_121};
  wire [7:0]    dataGroup_9_7 = dataGroup_lo_121[303:296];
  wire [511:0]  dataGroup_lo_122 = {dataGroup_lo_hi_122, dataGroup_lo_lo_122};
  wire [511:0]  dataGroup_hi_122 = {dataGroup_hi_hi_122, dataGroup_hi_lo_122};
  wire [7:0]    dataGroup_10_7 = dataGroup_lo_122[335:328];
  wire [511:0]  dataGroup_lo_123 = {dataGroup_lo_hi_123, dataGroup_lo_lo_123};
  wire [511:0]  dataGroup_hi_123 = {dataGroup_hi_hi_123, dataGroup_hi_lo_123};
  wire [7:0]    dataGroup_11_7 = dataGroup_lo_123[367:360];
  wire [511:0]  dataGroup_lo_124 = {dataGroup_lo_hi_124, dataGroup_lo_lo_124};
  wire [511:0]  dataGroup_hi_124 = {dataGroup_hi_hi_124, dataGroup_hi_lo_124};
  wire [7:0]    dataGroup_12_7 = dataGroup_lo_124[399:392];
  wire [511:0]  dataGroup_lo_125 = {dataGroup_lo_hi_125, dataGroup_lo_lo_125};
  wire [511:0]  dataGroup_hi_125 = {dataGroup_hi_hi_125, dataGroup_hi_lo_125};
  wire [7:0]    dataGroup_13_7 = dataGroup_lo_125[431:424];
  wire [511:0]  dataGroup_lo_126 = {dataGroup_lo_hi_126, dataGroup_lo_lo_126};
  wire [511:0]  dataGroup_hi_126 = {dataGroup_hi_hi_126, dataGroup_hi_lo_126};
  wire [7:0]    dataGroup_14_7 = dataGroup_lo_126[463:456];
  wire [511:0]  dataGroup_lo_127 = {dataGroup_lo_hi_127, dataGroup_lo_lo_127};
  wire [511:0]  dataGroup_hi_127 = {dataGroup_hi_hi_127, dataGroup_hi_lo_127};
  wire [7:0]    dataGroup_15_7 = dataGroup_lo_127[495:488];
  wire [15:0]   res_lo_lo_lo_7 = {dataGroup_1_7, dataGroup_0_7};
  wire [15:0]   res_lo_lo_hi_7 = {dataGroup_3_7, dataGroup_2_7};
  wire [31:0]   res_lo_lo_7 = {res_lo_lo_hi_7, res_lo_lo_lo_7};
  wire [15:0]   res_lo_hi_lo_7 = {dataGroup_5_7, dataGroup_4_7};
  wire [15:0]   res_lo_hi_hi_7 = {dataGroup_7_7, dataGroup_6_7};
  wire [31:0]   res_lo_hi_7 = {res_lo_hi_hi_7, res_lo_hi_lo_7};
  wire [63:0]   res_lo_7 = {res_lo_hi_7, res_lo_lo_7};
  wire [15:0]   res_hi_lo_lo_7 = {dataGroup_9_7, dataGroup_8_7};
  wire [15:0]   res_hi_lo_hi_7 = {dataGroup_11_7, dataGroup_10_7};
  wire [31:0]   res_hi_lo_7 = {res_hi_lo_hi_7, res_hi_lo_lo_7};
  wire [15:0]   res_hi_hi_lo_7 = {dataGroup_13_7, dataGroup_12_7};
  wire [15:0]   res_hi_hi_hi_7 = {dataGroup_15_7, dataGroup_14_7};
  wire [31:0]   res_hi_hi_7 = {res_hi_hi_hi_7, res_hi_hi_lo_7};
  wire [63:0]   res_hi_7 = {res_hi_hi_7, res_hi_lo_7};
  wire [127:0]  res_25 = {res_hi_7, res_lo_7};
  wire [511:0]  dataGroup_lo_128 = {dataGroup_lo_hi_128, dataGroup_lo_lo_128};
  wire [511:0]  dataGroup_hi_128 = {dataGroup_hi_hi_128, dataGroup_hi_lo_128};
  wire [7:0]    dataGroup_0_8 = dataGroup_lo_128[23:16];
  wire [511:0]  dataGroup_lo_129 = {dataGroup_lo_hi_129, dataGroup_lo_lo_129};
  wire [511:0]  dataGroup_hi_129 = {dataGroup_hi_hi_129, dataGroup_hi_lo_129};
  wire [7:0]    dataGroup_1_8 = dataGroup_lo_129[55:48];
  wire [511:0]  dataGroup_lo_130 = {dataGroup_lo_hi_130, dataGroup_lo_lo_130};
  wire [511:0]  dataGroup_hi_130 = {dataGroup_hi_hi_130, dataGroup_hi_lo_130};
  wire [7:0]    dataGroup_2_8 = dataGroup_lo_130[87:80];
  wire [511:0]  dataGroup_lo_131 = {dataGroup_lo_hi_131, dataGroup_lo_lo_131};
  wire [511:0]  dataGroup_hi_131 = {dataGroup_hi_hi_131, dataGroup_hi_lo_131};
  wire [7:0]    dataGroup_3_8 = dataGroup_lo_131[119:112];
  wire [511:0]  dataGroup_lo_132 = {dataGroup_lo_hi_132, dataGroup_lo_lo_132};
  wire [511:0]  dataGroup_hi_132 = {dataGroup_hi_hi_132, dataGroup_hi_lo_132};
  wire [7:0]    dataGroup_4_8 = dataGroup_lo_132[151:144];
  wire [511:0]  dataGroup_lo_133 = {dataGroup_lo_hi_133, dataGroup_lo_lo_133};
  wire [511:0]  dataGroup_hi_133 = {dataGroup_hi_hi_133, dataGroup_hi_lo_133};
  wire [7:0]    dataGroup_5_8 = dataGroup_lo_133[183:176];
  wire [511:0]  dataGroup_lo_134 = {dataGroup_lo_hi_134, dataGroup_lo_lo_134};
  wire [511:0]  dataGroup_hi_134 = {dataGroup_hi_hi_134, dataGroup_hi_lo_134};
  wire [7:0]    dataGroup_6_8 = dataGroup_lo_134[215:208];
  wire [511:0]  dataGroup_lo_135 = {dataGroup_lo_hi_135, dataGroup_lo_lo_135};
  wire [511:0]  dataGroup_hi_135 = {dataGroup_hi_hi_135, dataGroup_hi_lo_135};
  wire [7:0]    dataGroup_7_8 = dataGroup_lo_135[247:240];
  wire [511:0]  dataGroup_lo_136 = {dataGroup_lo_hi_136, dataGroup_lo_lo_136};
  wire [511:0]  dataGroup_hi_136 = {dataGroup_hi_hi_136, dataGroup_hi_lo_136};
  wire [7:0]    dataGroup_8_8 = dataGroup_lo_136[279:272];
  wire [511:0]  dataGroup_lo_137 = {dataGroup_lo_hi_137, dataGroup_lo_lo_137};
  wire [511:0]  dataGroup_hi_137 = {dataGroup_hi_hi_137, dataGroup_hi_lo_137};
  wire [7:0]    dataGroup_9_8 = dataGroup_lo_137[311:304];
  wire [511:0]  dataGroup_lo_138 = {dataGroup_lo_hi_138, dataGroup_lo_lo_138};
  wire [511:0]  dataGroup_hi_138 = {dataGroup_hi_hi_138, dataGroup_hi_lo_138};
  wire [7:0]    dataGroup_10_8 = dataGroup_lo_138[343:336];
  wire [511:0]  dataGroup_lo_139 = {dataGroup_lo_hi_139, dataGroup_lo_lo_139};
  wire [511:0]  dataGroup_hi_139 = {dataGroup_hi_hi_139, dataGroup_hi_lo_139};
  wire [7:0]    dataGroup_11_8 = dataGroup_lo_139[375:368];
  wire [511:0]  dataGroup_lo_140 = {dataGroup_lo_hi_140, dataGroup_lo_lo_140};
  wire [511:0]  dataGroup_hi_140 = {dataGroup_hi_hi_140, dataGroup_hi_lo_140};
  wire [7:0]    dataGroup_12_8 = dataGroup_lo_140[407:400];
  wire [511:0]  dataGroup_lo_141 = {dataGroup_lo_hi_141, dataGroup_lo_lo_141};
  wire [511:0]  dataGroup_hi_141 = {dataGroup_hi_hi_141, dataGroup_hi_lo_141};
  wire [7:0]    dataGroup_13_8 = dataGroup_lo_141[439:432];
  wire [511:0]  dataGroup_lo_142 = {dataGroup_lo_hi_142, dataGroup_lo_lo_142};
  wire [511:0]  dataGroup_hi_142 = {dataGroup_hi_hi_142, dataGroup_hi_lo_142};
  wire [7:0]    dataGroup_14_8 = dataGroup_lo_142[471:464];
  wire [511:0]  dataGroup_lo_143 = {dataGroup_lo_hi_143, dataGroup_lo_lo_143};
  wire [511:0]  dataGroup_hi_143 = {dataGroup_hi_hi_143, dataGroup_hi_lo_143};
  wire [7:0]    dataGroup_15_8 = dataGroup_lo_143[503:496];
  wire [15:0]   res_lo_lo_lo_8 = {dataGroup_1_8, dataGroup_0_8};
  wire [15:0]   res_lo_lo_hi_8 = {dataGroup_3_8, dataGroup_2_8};
  wire [31:0]   res_lo_lo_8 = {res_lo_lo_hi_8, res_lo_lo_lo_8};
  wire [15:0]   res_lo_hi_lo_8 = {dataGroup_5_8, dataGroup_4_8};
  wire [15:0]   res_lo_hi_hi_8 = {dataGroup_7_8, dataGroup_6_8};
  wire [31:0]   res_lo_hi_8 = {res_lo_hi_hi_8, res_lo_hi_lo_8};
  wire [63:0]   res_lo_8 = {res_lo_hi_8, res_lo_lo_8};
  wire [15:0]   res_hi_lo_lo_8 = {dataGroup_9_8, dataGroup_8_8};
  wire [15:0]   res_hi_lo_hi_8 = {dataGroup_11_8, dataGroup_10_8};
  wire [31:0]   res_hi_lo_8 = {res_hi_lo_hi_8, res_hi_lo_lo_8};
  wire [15:0]   res_hi_hi_lo_8 = {dataGroup_13_8, dataGroup_12_8};
  wire [15:0]   res_hi_hi_hi_8 = {dataGroup_15_8, dataGroup_14_8};
  wire [31:0]   res_hi_hi_8 = {res_hi_hi_hi_8, res_hi_hi_lo_8};
  wire [63:0]   res_hi_8 = {res_hi_hi_8, res_hi_lo_8};
  wire [127:0]  res_26 = {res_hi_8, res_lo_8};
  wire [511:0]  dataGroup_lo_144 = {dataGroup_lo_hi_144, dataGroup_lo_lo_144};
  wire [511:0]  dataGroup_hi_144 = {dataGroup_hi_hi_144, dataGroup_hi_lo_144};
  wire [7:0]    dataGroup_0_9 = dataGroup_lo_144[31:24];
  wire [511:0]  dataGroup_lo_145 = {dataGroup_lo_hi_145, dataGroup_lo_lo_145};
  wire [511:0]  dataGroup_hi_145 = {dataGroup_hi_hi_145, dataGroup_hi_lo_145};
  wire [7:0]    dataGroup_1_9 = dataGroup_lo_145[63:56];
  wire [511:0]  dataGroup_lo_146 = {dataGroup_lo_hi_146, dataGroup_lo_lo_146};
  wire [511:0]  dataGroup_hi_146 = {dataGroup_hi_hi_146, dataGroup_hi_lo_146};
  wire [7:0]    dataGroup_2_9 = dataGroup_lo_146[95:88];
  wire [511:0]  dataGroup_lo_147 = {dataGroup_lo_hi_147, dataGroup_lo_lo_147};
  wire [511:0]  dataGroup_hi_147 = {dataGroup_hi_hi_147, dataGroup_hi_lo_147};
  wire [7:0]    dataGroup_3_9 = dataGroup_lo_147[127:120];
  wire [511:0]  dataGroup_lo_148 = {dataGroup_lo_hi_148, dataGroup_lo_lo_148};
  wire [511:0]  dataGroup_hi_148 = {dataGroup_hi_hi_148, dataGroup_hi_lo_148};
  wire [7:0]    dataGroup_4_9 = dataGroup_lo_148[159:152];
  wire [511:0]  dataGroup_lo_149 = {dataGroup_lo_hi_149, dataGroup_lo_lo_149};
  wire [511:0]  dataGroup_hi_149 = {dataGroup_hi_hi_149, dataGroup_hi_lo_149};
  wire [7:0]    dataGroup_5_9 = dataGroup_lo_149[191:184];
  wire [511:0]  dataGroup_lo_150 = {dataGroup_lo_hi_150, dataGroup_lo_lo_150};
  wire [511:0]  dataGroup_hi_150 = {dataGroup_hi_hi_150, dataGroup_hi_lo_150};
  wire [7:0]    dataGroup_6_9 = dataGroup_lo_150[223:216];
  wire [511:0]  dataGroup_lo_151 = {dataGroup_lo_hi_151, dataGroup_lo_lo_151};
  wire [511:0]  dataGroup_hi_151 = {dataGroup_hi_hi_151, dataGroup_hi_lo_151};
  wire [7:0]    dataGroup_7_9 = dataGroup_lo_151[255:248];
  wire [511:0]  dataGroup_lo_152 = {dataGroup_lo_hi_152, dataGroup_lo_lo_152};
  wire [511:0]  dataGroup_hi_152 = {dataGroup_hi_hi_152, dataGroup_hi_lo_152};
  wire [7:0]    dataGroup_8_9 = dataGroup_lo_152[287:280];
  wire [511:0]  dataGroup_lo_153 = {dataGroup_lo_hi_153, dataGroup_lo_lo_153};
  wire [511:0]  dataGroup_hi_153 = {dataGroup_hi_hi_153, dataGroup_hi_lo_153};
  wire [7:0]    dataGroup_9_9 = dataGroup_lo_153[319:312];
  wire [511:0]  dataGroup_lo_154 = {dataGroup_lo_hi_154, dataGroup_lo_lo_154};
  wire [511:0]  dataGroup_hi_154 = {dataGroup_hi_hi_154, dataGroup_hi_lo_154};
  wire [7:0]    dataGroup_10_9 = dataGroup_lo_154[351:344];
  wire [511:0]  dataGroup_lo_155 = {dataGroup_lo_hi_155, dataGroup_lo_lo_155};
  wire [511:0]  dataGroup_hi_155 = {dataGroup_hi_hi_155, dataGroup_hi_lo_155};
  wire [7:0]    dataGroup_11_9 = dataGroup_lo_155[383:376];
  wire [511:0]  dataGroup_lo_156 = {dataGroup_lo_hi_156, dataGroup_lo_lo_156};
  wire [511:0]  dataGroup_hi_156 = {dataGroup_hi_hi_156, dataGroup_hi_lo_156};
  wire [7:0]    dataGroup_12_9 = dataGroup_lo_156[415:408];
  wire [511:0]  dataGroup_lo_157 = {dataGroup_lo_hi_157, dataGroup_lo_lo_157};
  wire [511:0]  dataGroup_hi_157 = {dataGroup_hi_hi_157, dataGroup_hi_lo_157};
  wire [7:0]    dataGroup_13_9 = dataGroup_lo_157[447:440];
  wire [511:0]  dataGroup_lo_158 = {dataGroup_lo_hi_158, dataGroup_lo_lo_158};
  wire [511:0]  dataGroup_hi_158 = {dataGroup_hi_hi_158, dataGroup_hi_lo_158};
  wire [7:0]    dataGroup_14_9 = dataGroup_lo_158[479:472];
  wire [511:0]  dataGroup_lo_159 = {dataGroup_lo_hi_159, dataGroup_lo_lo_159};
  wire [511:0]  dataGroup_hi_159 = {dataGroup_hi_hi_159, dataGroup_hi_lo_159};
  wire [7:0]    dataGroup_15_9 = dataGroup_lo_159[511:504];
  wire [15:0]   res_lo_lo_lo_9 = {dataGroup_1_9, dataGroup_0_9};
  wire [15:0]   res_lo_lo_hi_9 = {dataGroup_3_9, dataGroup_2_9};
  wire [31:0]   res_lo_lo_9 = {res_lo_lo_hi_9, res_lo_lo_lo_9};
  wire [15:0]   res_lo_hi_lo_9 = {dataGroup_5_9, dataGroup_4_9};
  wire [15:0]   res_lo_hi_hi_9 = {dataGroup_7_9, dataGroup_6_9};
  wire [31:0]   res_lo_hi_9 = {res_lo_hi_hi_9, res_lo_hi_lo_9};
  wire [63:0]   res_lo_9 = {res_lo_hi_9, res_lo_lo_9};
  wire [15:0]   res_hi_lo_lo_9 = {dataGroup_9_9, dataGroup_8_9};
  wire [15:0]   res_hi_lo_hi_9 = {dataGroup_11_9, dataGroup_10_9};
  wire [31:0]   res_hi_lo_9 = {res_hi_lo_hi_9, res_hi_lo_lo_9};
  wire [15:0]   res_hi_hi_lo_9 = {dataGroup_13_9, dataGroup_12_9};
  wire [15:0]   res_hi_hi_hi_9 = {dataGroup_15_9, dataGroup_14_9};
  wire [31:0]   res_hi_hi_9 = {res_hi_hi_hi_9, res_hi_hi_lo_9};
  wire [63:0]   res_hi_9 = {res_hi_hi_9, res_hi_lo_9};
  wire [127:0]  res_27 = {res_hi_9, res_lo_9};
  wire [255:0]  lo_lo_3 = {res_25, res_24};
  wire [255:0]  lo_hi_3 = {res_27, res_26};
  wire [511:0]  lo_3 = {lo_hi_3, lo_lo_3};
  wire [1023:0] regroupLoadData_0_3 = {512'h0, lo_3};
  wire [511:0]  dataGroup_lo_160 = {dataGroup_lo_hi_160, dataGroup_lo_lo_160};
  wire [511:0]  dataGroup_hi_160 = {dataGroup_hi_hi_160, dataGroup_hi_lo_160};
  wire [7:0]    dataGroup_0_10 = dataGroup_lo_160[7:0];
  wire [511:0]  dataGroup_lo_161 = {dataGroup_lo_hi_161, dataGroup_lo_lo_161};
  wire [511:0]  dataGroup_hi_161 = {dataGroup_hi_hi_161, dataGroup_hi_lo_161};
  wire [7:0]    dataGroup_1_10 = dataGroup_lo_161[47:40];
  wire [511:0]  dataGroup_lo_162 = {dataGroup_lo_hi_162, dataGroup_lo_lo_162};
  wire [511:0]  dataGroup_hi_162 = {dataGroup_hi_hi_162, dataGroup_hi_lo_162};
  wire [7:0]    dataGroup_2_10 = dataGroup_lo_162[87:80];
  wire [511:0]  dataGroup_lo_163 = {dataGroup_lo_hi_163, dataGroup_lo_lo_163};
  wire [511:0]  dataGroup_hi_163 = {dataGroup_hi_hi_163, dataGroup_hi_lo_163};
  wire [7:0]    dataGroup_3_10 = dataGroup_lo_163[127:120];
  wire [511:0]  dataGroup_lo_164 = {dataGroup_lo_hi_164, dataGroup_lo_lo_164};
  wire [511:0]  dataGroup_hi_164 = {dataGroup_hi_hi_164, dataGroup_hi_lo_164};
  wire [7:0]    dataGroup_4_10 = dataGroup_lo_164[167:160];
  wire [511:0]  dataGroup_lo_165 = {dataGroup_lo_hi_165, dataGroup_lo_lo_165};
  wire [511:0]  dataGroup_hi_165 = {dataGroup_hi_hi_165, dataGroup_hi_lo_165};
  wire [7:0]    dataGroup_5_10 = dataGroup_lo_165[207:200];
  wire [511:0]  dataGroup_lo_166 = {dataGroup_lo_hi_166, dataGroup_lo_lo_166};
  wire [511:0]  dataGroup_hi_166 = {dataGroup_hi_hi_166, dataGroup_hi_lo_166};
  wire [7:0]    dataGroup_6_10 = dataGroup_lo_166[247:240];
  wire [511:0]  dataGroup_lo_167 = {dataGroup_lo_hi_167, dataGroup_lo_lo_167};
  wire [511:0]  dataGroup_hi_167 = {dataGroup_hi_hi_167, dataGroup_hi_lo_167};
  wire [7:0]    dataGroup_7_10 = dataGroup_lo_167[287:280];
  wire [511:0]  dataGroup_lo_168 = {dataGroup_lo_hi_168, dataGroup_lo_lo_168};
  wire [511:0]  dataGroup_hi_168 = {dataGroup_hi_hi_168, dataGroup_hi_lo_168};
  wire [7:0]    dataGroup_8_10 = dataGroup_lo_168[327:320];
  wire [511:0]  dataGroup_lo_169 = {dataGroup_lo_hi_169, dataGroup_lo_lo_169};
  wire [511:0]  dataGroup_hi_169 = {dataGroup_hi_hi_169, dataGroup_hi_lo_169};
  wire [7:0]    dataGroup_9_10 = dataGroup_lo_169[367:360];
  wire [511:0]  dataGroup_lo_170 = {dataGroup_lo_hi_170, dataGroup_lo_lo_170};
  wire [511:0]  dataGroup_hi_170 = {dataGroup_hi_hi_170, dataGroup_hi_lo_170};
  wire [7:0]    dataGroup_10_10 = dataGroup_lo_170[407:400];
  wire [511:0]  dataGroup_lo_171 = {dataGroup_lo_hi_171, dataGroup_lo_lo_171};
  wire [511:0]  dataGroup_hi_171 = {dataGroup_hi_hi_171, dataGroup_hi_lo_171};
  wire [7:0]    dataGroup_11_10 = dataGroup_lo_171[447:440];
  wire [511:0]  dataGroup_lo_172 = {dataGroup_lo_hi_172, dataGroup_lo_lo_172};
  wire [511:0]  dataGroup_hi_172 = {dataGroup_hi_hi_172, dataGroup_hi_lo_172};
  wire [7:0]    dataGroup_12_10 = dataGroup_lo_172[487:480];
  wire [511:0]  dataGroup_lo_173 = {dataGroup_lo_hi_173, dataGroup_lo_lo_173};
  wire [511:0]  dataGroup_hi_173 = {dataGroup_hi_hi_173, dataGroup_hi_lo_173};
  wire [7:0]    dataGroup_13_10 = dataGroup_hi_173[15:8];
  wire [511:0]  dataGroup_lo_174 = {dataGroup_lo_hi_174, dataGroup_lo_lo_174};
  wire [511:0]  dataGroup_hi_174 = {dataGroup_hi_hi_174, dataGroup_hi_lo_174};
  wire [7:0]    dataGroup_14_10 = dataGroup_hi_174[55:48];
  wire [511:0]  dataGroup_lo_175 = {dataGroup_lo_hi_175, dataGroup_lo_lo_175};
  wire [511:0]  dataGroup_hi_175 = {dataGroup_hi_hi_175, dataGroup_hi_lo_175};
  wire [7:0]    dataGroup_15_10 = dataGroup_hi_175[95:88];
  wire [15:0]   res_lo_lo_lo_10 = {dataGroup_1_10, dataGroup_0_10};
  wire [15:0]   res_lo_lo_hi_10 = {dataGroup_3_10, dataGroup_2_10};
  wire [31:0]   res_lo_lo_10 = {res_lo_lo_hi_10, res_lo_lo_lo_10};
  wire [15:0]   res_lo_hi_lo_10 = {dataGroup_5_10, dataGroup_4_10};
  wire [15:0]   res_lo_hi_hi_10 = {dataGroup_7_10, dataGroup_6_10};
  wire [31:0]   res_lo_hi_10 = {res_lo_hi_hi_10, res_lo_hi_lo_10};
  wire [63:0]   res_lo_10 = {res_lo_hi_10, res_lo_lo_10};
  wire [15:0]   res_hi_lo_lo_10 = {dataGroup_9_10, dataGroup_8_10};
  wire [15:0]   res_hi_lo_hi_10 = {dataGroup_11_10, dataGroup_10_10};
  wire [31:0]   res_hi_lo_10 = {res_hi_lo_hi_10, res_hi_lo_lo_10};
  wire [15:0]   res_hi_hi_lo_10 = {dataGroup_13_10, dataGroup_12_10};
  wire [15:0]   res_hi_hi_hi_10 = {dataGroup_15_10, dataGroup_14_10};
  wire [31:0]   res_hi_hi_10 = {res_hi_hi_hi_10, res_hi_hi_lo_10};
  wire [63:0]   res_hi_10 = {res_hi_hi_10, res_hi_lo_10};
  wire [127:0]  res_32 = {res_hi_10, res_lo_10};
  wire [511:0]  dataGroup_lo_176 = {dataGroup_lo_hi_176, dataGroup_lo_lo_176};
  wire [511:0]  dataGroup_hi_176 = {dataGroup_hi_hi_176, dataGroup_hi_lo_176};
  wire [7:0]    dataGroup_0_11 = dataGroup_lo_176[15:8];
  wire [511:0]  dataGroup_lo_177 = {dataGroup_lo_hi_177, dataGroup_lo_lo_177};
  wire [511:0]  dataGroup_hi_177 = {dataGroup_hi_hi_177, dataGroup_hi_lo_177};
  wire [7:0]    dataGroup_1_11 = dataGroup_lo_177[55:48];
  wire [511:0]  dataGroup_lo_178 = {dataGroup_lo_hi_178, dataGroup_lo_lo_178};
  wire [511:0]  dataGroup_hi_178 = {dataGroup_hi_hi_178, dataGroup_hi_lo_178};
  wire [7:0]    dataGroup_2_11 = dataGroup_lo_178[95:88];
  wire [511:0]  dataGroup_lo_179 = {dataGroup_lo_hi_179, dataGroup_lo_lo_179};
  wire [511:0]  dataGroup_hi_179 = {dataGroup_hi_hi_179, dataGroup_hi_lo_179};
  wire [7:0]    dataGroup_3_11 = dataGroup_lo_179[135:128];
  wire [511:0]  dataGroup_lo_180 = {dataGroup_lo_hi_180, dataGroup_lo_lo_180};
  wire [511:0]  dataGroup_hi_180 = {dataGroup_hi_hi_180, dataGroup_hi_lo_180};
  wire [7:0]    dataGroup_4_11 = dataGroup_lo_180[175:168];
  wire [511:0]  dataGroup_lo_181 = {dataGroup_lo_hi_181, dataGroup_lo_lo_181};
  wire [511:0]  dataGroup_hi_181 = {dataGroup_hi_hi_181, dataGroup_hi_lo_181};
  wire [7:0]    dataGroup_5_11 = dataGroup_lo_181[215:208];
  wire [511:0]  dataGroup_lo_182 = {dataGroup_lo_hi_182, dataGroup_lo_lo_182};
  wire [511:0]  dataGroup_hi_182 = {dataGroup_hi_hi_182, dataGroup_hi_lo_182};
  wire [7:0]    dataGroup_6_11 = dataGroup_lo_182[255:248];
  wire [511:0]  dataGroup_lo_183 = {dataGroup_lo_hi_183, dataGroup_lo_lo_183};
  wire [511:0]  dataGroup_hi_183 = {dataGroup_hi_hi_183, dataGroup_hi_lo_183};
  wire [7:0]    dataGroup_7_11 = dataGroup_lo_183[295:288];
  wire [511:0]  dataGroup_lo_184 = {dataGroup_lo_hi_184, dataGroup_lo_lo_184};
  wire [511:0]  dataGroup_hi_184 = {dataGroup_hi_hi_184, dataGroup_hi_lo_184};
  wire [7:0]    dataGroup_8_11 = dataGroup_lo_184[335:328];
  wire [511:0]  dataGroup_lo_185 = {dataGroup_lo_hi_185, dataGroup_lo_lo_185};
  wire [511:0]  dataGroup_hi_185 = {dataGroup_hi_hi_185, dataGroup_hi_lo_185};
  wire [7:0]    dataGroup_9_11 = dataGroup_lo_185[375:368];
  wire [511:0]  dataGroup_lo_186 = {dataGroup_lo_hi_186, dataGroup_lo_lo_186};
  wire [511:0]  dataGroup_hi_186 = {dataGroup_hi_hi_186, dataGroup_hi_lo_186};
  wire [7:0]    dataGroup_10_11 = dataGroup_lo_186[415:408];
  wire [511:0]  dataGroup_lo_187 = {dataGroup_lo_hi_187, dataGroup_lo_lo_187};
  wire [511:0]  dataGroup_hi_187 = {dataGroup_hi_hi_187, dataGroup_hi_lo_187};
  wire [7:0]    dataGroup_11_11 = dataGroup_lo_187[455:448];
  wire [511:0]  dataGroup_lo_188 = {dataGroup_lo_hi_188, dataGroup_lo_lo_188};
  wire [511:0]  dataGroup_hi_188 = {dataGroup_hi_hi_188, dataGroup_hi_lo_188};
  wire [7:0]    dataGroup_12_11 = dataGroup_lo_188[495:488];
  wire [511:0]  dataGroup_lo_189 = {dataGroup_lo_hi_189, dataGroup_lo_lo_189};
  wire [511:0]  dataGroup_hi_189 = {dataGroup_hi_hi_189, dataGroup_hi_lo_189};
  wire [7:0]    dataGroup_13_11 = dataGroup_hi_189[23:16];
  wire [511:0]  dataGroup_lo_190 = {dataGroup_lo_hi_190, dataGroup_lo_lo_190};
  wire [511:0]  dataGroup_hi_190 = {dataGroup_hi_hi_190, dataGroup_hi_lo_190};
  wire [7:0]    dataGroup_14_11 = dataGroup_hi_190[63:56];
  wire [511:0]  dataGroup_lo_191 = {dataGroup_lo_hi_191, dataGroup_lo_lo_191};
  wire [511:0]  dataGroup_hi_191 = {dataGroup_hi_hi_191, dataGroup_hi_lo_191};
  wire [7:0]    dataGroup_15_11 = dataGroup_hi_191[103:96];
  wire [15:0]   res_lo_lo_lo_11 = {dataGroup_1_11, dataGroup_0_11};
  wire [15:0]   res_lo_lo_hi_11 = {dataGroup_3_11, dataGroup_2_11};
  wire [31:0]   res_lo_lo_11 = {res_lo_lo_hi_11, res_lo_lo_lo_11};
  wire [15:0]   res_lo_hi_lo_11 = {dataGroup_5_11, dataGroup_4_11};
  wire [15:0]   res_lo_hi_hi_11 = {dataGroup_7_11, dataGroup_6_11};
  wire [31:0]   res_lo_hi_11 = {res_lo_hi_hi_11, res_lo_hi_lo_11};
  wire [63:0]   res_lo_11 = {res_lo_hi_11, res_lo_lo_11};
  wire [15:0]   res_hi_lo_lo_11 = {dataGroup_9_11, dataGroup_8_11};
  wire [15:0]   res_hi_lo_hi_11 = {dataGroup_11_11, dataGroup_10_11};
  wire [31:0]   res_hi_lo_11 = {res_hi_lo_hi_11, res_hi_lo_lo_11};
  wire [15:0]   res_hi_hi_lo_11 = {dataGroup_13_11, dataGroup_12_11};
  wire [15:0]   res_hi_hi_hi_11 = {dataGroup_15_11, dataGroup_14_11};
  wire [31:0]   res_hi_hi_11 = {res_hi_hi_hi_11, res_hi_hi_lo_11};
  wire [63:0]   res_hi_11 = {res_hi_hi_11, res_hi_lo_11};
  wire [127:0]  res_33 = {res_hi_11, res_lo_11};
  wire [511:0]  dataGroup_lo_192 = {dataGroup_lo_hi_192, dataGroup_lo_lo_192};
  wire [511:0]  dataGroup_hi_192 = {dataGroup_hi_hi_192, dataGroup_hi_lo_192};
  wire [7:0]    dataGroup_0_12 = dataGroup_lo_192[23:16];
  wire [511:0]  dataGroup_lo_193 = {dataGroup_lo_hi_193, dataGroup_lo_lo_193};
  wire [511:0]  dataGroup_hi_193 = {dataGroup_hi_hi_193, dataGroup_hi_lo_193};
  wire [7:0]    dataGroup_1_12 = dataGroup_lo_193[63:56];
  wire [511:0]  dataGroup_lo_194 = {dataGroup_lo_hi_194, dataGroup_lo_lo_194};
  wire [511:0]  dataGroup_hi_194 = {dataGroup_hi_hi_194, dataGroup_hi_lo_194};
  wire [7:0]    dataGroup_2_12 = dataGroup_lo_194[103:96];
  wire [511:0]  dataGroup_lo_195 = {dataGroup_lo_hi_195, dataGroup_lo_lo_195};
  wire [511:0]  dataGroup_hi_195 = {dataGroup_hi_hi_195, dataGroup_hi_lo_195};
  wire [7:0]    dataGroup_3_12 = dataGroup_lo_195[143:136];
  wire [511:0]  dataGroup_lo_196 = {dataGroup_lo_hi_196, dataGroup_lo_lo_196};
  wire [511:0]  dataGroup_hi_196 = {dataGroup_hi_hi_196, dataGroup_hi_lo_196};
  wire [7:0]    dataGroup_4_12 = dataGroup_lo_196[183:176];
  wire [511:0]  dataGroup_lo_197 = {dataGroup_lo_hi_197, dataGroup_lo_lo_197};
  wire [511:0]  dataGroup_hi_197 = {dataGroup_hi_hi_197, dataGroup_hi_lo_197};
  wire [7:0]    dataGroup_5_12 = dataGroup_lo_197[223:216];
  wire [511:0]  dataGroup_lo_198 = {dataGroup_lo_hi_198, dataGroup_lo_lo_198};
  wire [511:0]  dataGroup_hi_198 = {dataGroup_hi_hi_198, dataGroup_hi_lo_198};
  wire [7:0]    dataGroup_6_12 = dataGroup_lo_198[263:256];
  wire [511:0]  dataGroup_lo_199 = {dataGroup_lo_hi_199, dataGroup_lo_lo_199};
  wire [511:0]  dataGroup_hi_199 = {dataGroup_hi_hi_199, dataGroup_hi_lo_199};
  wire [7:0]    dataGroup_7_12 = dataGroup_lo_199[303:296];
  wire [511:0]  dataGroup_lo_200 = {dataGroup_lo_hi_200, dataGroup_lo_lo_200};
  wire [511:0]  dataGroup_hi_200 = {dataGroup_hi_hi_200, dataGroup_hi_lo_200};
  wire [7:0]    dataGroup_8_12 = dataGroup_lo_200[343:336];
  wire [511:0]  dataGroup_lo_201 = {dataGroup_lo_hi_201, dataGroup_lo_lo_201};
  wire [511:0]  dataGroup_hi_201 = {dataGroup_hi_hi_201, dataGroup_hi_lo_201};
  wire [7:0]    dataGroup_9_12 = dataGroup_lo_201[383:376];
  wire [511:0]  dataGroup_lo_202 = {dataGroup_lo_hi_202, dataGroup_lo_lo_202};
  wire [511:0]  dataGroup_hi_202 = {dataGroup_hi_hi_202, dataGroup_hi_lo_202};
  wire [7:0]    dataGroup_10_12 = dataGroup_lo_202[423:416];
  wire [511:0]  dataGroup_lo_203 = {dataGroup_lo_hi_203, dataGroup_lo_lo_203};
  wire [511:0]  dataGroup_hi_203 = {dataGroup_hi_hi_203, dataGroup_hi_lo_203};
  wire [7:0]    dataGroup_11_12 = dataGroup_lo_203[463:456];
  wire [511:0]  dataGroup_lo_204 = {dataGroup_lo_hi_204, dataGroup_lo_lo_204};
  wire [511:0]  dataGroup_hi_204 = {dataGroup_hi_hi_204, dataGroup_hi_lo_204};
  wire [7:0]    dataGroup_12_12 = dataGroup_lo_204[503:496];
  wire [511:0]  dataGroup_lo_205 = {dataGroup_lo_hi_205, dataGroup_lo_lo_205};
  wire [511:0]  dataGroup_hi_205 = {dataGroup_hi_hi_205, dataGroup_hi_lo_205};
  wire [7:0]    dataGroup_13_12 = dataGroup_hi_205[31:24];
  wire [511:0]  dataGroup_lo_206 = {dataGroup_lo_hi_206, dataGroup_lo_lo_206};
  wire [511:0]  dataGroup_hi_206 = {dataGroup_hi_hi_206, dataGroup_hi_lo_206};
  wire [7:0]    dataGroup_14_12 = dataGroup_hi_206[71:64];
  wire [511:0]  dataGroup_lo_207 = {dataGroup_lo_hi_207, dataGroup_lo_lo_207};
  wire [511:0]  dataGroup_hi_207 = {dataGroup_hi_hi_207, dataGroup_hi_lo_207};
  wire [7:0]    dataGroup_15_12 = dataGroup_hi_207[111:104];
  wire [15:0]   res_lo_lo_lo_12 = {dataGroup_1_12, dataGroup_0_12};
  wire [15:0]   res_lo_lo_hi_12 = {dataGroup_3_12, dataGroup_2_12};
  wire [31:0]   res_lo_lo_12 = {res_lo_lo_hi_12, res_lo_lo_lo_12};
  wire [15:0]   res_lo_hi_lo_12 = {dataGroup_5_12, dataGroup_4_12};
  wire [15:0]   res_lo_hi_hi_12 = {dataGroup_7_12, dataGroup_6_12};
  wire [31:0]   res_lo_hi_12 = {res_lo_hi_hi_12, res_lo_hi_lo_12};
  wire [63:0]   res_lo_12 = {res_lo_hi_12, res_lo_lo_12};
  wire [15:0]   res_hi_lo_lo_12 = {dataGroup_9_12, dataGroup_8_12};
  wire [15:0]   res_hi_lo_hi_12 = {dataGroup_11_12, dataGroup_10_12};
  wire [31:0]   res_hi_lo_12 = {res_hi_lo_hi_12, res_hi_lo_lo_12};
  wire [15:0]   res_hi_hi_lo_12 = {dataGroup_13_12, dataGroup_12_12};
  wire [15:0]   res_hi_hi_hi_12 = {dataGroup_15_12, dataGroup_14_12};
  wire [31:0]   res_hi_hi_12 = {res_hi_hi_hi_12, res_hi_hi_lo_12};
  wire [63:0]   res_hi_12 = {res_hi_hi_12, res_hi_lo_12};
  wire [127:0]  res_34 = {res_hi_12, res_lo_12};
  wire [511:0]  dataGroup_lo_208 = {dataGroup_lo_hi_208, dataGroup_lo_lo_208};
  wire [511:0]  dataGroup_hi_208 = {dataGroup_hi_hi_208, dataGroup_hi_lo_208};
  wire [7:0]    dataGroup_0_13 = dataGroup_lo_208[31:24];
  wire [511:0]  dataGroup_lo_209 = {dataGroup_lo_hi_209, dataGroup_lo_lo_209};
  wire [511:0]  dataGroup_hi_209 = {dataGroup_hi_hi_209, dataGroup_hi_lo_209};
  wire [7:0]    dataGroup_1_13 = dataGroup_lo_209[71:64];
  wire [511:0]  dataGroup_lo_210 = {dataGroup_lo_hi_210, dataGroup_lo_lo_210};
  wire [511:0]  dataGroup_hi_210 = {dataGroup_hi_hi_210, dataGroup_hi_lo_210};
  wire [7:0]    dataGroup_2_13 = dataGroup_lo_210[111:104];
  wire [511:0]  dataGroup_lo_211 = {dataGroup_lo_hi_211, dataGroup_lo_lo_211};
  wire [511:0]  dataGroup_hi_211 = {dataGroup_hi_hi_211, dataGroup_hi_lo_211};
  wire [7:0]    dataGroup_3_13 = dataGroup_lo_211[151:144];
  wire [511:0]  dataGroup_lo_212 = {dataGroup_lo_hi_212, dataGroup_lo_lo_212};
  wire [511:0]  dataGroup_hi_212 = {dataGroup_hi_hi_212, dataGroup_hi_lo_212};
  wire [7:0]    dataGroup_4_13 = dataGroup_lo_212[191:184];
  wire [511:0]  dataGroup_lo_213 = {dataGroup_lo_hi_213, dataGroup_lo_lo_213};
  wire [511:0]  dataGroup_hi_213 = {dataGroup_hi_hi_213, dataGroup_hi_lo_213};
  wire [7:0]    dataGroup_5_13 = dataGroup_lo_213[231:224];
  wire [511:0]  dataGroup_lo_214 = {dataGroup_lo_hi_214, dataGroup_lo_lo_214};
  wire [511:0]  dataGroup_hi_214 = {dataGroup_hi_hi_214, dataGroup_hi_lo_214};
  wire [7:0]    dataGroup_6_13 = dataGroup_lo_214[271:264];
  wire [511:0]  dataGroup_lo_215 = {dataGroup_lo_hi_215, dataGroup_lo_lo_215};
  wire [511:0]  dataGroup_hi_215 = {dataGroup_hi_hi_215, dataGroup_hi_lo_215};
  wire [7:0]    dataGroup_7_13 = dataGroup_lo_215[311:304];
  wire [511:0]  dataGroup_lo_216 = {dataGroup_lo_hi_216, dataGroup_lo_lo_216};
  wire [511:0]  dataGroup_hi_216 = {dataGroup_hi_hi_216, dataGroup_hi_lo_216};
  wire [7:0]    dataGroup_8_13 = dataGroup_lo_216[351:344];
  wire [511:0]  dataGroup_lo_217 = {dataGroup_lo_hi_217, dataGroup_lo_lo_217};
  wire [511:0]  dataGroup_hi_217 = {dataGroup_hi_hi_217, dataGroup_hi_lo_217};
  wire [7:0]    dataGroup_9_13 = dataGroup_lo_217[391:384];
  wire [511:0]  dataGroup_lo_218 = {dataGroup_lo_hi_218, dataGroup_lo_lo_218};
  wire [511:0]  dataGroup_hi_218 = {dataGroup_hi_hi_218, dataGroup_hi_lo_218};
  wire [7:0]    dataGroup_10_13 = dataGroup_lo_218[431:424];
  wire [511:0]  dataGroup_lo_219 = {dataGroup_lo_hi_219, dataGroup_lo_lo_219};
  wire [511:0]  dataGroup_hi_219 = {dataGroup_hi_hi_219, dataGroup_hi_lo_219};
  wire [7:0]    dataGroup_11_13 = dataGroup_lo_219[471:464];
  wire [511:0]  dataGroup_lo_220 = {dataGroup_lo_hi_220, dataGroup_lo_lo_220};
  wire [511:0]  dataGroup_hi_220 = {dataGroup_hi_hi_220, dataGroup_hi_lo_220};
  wire [7:0]    dataGroup_12_13 = dataGroup_lo_220[511:504];
  wire [511:0]  dataGroup_lo_221 = {dataGroup_lo_hi_221, dataGroup_lo_lo_221};
  wire [511:0]  dataGroup_hi_221 = {dataGroup_hi_hi_221, dataGroup_hi_lo_221};
  wire [7:0]    dataGroup_13_13 = dataGroup_hi_221[39:32];
  wire [511:0]  dataGroup_lo_222 = {dataGroup_lo_hi_222, dataGroup_lo_lo_222};
  wire [511:0]  dataGroup_hi_222 = {dataGroup_hi_hi_222, dataGroup_hi_lo_222};
  wire [7:0]    dataGroup_14_13 = dataGroup_hi_222[79:72];
  wire [511:0]  dataGroup_lo_223 = {dataGroup_lo_hi_223, dataGroup_lo_lo_223};
  wire [511:0]  dataGroup_hi_223 = {dataGroup_hi_hi_223, dataGroup_hi_lo_223};
  wire [7:0]    dataGroup_15_13 = dataGroup_hi_223[119:112];
  wire [15:0]   res_lo_lo_lo_13 = {dataGroup_1_13, dataGroup_0_13};
  wire [15:0]   res_lo_lo_hi_13 = {dataGroup_3_13, dataGroup_2_13};
  wire [31:0]   res_lo_lo_13 = {res_lo_lo_hi_13, res_lo_lo_lo_13};
  wire [15:0]   res_lo_hi_lo_13 = {dataGroup_5_13, dataGroup_4_13};
  wire [15:0]   res_lo_hi_hi_13 = {dataGroup_7_13, dataGroup_6_13};
  wire [31:0]   res_lo_hi_13 = {res_lo_hi_hi_13, res_lo_hi_lo_13};
  wire [63:0]   res_lo_13 = {res_lo_hi_13, res_lo_lo_13};
  wire [15:0]   res_hi_lo_lo_13 = {dataGroup_9_13, dataGroup_8_13};
  wire [15:0]   res_hi_lo_hi_13 = {dataGroup_11_13, dataGroup_10_13};
  wire [31:0]   res_hi_lo_13 = {res_hi_lo_hi_13, res_hi_lo_lo_13};
  wire [15:0]   res_hi_hi_lo_13 = {dataGroup_13_13, dataGroup_12_13};
  wire [15:0]   res_hi_hi_hi_13 = {dataGroup_15_13, dataGroup_14_13};
  wire [31:0]   res_hi_hi_13 = {res_hi_hi_hi_13, res_hi_hi_lo_13};
  wire [63:0]   res_hi_13 = {res_hi_hi_13, res_hi_lo_13};
  wire [127:0]  res_35 = {res_hi_13, res_lo_13};
  wire [511:0]  dataGroup_lo_224 = {dataGroup_lo_hi_224, dataGroup_lo_lo_224};
  wire [511:0]  dataGroup_hi_224 = {dataGroup_hi_hi_224, dataGroup_hi_lo_224};
  wire [7:0]    dataGroup_0_14 = dataGroup_lo_224[39:32];
  wire [511:0]  dataGroup_lo_225 = {dataGroup_lo_hi_225, dataGroup_lo_lo_225};
  wire [511:0]  dataGroup_hi_225 = {dataGroup_hi_hi_225, dataGroup_hi_lo_225};
  wire [7:0]    dataGroup_1_14 = dataGroup_lo_225[79:72];
  wire [511:0]  dataGroup_lo_226 = {dataGroup_lo_hi_226, dataGroup_lo_lo_226};
  wire [511:0]  dataGroup_hi_226 = {dataGroup_hi_hi_226, dataGroup_hi_lo_226};
  wire [7:0]    dataGroup_2_14 = dataGroup_lo_226[119:112];
  wire [511:0]  dataGroup_lo_227 = {dataGroup_lo_hi_227, dataGroup_lo_lo_227};
  wire [511:0]  dataGroup_hi_227 = {dataGroup_hi_hi_227, dataGroup_hi_lo_227};
  wire [7:0]    dataGroup_3_14 = dataGroup_lo_227[159:152];
  wire [511:0]  dataGroup_lo_228 = {dataGroup_lo_hi_228, dataGroup_lo_lo_228};
  wire [511:0]  dataGroup_hi_228 = {dataGroup_hi_hi_228, dataGroup_hi_lo_228};
  wire [7:0]    dataGroup_4_14 = dataGroup_lo_228[199:192];
  wire [511:0]  dataGroup_lo_229 = {dataGroup_lo_hi_229, dataGroup_lo_lo_229};
  wire [511:0]  dataGroup_hi_229 = {dataGroup_hi_hi_229, dataGroup_hi_lo_229};
  wire [7:0]    dataGroup_5_14 = dataGroup_lo_229[239:232];
  wire [511:0]  dataGroup_lo_230 = {dataGroup_lo_hi_230, dataGroup_lo_lo_230};
  wire [511:0]  dataGroup_hi_230 = {dataGroup_hi_hi_230, dataGroup_hi_lo_230};
  wire [7:0]    dataGroup_6_14 = dataGroup_lo_230[279:272];
  wire [511:0]  dataGroup_lo_231 = {dataGroup_lo_hi_231, dataGroup_lo_lo_231};
  wire [511:0]  dataGroup_hi_231 = {dataGroup_hi_hi_231, dataGroup_hi_lo_231};
  wire [7:0]    dataGroup_7_14 = dataGroup_lo_231[319:312];
  wire [511:0]  dataGroup_lo_232 = {dataGroup_lo_hi_232, dataGroup_lo_lo_232};
  wire [511:0]  dataGroup_hi_232 = {dataGroup_hi_hi_232, dataGroup_hi_lo_232};
  wire [7:0]    dataGroup_8_14 = dataGroup_lo_232[359:352];
  wire [511:0]  dataGroup_lo_233 = {dataGroup_lo_hi_233, dataGroup_lo_lo_233};
  wire [511:0]  dataGroup_hi_233 = {dataGroup_hi_hi_233, dataGroup_hi_lo_233};
  wire [7:0]    dataGroup_9_14 = dataGroup_lo_233[399:392];
  wire [511:0]  dataGroup_lo_234 = {dataGroup_lo_hi_234, dataGroup_lo_lo_234};
  wire [511:0]  dataGroup_hi_234 = {dataGroup_hi_hi_234, dataGroup_hi_lo_234};
  wire [7:0]    dataGroup_10_14 = dataGroup_lo_234[439:432];
  wire [511:0]  dataGroup_lo_235 = {dataGroup_lo_hi_235, dataGroup_lo_lo_235};
  wire [511:0]  dataGroup_hi_235 = {dataGroup_hi_hi_235, dataGroup_hi_lo_235};
  wire [7:0]    dataGroup_11_14 = dataGroup_lo_235[479:472];
  wire [511:0]  dataGroup_lo_236 = {dataGroup_lo_hi_236, dataGroup_lo_lo_236};
  wire [511:0]  dataGroup_hi_236 = {dataGroup_hi_hi_236, dataGroup_hi_lo_236};
  wire [7:0]    dataGroup_12_14 = dataGroup_hi_236[7:0];
  wire [511:0]  dataGroup_lo_237 = {dataGroup_lo_hi_237, dataGroup_lo_lo_237};
  wire [511:0]  dataGroup_hi_237 = {dataGroup_hi_hi_237, dataGroup_hi_lo_237};
  wire [7:0]    dataGroup_13_14 = dataGroup_hi_237[47:40];
  wire [511:0]  dataGroup_lo_238 = {dataGroup_lo_hi_238, dataGroup_lo_lo_238};
  wire [511:0]  dataGroup_hi_238 = {dataGroup_hi_hi_238, dataGroup_hi_lo_238};
  wire [7:0]    dataGroup_14_14 = dataGroup_hi_238[87:80];
  wire [511:0]  dataGroup_lo_239 = {dataGroup_lo_hi_239, dataGroup_lo_lo_239};
  wire [511:0]  dataGroup_hi_239 = {dataGroup_hi_hi_239, dataGroup_hi_lo_239};
  wire [7:0]    dataGroup_15_14 = dataGroup_hi_239[127:120];
  wire [15:0]   res_lo_lo_lo_14 = {dataGroup_1_14, dataGroup_0_14};
  wire [15:0]   res_lo_lo_hi_14 = {dataGroup_3_14, dataGroup_2_14};
  wire [31:0]   res_lo_lo_14 = {res_lo_lo_hi_14, res_lo_lo_lo_14};
  wire [15:0]   res_lo_hi_lo_14 = {dataGroup_5_14, dataGroup_4_14};
  wire [15:0]   res_lo_hi_hi_14 = {dataGroup_7_14, dataGroup_6_14};
  wire [31:0]   res_lo_hi_14 = {res_lo_hi_hi_14, res_lo_hi_lo_14};
  wire [63:0]   res_lo_14 = {res_lo_hi_14, res_lo_lo_14};
  wire [15:0]   res_hi_lo_lo_14 = {dataGroup_9_14, dataGroup_8_14};
  wire [15:0]   res_hi_lo_hi_14 = {dataGroup_11_14, dataGroup_10_14};
  wire [31:0]   res_hi_lo_14 = {res_hi_lo_hi_14, res_hi_lo_lo_14};
  wire [15:0]   res_hi_hi_lo_14 = {dataGroup_13_14, dataGroup_12_14};
  wire [15:0]   res_hi_hi_hi_14 = {dataGroup_15_14, dataGroup_14_14};
  wire [31:0]   res_hi_hi_14 = {res_hi_hi_hi_14, res_hi_hi_lo_14};
  wire [63:0]   res_hi_14 = {res_hi_hi_14, res_hi_lo_14};
  wire [127:0]  res_36 = {res_hi_14, res_lo_14};
  wire [255:0]  lo_lo_4 = {res_33, res_32};
  wire [255:0]  lo_hi_4 = {res_35, res_34};
  wire [511:0]  lo_4 = {lo_hi_4, lo_lo_4};
  wire [255:0]  hi_lo_4 = {128'h0, res_36};
  wire [511:0]  hi_4 = {256'h0, hi_lo_4};
  wire [1023:0] regroupLoadData_0_4 = {hi_4, lo_4};
  wire [511:0]  dataGroup_lo_240 = {dataGroup_lo_hi_240, dataGroup_lo_lo_240};
  wire [511:0]  dataGroup_hi_240 = {dataGroup_hi_hi_240, dataGroup_hi_lo_240};
  wire [7:0]    dataGroup_0_15 = dataGroup_lo_240[7:0];
  wire [511:0]  dataGroup_lo_241 = {dataGroup_lo_hi_241, dataGroup_lo_lo_241};
  wire [511:0]  dataGroup_hi_241 = {dataGroup_hi_hi_241, dataGroup_hi_lo_241};
  wire [7:0]    dataGroup_1_15 = dataGroup_lo_241[55:48];
  wire [511:0]  dataGroup_lo_242 = {dataGroup_lo_hi_242, dataGroup_lo_lo_242};
  wire [511:0]  dataGroup_hi_242 = {dataGroup_hi_hi_242, dataGroup_hi_lo_242};
  wire [7:0]    dataGroup_2_15 = dataGroup_lo_242[103:96];
  wire [511:0]  dataGroup_lo_243 = {dataGroup_lo_hi_243, dataGroup_lo_lo_243};
  wire [511:0]  dataGroup_hi_243 = {dataGroup_hi_hi_243, dataGroup_hi_lo_243};
  wire [7:0]    dataGroup_3_15 = dataGroup_lo_243[151:144];
  wire [511:0]  dataGroup_lo_244 = {dataGroup_lo_hi_244, dataGroup_lo_lo_244};
  wire [511:0]  dataGroup_hi_244 = {dataGroup_hi_hi_244, dataGroup_hi_lo_244};
  wire [7:0]    dataGroup_4_15 = dataGroup_lo_244[199:192];
  wire [511:0]  dataGroup_lo_245 = {dataGroup_lo_hi_245, dataGroup_lo_lo_245};
  wire [511:0]  dataGroup_hi_245 = {dataGroup_hi_hi_245, dataGroup_hi_lo_245};
  wire [7:0]    dataGroup_5_15 = dataGroup_lo_245[247:240];
  wire [511:0]  dataGroup_lo_246 = {dataGroup_lo_hi_246, dataGroup_lo_lo_246};
  wire [511:0]  dataGroup_hi_246 = {dataGroup_hi_hi_246, dataGroup_hi_lo_246};
  wire [7:0]    dataGroup_6_15 = dataGroup_lo_246[295:288];
  wire [511:0]  dataGroup_lo_247 = {dataGroup_lo_hi_247, dataGroup_lo_lo_247};
  wire [511:0]  dataGroup_hi_247 = {dataGroup_hi_hi_247, dataGroup_hi_lo_247};
  wire [7:0]    dataGroup_7_15 = dataGroup_lo_247[343:336];
  wire [511:0]  dataGroup_lo_248 = {dataGroup_lo_hi_248, dataGroup_lo_lo_248};
  wire [511:0]  dataGroup_hi_248 = {dataGroup_hi_hi_248, dataGroup_hi_lo_248};
  wire [7:0]    dataGroup_8_15 = dataGroup_lo_248[391:384];
  wire [511:0]  dataGroup_lo_249 = {dataGroup_lo_hi_249, dataGroup_lo_lo_249};
  wire [511:0]  dataGroup_hi_249 = {dataGroup_hi_hi_249, dataGroup_hi_lo_249};
  wire [7:0]    dataGroup_9_15 = dataGroup_lo_249[439:432];
  wire [511:0]  dataGroup_lo_250 = {dataGroup_lo_hi_250, dataGroup_lo_lo_250};
  wire [511:0]  dataGroup_hi_250 = {dataGroup_hi_hi_250, dataGroup_hi_lo_250};
  wire [7:0]    dataGroup_10_15 = dataGroup_lo_250[487:480];
  wire [511:0]  dataGroup_lo_251 = {dataGroup_lo_hi_251, dataGroup_lo_lo_251};
  wire [511:0]  dataGroup_hi_251 = {dataGroup_hi_hi_251, dataGroup_hi_lo_251};
  wire [7:0]    dataGroup_11_15 = dataGroup_hi_251[23:16];
  wire [511:0]  dataGroup_lo_252 = {dataGroup_lo_hi_252, dataGroup_lo_lo_252};
  wire [511:0]  dataGroup_hi_252 = {dataGroup_hi_hi_252, dataGroup_hi_lo_252};
  wire [7:0]    dataGroup_12_15 = dataGroup_hi_252[71:64];
  wire [511:0]  dataGroup_lo_253 = {dataGroup_lo_hi_253, dataGroup_lo_lo_253};
  wire [511:0]  dataGroup_hi_253 = {dataGroup_hi_hi_253, dataGroup_hi_lo_253};
  wire [7:0]    dataGroup_13_15 = dataGroup_hi_253[119:112];
  wire [511:0]  dataGroup_lo_254 = {dataGroup_lo_hi_254, dataGroup_lo_lo_254};
  wire [511:0]  dataGroup_hi_254 = {dataGroup_hi_hi_254, dataGroup_hi_lo_254};
  wire [7:0]    dataGroup_14_15 = dataGroup_hi_254[167:160];
  wire [511:0]  dataGroup_lo_255 = {dataGroup_lo_hi_255, dataGroup_lo_lo_255};
  wire [511:0]  dataGroup_hi_255 = {dataGroup_hi_hi_255, dataGroup_hi_lo_255};
  wire [7:0]    dataGroup_15_15 = dataGroup_hi_255[215:208];
  wire [15:0]   res_lo_lo_lo_15 = {dataGroup_1_15, dataGroup_0_15};
  wire [15:0]   res_lo_lo_hi_15 = {dataGroup_3_15, dataGroup_2_15};
  wire [31:0]   res_lo_lo_15 = {res_lo_lo_hi_15, res_lo_lo_lo_15};
  wire [15:0]   res_lo_hi_lo_15 = {dataGroup_5_15, dataGroup_4_15};
  wire [15:0]   res_lo_hi_hi_15 = {dataGroup_7_15, dataGroup_6_15};
  wire [31:0]   res_lo_hi_15 = {res_lo_hi_hi_15, res_lo_hi_lo_15};
  wire [63:0]   res_lo_15 = {res_lo_hi_15, res_lo_lo_15};
  wire [15:0]   res_hi_lo_lo_15 = {dataGroup_9_15, dataGroup_8_15};
  wire [15:0]   res_hi_lo_hi_15 = {dataGroup_11_15, dataGroup_10_15};
  wire [31:0]   res_hi_lo_15 = {res_hi_lo_hi_15, res_hi_lo_lo_15};
  wire [15:0]   res_hi_hi_lo_15 = {dataGroup_13_15, dataGroup_12_15};
  wire [15:0]   res_hi_hi_hi_15 = {dataGroup_15_15, dataGroup_14_15};
  wire [31:0]   res_hi_hi_15 = {res_hi_hi_hi_15, res_hi_hi_lo_15};
  wire [63:0]   res_hi_15 = {res_hi_hi_15, res_hi_lo_15};
  wire [127:0]  res_40 = {res_hi_15, res_lo_15};
  wire [511:0]  dataGroup_lo_256 = {dataGroup_lo_hi_256, dataGroup_lo_lo_256};
  wire [511:0]  dataGroup_hi_256 = {dataGroup_hi_hi_256, dataGroup_hi_lo_256};
  wire [7:0]    dataGroup_0_16 = dataGroup_lo_256[15:8];
  wire [511:0]  dataGroup_lo_257 = {dataGroup_lo_hi_257, dataGroup_lo_lo_257};
  wire [511:0]  dataGroup_hi_257 = {dataGroup_hi_hi_257, dataGroup_hi_lo_257};
  wire [7:0]    dataGroup_1_16 = dataGroup_lo_257[63:56];
  wire [511:0]  dataGroup_lo_258 = {dataGroup_lo_hi_258, dataGroup_lo_lo_258};
  wire [511:0]  dataGroup_hi_258 = {dataGroup_hi_hi_258, dataGroup_hi_lo_258};
  wire [7:0]    dataGroup_2_16 = dataGroup_lo_258[111:104];
  wire [511:0]  dataGroup_lo_259 = {dataGroup_lo_hi_259, dataGroup_lo_lo_259};
  wire [511:0]  dataGroup_hi_259 = {dataGroup_hi_hi_259, dataGroup_hi_lo_259};
  wire [7:0]    dataGroup_3_16 = dataGroup_lo_259[159:152];
  wire [511:0]  dataGroup_lo_260 = {dataGroup_lo_hi_260, dataGroup_lo_lo_260};
  wire [511:0]  dataGroup_hi_260 = {dataGroup_hi_hi_260, dataGroup_hi_lo_260};
  wire [7:0]    dataGroup_4_16 = dataGroup_lo_260[207:200];
  wire [511:0]  dataGroup_lo_261 = {dataGroup_lo_hi_261, dataGroup_lo_lo_261};
  wire [511:0]  dataGroup_hi_261 = {dataGroup_hi_hi_261, dataGroup_hi_lo_261};
  wire [7:0]    dataGroup_5_16 = dataGroup_lo_261[255:248];
  wire [511:0]  dataGroup_lo_262 = {dataGroup_lo_hi_262, dataGroup_lo_lo_262};
  wire [511:0]  dataGroup_hi_262 = {dataGroup_hi_hi_262, dataGroup_hi_lo_262};
  wire [7:0]    dataGroup_6_16 = dataGroup_lo_262[303:296];
  wire [511:0]  dataGroup_lo_263 = {dataGroup_lo_hi_263, dataGroup_lo_lo_263};
  wire [511:0]  dataGroup_hi_263 = {dataGroup_hi_hi_263, dataGroup_hi_lo_263};
  wire [7:0]    dataGroup_7_16 = dataGroup_lo_263[351:344];
  wire [511:0]  dataGroup_lo_264 = {dataGroup_lo_hi_264, dataGroup_lo_lo_264};
  wire [511:0]  dataGroup_hi_264 = {dataGroup_hi_hi_264, dataGroup_hi_lo_264};
  wire [7:0]    dataGroup_8_16 = dataGroup_lo_264[399:392];
  wire [511:0]  dataGroup_lo_265 = {dataGroup_lo_hi_265, dataGroup_lo_lo_265};
  wire [511:0]  dataGroup_hi_265 = {dataGroup_hi_hi_265, dataGroup_hi_lo_265};
  wire [7:0]    dataGroup_9_16 = dataGroup_lo_265[447:440];
  wire [511:0]  dataGroup_lo_266 = {dataGroup_lo_hi_266, dataGroup_lo_lo_266};
  wire [511:0]  dataGroup_hi_266 = {dataGroup_hi_hi_266, dataGroup_hi_lo_266};
  wire [7:0]    dataGroup_10_16 = dataGroup_lo_266[495:488];
  wire [511:0]  dataGroup_lo_267 = {dataGroup_lo_hi_267, dataGroup_lo_lo_267};
  wire [511:0]  dataGroup_hi_267 = {dataGroup_hi_hi_267, dataGroup_hi_lo_267};
  wire [7:0]    dataGroup_11_16 = dataGroup_hi_267[31:24];
  wire [511:0]  dataGroup_lo_268 = {dataGroup_lo_hi_268, dataGroup_lo_lo_268};
  wire [511:0]  dataGroup_hi_268 = {dataGroup_hi_hi_268, dataGroup_hi_lo_268};
  wire [7:0]    dataGroup_12_16 = dataGroup_hi_268[79:72];
  wire [511:0]  dataGroup_lo_269 = {dataGroup_lo_hi_269, dataGroup_lo_lo_269};
  wire [511:0]  dataGroup_hi_269 = {dataGroup_hi_hi_269, dataGroup_hi_lo_269};
  wire [7:0]    dataGroup_13_16 = dataGroup_hi_269[127:120];
  wire [511:0]  dataGroup_lo_270 = {dataGroup_lo_hi_270, dataGroup_lo_lo_270};
  wire [511:0]  dataGroup_hi_270 = {dataGroup_hi_hi_270, dataGroup_hi_lo_270};
  wire [7:0]    dataGroup_14_16 = dataGroup_hi_270[175:168];
  wire [511:0]  dataGroup_lo_271 = {dataGroup_lo_hi_271, dataGroup_lo_lo_271};
  wire [511:0]  dataGroup_hi_271 = {dataGroup_hi_hi_271, dataGroup_hi_lo_271};
  wire [7:0]    dataGroup_15_16 = dataGroup_hi_271[223:216];
  wire [15:0]   res_lo_lo_lo_16 = {dataGroup_1_16, dataGroup_0_16};
  wire [15:0]   res_lo_lo_hi_16 = {dataGroup_3_16, dataGroup_2_16};
  wire [31:0]   res_lo_lo_16 = {res_lo_lo_hi_16, res_lo_lo_lo_16};
  wire [15:0]   res_lo_hi_lo_16 = {dataGroup_5_16, dataGroup_4_16};
  wire [15:0]   res_lo_hi_hi_16 = {dataGroup_7_16, dataGroup_6_16};
  wire [31:0]   res_lo_hi_16 = {res_lo_hi_hi_16, res_lo_hi_lo_16};
  wire [63:0]   res_lo_16 = {res_lo_hi_16, res_lo_lo_16};
  wire [15:0]   res_hi_lo_lo_16 = {dataGroup_9_16, dataGroup_8_16};
  wire [15:0]   res_hi_lo_hi_16 = {dataGroup_11_16, dataGroup_10_16};
  wire [31:0]   res_hi_lo_16 = {res_hi_lo_hi_16, res_hi_lo_lo_16};
  wire [15:0]   res_hi_hi_lo_16 = {dataGroup_13_16, dataGroup_12_16};
  wire [15:0]   res_hi_hi_hi_16 = {dataGroup_15_16, dataGroup_14_16};
  wire [31:0]   res_hi_hi_16 = {res_hi_hi_hi_16, res_hi_hi_lo_16};
  wire [63:0]   res_hi_16 = {res_hi_hi_16, res_hi_lo_16};
  wire [127:0]  res_41 = {res_hi_16, res_lo_16};
  wire [511:0]  dataGroup_lo_272 = {dataGroup_lo_hi_272, dataGroup_lo_lo_272};
  wire [511:0]  dataGroup_hi_272 = {dataGroup_hi_hi_272, dataGroup_hi_lo_272};
  wire [7:0]    dataGroup_0_17 = dataGroup_lo_272[23:16];
  wire [511:0]  dataGroup_lo_273 = {dataGroup_lo_hi_273, dataGroup_lo_lo_273};
  wire [511:0]  dataGroup_hi_273 = {dataGroup_hi_hi_273, dataGroup_hi_lo_273};
  wire [7:0]    dataGroup_1_17 = dataGroup_lo_273[71:64];
  wire [511:0]  dataGroup_lo_274 = {dataGroup_lo_hi_274, dataGroup_lo_lo_274};
  wire [511:0]  dataGroup_hi_274 = {dataGroup_hi_hi_274, dataGroup_hi_lo_274};
  wire [7:0]    dataGroup_2_17 = dataGroup_lo_274[119:112];
  wire [511:0]  dataGroup_lo_275 = {dataGroup_lo_hi_275, dataGroup_lo_lo_275};
  wire [511:0]  dataGroup_hi_275 = {dataGroup_hi_hi_275, dataGroup_hi_lo_275};
  wire [7:0]    dataGroup_3_17 = dataGroup_lo_275[167:160];
  wire [511:0]  dataGroup_lo_276 = {dataGroup_lo_hi_276, dataGroup_lo_lo_276};
  wire [511:0]  dataGroup_hi_276 = {dataGroup_hi_hi_276, dataGroup_hi_lo_276};
  wire [7:0]    dataGroup_4_17 = dataGroup_lo_276[215:208];
  wire [511:0]  dataGroup_lo_277 = {dataGroup_lo_hi_277, dataGroup_lo_lo_277};
  wire [511:0]  dataGroup_hi_277 = {dataGroup_hi_hi_277, dataGroup_hi_lo_277};
  wire [7:0]    dataGroup_5_17 = dataGroup_lo_277[263:256];
  wire [511:0]  dataGroup_lo_278 = {dataGroup_lo_hi_278, dataGroup_lo_lo_278};
  wire [511:0]  dataGroup_hi_278 = {dataGroup_hi_hi_278, dataGroup_hi_lo_278};
  wire [7:0]    dataGroup_6_17 = dataGroup_lo_278[311:304];
  wire [511:0]  dataGroup_lo_279 = {dataGroup_lo_hi_279, dataGroup_lo_lo_279};
  wire [511:0]  dataGroup_hi_279 = {dataGroup_hi_hi_279, dataGroup_hi_lo_279};
  wire [7:0]    dataGroup_7_17 = dataGroup_lo_279[359:352];
  wire [511:0]  dataGroup_lo_280 = {dataGroup_lo_hi_280, dataGroup_lo_lo_280};
  wire [511:0]  dataGroup_hi_280 = {dataGroup_hi_hi_280, dataGroup_hi_lo_280};
  wire [7:0]    dataGroup_8_17 = dataGroup_lo_280[407:400];
  wire [511:0]  dataGroup_lo_281 = {dataGroup_lo_hi_281, dataGroup_lo_lo_281};
  wire [511:0]  dataGroup_hi_281 = {dataGroup_hi_hi_281, dataGroup_hi_lo_281};
  wire [7:0]    dataGroup_9_17 = dataGroup_lo_281[455:448];
  wire [511:0]  dataGroup_lo_282 = {dataGroup_lo_hi_282, dataGroup_lo_lo_282};
  wire [511:0]  dataGroup_hi_282 = {dataGroup_hi_hi_282, dataGroup_hi_lo_282};
  wire [7:0]    dataGroup_10_17 = dataGroup_lo_282[503:496];
  wire [511:0]  dataGroup_lo_283 = {dataGroup_lo_hi_283, dataGroup_lo_lo_283};
  wire [511:0]  dataGroup_hi_283 = {dataGroup_hi_hi_283, dataGroup_hi_lo_283};
  wire [7:0]    dataGroup_11_17 = dataGroup_hi_283[39:32];
  wire [511:0]  dataGroup_lo_284 = {dataGroup_lo_hi_284, dataGroup_lo_lo_284};
  wire [511:0]  dataGroup_hi_284 = {dataGroup_hi_hi_284, dataGroup_hi_lo_284};
  wire [7:0]    dataGroup_12_17 = dataGroup_hi_284[87:80];
  wire [511:0]  dataGroup_lo_285 = {dataGroup_lo_hi_285, dataGroup_lo_lo_285};
  wire [511:0]  dataGroup_hi_285 = {dataGroup_hi_hi_285, dataGroup_hi_lo_285};
  wire [7:0]    dataGroup_13_17 = dataGroup_hi_285[135:128];
  wire [511:0]  dataGroup_lo_286 = {dataGroup_lo_hi_286, dataGroup_lo_lo_286};
  wire [511:0]  dataGroup_hi_286 = {dataGroup_hi_hi_286, dataGroup_hi_lo_286};
  wire [7:0]    dataGroup_14_17 = dataGroup_hi_286[183:176];
  wire [511:0]  dataGroup_lo_287 = {dataGroup_lo_hi_287, dataGroup_lo_lo_287};
  wire [511:0]  dataGroup_hi_287 = {dataGroup_hi_hi_287, dataGroup_hi_lo_287};
  wire [7:0]    dataGroup_15_17 = dataGroup_hi_287[231:224];
  wire [15:0]   res_lo_lo_lo_17 = {dataGroup_1_17, dataGroup_0_17};
  wire [15:0]   res_lo_lo_hi_17 = {dataGroup_3_17, dataGroup_2_17};
  wire [31:0]   res_lo_lo_17 = {res_lo_lo_hi_17, res_lo_lo_lo_17};
  wire [15:0]   res_lo_hi_lo_17 = {dataGroup_5_17, dataGroup_4_17};
  wire [15:0]   res_lo_hi_hi_17 = {dataGroup_7_17, dataGroup_6_17};
  wire [31:0]   res_lo_hi_17 = {res_lo_hi_hi_17, res_lo_hi_lo_17};
  wire [63:0]   res_lo_17 = {res_lo_hi_17, res_lo_lo_17};
  wire [15:0]   res_hi_lo_lo_17 = {dataGroup_9_17, dataGroup_8_17};
  wire [15:0]   res_hi_lo_hi_17 = {dataGroup_11_17, dataGroup_10_17};
  wire [31:0]   res_hi_lo_17 = {res_hi_lo_hi_17, res_hi_lo_lo_17};
  wire [15:0]   res_hi_hi_lo_17 = {dataGroup_13_17, dataGroup_12_17};
  wire [15:0]   res_hi_hi_hi_17 = {dataGroup_15_17, dataGroup_14_17};
  wire [31:0]   res_hi_hi_17 = {res_hi_hi_hi_17, res_hi_hi_lo_17};
  wire [63:0]   res_hi_17 = {res_hi_hi_17, res_hi_lo_17};
  wire [127:0]  res_42 = {res_hi_17, res_lo_17};
  wire [511:0]  dataGroup_lo_288 = {dataGroup_lo_hi_288, dataGroup_lo_lo_288};
  wire [511:0]  dataGroup_hi_288 = {dataGroup_hi_hi_288, dataGroup_hi_lo_288};
  wire [7:0]    dataGroup_0_18 = dataGroup_lo_288[31:24];
  wire [511:0]  dataGroup_lo_289 = {dataGroup_lo_hi_289, dataGroup_lo_lo_289};
  wire [511:0]  dataGroup_hi_289 = {dataGroup_hi_hi_289, dataGroup_hi_lo_289};
  wire [7:0]    dataGroup_1_18 = dataGroup_lo_289[79:72];
  wire [511:0]  dataGroup_lo_290 = {dataGroup_lo_hi_290, dataGroup_lo_lo_290};
  wire [511:0]  dataGroup_hi_290 = {dataGroup_hi_hi_290, dataGroup_hi_lo_290};
  wire [7:0]    dataGroup_2_18 = dataGroup_lo_290[127:120];
  wire [511:0]  dataGroup_lo_291 = {dataGroup_lo_hi_291, dataGroup_lo_lo_291};
  wire [511:0]  dataGroup_hi_291 = {dataGroup_hi_hi_291, dataGroup_hi_lo_291};
  wire [7:0]    dataGroup_3_18 = dataGroup_lo_291[175:168];
  wire [511:0]  dataGroup_lo_292 = {dataGroup_lo_hi_292, dataGroup_lo_lo_292};
  wire [511:0]  dataGroup_hi_292 = {dataGroup_hi_hi_292, dataGroup_hi_lo_292};
  wire [7:0]    dataGroup_4_18 = dataGroup_lo_292[223:216];
  wire [511:0]  dataGroup_lo_293 = {dataGroup_lo_hi_293, dataGroup_lo_lo_293};
  wire [511:0]  dataGroup_hi_293 = {dataGroup_hi_hi_293, dataGroup_hi_lo_293};
  wire [7:0]    dataGroup_5_18 = dataGroup_lo_293[271:264];
  wire [511:0]  dataGroup_lo_294 = {dataGroup_lo_hi_294, dataGroup_lo_lo_294};
  wire [511:0]  dataGroup_hi_294 = {dataGroup_hi_hi_294, dataGroup_hi_lo_294};
  wire [7:0]    dataGroup_6_18 = dataGroup_lo_294[319:312];
  wire [511:0]  dataGroup_lo_295 = {dataGroup_lo_hi_295, dataGroup_lo_lo_295};
  wire [511:0]  dataGroup_hi_295 = {dataGroup_hi_hi_295, dataGroup_hi_lo_295};
  wire [7:0]    dataGroup_7_18 = dataGroup_lo_295[367:360];
  wire [511:0]  dataGroup_lo_296 = {dataGroup_lo_hi_296, dataGroup_lo_lo_296};
  wire [511:0]  dataGroup_hi_296 = {dataGroup_hi_hi_296, dataGroup_hi_lo_296};
  wire [7:0]    dataGroup_8_18 = dataGroup_lo_296[415:408];
  wire [511:0]  dataGroup_lo_297 = {dataGroup_lo_hi_297, dataGroup_lo_lo_297};
  wire [511:0]  dataGroup_hi_297 = {dataGroup_hi_hi_297, dataGroup_hi_lo_297};
  wire [7:0]    dataGroup_9_18 = dataGroup_lo_297[463:456];
  wire [511:0]  dataGroup_lo_298 = {dataGroup_lo_hi_298, dataGroup_lo_lo_298};
  wire [511:0]  dataGroup_hi_298 = {dataGroup_hi_hi_298, dataGroup_hi_lo_298};
  wire [7:0]    dataGroup_10_18 = dataGroup_lo_298[511:504];
  wire [511:0]  dataGroup_lo_299 = {dataGroup_lo_hi_299, dataGroup_lo_lo_299};
  wire [511:0]  dataGroup_hi_299 = {dataGroup_hi_hi_299, dataGroup_hi_lo_299};
  wire [7:0]    dataGroup_11_18 = dataGroup_hi_299[47:40];
  wire [511:0]  dataGroup_lo_300 = {dataGroup_lo_hi_300, dataGroup_lo_lo_300};
  wire [511:0]  dataGroup_hi_300 = {dataGroup_hi_hi_300, dataGroup_hi_lo_300};
  wire [7:0]    dataGroup_12_18 = dataGroup_hi_300[95:88];
  wire [511:0]  dataGroup_lo_301 = {dataGroup_lo_hi_301, dataGroup_lo_lo_301};
  wire [511:0]  dataGroup_hi_301 = {dataGroup_hi_hi_301, dataGroup_hi_lo_301};
  wire [7:0]    dataGroup_13_18 = dataGroup_hi_301[143:136];
  wire [511:0]  dataGroup_lo_302 = {dataGroup_lo_hi_302, dataGroup_lo_lo_302};
  wire [511:0]  dataGroup_hi_302 = {dataGroup_hi_hi_302, dataGroup_hi_lo_302};
  wire [7:0]    dataGroup_14_18 = dataGroup_hi_302[191:184];
  wire [511:0]  dataGroup_lo_303 = {dataGroup_lo_hi_303, dataGroup_lo_lo_303};
  wire [511:0]  dataGroup_hi_303 = {dataGroup_hi_hi_303, dataGroup_hi_lo_303};
  wire [7:0]    dataGroup_15_18 = dataGroup_hi_303[239:232];
  wire [15:0]   res_lo_lo_lo_18 = {dataGroup_1_18, dataGroup_0_18};
  wire [15:0]   res_lo_lo_hi_18 = {dataGroup_3_18, dataGroup_2_18};
  wire [31:0]   res_lo_lo_18 = {res_lo_lo_hi_18, res_lo_lo_lo_18};
  wire [15:0]   res_lo_hi_lo_18 = {dataGroup_5_18, dataGroup_4_18};
  wire [15:0]   res_lo_hi_hi_18 = {dataGroup_7_18, dataGroup_6_18};
  wire [31:0]   res_lo_hi_18 = {res_lo_hi_hi_18, res_lo_hi_lo_18};
  wire [63:0]   res_lo_18 = {res_lo_hi_18, res_lo_lo_18};
  wire [15:0]   res_hi_lo_lo_18 = {dataGroup_9_18, dataGroup_8_18};
  wire [15:0]   res_hi_lo_hi_18 = {dataGroup_11_18, dataGroup_10_18};
  wire [31:0]   res_hi_lo_18 = {res_hi_lo_hi_18, res_hi_lo_lo_18};
  wire [15:0]   res_hi_hi_lo_18 = {dataGroup_13_18, dataGroup_12_18};
  wire [15:0]   res_hi_hi_hi_18 = {dataGroup_15_18, dataGroup_14_18};
  wire [31:0]   res_hi_hi_18 = {res_hi_hi_hi_18, res_hi_hi_lo_18};
  wire [63:0]   res_hi_18 = {res_hi_hi_18, res_hi_lo_18};
  wire [127:0]  res_43 = {res_hi_18, res_lo_18};
  wire [511:0]  dataGroup_lo_304 = {dataGroup_lo_hi_304, dataGroup_lo_lo_304};
  wire [511:0]  dataGroup_hi_304 = {dataGroup_hi_hi_304, dataGroup_hi_lo_304};
  wire [7:0]    dataGroup_0_19 = dataGroup_lo_304[39:32];
  wire [511:0]  dataGroup_lo_305 = {dataGroup_lo_hi_305, dataGroup_lo_lo_305};
  wire [511:0]  dataGroup_hi_305 = {dataGroup_hi_hi_305, dataGroup_hi_lo_305};
  wire [7:0]    dataGroup_1_19 = dataGroup_lo_305[87:80];
  wire [511:0]  dataGroup_lo_306 = {dataGroup_lo_hi_306, dataGroup_lo_lo_306};
  wire [511:0]  dataGroup_hi_306 = {dataGroup_hi_hi_306, dataGroup_hi_lo_306};
  wire [7:0]    dataGroup_2_19 = dataGroup_lo_306[135:128];
  wire [511:0]  dataGroup_lo_307 = {dataGroup_lo_hi_307, dataGroup_lo_lo_307};
  wire [511:0]  dataGroup_hi_307 = {dataGroup_hi_hi_307, dataGroup_hi_lo_307};
  wire [7:0]    dataGroup_3_19 = dataGroup_lo_307[183:176];
  wire [511:0]  dataGroup_lo_308 = {dataGroup_lo_hi_308, dataGroup_lo_lo_308};
  wire [511:0]  dataGroup_hi_308 = {dataGroup_hi_hi_308, dataGroup_hi_lo_308};
  wire [7:0]    dataGroup_4_19 = dataGroup_lo_308[231:224];
  wire [511:0]  dataGroup_lo_309 = {dataGroup_lo_hi_309, dataGroup_lo_lo_309};
  wire [511:0]  dataGroup_hi_309 = {dataGroup_hi_hi_309, dataGroup_hi_lo_309};
  wire [7:0]    dataGroup_5_19 = dataGroup_lo_309[279:272];
  wire [511:0]  dataGroup_lo_310 = {dataGroup_lo_hi_310, dataGroup_lo_lo_310};
  wire [511:0]  dataGroup_hi_310 = {dataGroup_hi_hi_310, dataGroup_hi_lo_310};
  wire [7:0]    dataGroup_6_19 = dataGroup_lo_310[327:320];
  wire [511:0]  dataGroup_lo_311 = {dataGroup_lo_hi_311, dataGroup_lo_lo_311};
  wire [511:0]  dataGroup_hi_311 = {dataGroup_hi_hi_311, dataGroup_hi_lo_311};
  wire [7:0]    dataGroup_7_19 = dataGroup_lo_311[375:368];
  wire [511:0]  dataGroup_lo_312 = {dataGroup_lo_hi_312, dataGroup_lo_lo_312};
  wire [511:0]  dataGroup_hi_312 = {dataGroup_hi_hi_312, dataGroup_hi_lo_312};
  wire [7:0]    dataGroup_8_19 = dataGroup_lo_312[423:416];
  wire [511:0]  dataGroup_lo_313 = {dataGroup_lo_hi_313, dataGroup_lo_lo_313};
  wire [511:0]  dataGroup_hi_313 = {dataGroup_hi_hi_313, dataGroup_hi_lo_313};
  wire [7:0]    dataGroup_9_19 = dataGroup_lo_313[471:464];
  wire [511:0]  dataGroup_lo_314 = {dataGroup_lo_hi_314, dataGroup_lo_lo_314};
  wire [511:0]  dataGroup_hi_314 = {dataGroup_hi_hi_314, dataGroup_hi_lo_314};
  wire [7:0]    dataGroup_10_19 = dataGroup_hi_314[7:0];
  wire [511:0]  dataGroup_lo_315 = {dataGroup_lo_hi_315, dataGroup_lo_lo_315};
  wire [511:0]  dataGroup_hi_315 = {dataGroup_hi_hi_315, dataGroup_hi_lo_315};
  wire [7:0]    dataGroup_11_19 = dataGroup_hi_315[55:48];
  wire [511:0]  dataGroup_lo_316 = {dataGroup_lo_hi_316, dataGroup_lo_lo_316};
  wire [511:0]  dataGroup_hi_316 = {dataGroup_hi_hi_316, dataGroup_hi_lo_316};
  wire [7:0]    dataGroup_12_19 = dataGroup_hi_316[103:96];
  wire [511:0]  dataGroup_lo_317 = {dataGroup_lo_hi_317, dataGroup_lo_lo_317};
  wire [511:0]  dataGroup_hi_317 = {dataGroup_hi_hi_317, dataGroup_hi_lo_317};
  wire [7:0]    dataGroup_13_19 = dataGroup_hi_317[151:144];
  wire [511:0]  dataGroup_lo_318 = {dataGroup_lo_hi_318, dataGroup_lo_lo_318};
  wire [511:0]  dataGroup_hi_318 = {dataGroup_hi_hi_318, dataGroup_hi_lo_318};
  wire [7:0]    dataGroup_14_19 = dataGroup_hi_318[199:192];
  wire [511:0]  dataGroup_lo_319 = {dataGroup_lo_hi_319, dataGroup_lo_lo_319};
  wire [511:0]  dataGroup_hi_319 = {dataGroup_hi_hi_319, dataGroup_hi_lo_319};
  wire [7:0]    dataGroup_15_19 = dataGroup_hi_319[247:240];
  wire [15:0]   res_lo_lo_lo_19 = {dataGroup_1_19, dataGroup_0_19};
  wire [15:0]   res_lo_lo_hi_19 = {dataGroup_3_19, dataGroup_2_19};
  wire [31:0]   res_lo_lo_19 = {res_lo_lo_hi_19, res_lo_lo_lo_19};
  wire [15:0]   res_lo_hi_lo_19 = {dataGroup_5_19, dataGroup_4_19};
  wire [15:0]   res_lo_hi_hi_19 = {dataGroup_7_19, dataGroup_6_19};
  wire [31:0]   res_lo_hi_19 = {res_lo_hi_hi_19, res_lo_hi_lo_19};
  wire [63:0]   res_lo_19 = {res_lo_hi_19, res_lo_lo_19};
  wire [15:0]   res_hi_lo_lo_19 = {dataGroup_9_19, dataGroup_8_19};
  wire [15:0]   res_hi_lo_hi_19 = {dataGroup_11_19, dataGroup_10_19};
  wire [31:0]   res_hi_lo_19 = {res_hi_lo_hi_19, res_hi_lo_lo_19};
  wire [15:0]   res_hi_hi_lo_19 = {dataGroup_13_19, dataGroup_12_19};
  wire [15:0]   res_hi_hi_hi_19 = {dataGroup_15_19, dataGroup_14_19};
  wire [31:0]   res_hi_hi_19 = {res_hi_hi_hi_19, res_hi_hi_lo_19};
  wire [63:0]   res_hi_19 = {res_hi_hi_19, res_hi_lo_19};
  wire [127:0]  res_44 = {res_hi_19, res_lo_19};
  wire [511:0]  dataGroup_lo_320 = {dataGroup_lo_hi_320, dataGroup_lo_lo_320};
  wire [511:0]  dataGroup_hi_320 = {dataGroup_hi_hi_320, dataGroup_hi_lo_320};
  wire [7:0]    dataGroup_0_20 = dataGroup_lo_320[47:40];
  wire [511:0]  dataGroup_lo_321 = {dataGroup_lo_hi_321, dataGroup_lo_lo_321};
  wire [511:0]  dataGroup_hi_321 = {dataGroup_hi_hi_321, dataGroup_hi_lo_321};
  wire [7:0]    dataGroup_1_20 = dataGroup_lo_321[95:88];
  wire [511:0]  dataGroup_lo_322 = {dataGroup_lo_hi_322, dataGroup_lo_lo_322};
  wire [511:0]  dataGroup_hi_322 = {dataGroup_hi_hi_322, dataGroup_hi_lo_322};
  wire [7:0]    dataGroup_2_20 = dataGroup_lo_322[143:136];
  wire [511:0]  dataGroup_lo_323 = {dataGroup_lo_hi_323, dataGroup_lo_lo_323};
  wire [511:0]  dataGroup_hi_323 = {dataGroup_hi_hi_323, dataGroup_hi_lo_323};
  wire [7:0]    dataGroup_3_20 = dataGroup_lo_323[191:184];
  wire [511:0]  dataGroup_lo_324 = {dataGroup_lo_hi_324, dataGroup_lo_lo_324};
  wire [511:0]  dataGroup_hi_324 = {dataGroup_hi_hi_324, dataGroup_hi_lo_324};
  wire [7:0]    dataGroup_4_20 = dataGroup_lo_324[239:232];
  wire [511:0]  dataGroup_lo_325 = {dataGroup_lo_hi_325, dataGroup_lo_lo_325};
  wire [511:0]  dataGroup_hi_325 = {dataGroup_hi_hi_325, dataGroup_hi_lo_325};
  wire [7:0]    dataGroup_5_20 = dataGroup_lo_325[287:280];
  wire [511:0]  dataGroup_lo_326 = {dataGroup_lo_hi_326, dataGroup_lo_lo_326};
  wire [511:0]  dataGroup_hi_326 = {dataGroup_hi_hi_326, dataGroup_hi_lo_326};
  wire [7:0]    dataGroup_6_20 = dataGroup_lo_326[335:328];
  wire [511:0]  dataGroup_lo_327 = {dataGroup_lo_hi_327, dataGroup_lo_lo_327};
  wire [511:0]  dataGroup_hi_327 = {dataGroup_hi_hi_327, dataGroup_hi_lo_327};
  wire [7:0]    dataGroup_7_20 = dataGroup_lo_327[383:376];
  wire [511:0]  dataGroup_lo_328 = {dataGroup_lo_hi_328, dataGroup_lo_lo_328};
  wire [511:0]  dataGroup_hi_328 = {dataGroup_hi_hi_328, dataGroup_hi_lo_328};
  wire [7:0]    dataGroup_8_20 = dataGroup_lo_328[431:424];
  wire [511:0]  dataGroup_lo_329 = {dataGroup_lo_hi_329, dataGroup_lo_lo_329};
  wire [511:0]  dataGroup_hi_329 = {dataGroup_hi_hi_329, dataGroup_hi_lo_329};
  wire [7:0]    dataGroup_9_20 = dataGroup_lo_329[479:472];
  wire [511:0]  dataGroup_lo_330 = {dataGroup_lo_hi_330, dataGroup_lo_lo_330};
  wire [511:0]  dataGroup_hi_330 = {dataGroup_hi_hi_330, dataGroup_hi_lo_330};
  wire [7:0]    dataGroup_10_20 = dataGroup_hi_330[15:8];
  wire [511:0]  dataGroup_lo_331 = {dataGroup_lo_hi_331, dataGroup_lo_lo_331};
  wire [511:0]  dataGroup_hi_331 = {dataGroup_hi_hi_331, dataGroup_hi_lo_331};
  wire [7:0]    dataGroup_11_20 = dataGroup_hi_331[63:56];
  wire [511:0]  dataGroup_lo_332 = {dataGroup_lo_hi_332, dataGroup_lo_lo_332};
  wire [511:0]  dataGroup_hi_332 = {dataGroup_hi_hi_332, dataGroup_hi_lo_332};
  wire [7:0]    dataGroup_12_20 = dataGroup_hi_332[111:104];
  wire [511:0]  dataGroup_lo_333 = {dataGroup_lo_hi_333, dataGroup_lo_lo_333};
  wire [511:0]  dataGroup_hi_333 = {dataGroup_hi_hi_333, dataGroup_hi_lo_333};
  wire [7:0]    dataGroup_13_20 = dataGroup_hi_333[159:152];
  wire [511:0]  dataGroup_lo_334 = {dataGroup_lo_hi_334, dataGroup_lo_lo_334};
  wire [511:0]  dataGroup_hi_334 = {dataGroup_hi_hi_334, dataGroup_hi_lo_334};
  wire [7:0]    dataGroup_14_20 = dataGroup_hi_334[207:200];
  wire [511:0]  dataGroup_lo_335 = {dataGroup_lo_hi_335, dataGroup_lo_lo_335};
  wire [511:0]  dataGroup_hi_335 = {dataGroup_hi_hi_335, dataGroup_hi_lo_335};
  wire [7:0]    dataGroup_15_20 = dataGroup_hi_335[255:248];
  wire [15:0]   res_lo_lo_lo_20 = {dataGroup_1_20, dataGroup_0_20};
  wire [15:0]   res_lo_lo_hi_20 = {dataGroup_3_20, dataGroup_2_20};
  wire [31:0]   res_lo_lo_20 = {res_lo_lo_hi_20, res_lo_lo_lo_20};
  wire [15:0]   res_lo_hi_lo_20 = {dataGroup_5_20, dataGroup_4_20};
  wire [15:0]   res_lo_hi_hi_20 = {dataGroup_7_20, dataGroup_6_20};
  wire [31:0]   res_lo_hi_20 = {res_lo_hi_hi_20, res_lo_hi_lo_20};
  wire [63:0]   res_lo_20 = {res_lo_hi_20, res_lo_lo_20};
  wire [15:0]   res_hi_lo_lo_20 = {dataGroup_9_20, dataGroup_8_20};
  wire [15:0]   res_hi_lo_hi_20 = {dataGroup_11_20, dataGroup_10_20};
  wire [31:0]   res_hi_lo_20 = {res_hi_lo_hi_20, res_hi_lo_lo_20};
  wire [15:0]   res_hi_hi_lo_20 = {dataGroup_13_20, dataGroup_12_20};
  wire [15:0]   res_hi_hi_hi_20 = {dataGroup_15_20, dataGroup_14_20};
  wire [31:0]   res_hi_hi_20 = {res_hi_hi_hi_20, res_hi_hi_lo_20};
  wire [63:0]   res_hi_20 = {res_hi_hi_20, res_hi_lo_20};
  wire [127:0]  res_45 = {res_hi_20, res_lo_20};
  wire [255:0]  lo_lo_5 = {res_41, res_40};
  wire [255:0]  lo_hi_5 = {res_43, res_42};
  wire [511:0]  lo_5 = {lo_hi_5, lo_lo_5};
  wire [255:0]  hi_lo_5 = {res_45, res_44};
  wire [511:0]  hi_5 = {256'h0, hi_lo_5};
  wire [1023:0] regroupLoadData_0_5 = {hi_5, lo_5};
  wire [511:0]  dataGroup_lo_336 = {dataGroup_lo_hi_336, dataGroup_lo_lo_336};
  wire [511:0]  dataGroup_hi_336 = {dataGroup_hi_hi_336, dataGroup_hi_lo_336};
  wire [7:0]    dataGroup_0_21 = dataGroup_lo_336[7:0];
  wire [511:0]  dataGroup_lo_337 = {dataGroup_lo_hi_337, dataGroup_lo_lo_337};
  wire [511:0]  dataGroup_hi_337 = {dataGroup_hi_hi_337, dataGroup_hi_lo_337};
  wire [7:0]    dataGroup_1_21 = dataGroup_lo_337[63:56];
  wire [511:0]  dataGroup_lo_338 = {dataGroup_lo_hi_338, dataGroup_lo_lo_338};
  wire [511:0]  dataGroup_hi_338 = {dataGroup_hi_hi_338, dataGroup_hi_lo_338};
  wire [7:0]    dataGroup_2_21 = dataGroup_lo_338[119:112];
  wire [511:0]  dataGroup_lo_339 = {dataGroup_lo_hi_339, dataGroup_lo_lo_339};
  wire [511:0]  dataGroup_hi_339 = {dataGroup_hi_hi_339, dataGroup_hi_lo_339};
  wire [7:0]    dataGroup_3_21 = dataGroup_lo_339[175:168];
  wire [511:0]  dataGroup_lo_340 = {dataGroup_lo_hi_340, dataGroup_lo_lo_340};
  wire [511:0]  dataGroup_hi_340 = {dataGroup_hi_hi_340, dataGroup_hi_lo_340};
  wire [7:0]    dataGroup_4_21 = dataGroup_lo_340[231:224];
  wire [511:0]  dataGroup_lo_341 = {dataGroup_lo_hi_341, dataGroup_lo_lo_341};
  wire [511:0]  dataGroup_hi_341 = {dataGroup_hi_hi_341, dataGroup_hi_lo_341};
  wire [7:0]    dataGroup_5_21 = dataGroup_lo_341[287:280];
  wire [511:0]  dataGroup_lo_342 = {dataGroup_lo_hi_342, dataGroup_lo_lo_342};
  wire [511:0]  dataGroup_hi_342 = {dataGroup_hi_hi_342, dataGroup_hi_lo_342};
  wire [7:0]    dataGroup_6_21 = dataGroup_lo_342[343:336];
  wire [511:0]  dataGroup_lo_343 = {dataGroup_lo_hi_343, dataGroup_lo_lo_343};
  wire [511:0]  dataGroup_hi_343 = {dataGroup_hi_hi_343, dataGroup_hi_lo_343};
  wire [7:0]    dataGroup_7_21 = dataGroup_lo_343[399:392];
  wire [511:0]  dataGroup_lo_344 = {dataGroup_lo_hi_344, dataGroup_lo_lo_344};
  wire [511:0]  dataGroup_hi_344 = {dataGroup_hi_hi_344, dataGroup_hi_lo_344};
  wire [7:0]    dataGroup_8_21 = dataGroup_lo_344[455:448];
  wire [511:0]  dataGroup_lo_345 = {dataGroup_lo_hi_345, dataGroup_lo_lo_345};
  wire [511:0]  dataGroup_hi_345 = {dataGroup_hi_hi_345, dataGroup_hi_lo_345};
  wire [7:0]    dataGroup_9_21 = dataGroup_lo_345[511:504];
  wire [511:0]  dataGroup_lo_346 = {dataGroup_lo_hi_346, dataGroup_lo_lo_346};
  wire [511:0]  dataGroup_hi_346 = {dataGroup_hi_hi_346, dataGroup_hi_lo_346};
  wire [7:0]    dataGroup_10_21 = dataGroup_hi_346[55:48];
  wire [511:0]  dataGroup_lo_347 = {dataGroup_lo_hi_347, dataGroup_lo_lo_347};
  wire [511:0]  dataGroup_hi_347 = {dataGroup_hi_hi_347, dataGroup_hi_lo_347};
  wire [7:0]    dataGroup_11_21 = dataGroup_hi_347[111:104];
  wire [511:0]  dataGroup_lo_348 = {dataGroup_lo_hi_348, dataGroup_lo_lo_348};
  wire [511:0]  dataGroup_hi_348 = {dataGroup_hi_hi_348, dataGroup_hi_lo_348};
  wire [7:0]    dataGroup_12_21 = dataGroup_hi_348[167:160];
  wire [511:0]  dataGroup_lo_349 = {dataGroup_lo_hi_349, dataGroup_lo_lo_349};
  wire [511:0]  dataGroup_hi_349 = {dataGroup_hi_hi_349, dataGroup_hi_lo_349};
  wire [7:0]    dataGroup_13_21 = dataGroup_hi_349[223:216];
  wire [511:0]  dataGroup_lo_350 = {dataGroup_lo_hi_350, dataGroup_lo_lo_350};
  wire [511:0]  dataGroup_hi_350 = {dataGroup_hi_hi_350, dataGroup_hi_lo_350};
  wire [7:0]    dataGroup_14_21 = dataGroup_hi_350[279:272];
  wire [511:0]  dataGroup_lo_351 = {dataGroup_lo_hi_351, dataGroup_lo_lo_351};
  wire [511:0]  dataGroup_hi_351 = {dataGroup_hi_hi_351, dataGroup_hi_lo_351};
  wire [7:0]    dataGroup_15_21 = dataGroup_hi_351[335:328];
  wire [15:0]   res_lo_lo_lo_21 = {dataGroup_1_21, dataGroup_0_21};
  wire [15:0]   res_lo_lo_hi_21 = {dataGroup_3_21, dataGroup_2_21};
  wire [31:0]   res_lo_lo_21 = {res_lo_lo_hi_21, res_lo_lo_lo_21};
  wire [15:0]   res_lo_hi_lo_21 = {dataGroup_5_21, dataGroup_4_21};
  wire [15:0]   res_lo_hi_hi_21 = {dataGroup_7_21, dataGroup_6_21};
  wire [31:0]   res_lo_hi_21 = {res_lo_hi_hi_21, res_lo_hi_lo_21};
  wire [63:0]   res_lo_21 = {res_lo_hi_21, res_lo_lo_21};
  wire [15:0]   res_hi_lo_lo_21 = {dataGroup_9_21, dataGroup_8_21};
  wire [15:0]   res_hi_lo_hi_21 = {dataGroup_11_21, dataGroup_10_21};
  wire [31:0]   res_hi_lo_21 = {res_hi_lo_hi_21, res_hi_lo_lo_21};
  wire [15:0]   res_hi_hi_lo_21 = {dataGroup_13_21, dataGroup_12_21};
  wire [15:0]   res_hi_hi_hi_21 = {dataGroup_15_21, dataGroup_14_21};
  wire [31:0]   res_hi_hi_21 = {res_hi_hi_hi_21, res_hi_hi_lo_21};
  wire [63:0]   res_hi_21 = {res_hi_hi_21, res_hi_lo_21};
  wire [127:0]  res_48 = {res_hi_21, res_lo_21};
  wire [511:0]  dataGroup_lo_352 = {dataGroup_lo_hi_352, dataGroup_lo_lo_352};
  wire [511:0]  dataGroup_hi_352 = {dataGroup_hi_hi_352, dataGroup_hi_lo_352};
  wire [7:0]    dataGroup_0_22 = dataGroup_lo_352[15:8];
  wire [511:0]  dataGroup_lo_353 = {dataGroup_lo_hi_353, dataGroup_lo_lo_353};
  wire [511:0]  dataGroup_hi_353 = {dataGroup_hi_hi_353, dataGroup_hi_lo_353};
  wire [7:0]    dataGroup_1_22 = dataGroup_lo_353[71:64];
  wire [511:0]  dataGroup_lo_354 = {dataGroup_lo_hi_354, dataGroup_lo_lo_354};
  wire [511:0]  dataGroup_hi_354 = {dataGroup_hi_hi_354, dataGroup_hi_lo_354};
  wire [7:0]    dataGroup_2_22 = dataGroup_lo_354[127:120];
  wire [511:0]  dataGroup_lo_355 = {dataGroup_lo_hi_355, dataGroup_lo_lo_355};
  wire [511:0]  dataGroup_hi_355 = {dataGroup_hi_hi_355, dataGroup_hi_lo_355};
  wire [7:0]    dataGroup_3_22 = dataGroup_lo_355[183:176];
  wire [511:0]  dataGroup_lo_356 = {dataGroup_lo_hi_356, dataGroup_lo_lo_356};
  wire [511:0]  dataGroup_hi_356 = {dataGroup_hi_hi_356, dataGroup_hi_lo_356};
  wire [7:0]    dataGroup_4_22 = dataGroup_lo_356[239:232];
  wire [511:0]  dataGroup_lo_357 = {dataGroup_lo_hi_357, dataGroup_lo_lo_357};
  wire [511:0]  dataGroup_hi_357 = {dataGroup_hi_hi_357, dataGroup_hi_lo_357};
  wire [7:0]    dataGroup_5_22 = dataGroup_lo_357[295:288];
  wire [511:0]  dataGroup_lo_358 = {dataGroup_lo_hi_358, dataGroup_lo_lo_358};
  wire [511:0]  dataGroup_hi_358 = {dataGroup_hi_hi_358, dataGroup_hi_lo_358};
  wire [7:0]    dataGroup_6_22 = dataGroup_lo_358[351:344];
  wire [511:0]  dataGroup_lo_359 = {dataGroup_lo_hi_359, dataGroup_lo_lo_359};
  wire [511:0]  dataGroup_hi_359 = {dataGroup_hi_hi_359, dataGroup_hi_lo_359};
  wire [7:0]    dataGroup_7_22 = dataGroup_lo_359[407:400];
  wire [511:0]  dataGroup_lo_360 = {dataGroup_lo_hi_360, dataGroup_lo_lo_360};
  wire [511:0]  dataGroup_hi_360 = {dataGroup_hi_hi_360, dataGroup_hi_lo_360};
  wire [7:0]    dataGroup_8_22 = dataGroup_lo_360[463:456];
  wire [511:0]  dataGroup_lo_361 = {dataGroup_lo_hi_361, dataGroup_lo_lo_361};
  wire [511:0]  dataGroup_hi_361 = {dataGroup_hi_hi_361, dataGroup_hi_lo_361};
  wire [7:0]    dataGroup_9_22 = dataGroup_hi_361[7:0];
  wire [511:0]  dataGroup_lo_362 = {dataGroup_lo_hi_362, dataGroup_lo_lo_362};
  wire [511:0]  dataGroup_hi_362 = {dataGroup_hi_hi_362, dataGroup_hi_lo_362};
  wire [7:0]    dataGroup_10_22 = dataGroup_hi_362[63:56];
  wire [511:0]  dataGroup_lo_363 = {dataGroup_lo_hi_363, dataGroup_lo_lo_363};
  wire [511:0]  dataGroup_hi_363 = {dataGroup_hi_hi_363, dataGroup_hi_lo_363};
  wire [7:0]    dataGroup_11_22 = dataGroup_hi_363[119:112];
  wire [511:0]  dataGroup_lo_364 = {dataGroup_lo_hi_364, dataGroup_lo_lo_364};
  wire [511:0]  dataGroup_hi_364 = {dataGroup_hi_hi_364, dataGroup_hi_lo_364};
  wire [7:0]    dataGroup_12_22 = dataGroup_hi_364[175:168];
  wire [511:0]  dataGroup_lo_365 = {dataGroup_lo_hi_365, dataGroup_lo_lo_365};
  wire [511:0]  dataGroup_hi_365 = {dataGroup_hi_hi_365, dataGroup_hi_lo_365};
  wire [7:0]    dataGroup_13_22 = dataGroup_hi_365[231:224];
  wire [511:0]  dataGroup_lo_366 = {dataGroup_lo_hi_366, dataGroup_lo_lo_366};
  wire [511:0]  dataGroup_hi_366 = {dataGroup_hi_hi_366, dataGroup_hi_lo_366};
  wire [7:0]    dataGroup_14_22 = dataGroup_hi_366[287:280];
  wire [511:0]  dataGroup_lo_367 = {dataGroup_lo_hi_367, dataGroup_lo_lo_367};
  wire [511:0]  dataGroup_hi_367 = {dataGroup_hi_hi_367, dataGroup_hi_lo_367};
  wire [7:0]    dataGroup_15_22 = dataGroup_hi_367[343:336];
  wire [15:0]   res_lo_lo_lo_22 = {dataGroup_1_22, dataGroup_0_22};
  wire [15:0]   res_lo_lo_hi_22 = {dataGroup_3_22, dataGroup_2_22};
  wire [31:0]   res_lo_lo_22 = {res_lo_lo_hi_22, res_lo_lo_lo_22};
  wire [15:0]   res_lo_hi_lo_22 = {dataGroup_5_22, dataGroup_4_22};
  wire [15:0]   res_lo_hi_hi_22 = {dataGroup_7_22, dataGroup_6_22};
  wire [31:0]   res_lo_hi_22 = {res_lo_hi_hi_22, res_lo_hi_lo_22};
  wire [63:0]   res_lo_22 = {res_lo_hi_22, res_lo_lo_22};
  wire [15:0]   res_hi_lo_lo_22 = {dataGroup_9_22, dataGroup_8_22};
  wire [15:0]   res_hi_lo_hi_22 = {dataGroup_11_22, dataGroup_10_22};
  wire [31:0]   res_hi_lo_22 = {res_hi_lo_hi_22, res_hi_lo_lo_22};
  wire [15:0]   res_hi_hi_lo_22 = {dataGroup_13_22, dataGroup_12_22};
  wire [15:0]   res_hi_hi_hi_22 = {dataGroup_15_22, dataGroup_14_22};
  wire [31:0]   res_hi_hi_22 = {res_hi_hi_hi_22, res_hi_hi_lo_22};
  wire [63:0]   res_hi_22 = {res_hi_hi_22, res_hi_lo_22};
  wire [127:0]  res_49 = {res_hi_22, res_lo_22};
  wire [511:0]  dataGroup_lo_368 = {dataGroup_lo_hi_368, dataGroup_lo_lo_368};
  wire [511:0]  dataGroup_hi_368 = {dataGroup_hi_hi_368, dataGroup_hi_lo_368};
  wire [7:0]    dataGroup_0_23 = dataGroup_lo_368[23:16];
  wire [511:0]  dataGroup_lo_369 = {dataGroup_lo_hi_369, dataGroup_lo_lo_369};
  wire [511:0]  dataGroup_hi_369 = {dataGroup_hi_hi_369, dataGroup_hi_lo_369};
  wire [7:0]    dataGroup_1_23 = dataGroup_lo_369[79:72];
  wire [511:0]  dataGroup_lo_370 = {dataGroup_lo_hi_370, dataGroup_lo_lo_370};
  wire [511:0]  dataGroup_hi_370 = {dataGroup_hi_hi_370, dataGroup_hi_lo_370};
  wire [7:0]    dataGroup_2_23 = dataGroup_lo_370[135:128];
  wire [511:0]  dataGroup_lo_371 = {dataGroup_lo_hi_371, dataGroup_lo_lo_371};
  wire [511:0]  dataGroup_hi_371 = {dataGroup_hi_hi_371, dataGroup_hi_lo_371};
  wire [7:0]    dataGroup_3_23 = dataGroup_lo_371[191:184];
  wire [511:0]  dataGroup_lo_372 = {dataGroup_lo_hi_372, dataGroup_lo_lo_372};
  wire [511:0]  dataGroup_hi_372 = {dataGroup_hi_hi_372, dataGroup_hi_lo_372};
  wire [7:0]    dataGroup_4_23 = dataGroup_lo_372[247:240];
  wire [511:0]  dataGroup_lo_373 = {dataGroup_lo_hi_373, dataGroup_lo_lo_373};
  wire [511:0]  dataGroup_hi_373 = {dataGroup_hi_hi_373, dataGroup_hi_lo_373};
  wire [7:0]    dataGroup_5_23 = dataGroup_lo_373[303:296];
  wire [511:0]  dataGroup_lo_374 = {dataGroup_lo_hi_374, dataGroup_lo_lo_374};
  wire [511:0]  dataGroup_hi_374 = {dataGroup_hi_hi_374, dataGroup_hi_lo_374};
  wire [7:0]    dataGroup_6_23 = dataGroup_lo_374[359:352];
  wire [511:0]  dataGroup_lo_375 = {dataGroup_lo_hi_375, dataGroup_lo_lo_375};
  wire [511:0]  dataGroup_hi_375 = {dataGroup_hi_hi_375, dataGroup_hi_lo_375};
  wire [7:0]    dataGroup_7_23 = dataGroup_lo_375[415:408];
  wire [511:0]  dataGroup_lo_376 = {dataGroup_lo_hi_376, dataGroup_lo_lo_376};
  wire [511:0]  dataGroup_hi_376 = {dataGroup_hi_hi_376, dataGroup_hi_lo_376};
  wire [7:0]    dataGroup_8_23 = dataGroup_lo_376[471:464];
  wire [511:0]  dataGroup_lo_377 = {dataGroup_lo_hi_377, dataGroup_lo_lo_377};
  wire [511:0]  dataGroup_hi_377 = {dataGroup_hi_hi_377, dataGroup_hi_lo_377};
  wire [7:0]    dataGroup_9_23 = dataGroup_hi_377[15:8];
  wire [511:0]  dataGroup_lo_378 = {dataGroup_lo_hi_378, dataGroup_lo_lo_378};
  wire [511:0]  dataGroup_hi_378 = {dataGroup_hi_hi_378, dataGroup_hi_lo_378};
  wire [7:0]    dataGroup_10_23 = dataGroup_hi_378[71:64];
  wire [511:0]  dataGroup_lo_379 = {dataGroup_lo_hi_379, dataGroup_lo_lo_379};
  wire [511:0]  dataGroup_hi_379 = {dataGroup_hi_hi_379, dataGroup_hi_lo_379};
  wire [7:0]    dataGroup_11_23 = dataGroup_hi_379[127:120];
  wire [511:0]  dataGroup_lo_380 = {dataGroup_lo_hi_380, dataGroup_lo_lo_380};
  wire [511:0]  dataGroup_hi_380 = {dataGroup_hi_hi_380, dataGroup_hi_lo_380};
  wire [7:0]    dataGroup_12_23 = dataGroup_hi_380[183:176];
  wire [511:0]  dataGroup_lo_381 = {dataGroup_lo_hi_381, dataGroup_lo_lo_381};
  wire [511:0]  dataGroup_hi_381 = {dataGroup_hi_hi_381, dataGroup_hi_lo_381};
  wire [7:0]    dataGroup_13_23 = dataGroup_hi_381[239:232];
  wire [511:0]  dataGroup_lo_382 = {dataGroup_lo_hi_382, dataGroup_lo_lo_382};
  wire [511:0]  dataGroup_hi_382 = {dataGroup_hi_hi_382, dataGroup_hi_lo_382};
  wire [7:0]    dataGroup_14_23 = dataGroup_hi_382[295:288];
  wire [511:0]  dataGroup_lo_383 = {dataGroup_lo_hi_383, dataGroup_lo_lo_383};
  wire [511:0]  dataGroup_hi_383 = {dataGroup_hi_hi_383, dataGroup_hi_lo_383};
  wire [7:0]    dataGroup_15_23 = dataGroup_hi_383[351:344];
  wire [15:0]   res_lo_lo_lo_23 = {dataGroup_1_23, dataGroup_0_23};
  wire [15:0]   res_lo_lo_hi_23 = {dataGroup_3_23, dataGroup_2_23};
  wire [31:0]   res_lo_lo_23 = {res_lo_lo_hi_23, res_lo_lo_lo_23};
  wire [15:0]   res_lo_hi_lo_23 = {dataGroup_5_23, dataGroup_4_23};
  wire [15:0]   res_lo_hi_hi_23 = {dataGroup_7_23, dataGroup_6_23};
  wire [31:0]   res_lo_hi_23 = {res_lo_hi_hi_23, res_lo_hi_lo_23};
  wire [63:0]   res_lo_23 = {res_lo_hi_23, res_lo_lo_23};
  wire [15:0]   res_hi_lo_lo_23 = {dataGroup_9_23, dataGroup_8_23};
  wire [15:0]   res_hi_lo_hi_23 = {dataGroup_11_23, dataGroup_10_23};
  wire [31:0]   res_hi_lo_23 = {res_hi_lo_hi_23, res_hi_lo_lo_23};
  wire [15:0]   res_hi_hi_lo_23 = {dataGroup_13_23, dataGroup_12_23};
  wire [15:0]   res_hi_hi_hi_23 = {dataGroup_15_23, dataGroup_14_23};
  wire [31:0]   res_hi_hi_23 = {res_hi_hi_hi_23, res_hi_hi_lo_23};
  wire [63:0]   res_hi_23 = {res_hi_hi_23, res_hi_lo_23};
  wire [127:0]  res_50 = {res_hi_23, res_lo_23};
  wire [511:0]  dataGroup_lo_384 = {dataGroup_lo_hi_384, dataGroup_lo_lo_384};
  wire [511:0]  dataGroup_hi_384 = {dataGroup_hi_hi_384, dataGroup_hi_lo_384};
  wire [7:0]    dataGroup_0_24 = dataGroup_lo_384[31:24];
  wire [511:0]  dataGroup_lo_385 = {dataGroup_lo_hi_385, dataGroup_lo_lo_385};
  wire [511:0]  dataGroup_hi_385 = {dataGroup_hi_hi_385, dataGroup_hi_lo_385};
  wire [7:0]    dataGroup_1_24 = dataGroup_lo_385[87:80];
  wire [511:0]  dataGroup_lo_386 = {dataGroup_lo_hi_386, dataGroup_lo_lo_386};
  wire [511:0]  dataGroup_hi_386 = {dataGroup_hi_hi_386, dataGroup_hi_lo_386};
  wire [7:0]    dataGroup_2_24 = dataGroup_lo_386[143:136];
  wire [511:0]  dataGroup_lo_387 = {dataGroup_lo_hi_387, dataGroup_lo_lo_387};
  wire [511:0]  dataGroup_hi_387 = {dataGroup_hi_hi_387, dataGroup_hi_lo_387};
  wire [7:0]    dataGroup_3_24 = dataGroup_lo_387[199:192];
  wire [511:0]  dataGroup_lo_388 = {dataGroup_lo_hi_388, dataGroup_lo_lo_388};
  wire [511:0]  dataGroup_hi_388 = {dataGroup_hi_hi_388, dataGroup_hi_lo_388};
  wire [7:0]    dataGroup_4_24 = dataGroup_lo_388[255:248];
  wire [511:0]  dataGroup_lo_389 = {dataGroup_lo_hi_389, dataGroup_lo_lo_389};
  wire [511:0]  dataGroup_hi_389 = {dataGroup_hi_hi_389, dataGroup_hi_lo_389};
  wire [7:0]    dataGroup_5_24 = dataGroup_lo_389[311:304];
  wire [511:0]  dataGroup_lo_390 = {dataGroup_lo_hi_390, dataGroup_lo_lo_390};
  wire [511:0]  dataGroup_hi_390 = {dataGroup_hi_hi_390, dataGroup_hi_lo_390};
  wire [7:0]    dataGroup_6_24 = dataGroup_lo_390[367:360];
  wire [511:0]  dataGroup_lo_391 = {dataGroup_lo_hi_391, dataGroup_lo_lo_391};
  wire [511:0]  dataGroup_hi_391 = {dataGroup_hi_hi_391, dataGroup_hi_lo_391};
  wire [7:0]    dataGroup_7_24 = dataGroup_lo_391[423:416];
  wire [511:0]  dataGroup_lo_392 = {dataGroup_lo_hi_392, dataGroup_lo_lo_392};
  wire [511:0]  dataGroup_hi_392 = {dataGroup_hi_hi_392, dataGroup_hi_lo_392};
  wire [7:0]    dataGroup_8_24 = dataGroup_lo_392[479:472];
  wire [511:0]  dataGroup_lo_393 = {dataGroup_lo_hi_393, dataGroup_lo_lo_393};
  wire [511:0]  dataGroup_hi_393 = {dataGroup_hi_hi_393, dataGroup_hi_lo_393};
  wire [7:0]    dataGroup_9_24 = dataGroup_hi_393[23:16];
  wire [511:0]  dataGroup_lo_394 = {dataGroup_lo_hi_394, dataGroup_lo_lo_394};
  wire [511:0]  dataGroup_hi_394 = {dataGroup_hi_hi_394, dataGroup_hi_lo_394};
  wire [7:0]    dataGroup_10_24 = dataGroup_hi_394[79:72];
  wire [511:0]  dataGroup_lo_395 = {dataGroup_lo_hi_395, dataGroup_lo_lo_395};
  wire [511:0]  dataGroup_hi_395 = {dataGroup_hi_hi_395, dataGroup_hi_lo_395};
  wire [7:0]    dataGroup_11_24 = dataGroup_hi_395[135:128];
  wire [511:0]  dataGroup_lo_396 = {dataGroup_lo_hi_396, dataGroup_lo_lo_396};
  wire [511:0]  dataGroup_hi_396 = {dataGroup_hi_hi_396, dataGroup_hi_lo_396};
  wire [7:0]    dataGroup_12_24 = dataGroup_hi_396[191:184];
  wire [511:0]  dataGroup_lo_397 = {dataGroup_lo_hi_397, dataGroup_lo_lo_397};
  wire [511:0]  dataGroup_hi_397 = {dataGroup_hi_hi_397, dataGroup_hi_lo_397};
  wire [7:0]    dataGroup_13_24 = dataGroup_hi_397[247:240];
  wire [511:0]  dataGroup_lo_398 = {dataGroup_lo_hi_398, dataGroup_lo_lo_398};
  wire [511:0]  dataGroup_hi_398 = {dataGroup_hi_hi_398, dataGroup_hi_lo_398};
  wire [7:0]    dataGroup_14_24 = dataGroup_hi_398[303:296];
  wire [511:0]  dataGroup_lo_399 = {dataGroup_lo_hi_399, dataGroup_lo_lo_399};
  wire [511:0]  dataGroup_hi_399 = {dataGroup_hi_hi_399, dataGroup_hi_lo_399};
  wire [7:0]    dataGroup_15_24 = dataGroup_hi_399[359:352];
  wire [15:0]   res_lo_lo_lo_24 = {dataGroup_1_24, dataGroup_0_24};
  wire [15:0]   res_lo_lo_hi_24 = {dataGroup_3_24, dataGroup_2_24};
  wire [31:0]   res_lo_lo_24 = {res_lo_lo_hi_24, res_lo_lo_lo_24};
  wire [15:0]   res_lo_hi_lo_24 = {dataGroup_5_24, dataGroup_4_24};
  wire [15:0]   res_lo_hi_hi_24 = {dataGroup_7_24, dataGroup_6_24};
  wire [31:0]   res_lo_hi_24 = {res_lo_hi_hi_24, res_lo_hi_lo_24};
  wire [63:0]   res_lo_24 = {res_lo_hi_24, res_lo_lo_24};
  wire [15:0]   res_hi_lo_lo_24 = {dataGroup_9_24, dataGroup_8_24};
  wire [15:0]   res_hi_lo_hi_24 = {dataGroup_11_24, dataGroup_10_24};
  wire [31:0]   res_hi_lo_24 = {res_hi_lo_hi_24, res_hi_lo_lo_24};
  wire [15:0]   res_hi_hi_lo_24 = {dataGroup_13_24, dataGroup_12_24};
  wire [15:0]   res_hi_hi_hi_24 = {dataGroup_15_24, dataGroup_14_24};
  wire [31:0]   res_hi_hi_24 = {res_hi_hi_hi_24, res_hi_hi_lo_24};
  wire [63:0]   res_hi_24 = {res_hi_hi_24, res_hi_lo_24};
  wire [127:0]  res_51 = {res_hi_24, res_lo_24};
  wire [511:0]  dataGroup_lo_400 = {dataGroup_lo_hi_400, dataGroup_lo_lo_400};
  wire [511:0]  dataGroup_hi_400 = {dataGroup_hi_hi_400, dataGroup_hi_lo_400};
  wire [7:0]    dataGroup_0_25 = dataGroup_lo_400[39:32];
  wire [511:0]  dataGroup_lo_401 = {dataGroup_lo_hi_401, dataGroup_lo_lo_401};
  wire [511:0]  dataGroup_hi_401 = {dataGroup_hi_hi_401, dataGroup_hi_lo_401};
  wire [7:0]    dataGroup_1_25 = dataGroup_lo_401[95:88];
  wire [511:0]  dataGroup_lo_402 = {dataGroup_lo_hi_402, dataGroup_lo_lo_402};
  wire [511:0]  dataGroup_hi_402 = {dataGroup_hi_hi_402, dataGroup_hi_lo_402};
  wire [7:0]    dataGroup_2_25 = dataGroup_lo_402[151:144];
  wire [511:0]  dataGroup_lo_403 = {dataGroup_lo_hi_403, dataGroup_lo_lo_403};
  wire [511:0]  dataGroup_hi_403 = {dataGroup_hi_hi_403, dataGroup_hi_lo_403};
  wire [7:0]    dataGroup_3_25 = dataGroup_lo_403[207:200];
  wire [511:0]  dataGroup_lo_404 = {dataGroup_lo_hi_404, dataGroup_lo_lo_404};
  wire [511:0]  dataGroup_hi_404 = {dataGroup_hi_hi_404, dataGroup_hi_lo_404};
  wire [7:0]    dataGroup_4_25 = dataGroup_lo_404[263:256];
  wire [511:0]  dataGroup_lo_405 = {dataGroup_lo_hi_405, dataGroup_lo_lo_405};
  wire [511:0]  dataGroup_hi_405 = {dataGroup_hi_hi_405, dataGroup_hi_lo_405};
  wire [7:0]    dataGroup_5_25 = dataGroup_lo_405[319:312];
  wire [511:0]  dataGroup_lo_406 = {dataGroup_lo_hi_406, dataGroup_lo_lo_406};
  wire [511:0]  dataGroup_hi_406 = {dataGroup_hi_hi_406, dataGroup_hi_lo_406};
  wire [7:0]    dataGroup_6_25 = dataGroup_lo_406[375:368];
  wire [511:0]  dataGroup_lo_407 = {dataGroup_lo_hi_407, dataGroup_lo_lo_407};
  wire [511:0]  dataGroup_hi_407 = {dataGroup_hi_hi_407, dataGroup_hi_lo_407};
  wire [7:0]    dataGroup_7_25 = dataGroup_lo_407[431:424];
  wire [511:0]  dataGroup_lo_408 = {dataGroup_lo_hi_408, dataGroup_lo_lo_408};
  wire [511:0]  dataGroup_hi_408 = {dataGroup_hi_hi_408, dataGroup_hi_lo_408};
  wire [7:0]    dataGroup_8_25 = dataGroup_lo_408[487:480];
  wire [511:0]  dataGroup_lo_409 = {dataGroup_lo_hi_409, dataGroup_lo_lo_409};
  wire [511:0]  dataGroup_hi_409 = {dataGroup_hi_hi_409, dataGroup_hi_lo_409};
  wire [7:0]    dataGroup_9_25 = dataGroup_hi_409[31:24];
  wire [511:0]  dataGroup_lo_410 = {dataGroup_lo_hi_410, dataGroup_lo_lo_410};
  wire [511:0]  dataGroup_hi_410 = {dataGroup_hi_hi_410, dataGroup_hi_lo_410};
  wire [7:0]    dataGroup_10_25 = dataGroup_hi_410[87:80];
  wire [511:0]  dataGroup_lo_411 = {dataGroup_lo_hi_411, dataGroup_lo_lo_411};
  wire [511:0]  dataGroup_hi_411 = {dataGroup_hi_hi_411, dataGroup_hi_lo_411};
  wire [7:0]    dataGroup_11_25 = dataGroup_hi_411[143:136];
  wire [511:0]  dataGroup_lo_412 = {dataGroup_lo_hi_412, dataGroup_lo_lo_412};
  wire [511:0]  dataGroup_hi_412 = {dataGroup_hi_hi_412, dataGroup_hi_lo_412};
  wire [7:0]    dataGroup_12_25 = dataGroup_hi_412[199:192];
  wire [511:0]  dataGroup_lo_413 = {dataGroup_lo_hi_413, dataGroup_lo_lo_413};
  wire [511:0]  dataGroup_hi_413 = {dataGroup_hi_hi_413, dataGroup_hi_lo_413};
  wire [7:0]    dataGroup_13_25 = dataGroup_hi_413[255:248];
  wire [511:0]  dataGroup_lo_414 = {dataGroup_lo_hi_414, dataGroup_lo_lo_414};
  wire [511:0]  dataGroup_hi_414 = {dataGroup_hi_hi_414, dataGroup_hi_lo_414};
  wire [7:0]    dataGroup_14_25 = dataGroup_hi_414[311:304];
  wire [511:0]  dataGroup_lo_415 = {dataGroup_lo_hi_415, dataGroup_lo_lo_415};
  wire [511:0]  dataGroup_hi_415 = {dataGroup_hi_hi_415, dataGroup_hi_lo_415};
  wire [7:0]    dataGroup_15_25 = dataGroup_hi_415[367:360];
  wire [15:0]   res_lo_lo_lo_25 = {dataGroup_1_25, dataGroup_0_25};
  wire [15:0]   res_lo_lo_hi_25 = {dataGroup_3_25, dataGroup_2_25};
  wire [31:0]   res_lo_lo_25 = {res_lo_lo_hi_25, res_lo_lo_lo_25};
  wire [15:0]   res_lo_hi_lo_25 = {dataGroup_5_25, dataGroup_4_25};
  wire [15:0]   res_lo_hi_hi_25 = {dataGroup_7_25, dataGroup_6_25};
  wire [31:0]   res_lo_hi_25 = {res_lo_hi_hi_25, res_lo_hi_lo_25};
  wire [63:0]   res_lo_25 = {res_lo_hi_25, res_lo_lo_25};
  wire [15:0]   res_hi_lo_lo_25 = {dataGroup_9_25, dataGroup_8_25};
  wire [15:0]   res_hi_lo_hi_25 = {dataGroup_11_25, dataGroup_10_25};
  wire [31:0]   res_hi_lo_25 = {res_hi_lo_hi_25, res_hi_lo_lo_25};
  wire [15:0]   res_hi_hi_lo_25 = {dataGroup_13_25, dataGroup_12_25};
  wire [15:0]   res_hi_hi_hi_25 = {dataGroup_15_25, dataGroup_14_25};
  wire [31:0]   res_hi_hi_25 = {res_hi_hi_hi_25, res_hi_hi_lo_25};
  wire [63:0]   res_hi_25 = {res_hi_hi_25, res_hi_lo_25};
  wire [127:0]  res_52 = {res_hi_25, res_lo_25};
  wire [511:0]  dataGroup_lo_416 = {dataGroup_lo_hi_416, dataGroup_lo_lo_416};
  wire [511:0]  dataGroup_hi_416 = {dataGroup_hi_hi_416, dataGroup_hi_lo_416};
  wire [7:0]    dataGroup_0_26 = dataGroup_lo_416[47:40];
  wire [511:0]  dataGroup_lo_417 = {dataGroup_lo_hi_417, dataGroup_lo_lo_417};
  wire [511:0]  dataGroup_hi_417 = {dataGroup_hi_hi_417, dataGroup_hi_lo_417};
  wire [7:0]    dataGroup_1_26 = dataGroup_lo_417[103:96];
  wire [511:0]  dataGroup_lo_418 = {dataGroup_lo_hi_418, dataGroup_lo_lo_418};
  wire [511:0]  dataGroup_hi_418 = {dataGroup_hi_hi_418, dataGroup_hi_lo_418};
  wire [7:0]    dataGroup_2_26 = dataGroup_lo_418[159:152];
  wire [511:0]  dataGroup_lo_419 = {dataGroup_lo_hi_419, dataGroup_lo_lo_419};
  wire [511:0]  dataGroup_hi_419 = {dataGroup_hi_hi_419, dataGroup_hi_lo_419};
  wire [7:0]    dataGroup_3_26 = dataGroup_lo_419[215:208];
  wire [511:0]  dataGroup_lo_420 = {dataGroup_lo_hi_420, dataGroup_lo_lo_420};
  wire [511:0]  dataGroup_hi_420 = {dataGroup_hi_hi_420, dataGroup_hi_lo_420};
  wire [7:0]    dataGroup_4_26 = dataGroup_lo_420[271:264];
  wire [511:0]  dataGroup_lo_421 = {dataGroup_lo_hi_421, dataGroup_lo_lo_421};
  wire [511:0]  dataGroup_hi_421 = {dataGroup_hi_hi_421, dataGroup_hi_lo_421};
  wire [7:0]    dataGroup_5_26 = dataGroup_lo_421[327:320];
  wire [511:0]  dataGroup_lo_422 = {dataGroup_lo_hi_422, dataGroup_lo_lo_422};
  wire [511:0]  dataGroup_hi_422 = {dataGroup_hi_hi_422, dataGroup_hi_lo_422};
  wire [7:0]    dataGroup_6_26 = dataGroup_lo_422[383:376];
  wire [511:0]  dataGroup_lo_423 = {dataGroup_lo_hi_423, dataGroup_lo_lo_423};
  wire [511:0]  dataGroup_hi_423 = {dataGroup_hi_hi_423, dataGroup_hi_lo_423};
  wire [7:0]    dataGroup_7_26 = dataGroup_lo_423[439:432];
  wire [511:0]  dataGroup_lo_424 = {dataGroup_lo_hi_424, dataGroup_lo_lo_424};
  wire [511:0]  dataGroup_hi_424 = {dataGroup_hi_hi_424, dataGroup_hi_lo_424};
  wire [7:0]    dataGroup_8_26 = dataGroup_lo_424[495:488];
  wire [511:0]  dataGroup_lo_425 = {dataGroup_lo_hi_425, dataGroup_lo_lo_425};
  wire [511:0]  dataGroup_hi_425 = {dataGroup_hi_hi_425, dataGroup_hi_lo_425};
  wire [7:0]    dataGroup_9_26 = dataGroup_hi_425[39:32];
  wire [511:0]  dataGroup_lo_426 = {dataGroup_lo_hi_426, dataGroup_lo_lo_426};
  wire [511:0]  dataGroup_hi_426 = {dataGroup_hi_hi_426, dataGroup_hi_lo_426};
  wire [7:0]    dataGroup_10_26 = dataGroup_hi_426[95:88];
  wire [511:0]  dataGroup_lo_427 = {dataGroup_lo_hi_427, dataGroup_lo_lo_427};
  wire [511:0]  dataGroup_hi_427 = {dataGroup_hi_hi_427, dataGroup_hi_lo_427};
  wire [7:0]    dataGroup_11_26 = dataGroup_hi_427[151:144];
  wire [511:0]  dataGroup_lo_428 = {dataGroup_lo_hi_428, dataGroup_lo_lo_428};
  wire [511:0]  dataGroup_hi_428 = {dataGroup_hi_hi_428, dataGroup_hi_lo_428};
  wire [7:0]    dataGroup_12_26 = dataGroup_hi_428[207:200];
  wire [511:0]  dataGroup_lo_429 = {dataGroup_lo_hi_429, dataGroup_lo_lo_429};
  wire [511:0]  dataGroup_hi_429 = {dataGroup_hi_hi_429, dataGroup_hi_lo_429};
  wire [7:0]    dataGroup_13_26 = dataGroup_hi_429[263:256];
  wire [511:0]  dataGroup_lo_430 = {dataGroup_lo_hi_430, dataGroup_lo_lo_430};
  wire [511:0]  dataGroup_hi_430 = {dataGroup_hi_hi_430, dataGroup_hi_lo_430};
  wire [7:0]    dataGroup_14_26 = dataGroup_hi_430[319:312];
  wire [511:0]  dataGroup_lo_431 = {dataGroup_lo_hi_431, dataGroup_lo_lo_431};
  wire [511:0]  dataGroup_hi_431 = {dataGroup_hi_hi_431, dataGroup_hi_lo_431};
  wire [7:0]    dataGroup_15_26 = dataGroup_hi_431[375:368];
  wire [15:0]   res_lo_lo_lo_26 = {dataGroup_1_26, dataGroup_0_26};
  wire [15:0]   res_lo_lo_hi_26 = {dataGroup_3_26, dataGroup_2_26};
  wire [31:0]   res_lo_lo_26 = {res_lo_lo_hi_26, res_lo_lo_lo_26};
  wire [15:0]   res_lo_hi_lo_26 = {dataGroup_5_26, dataGroup_4_26};
  wire [15:0]   res_lo_hi_hi_26 = {dataGroup_7_26, dataGroup_6_26};
  wire [31:0]   res_lo_hi_26 = {res_lo_hi_hi_26, res_lo_hi_lo_26};
  wire [63:0]   res_lo_26 = {res_lo_hi_26, res_lo_lo_26};
  wire [15:0]   res_hi_lo_lo_26 = {dataGroup_9_26, dataGroup_8_26};
  wire [15:0]   res_hi_lo_hi_26 = {dataGroup_11_26, dataGroup_10_26};
  wire [31:0]   res_hi_lo_26 = {res_hi_lo_hi_26, res_hi_lo_lo_26};
  wire [15:0]   res_hi_hi_lo_26 = {dataGroup_13_26, dataGroup_12_26};
  wire [15:0]   res_hi_hi_hi_26 = {dataGroup_15_26, dataGroup_14_26};
  wire [31:0]   res_hi_hi_26 = {res_hi_hi_hi_26, res_hi_hi_lo_26};
  wire [63:0]   res_hi_26 = {res_hi_hi_26, res_hi_lo_26};
  wire [127:0]  res_53 = {res_hi_26, res_lo_26};
  wire [511:0]  dataGroup_lo_432 = {dataGroup_lo_hi_432, dataGroup_lo_lo_432};
  wire [511:0]  dataGroup_hi_432 = {dataGroup_hi_hi_432, dataGroup_hi_lo_432};
  wire [7:0]    dataGroup_0_27 = dataGroup_lo_432[55:48];
  wire [511:0]  dataGroup_lo_433 = {dataGroup_lo_hi_433, dataGroup_lo_lo_433};
  wire [511:0]  dataGroup_hi_433 = {dataGroup_hi_hi_433, dataGroup_hi_lo_433};
  wire [7:0]    dataGroup_1_27 = dataGroup_lo_433[111:104];
  wire [511:0]  dataGroup_lo_434 = {dataGroup_lo_hi_434, dataGroup_lo_lo_434};
  wire [511:0]  dataGroup_hi_434 = {dataGroup_hi_hi_434, dataGroup_hi_lo_434};
  wire [7:0]    dataGroup_2_27 = dataGroup_lo_434[167:160];
  wire [511:0]  dataGroup_lo_435 = {dataGroup_lo_hi_435, dataGroup_lo_lo_435};
  wire [511:0]  dataGroup_hi_435 = {dataGroup_hi_hi_435, dataGroup_hi_lo_435};
  wire [7:0]    dataGroup_3_27 = dataGroup_lo_435[223:216];
  wire [511:0]  dataGroup_lo_436 = {dataGroup_lo_hi_436, dataGroup_lo_lo_436};
  wire [511:0]  dataGroup_hi_436 = {dataGroup_hi_hi_436, dataGroup_hi_lo_436};
  wire [7:0]    dataGroup_4_27 = dataGroup_lo_436[279:272];
  wire [511:0]  dataGroup_lo_437 = {dataGroup_lo_hi_437, dataGroup_lo_lo_437};
  wire [511:0]  dataGroup_hi_437 = {dataGroup_hi_hi_437, dataGroup_hi_lo_437};
  wire [7:0]    dataGroup_5_27 = dataGroup_lo_437[335:328];
  wire [511:0]  dataGroup_lo_438 = {dataGroup_lo_hi_438, dataGroup_lo_lo_438};
  wire [511:0]  dataGroup_hi_438 = {dataGroup_hi_hi_438, dataGroup_hi_lo_438};
  wire [7:0]    dataGroup_6_27 = dataGroup_lo_438[391:384];
  wire [511:0]  dataGroup_lo_439 = {dataGroup_lo_hi_439, dataGroup_lo_lo_439};
  wire [511:0]  dataGroup_hi_439 = {dataGroup_hi_hi_439, dataGroup_hi_lo_439};
  wire [7:0]    dataGroup_7_27 = dataGroup_lo_439[447:440];
  wire [511:0]  dataGroup_lo_440 = {dataGroup_lo_hi_440, dataGroup_lo_lo_440};
  wire [511:0]  dataGroup_hi_440 = {dataGroup_hi_hi_440, dataGroup_hi_lo_440};
  wire [7:0]    dataGroup_8_27 = dataGroup_lo_440[503:496];
  wire [511:0]  dataGroup_lo_441 = {dataGroup_lo_hi_441, dataGroup_lo_lo_441};
  wire [511:0]  dataGroup_hi_441 = {dataGroup_hi_hi_441, dataGroup_hi_lo_441};
  wire [7:0]    dataGroup_9_27 = dataGroup_hi_441[47:40];
  wire [511:0]  dataGroup_lo_442 = {dataGroup_lo_hi_442, dataGroup_lo_lo_442};
  wire [511:0]  dataGroup_hi_442 = {dataGroup_hi_hi_442, dataGroup_hi_lo_442};
  wire [7:0]    dataGroup_10_27 = dataGroup_hi_442[103:96];
  wire [511:0]  dataGroup_lo_443 = {dataGroup_lo_hi_443, dataGroup_lo_lo_443};
  wire [511:0]  dataGroup_hi_443 = {dataGroup_hi_hi_443, dataGroup_hi_lo_443};
  wire [7:0]    dataGroup_11_27 = dataGroup_hi_443[159:152];
  wire [511:0]  dataGroup_lo_444 = {dataGroup_lo_hi_444, dataGroup_lo_lo_444};
  wire [511:0]  dataGroup_hi_444 = {dataGroup_hi_hi_444, dataGroup_hi_lo_444};
  wire [7:0]    dataGroup_12_27 = dataGroup_hi_444[215:208];
  wire [511:0]  dataGroup_lo_445 = {dataGroup_lo_hi_445, dataGroup_lo_lo_445};
  wire [511:0]  dataGroup_hi_445 = {dataGroup_hi_hi_445, dataGroup_hi_lo_445};
  wire [7:0]    dataGroup_13_27 = dataGroup_hi_445[271:264];
  wire [511:0]  dataGroup_lo_446 = {dataGroup_lo_hi_446, dataGroup_lo_lo_446};
  wire [511:0]  dataGroup_hi_446 = {dataGroup_hi_hi_446, dataGroup_hi_lo_446};
  wire [7:0]    dataGroup_14_27 = dataGroup_hi_446[327:320];
  wire [511:0]  dataGroup_lo_447 = {dataGroup_lo_hi_447, dataGroup_lo_lo_447};
  wire [511:0]  dataGroup_hi_447 = {dataGroup_hi_hi_447, dataGroup_hi_lo_447};
  wire [7:0]    dataGroup_15_27 = dataGroup_hi_447[383:376];
  wire [15:0]   res_lo_lo_lo_27 = {dataGroup_1_27, dataGroup_0_27};
  wire [15:0]   res_lo_lo_hi_27 = {dataGroup_3_27, dataGroup_2_27};
  wire [31:0]   res_lo_lo_27 = {res_lo_lo_hi_27, res_lo_lo_lo_27};
  wire [15:0]   res_lo_hi_lo_27 = {dataGroup_5_27, dataGroup_4_27};
  wire [15:0]   res_lo_hi_hi_27 = {dataGroup_7_27, dataGroup_6_27};
  wire [31:0]   res_lo_hi_27 = {res_lo_hi_hi_27, res_lo_hi_lo_27};
  wire [63:0]   res_lo_27 = {res_lo_hi_27, res_lo_lo_27};
  wire [15:0]   res_hi_lo_lo_27 = {dataGroup_9_27, dataGroup_8_27};
  wire [15:0]   res_hi_lo_hi_27 = {dataGroup_11_27, dataGroup_10_27};
  wire [31:0]   res_hi_lo_27 = {res_hi_lo_hi_27, res_hi_lo_lo_27};
  wire [15:0]   res_hi_hi_lo_27 = {dataGroup_13_27, dataGroup_12_27};
  wire [15:0]   res_hi_hi_hi_27 = {dataGroup_15_27, dataGroup_14_27};
  wire [31:0]   res_hi_hi_27 = {res_hi_hi_hi_27, res_hi_hi_lo_27};
  wire [63:0]   res_hi_27 = {res_hi_hi_27, res_hi_lo_27};
  wire [127:0]  res_54 = {res_hi_27, res_lo_27};
  wire [255:0]  lo_lo_6 = {res_49, res_48};
  wire [255:0]  lo_hi_6 = {res_51, res_50};
  wire [511:0]  lo_6 = {lo_hi_6, lo_lo_6};
  wire [255:0]  hi_lo_6 = {res_53, res_52};
  wire [255:0]  hi_hi_6 = {128'h0, res_54};
  wire [511:0]  hi_6 = {hi_hi_6, hi_lo_6};
  wire [1023:0] regroupLoadData_0_6 = {hi_6, lo_6};
  wire [511:0]  dataGroup_lo_448 = {dataGroup_lo_hi_448, dataGroup_lo_lo_448};
  wire [511:0]  dataGroup_hi_448 = {dataGroup_hi_hi_448, dataGroup_hi_lo_448};
  wire [7:0]    dataGroup_0_28 = dataGroup_lo_448[7:0];
  wire [511:0]  dataGroup_lo_449 = {dataGroup_lo_hi_449, dataGroup_lo_lo_449};
  wire [511:0]  dataGroup_hi_449 = {dataGroup_hi_hi_449, dataGroup_hi_lo_449};
  wire [7:0]    dataGroup_1_28 = dataGroup_lo_449[71:64];
  wire [511:0]  dataGroup_lo_450 = {dataGroup_lo_hi_450, dataGroup_lo_lo_450};
  wire [511:0]  dataGroup_hi_450 = {dataGroup_hi_hi_450, dataGroup_hi_lo_450};
  wire [7:0]    dataGroup_2_28 = dataGroup_lo_450[135:128];
  wire [511:0]  dataGroup_lo_451 = {dataGroup_lo_hi_451, dataGroup_lo_lo_451};
  wire [511:0]  dataGroup_hi_451 = {dataGroup_hi_hi_451, dataGroup_hi_lo_451};
  wire [7:0]    dataGroup_3_28 = dataGroup_lo_451[199:192];
  wire [511:0]  dataGroup_lo_452 = {dataGroup_lo_hi_452, dataGroup_lo_lo_452};
  wire [511:0]  dataGroup_hi_452 = {dataGroup_hi_hi_452, dataGroup_hi_lo_452};
  wire [7:0]    dataGroup_4_28 = dataGroup_lo_452[263:256];
  wire [511:0]  dataGroup_lo_453 = {dataGroup_lo_hi_453, dataGroup_lo_lo_453};
  wire [511:0]  dataGroup_hi_453 = {dataGroup_hi_hi_453, dataGroup_hi_lo_453};
  wire [7:0]    dataGroup_5_28 = dataGroup_lo_453[327:320];
  wire [511:0]  dataGroup_lo_454 = {dataGroup_lo_hi_454, dataGroup_lo_lo_454};
  wire [511:0]  dataGroup_hi_454 = {dataGroup_hi_hi_454, dataGroup_hi_lo_454};
  wire [7:0]    dataGroup_6_28 = dataGroup_lo_454[391:384];
  wire [511:0]  dataGroup_lo_455 = {dataGroup_lo_hi_455, dataGroup_lo_lo_455};
  wire [511:0]  dataGroup_hi_455 = {dataGroup_hi_hi_455, dataGroup_hi_lo_455};
  wire [7:0]    dataGroup_7_28 = dataGroup_lo_455[455:448];
  wire [511:0]  dataGroup_lo_456 = {dataGroup_lo_hi_456, dataGroup_lo_lo_456};
  wire [511:0]  dataGroup_hi_456 = {dataGroup_hi_hi_456, dataGroup_hi_lo_456};
  wire [7:0]    dataGroup_8_28 = dataGroup_hi_456[7:0];
  wire [511:0]  dataGroup_lo_457 = {dataGroup_lo_hi_457, dataGroup_lo_lo_457};
  wire [511:0]  dataGroup_hi_457 = {dataGroup_hi_hi_457, dataGroup_hi_lo_457};
  wire [7:0]    dataGroup_9_28 = dataGroup_hi_457[71:64];
  wire [511:0]  dataGroup_lo_458 = {dataGroup_lo_hi_458, dataGroup_lo_lo_458};
  wire [511:0]  dataGroup_hi_458 = {dataGroup_hi_hi_458, dataGroup_hi_lo_458};
  wire [7:0]    dataGroup_10_28 = dataGroup_hi_458[135:128];
  wire [511:0]  dataGroup_lo_459 = {dataGroup_lo_hi_459, dataGroup_lo_lo_459};
  wire [511:0]  dataGroup_hi_459 = {dataGroup_hi_hi_459, dataGroup_hi_lo_459};
  wire [7:0]    dataGroup_11_28 = dataGroup_hi_459[199:192];
  wire [511:0]  dataGroup_lo_460 = {dataGroup_lo_hi_460, dataGroup_lo_lo_460};
  wire [511:0]  dataGroup_hi_460 = {dataGroup_hi_hi_460, dataGroup_hi_lo_460};
  wire [7:0]    dataGroup_12_28 = dataGroup_hi_460[263:256];
  wire [511:0]  dataGroup_lo_461 = {dataGroup_lo_hi_461, dataGroup_lo_lo_461};
  wire [511:0]  dataGroup_hi_461 = {dataGroup_hi_hi_461, dataGroup_hi_lo_461};
  wire [7:0]    dataGroup_13_28 = dataGroup_hi_461[327:320];
  wire [511:0]  dataGroup_lo_462 = {dataGroup_lo_hi_462, dataGroup_lo_lo_462};
  wire [511:0]  dataGroup_hi_462 = {dataGroup_hi_hi_462, dataGroup_hi_lo_462};
  wire [7:0]    dataGroup_14_28 = dataGroup_hi_462[391:384];
  wire [511:0]  dataGroup_lo_463 = {dataGroup_lo_hi_463, dataGroup_lo_lo_463};
  wire [511:0]  dataGroup_hi_463 = {dataGroup_hi_hi_463, dataGroup_hi_lo_463};
  wire [7:0]    dataGroup_15_28 = dataGroup_hi_463[455:448];
  wire [15:0]   res_lo_lo_lo_28 = {dataGroup_1_28, dataGroup_0_28};
  wire [15:0]   res_lo_lo_hi_28 = {dataGroup_3_28, dataGroup_2_28};
  wire [31:0]   res_lo_lo_28 = {res_lo_lo_hi_28, res_lo_lo_lo_28};
  wire [15:0]   res_lo_hi_lo_28 = {dataGroup_5_28, dataGroup_4_28};
  wire [15:0]   res_lo_hi_hi_28 = {dataGroup_7_28, dataGroup_6_28};
  wire [31:0]   res_lo_hi_28 = {res_lo_hi_hi_28, res_lo_hi_lo_28};
  wire [63:0]   res_lo_28 = {res_lo_hi_28, res_lo_lo_28};
  wire [15:0]   res_hi_lo_lo_28 = {dataGroup_9_28, dataGroup_8_28};
  wire [15:0]   res_hi_lo_hi_28 = {dataGroup_11_28, dataGroup_10_28};
  wire [31:0]   res_hi_lo_28 = {res_hi_lo_hi_28, res_hi_lo_lo_28};
  wire [15:0]   res_hi_hi_lo_28 = {dataGroup_13_28, dataGroup_12_28};
  wire [15:0]   res_hi_hi_hi_28 = {dataGroup_15_28, dataGroup_14_28};
  wire [31:0]   res_hi_hi_28 = {res_hi_hi_hi_28, res_hi_hi_lo_28};
  wire [63:0]   res_hi_28 = {res_hi_hi_28, res_hi_lo_28};
  wire [127:0]  res_56 = {res_hi_28, res_lo_28};
  wire [511:0]  dataGroup_lo_464 = {dataGroup_lo_hi_464, dataGroup_lo_lo_464};
  wire [511:0]  dataGroup_hi_464 = {dataGroup_hi_hi_464, dataGroup_hi_lo_464};
  wire [7:0]    dataGroup_0_29 = dataGroup_lo_464[15:8];
  wire [511:0]  dataGroup_lo_465 = {dataGroup_lo_hi_465, dataGroup_lo_lo_465};
  wire [511:0]  dataGroup_hi_465 = {dataGroup_hi_hi_465, dataGroup_hi_lo_465};
  wire [7:0]    dataGroup_1_29 = dataGroup_lo_465[79:72];
  wire [511:0]  dataGroup_lo_466 = {dataGroup_lo_hi_466, dataGroup_lo_lo_466};
  wire [511:0]  dataGroup_hi_466 = {dataGroup_hi_hi_466, dataGroup_hi_lo_466};
  wire [7:0]    dataGroup_2_29 = dataGroup_lo_466[143:136];
  wire [511:0]  dataGroup_lo_467 = {dataGroup_lo_hi_467, dataGroup_lo_lo_467};
  wire [511:0]  dataGroup_hi_467 = {dataGroup_hi_hi_467, dataGroup_hi_lo_467};
  wire [7:0]    dataGroup_3_29 = dataGroup_lo_467[207:200];
  wire [511:0]  dataGroup_lo_468 = {dataGroup_lo_hi_468, dataGroup_lo_lo_468};
  wire [511:0]  dataGroup_hi_468 = {dataGroup_hi_hi_468, dataGroup_hi_lo_468};
  wire [7:0]    dataGroup_4_29 = dataGroup_lo_468[271:264];
  wire [511:0]  dataGroup_lo_469 = {dataGroup_lo_hi_469, dataGroup_lo_lo_469};
  wire [511:0]  dataGroup_hi_469 = {dataGroup_hi_hi_469, dataGroup_hi_lo_469};
  wire [7:0]    dataGroup_5_29 = dataGroup_lo_469[335:328];
  wire [511:0]  dataGroup_lo_470 = {dataGroup_lo_hi_470, dataGroup_lo_lo_470};
  wire [511:0]  dataGroup_hi_470 = {dataGroup_hi_hi_470, dataGroup_hi_lo_470};
  wire [7:0]    dataGroup_6_29 = dataGroup_lo_470[399:392];
  wire [511:0]  dataGroup_lo_471 = {dataGroup_lo_hi_471, dataGroup_lo_lo_471};
  wire [511:0]  dataGroup_hi_471 = {dataGroup_hi_hi_471, dataGroup_hi_lo_471};
  wire [7:0]    dataGroup_7_29 = dataGroup_lo_471[463:456];
  wire [511:0]  dataGroup_lo_472 = {dataGroup_lo_hi_472, dataGroup_lo_lo_472};
  wire [511:0]  dataGroup_hi_472 = {dataGroup_hi_hi_472, dataGroup_hi_lo_472};
  wire [7:0]    dataGroup_8_29 = dataGroup_hi_472[15:8];
  wire [511:0]  dataGroup_lo_473 = {dataGroup_lo_hi_473, dataGroup_lo_lo_473};
  wire [511:0]  dataGroup_hi_473 = {dataGroup_hi_hi_473, dataGroup_hi_lo_473};
  wire [7:0]    dataGroup_9_29 = dataGroup_hi_473[79:72];
  wire [511:0]  dataGroup_lo_474 = {dataGroup_lo_hi_474, dataGroup_lo_lo_474};
  wire [511:0]  dataGroup_hi_474 = {dataGroup_hi_hi_474, dataGroup_hi_lo_474};
  wire [7:0]    dataGroup_10_29 = dataGroup_hi_474[143:136];
  wire [511:0]  dataGroup_lo_475 = {dataGroup_lo_hi_475, dataGroup_lo_lo_475};
  wire [511:0]  dataGroup_hi_475 = {dataGroup_hi_hi_475, dataGroup_hi_lo_475};
  wire [7:0]    dataGroup_11_29 = dataGroup_hi_475[207:200];
  wire [511:0]  dataGroup_lo_476 = {dataGroup_lo_hi_476, dataGroup_lo_lo_476};
  wire [511:0]  dataGroup_hi_476 = {dataGroup_hi_hi_476, dataGroup_hi_lo_476};
  wire [7:0]    dataGroup_12_29 = dataGroup_hi_476[271:264];
  wire [511:0]  dataGroup_lo_477 = {dataGroup_lo_hi_477, dataGroup_lo_lo_477};
  wire [511:0]  dataGroup_hi_477 = {dataGroup_hi_hi_477, dataGroup_hi_lo_477};
  wire [7:0]    dataGroup_13_29 = dataGroup_hi_477[335:328];
  wire [511:0]  dataGroup_lo_478 = {dataGroup_lo_hi_478, dataGroup_lo_lo_478};
  wire [511:0]  dataGroup_hi_478 = {dataGroup_hi_hi_478, dataGroup_hi_lo_478};
  wire [7:0]    dataGroup_14_29 = dataGroup_hi_478[399:392];
  wire [511:0]  dataGroup_lo_479 = {dataGroup_lo_hi_479, dataGroup_lo_lo_479};
  wire [511:0]  dataGroup_hi_479 = {dataGroup_hi_hi_479, dataGroup_hi_lo_479};
  wire [7:0]    dataGroup_15_29 = dataGroup_hi_479[463:456];
  wire [15:0]   res_lo_lo_lo_29 = {dataGroup_1_29, dataGroup_0_29};
  wire [15:0]   res_lo_lo_hi_29 = {dataGroup_3_29, dataGroup_2_29};
  wire [31:0]   res_lo_lo_29 = {res_lo_lo_hi_29, res_lo_lo_lo_29};
  wire [15:0]   res_lo_hi_lo_29 = {dataGroup_5_29, dataGroup_4_29};
  wire [15:0]   res_lo_hi_hi_29 = {dataGroup_7_29, dataGroup_6_29};
  wire [31:0]   res_lo_hi_29 = {res_lo_hi_hi_29, res_lo_hi_lo_29};
  wire [63:0]   res_lo_29 = {res_lo_hi_29, res_lo_lo_29};
  wire [15:0]   res_hi_lo_lo_29 = {dataGroup_9_29, dataGroup_8_29};
  wire [15:0]   res_hi_lo_hi_29 = {dataGroup_11_29, dataGroup_10_29};
  wire [31:0]   res_hi_lo_29 = {res_hi_lo_hi_29, res_hi_lo_lo_29};
  wire [15:0]   res_hi_hi_lo_29 = {dataGroup_13_29, dataGroup_12_29};
  wire [15:0]   res_hi_hi_hi_29 = {dataGroup_15_29, dataGroup_14_29};
  wire [31:0]   res_hi_hi_29 = {res_hi_hi_hi_29, res_hi_hi_lo_29};
  wire [63:0]   res_hi_29 = {res_hi_hi_29, res_hi_lo_29};
  wire [127:0]  res_57 = {res_hi_29, res_lo_29};
  wire [511:0]  dataGroup_lo_480 = {dataGroup_lo_hi_480, dataGroup_lo_lo_480};
  wire [511:0]  dataGroup_hi_480 = {dataGroup_hi_hi_480, dataGroup_hi_lo_480};
  wire [7:0]    dataGroup_0_30 = dataGroup_lo_480[23:16];
  wire [511:0]  dataGroup_lo_481 = {dataGroup_lo_hi_481, dataGroup_lo_lo_481};
  wire [511:0]  dataGroup_hi_481 = {dataGroup_hi_hi_481, dataGroup_hi_lo_481};
  wire [7:0]    dataGroup_1_30 = dataGroup_lo_481[87:80];
  wire [511:0]  dataGroup_lo_482 = {dataGroup_lo_hi_482, dataGroup_lo_lo_482};
  wire [511:0]  dataGroup_hi_482 = {dataGroup_hi_hi_482, dataGroup_hi_lo_482};
  wire [7:0]    dataGroup_2_30 = dataGroup_lo_482[151:144];
  wire [511:0]  dataGroup_lo_483 = {dataGroup_lo_hi_483, dataGroup_lo_lo_483};
  wire [511:0]  dataGroup_hi_483 = {dataGroup_hi_hi_483, dataGroup_hi_lo_483};
  wire [7:0]    dataGroup_3_30 = dataGroup_lo_483[215:208];
  wire [511:0]  dataGroup_lo_484 = {dataGroup_lo_hi_484, dataGroup_lo_lo_484};
  wire [511:0]  dataGroup_hi_484 = {dataGroup_hi_hi_484, dataGroup_hi_lo_484};
  wire [7:0]    dataGroup_4_30 = dataGroup_lo_484[279:272];
  wire [511:0]  dataGroup_lo_485 = {dataGroup_lo_hi_485, dataGroup_lo_lo_485};
  wire [511:0]  dataGroup_hi_485 = {dataGroup_hi_hi_485, dataGroup_hi_lo_485};
  wire [7:0]    dataGroup_5_30 = dataGroup_lo_485[343:336];
  wire [511:0]  dataGroup_lo_486 = {dataGroup_lo_hi_486, dataGroup_lo_lo_486};
  wire [511:0]  dataGroup_hi_486 = {dataGroup_hi_hi_486, dataGroup_hi_lo_486};
  wire [7:0]    dataGroup_6_30 = dataGroup_lo_486[407:400];
  wire [511:0]  dataGroup_lo_487 = {dataGroup_lo_hi_487, dataGroup_lo_lo_487};
  wire [511:0]  dataGroup_hi_487 = {dataGroup_hi_hi_487, dataGroup_hi_lo_487};
  wire [7:0]    dataGroup_7_30 = dataGroup_lo_487[471:464];
  wire [511:0]  dataGroup_lo_488 = {dataGroup_lo_hi_488, dataGroup_lo_lo_488};
  wire [511:0]  dataGroup_hi_488 = {dataGroup_hi_hi_488, dataGroup_hi_lo_488};
  wire [7:0]    dataGroup_8_30 = dataGroup_hi_488[23:16];
  wire [511:0]  dataGroup_lo_489 = {dataGroup_lo_hi_489, dataGroup_lo_lo_489};
  wire [511:0]  dataGroup_hi_489 = {dataGroup_hi_hi_489, dataGroup_hi_lo_489};
  wire [7:0]    dataGroup_9_30 = dataGroup_hi_489[87:80];
  wire [511:0]  dataGroup_lo_490 = {dataGroup_lo_hi_490, dataGroup_lo_lo_490};
  wire [511:0]  dataGroup_hi_490 = {dataGroup_hi_hi_490, dataGroup_hi_lo_490};
  wire [7:0]    dataGroup_10_30 = dataGroup_hi_490[151:144];
  wire [511:0]  dataGroup_lo_491 = {dataGroup_lo_hi_491, dataGroup_lo_lo_491};
  wire [511:0]  dataGroup_hi_491 = {dataGroup_hi_hi_491, dataGroup_hi_lo_491};
  wire [7:0]    dataGroup_11_30 = dataGroup_hi_491[215:208];
  wire [511:0]  dataGroup_lo_492 = {dataGroup_lo_hi_492, dataGroup_lo_lo_492};
  wire [511:0]  dataGroup_hi_492 = {dataGroup_hi_hi_492, dataGroup_hi_lo_492};
  wire [7:0]    dataGroup_12_30 = dataGroup_hi_492[279:272];
  wire [511:0]  dataGroup_lo_493 = {dataGroup_lo_hi_493, dataGroup_lo_lo_493};
  wire [511:0]  dataGroup_hi_493 = {dataGroup_hi_hi_493, dataGroup_hi_lo_493};
  wire [7:0]    dataGroup_13_30 = dataGroup_hi_493[343:336];
  wire [511:0]  dataGroup_lo_494 = {dataGroup_lo_hi_494, dataGroup_lo_lo_494};
  wire [511:0]  dataGroup_hi_494 = {dataGroup_hi_hi_494, dataGroup_hi_lo_494};
  wire [7:0]    dataGroup_14_30 = dataGroup_hi_494[407:400];
  wire [511:0]  dataGroup_lo_495 = {dataGroup_lo_hi_495, dataGroup_lo_lo_495};
  wire [511:0]  dataGroup_hi_495 = {dataGroup_hi_hi_495, dataGroup_hi_lo_495};
  wire [7:0]    dataGroup_15_30 = dataGroup_hi_495[471:464];
  wire [15:0]   res_lo_lo_lo_30 = {dataGroup_1_30, dataGroup_0_30};
  wire [15:0]   res_lo_lo_hi_30 = {dataGroup_3_30, dataGroup_2_30};
  wire [31:0]   res_lo_lo_30 = {res_lo_lo_hi_30, res_lo_lo_lo_30};
  wire [15:0]   res_lo_hi_lo_30 = {dataGroup_5_30, dataGroup_4_30};
  wire [15:0]   res_lo_hi_hi_30 = {dataGroup_7_30, dataGroup_6_30};
  wire [31:0]   res_lo_hi_30 = {res_lo_hi_hi_30, res_lo_hi_lo_30};
  wire [63:0]   res_lo_30 = {res_lo_hi_30, res_lo_lo_30};
  wire [15:0]   res_hi_lo_lo_30 = {dataGroup_9_30, dataGroup_8_30};
  wire [15:0]   res_hi_lo_hi_30 = {dataGroup_11_30, dataGroup_10_30};
  wire [31:0]   res_hi_lo_30 = {res_hi_lo_hi_30, res_hi_lo_lo_30};
  wire [15:0]   res_hi_hi_lo_30 = {dataGroup_13_30, dataGroup_12_30};
  wire [15:0]   res_hi_hi_hi_30 = {dataGroup_15_30, dataGroup_14_30};
  wire [31:0]   res_hi_hi_30 = {res_hi_hi_hi_30, res_hi_hi_lo_30};
  wire [63:0]   res_hi_30 = {res_hi_hi_30, res_hi_lo_30};
  wire [127:0]  res_58 = {res_hi_30, res_lo_30};
  wire [511:0]  dataGroup_lo_496 = {dataGroup_lo_hi_496, dataGroup_lo_lo_496};
  wire [511:0]  dataGroup_hi_496 = {dataGroup_hi_hi_496, dataGroup_hi_lo_496};
  wire [7:0]    dataGroup_0_31 = dataGroup_lo_496[31:24];
  wire [511:0]  dataGroup_lo_497 = {dataGroup_lo_hi_497, dataGroup_lo_lo_497};
  wire [511:0]  dataGroup_hi_497 = {dataGroup_hi_hi_497, dataGroup_hi_lo_497};
  wire [7:0]    dataGroup_1_31 = dataGroup_lo_497[95:88];
  wire [511:0]  dataGroup_lo_498 = {dataGroup_lo_hi_498, dataGroup_lo_lo_498};
  wire [511:0]  dataGroup_hi_498 = {dataGroup_hi_hi_498, dataGroup_hi_lo_498};
  wire [7:0]    dataGroup_2_31 = dataGroup_lo_498[159:152];
  wire [511:0]  dataGroup_lo_499 = {dataGroup_lo_hi_499, dataGroup_lo_lo_499};
  wire [511:0]  dataGroup_hi_499 = {dataGroup_hi_hi_499, dataGroup_hi_lo_499};
  wire [7:0]    dataGroup_3_31 = dataGroup_lo_499[223:216];
  wire [511:0]  dataGroup_lo_500 = {dataGroup_lo_hi_500, dataGroup_lo_lo_500};
  wire [511:0]  dataGroup_hi_500 = {dataGroup_hi_hi_500, dataGroup_hi_lo_500};
  wire [7:0]    dataGroup_4_31 = dataGroup_lo_500[287:280];
  wire [511:0]  dataGroup_lo_501 = {dataGroup_lo_hi_501, dataGroup_lo_lo_501};
  wire [511:0]  dataGroup_hi_501 = {dataGroup_hi_hi_501, dataGroup_hi_lo_501};
  wire [7:0]    dataGroup_5_31 = dataGroup_lo_501[351:344];
  wire [511:0]  dataGroup_lo_502 = {dataGroup_lo_hi_502, dataGroup_lo_lo_502};
  wire [511:0]  dataGroup_hi_502 = {dataGroup_hi_hi_502, dataGroup_hi_lo_502};
  wire [7:0]    dataGroup_6_31 = dataGroup_lo_502[415:408];
  wire [511:0]  dataGroup_lo_503 = {dataGroup_lo_hi_503, dataGroup_lo_lo_503};
  wire [511:0]  dataGroup_hi_503 = {dataGroup_hi_hi_503, dataGroup_hi_lo_503};
  wire [7:0]    dataGroup_7_31 = dataGroup_lo_503[479:472];
  wire [511:0]  dataGroup_lo_504 = {dataGroup_lo_hi_504, dataGroup_lo_lo_504};
  wire [511:0]  dataGroup_hi_504 = {dataGroup_hi_hi_504, dataGroup_hi_lo_504};
  wire [7:0]    dataGroup_8_31 = dataGroup_hi_504[31:24];
  wire [511:0]  dataGroup_lo_505 = {dataGroup_lo_hi_505, dataGroup_lo_lo_505};
  wire [511:0]  dataGroup_hi_505 = {dataGroup_hi_hi_505, dataGroup_hi_lo_505};
  wire [7:0]    dataGroup_9_31 = dataGroup_hi_505[95:88];
  wire [511:0]  dataGroup_lo_506 = {dataGroup_lo_hi_506, dataGroup_lo_lo_506};
  wire [511:0]  dataGroup_hi_506 = {dataGroup_hi_hi_506, dataGroup_hi_lo_506};
  wire [7:0]    dataGroup_10_31 = dataGroup_hi_506[159:152];
  wire [511:0]  dataGroup_lo_507 = {dataGroup_lo_hi_507, dataGroup_lo_lo_507};
  wire [511:0]  dataGroup_hi_507 = {dataGroup_hi_hi_507, dataGroup_hi_lo_507};
  wire [7:0]    dataGroup_11_31 = dataGroup_hi_507[223:216];
  wire [511:0]  dataGroup_lo_508 = {dataGroup_lo_hi_508, dataGroup_lo_lo_508};
  wire [511:0]  dataGroup_hi_508 = {dataGroup_hi_hi_508, dataGroup_hi_lo_508};
  wire [7:0]    dataGroup_12_31 = dataGroup_hi_508[287:280];
  wire [511:0]  dataGroup_lo_509 = {dataGroup_lo_hi_509, dataGroup_lo_lo_509};
  wire [511:0]  dataGroup_hi_509 = {dataGroup_hi_hi_509, dataGroup_hi_lo_509};
  wire [7:0]    dataGroup_13_31 = dataGroup_hi_509[351:344];
  wire [511:0]  dataGroup_lo_510 = {dataGroup_lo_hi_510, dataGroup_lo_lo_510};
  wire [511:0]  dataGroup_hi_510 = {dataGroup_hi_hi_510, dataGroup_hi_lo_510};
  wire [7:0]    dataGroup_14_31 = dataGroup_hi_510[415:408];
  wire [511:0]  dataGroup_lo_511 = {dataGroup_lo_hi_511, dataGroup_lo_lo_511};
  wire [511:0]  dataGroup_hi_511 = {dataGroup_hi_hi_511, dataGroup_hi_lo_511};
  wire [7:0]    dataGroup_15_31 = dataGroup_hi_511[479:472];
  wire [15:0]   res_lo_lo_lo_31 = {dataGroup_1_31, dataGroup_0_31};
  wire [15:0]   res_lo_lo_hi_31 = {dataGroup_3_31, dataGroup_2_31};
  wire [31:0]   res_lo_lo_31 = {res_lo_lo_hi_31, res_lo_lo_lo_31};
  wire [15:0]   res_lo_hi_lo_31 = {dataGroup_5_31, dataGroup_4_31};
  wire [15:0]   res_lo_hi_hi_31 = {dataGroup_7_31, dataGroup_6_31};
  wire [31:0]   res_lo_hi_31 = {res_lo_hi_hi_31, res_lo_hi_lo_31};
  wire [63:0]   res_lo_31 = {res_lo_hi_31, res_lo_lo_31};
  wire [15:0]   res_hi_lo_lo_31 = {dataGroup_9_31, dataGroup_8_31};
  wire [15:0]   res_hi_lo_hi_31 = {dataGroup_11_31, dataGroup_10_31};
  wire [31:0]   res_hi_lo_31 = {res_hi_lo_hi_31, res_hi_lo_lo_31};
  wire [15:0]   res_hi_hi_lo_31 = {dataGroup_13_31, dataGroup_12_31};
  wire [15:0]   res_hi_hi_hi_31 = {dataGroup_15_31, dataGroup_14_31};
  wire [31:0]   res_hi_hi_31 = {res_hi_hi_hi_31, res_hi_hi_lo_31};
  wire [63:0]   res_hi_31 = {res_hi_hi_31, res_hi_lo_31};
  wire [127:0]  res_59 = {res_hi_31, res_lo_31};
  wire [511:0]  dataGroup_lo_512 = {dataGroup_lo_hi_512, dataGroup_lo_lo_512};
  wire [511:0]  dataGroup_hi_512 = {dataGroup_hi_hi_512, dataGroup_hi_lo_512};
  wire [7:0]    dataGroup_0_32 = dataGroup_lo_512[39:32];
  wire [511:0]  dataGroup_lo_513 = {dataGroup_lo_hi_513, dataGroup_lo_lo_513};
  wire [511:0]  dataGroup_hi_513 = {dataGroup_hi_hi_513, dataGroup_hi_lo_513};
  wire [7:0]    dataGroup_1_32 = dataGroup_lo_513[103:96];
  wire [511:0]  dataGroup_lo_514 = {dataGroup_lo_hi_514, dataGroup_lo_lo_514};
  wire [511:0]  dataGroup_hi_514 = {dataGroup_hi_hi_514, dataGroup_hi_lo_514};
  wire [7:0]    dataGroup_2_32 = dataGroup_lo_514[167:160];
  wire [511:0]  dataGroup_lo_515 = {dataGroup_lo_hi_515, dataGroup_lo_lo_515};
  wire [511:0]  dataGroup_hi_515 = {dataGroup_hi_hi_515, dataGroup_hi_lo_515};
  wire [7:0]    dataGroup_3_32 = dataGroup_lo_515[231:224];
  wire [511:0]  dataGroup_lo_516 = {dataGroup_lo_hi_516, dataGroup_lo_lo_516};
  wire [511:0]  dataGroup_hi_516 = {dataGroup_hi_hi_516, dataGroup_hi_lo_516};
  wire [7:0]    dataGroup_4_32 = dataGroup_lo_516[295:288];
  wire [511:0]  dataGroup_lo_517 = {dataGroup_lo_hi_517, dataGroup_lo_lo_517};
  wire [511:0]  dataGroup_hi_517 = {dataGroup_hi_hi_517, dataGroup_hi_lo_517};
  wire [7:0]    dataGroup_5_32 = dataGroup_lo_517[359:352];
  wire [511:0]  dataGroup_lo_518 = {dataGroup_lo_hi_518, dataGroup_lo_lo_518};
  wire [511:0]  dataGroup_hi_518 = {dataGroup_hi_hi_518, dataGroup_hi_lo_518};
  wire [7:0]    dataGroup_6_32 = dataGroup_lo_518[423:416];
  wire [511:0]  dataGroup_lo_519 = {dataGroup_lo_hi_519, dataGroup_lo_lo_519};
  wire [511:0]  dataGroup_hi_519 = {dataGroup_hi_hi_519, dataGroup_hi_lo_519};
  wire [7:0]    dataGroup_7_32 = dataGroup_lo_519[487:480];
  wire [511:0]  dataGroup_lo_520 = {dataGroup_lo_hi_520, dataGroup_lo_lo_520};
  wire [511:0]  dataGroup_hi_520 = {dataGroup_hi_hi_520, dataGroup_hi_lo_520};
  wire [7:0]    dataGroup_8_32 = dataGroup_hi_520[39:32];
  wire [511:0]  dataGroup_lo_521 = {dataGroup_lo_hi_521, dataGroup_lo_lo_521};
  wire [511:0]  dataGroup_hi_521 = {dataGroup_hi_hi_521, dataGroup_hi_lo_521};
  wire [7:0]    dataGroup_9_32 = dataGroup_hi_521[103:96];
  wire [511:0]  dataGroup_lo_522 = {dataGroup_lo_hi_522, dataGroup_lo_lo_522};
  wire [511:0]  dataGroup_hi_522 = {dataGroup_hi_hi_522, dataGroup_hi_lo_522};
  wire [7:0]    dataGroup_10_32 = dataGroup_hi_522[167:160];
  wire [511:0]  dataGroup_lo_523 = {dataGroup_lo_hi_523, dataGroup_lo_lo_523};
  wire [511:0]  dataGroup_hi_523 = {dataGroup_hi_hi_523, dataGroup_hi_lo_523};
  wire [7:0]    dataGroup_11_32 = dataGroup_hi_523[231:224];
  wire [511:0]  dataGroup_lo_524 = {dataGroup_lo_hi_524, dataGroup_lo_lo_524};
  wire [511:0]  dataGroup_hi_524 = {dataGroup_hi_hi_524, dataGroup_hi_lo_524};
  wire [7:0]    dataGroup_12_32 = dataGroup_hi_524[295:288];
  wire [511:0]  dataGroup_lo_525 = {dataGroup_lo_hi_525, dataGroup_lo_lo_525};
  wire [511:0]  dataGroup_hi_525 = {dataGroup_hi_hi_525, dataGroup_hi_lo_525};
  wire [7:0]    dataGroup_13_32 = dataGroup_hi_525[359:352];
  wire [511:0]  dataGroup_lo_526 = {dataGroup_lo_hi_526, dataGroup_lo_lo_526};
  wire [511:0]  dataGroup_hi_526 = {dataGroup_hi_hi_526, dataGroup_hi_lo_526};
  wire [7:0]    dataGroup_14_32 = dataGroup_hi_526[423:416];
  wire [511:0]  dataGroup_lo_527 = {dataGroup_lo_hi_527, dataGroup_lo_lo_527};
  wire [511:0]  dataGroup_hi_527 = {dataGroup_hi_hi_527, dataGroup_hi_lo_527};
  wire [7:0]    dataGroup_15_32 = dataGroup_hi_527[487:480];
  wire [15:0]   res_lo_lo_lo_32 = {dataGroup_1_32, dataGroup_0_32};
  wire [15:0]   res_lo_lo_hi_32 = {dataGroup_3_32, dataGroup_2_32};
  wire [31:0]   res_lo_lo_32 = {res_lo_lo_hi_32, res_lo_lo_lo_32};
  wire [15:0]   res_lo_hi_lo_32 = {dataGroup_5_32, dataGroup_4_32};
  wire [15:0]   res_lo_hi_hi_32 = {dataGroup_7_32, dataGroup_6_32};
  wire [31:0]   res_lo_hi_32 = {res_lo_hi_hi_32, res_lo_hi_lo_32};
  wire [63:0]   res_lo_32 = {res_lo_hi_32, res_lo_lo_32};
  wire [15:0]   res_hi_lo_lo_32 = {dataGroup_9_32, dataGroup_8_32};
  wire [15:0]   res_hi_lo_hi_32 = {dataGroup_11_32, dataGroup_10_32};
  wire [31:0]   res_hi_lo_32 = {res_hi_lo_hi_32, res_hi_lo_lo_32};
  wire [15:0]   res_hi_hi_lo_32 = {dataGroup_13_32, dataGroup_12_32};
  wire [15:0]   res_hi_hi_hi_32 = {dataGroup_15_32, dataGroup_14_32};
  wire [31:0]   res_hi_hi_32 = {res_hi_hi_hi_32, res_hi_hi_lo_32};
  wire [63:0]   res_hi_32 = {res_hi_hi_32, res_hi_lo_32};
  wire [127:0]  res_60 = {res_hi_32, res_lo_32};
  wire [511:0]  dataGroup_lo_528 = {dataGroup_lo_hi_528, dataGroup_lo_lo_528};
  wire [511:0]  dataGroup_hi_528 = {dataGroup_hi_hi_528, dataGroup_hi_lo_528};
  wire [7:0]    dataGroup_0_33 = dataGroup_lo_528[47:40];
  wire [511:0]  dataGroup_lo_529 = {dataGroup_lo_hi_529, dataGroup_lo_lo_529};
  wire [511:0]  dataGroup_hi_529 = {dataGroup_hi_hi_529, dataGroup_hi_lo_529};
  wire [7:0]    dataGroup_1_33 = dataGroup_lo_529[111:104];
  wire [511:0]  dataGroup_lo_530 = {dataGroup_lo_hi_530, dataGroup_lo_lo_530};
  wire [511:0]  dataGroup_hi_530 = {dataGroup_hi_hi_530, dataGroup_hi_lo_530};
  wire [7:0]    dataGroup_2_33 = dataGroup_lo_530[175:168];
  wire [511:0]  dataGroup_lo_531 = {dataGroup_lo_hi_531, dataGroup_lo_lo_531};
  wire [511:0]  dataGroup_hi_531 = {dataGroup_hi_hi_531, dataGroup_hi_lo_531};
  wire [7:0]    dataGroup_3_33 = dataGroup_lo_531[239:232];
  wire [511:0]  dataGroup_lo_532 = {dataGroup_lo_hi_532, dataGroup_lo_lo_532};
  wire [511:0]  dataGroup_hi_532 = {dataGroup_hi_hi_532, dataGroup_hi_lo_532};
  wire [7:0]    dataGroup_4_33 = dataGroup_lo_532[303:296];
  wire [511:0]  dataGroup_lo_533 = {dataGroup_lo_hi_533, dataGroup_lo_lo_533};
  wire [511:0]  dataGroup_hi_533 = {dataGroup_hi_hi_533, dataGroup_hi_lo_533};
  wire [7:0]    dataGroup_5_33 = dataGroup_lo_533[367:360];
  wire [511:0]  dataGroup_lo_534 = {dataGroup_lo_hi_534, dataGroup_lo_lo_534};
  wire [511:0]  dataGroup_hi_534 = {dataGroup_hi_hi_534, dataGroup_hi_lo_534};
  wire [7:0]    dataGroup_6_33 = dataGroup_lo_534[431:424];
  wire [511:0]  dataGroup_lo_535 = {dataGroup_lo_hi_535, dataGroup_lo_lo_535};
  wire [511:0]  dataGroup_hi_535 = {dataGroup_hi_hi_535, dataGroup_hi_lo_535};
  wire [7:0]    dataGroup_7_33 = dataGroup_lo_535[495:488];
  wire [511:0]  dataGroup_lo_536 = {dataGroup_lo_hi_536, dataGroup_lo_lo_536};
  wire [511:0]  dataGroup_hi_536 = {dataGroup_hi_hi_536, dataGroup_hi_lo_536};
  wire [7:0]    dataGroup_8_33 = dataGroup_hi_536[47:40];
  wire [511:0]  dataGroup_lo_537 = {dataGroup_lo_hi_537, dataGroup_lo_lo_537};
  wire [511:0]  dataGroup_hi_537 = {dataGroup_hi_hi_537, dataGroup_hi_lo_537};
  wire [7:0]    dataGroup_9_33 = dataGroup_hi_537[111:104];
  wire [511:0]  dataGroup_lo_538 = {dataGroup_lo_hi_538, dataGroup_lo_lo_538};
  wire [511:0]  dataGroup_hi_538 = {dataGroup_hi_hi_538, dataGroup_hi_lo_538};
  wire [7:0]    dataGroup_10_33 = dataGroup_hi_538[175:168];
  wire [511:0]  dataGroup_lo_539 = {dataGroup_lo_hi_539, dataGroup_lo_lo_539};
  wire [511:0]  dataGroup_hi_539 = {dataGroup_hi_hi_539, dataGroup_hi_lo_539};
  wire [7:0]    dataGroup_11_33 = dataGroup_hi_539[239:232];
  wire [511:0]  dataGroup_lo_540 = {dataGroup_lo_hi_540, dataGroup_lo_lo_540};
  wire [511:0]  dataGroup_hi_540 = {dataGroup_hi_hi_540, dataGroup_hi_lo_540};
  wire [7:0]    dataGroup_12_33 = dataGroup_hi_540[303:296];
  wire [511:0]  dataGroup_lo_541 = {dataGroup_lo_hi_541, dataGroup_lo_lo_541};
  wire [511:0]  dataGroup_hi_541 = {dataGroup_hi_hi_541, dataGroup_hi_lo_541};
  wire [7:0]    dataGroup_13_33 = dataGroup_hi_541[367:360];
  wire [511:0]  dataGroup_lo_542 = {dataGroup_lo_hi_542, dataGroup_lo_lo_542};
  wire [511:0]  dataGroup_hi_542 = {dataGroup_hi_hi_542, dataGroup_hi_lo_542};
  wire [7:0]    dataGroup_14_33 = dataGroup_hi_542[431:424];
  wire [511:0]  dataGroup_lo_543 = {dataGroup_lo_hi_543, dataGroup_lo_lo_543};
  wire [511:0]  dataGroup_hi_543 = {dataGroup_hi_hi_543, dataGroup_hi_lo_543};
  wire [7:0]    dataGroup_15_33 = dataGroup_hi_543[495:488];
  wire [15:0]   res_lo_lo_lo_33 = {dataGroup_1_33, dataGroup_0_33};
  wire [15:0]   res_lo_lo_hi_33 = {dataGroup_3_33, dataGroup_2_33};
  wire [31:0]   res_lo_lo_33 = {res_lo_lo_hi_33, res_lo_lo_lo_33};
  wire [15:0]   res_lo_hi_lo_33 = {dataGroup_5_33, dataGroup_4_33};
  wire [15:0]   res_lo_hi_hi_33 = {dataGroup_7_33, dataGroup_6_33};
  wire [31:0]   res_lo_hi_33 = {res_lo_hi_hi_33, res_lo_hi_lo_33};
  wire [63:0]   res_lo_33 = {res_lo_hi_33, res_lo_lo_33};
  wire [15:0]   res_hi_lo_lo_33 = {dataGroup_9_33, dataGroup_8_33};
  wire [15:0]   res_hi_lo_hi_33 = {dataGroup_11_33, dataGroup_10_33};
  wire [31:0]   res_hi_lo_33 = {res_hi_lo_hi_33, res_hi_lo_lo_33};
  wire [15:0]   res_hi_hi_lo_33 = {dataGroup_13_33, dataGroup_12_33};
  wire [15:0]   res_hi_hi_hi_33 = {dataGroup_15_33, dataGroup_14_33};
  wire [31:0]   res_hi_hi_33 = {res_hi_hi_hi_33, res_hi_hi_lo_33};
  wire [63:0]   res_hi_33 = {res_hi_hi_33, res_hi_lo_33};
  wire [127:0]  res_61 = {res_hi_33, res_lo_33};
  wire [511:0]  dataGroup_lo_544 = {dataGroup_lo_hi_544, dataGroup_lo_lo_544};
  wire [511:0]  dataGroup_hi_544 = {dataGroup_hi_hi_544, dataGroup_hi_lo_544};
  wire [7:0]    dataGroup_0_34 = dataGroup_lo_544[55:48];
  wire [511:0]  dataGroup_lo_545 = {dataGroup_lo_hi_545, dataGroup_lo_lo_545};
  wire [511:0]  dataGroup_hi_545 = {dataGroup_hi_hi_545, dataGroup_hi_lo_545};
  wire [7:0]    dataGroup_1_34 = dataGroup_lo_545[119:112];
  wire [511:0]  dataGroup_lo_546 = {dataGroup_lo_hi_546, dataGroup_lo_lo_546};
  wire [511:0]  dataGroup_hi_546 = {dataGroup_hi_hi_546, dataGroup_hi_lo_546};
  wire [7:0]    dataGroup_2_34 = dataGroup_lo_546[183:176];
  wire [511:0]  dataGroup_lo_547 = {dataGroup_lo_hi_547, dataGroup_lo_lo_547};
  wire [511:0]  dataGroup_hi_547 = {dataGroup_hi_hi_547, dataGroup_hi_lo_547};
  wire [7:0]    dataGroup_3_34 = dataGroup_lo_547[247:240];
  wire [511:0]  dataGroup_lo_548 = {dataGroup_lo_hi_548, dataGroup_lo_lo_548};
  wire [511:0]  dataGroup_hi_548 = {dataGroup_hi_hi_548, dataGroup_hi_lo_548};
  wire [7:0]    dataGroup_4_34 = dataGroup_lo_548[311:304];
  wire [511:0]  dataGroup_lo_549 = {dataGroup_lo_hi_549, dataGroup_lo_lo_549};
  wire [511:0]  dataGroup_hi_549 = {dataGroup_hi_hi_549, dataGroup_hi_lo_549};
  wire [7:0]    dataGroup_5_34 = dataGroup_lo_549[375:368];
  wire [511:0]  dataGroup_lo_550 = {dataGroup_lo_hi_550, dataGroup_lo_lo_550};
  wire [511:0]  dataGroup_hi_550 = {dataGroup_hi_hi_550, dataGroup_hi_lo_550};
  wire [7:0]    dataGroup_6_34 = dataGroup_lo_550[439:432];
  wire [511:0]  dataGroup_lo_551 = {dataGroup_lo_hi_551, dataGroup_lo_lo_551};
  wire [511:0]  dataGroup_hi_551 = {dataGroup_hi_hi_551, dataGroup_hi_lo_551};
  wire [7:0]    dataGroup_7_34 = dataGroup_lo_551[503:496];
  wire [511:0]  dataGroup_lo_552 = {dataGroup_lo_hi_552, dataGroup_lo_lo_552};
  wire [511:0]  dataGroup_hi_552 = {dataGroup_hi_hi_552, dataGroup_hi_lo_552};
  wire [7:0]    dataGroup_8_34 = dataGroup_hi_552[55:48];
  wire [511:0]  dataGroup_lo_553 = {dataGroup_lo_hi_553, dataGroup_lo_lo_553};
  wire [511:0]  dataGroup_hi_553 = {dataGroup_hi_hi_553, dataGroup_hi_lo_553};
  wire [7:0]    dataGroup_9_34 = dataGroup_hi_553[119:112];
  wire [511:0]  dataGroup_lo_554 = {dataGroup_lo_hi_554, dataGroup_lo_lo_554};
  wire [511:0]  dataGroup_hi_554 = {dataGroup_hi_hi_554, dataGroup_hi_lo_554};
  wire [7:0]    dataGroup_10_34 = dataGroup_hi_554[183:176];
  wire [511:0]  dataGroup_lo_555 = {dataGroup_lo_hi_555, dataGroup_lo_lo_555};
  wire [511:0]  dataGroup_hi_555 = {dataGroup_hi_hi_555, dataGroup_hi_lo_555};
  wire [7:0]    dataGroup_11_34 = dataGroup_hi_555[247:240];
  wire [511:0]  dataGroup_lo_556 = {dataGroup_lo_hi_556, dataGroup_lo_lo_556};
  wire [511:0]  dataGroup_hi_556 = {dataGroup_hi_hi_556, dataGroup_hi_lo_556};
  wire [7:0]    dataGroup_12_34 = dataGroup_hi_556[311:304];
  wire [511:0]  dataGroup_lo_557 = {dataGroup_lo_hi_557, dataGroup_lo_lo_557};
  wire [511:0]  dataGroup_hi_557 = {dataGroup_hi_hi_557, dataGroup_hi_lo_557};
  wire [7:0]    dataGroup_13_34 = dataGroup_hi_557[375:368];
  wire [511:0]  dataGroup_lo_558 = {dataGroup_lo_hi_558, dataGroup_lo_lo_558};
  wire [511:0]  dataGroup_hi_558 = {dataGroup_hi_hi_558, dataGroup_hi_lo_558};
  wire [7:0]    dataGroup_14_34 = dataGroup_hi_558[439:432];
  wire [511:0]  dataGroup_lo_559 = {dataGroup_lo_hi_559, dataGroup_lo_lo_559};
  wire [511:0]  dataGroup_hi_559 = {dataGroup_hi_hi_559, dataGroup_hi_lo_559};
  wire [7:0]    dataGroup_15_34 = dataGroup_hi_559[503:496];
  wire [15:0]   res_lo_lo_lo_34 = {dataGroup_1_34, dataGroup_0_34};
  wire [15:0]   res_lo_lo_hi_34 = {dataGroup_3_34, dataGroup_2_34};
  wire [31:0]   res_lo_lo_34 = {res_lo_lo_hi_34, res_lo_lo_lo_34};
  wire [15:0]   res_lo_hi_lo_34 = {dataGroup_5_34, dataGroup_4_34};
  wire [15:0]   res_lo_hi_hi_34 = {dataGroup_7_34, dataGroup_6_34};
  wire [31:0]   res_lo_hi_34 = {res_lo_hi_hi_34, res_lo_hi_lo_34};
  wire [63:0]   res_lo_34 = {res_lo_hi_34, res_lo_lo_34};
  wire [15:0]   res_hi_lo_lo_34 = {dataGroup_9_34, dataGroup_8_34};
  wire [15:0]   res_hi_lo_hi_34 = {dataGroup_11_34, dataGroup_10_34};
  wire [31:0]   res_hi_lo_34 = {res_hi_lo_hi_34, res_hi_lo_lo_34};
  wire [15:0]   res_hi_hi_lo_34 = {dataGroup_13_34, dataGroup_12_34};
  wire [15:0]   res_hi_hi_hi_34 = {dataGroup_15_34, dataGroup_14_34};
  wire [31:0]   res_hi_hi_34 = {res_hi_hi_hi_34, res_hi_hi_lo_34};
  wire [63:0]   res_hi_34 = {res_hi_hi_34, res_hi_lo_34};
  wire [127:0]  res_62 = {res_hi_34, res_lo_34};
  wire [511:0]  dataGroup_lo_560 = {dataGroup_lo_hi_560, dataGroup_lo_lo_560};
  wire [511:0]  dataGroup_hi_560 = {dataGroup_hi_hi_560, dataGroup_hi_lo_560};
  wire [7:0]    dataGroup_0_35 = dataGroup_lo_560[63:56];
  wire [511:0]  dataGroup_lo_561 = {dataGroup_lo_hi_561, dataGroup_lo_lo_561};
  wire [511:0]  dataGroup_hi_561 = {dataGroup_hi_hi_561, dataGroup_hi_lo_561};
  wire [7:0]    dataGroup_1_35 = dataGroup_lo_561[127:120];
  wire [511:0]  dataGroup_lo_562 = {dataGroup_lo_hi_562, dataGroup_lo_lo_562};
  wire [511:0]  dataGroup_hi_562 = {dataGroup_hi_hi_562, dataGroup_hi_lo_562};
  wire [7:0]    dataGroup_2_35 = dataGroup_lo_562[191:184];
  wire [511:0]  dataGroup_lo_563 = {dataGroup_lo_hi_563, dataGroup_lo_lo_563};
  wire [511:0]  dataGroup_hi_563 = {dataGroup_hi_hi_563, dataGroup_hi_lo_563};
  wire [7:0]    dataGroup_3_35 = dataGroup_lo_563[255:248];
  wire [511:0]  dataGroup_lo_564 = {dataGroup_lo_hi_564, dataGroup_lo_lo_564};
  wire [511:0]  dataGroup_hi_564 = {dataGroup_hi_hi_564, dataGroup_hi_lo_564};
  wire [7:0]    dataGroup_4_35 = dataGroup_lo_564[319:312];
  wire [511:0]  dataGroup_lo_565 = {dataGroup_lo_hi_565, dataGroup_lo_lo_565};
  wire [511:0]  dataGroup_hi_565 = {dataGroup_hi_hi_565, dataGroup_hi_lo_565};
  wire [7:0]    dataGroup_5_35 = dataGroup_lo_565[383:376];
  wire [511:0]  dataGroup_lo_566 = {dataGroup_lo_hi_566, dataGroup_lo_lo_566};
  wire [511:0]  dataGroup_hi_566 = {dataGroup_hi_hi_566, dataGroup_hi_lo_566};
  wire [7:0]    dataGroup_6_35 = dataGroup_lo_566[447:440];
  wire [511:0]  dataGroup_lo_567 = {dataGroup_lo_hi_567, dataGroup_lo_lo_567};
  wire [511:0]  dataGroup_hi_567 = {dataGroup_hi_hi_567, dataGroup_hi_lo_567};
  wire [7:0]    dataGroup_7_35 = dataGroup_lo_567[511:504];
  wire [511:0]  dataGroup_lo_568 = {dataGroup_lo_hi_568, dataGroup_lo_lo_568};
  wire [511:0]  dataGroup_hi_568 = {dataGroup_hi_hi_568, dataGroup_hi_lo_568};
  wire [7:0]    dataGroup_8_35 = dataGroup_hi_568[63:56];
  wire [511:0]  dataGroup_lo_569 = {dataGroup_lo_hi_569, dataGroup_lo_lo_569};
  wire [511:0]  dataGroup_hi_569 = {dataGroup_hi_hi_569, dataGroup_hi_lo_569};
  wire [7:0]    dataGroup_9_35 = dataGroup_hi_569[127:120];
  wire [511:0]  dataGroup_lo_570 = {dataGroup_lo_hi_570, dataGroup_lo_lo_570};
  wire [511:0]  dataGroup_hi_570 = {dataGroup_hi_hi_570, dataGroup_hi_lo_570};
  wire [7:0]    dataGroup_10_35 = dataGroup_hi_570[191:184];
  wire [511:0]  dataGroup_lo_571 = {dataGroup_lo_hi_571, dataGroup_lo_lo_571};
  wire [511:0]  dataGroup_hi_571 = {dataGroup_hi_hi_571, dataGroup_hi_lo_571};
  wire [7:0]    dataGroup_11_35 = dataGroup_hi_571[255:248];
  wire [511:0]  dataGroup_lo_572 = {dataGroup_lo_hi_572, dataGroup_lo_lo_572};
  wire [511:0]  dataGroup_hi_572 = {dataGroup_hi_hi_572, dataGroup_hi_lo_572};
  wire [7:0]    dataGroup_12_35 = dataGroup_hi_572[319:312];
  wire [511:0]  dataGroup_lo_573 = {dataGroup_lo_hi_573, dataGroup_lo_lo_573};
  wire [511:0]  dataGroup_hi_573 = {dataGroup_hi_hi_573, dataGroup_hi_lo_573};
  wire [7:0]    dataGroup_13_35 = dataGroup_hi_573[383:376];
  wire [511:0]  dataGroup_lo_574 = {dataGroup_lo_hi_574, dataGroup_lo_lo_574};
  wire [511:0]  dataGroup_hi_574 = {dataGroup_hi_hi_574, dataGroup_hi_lo_574};
  wire [7:0]    dataGroup_14_35 = dataGroup_hi_574[447:440];
  wire [511:0]  dataGroup_lo_575 = {dataGroup_lo_hi_575, dataGroup_lo_lo_575};
  wire [511:0]  dataGroup_hi_575 = {dataGroup_hi_hi_575, dataGroup_hi_lo_575};
  wire [7:0]    dataGroup_15_35 = dataGroup_hi_575[511:504];
  wire [15:0]   res_lo_lo_lo_35 = {dataGroup_1_35, dataGroup_0_35};
  wire [15:0]   res_lo_lo_hi_35 = {dataGroup_3_35, dataGroup_2_35};
  wire [31:0]   res_lo_lo_35 = {res_lo_lo_hi_35, res_lo_lo_lo_35};
  wire [15:0]   res_lo_hi_lo_35 = {dataGroup_5_35, dataGroup_4_35};
  wire [15:0]   res_lo_hi_hi_35 = {dataGroup_7_35, dataGroup_6_35};
  wire [31:0]   res_lo_hi_35 = {res_lo_hi_hi_35, res_lo_hi_lo_35};
  wire [63:0]   res_lo_35 = {res_lo_hi_35, res_lo_lo_35};
  wire [15:0]   res_hi_lo_lo_35 = {dataGroup_9_35, dataGroup_8_35};
  wire [15:0]   res_hi_lo_hi_35 = {dataGroup_11_35, dataGroup_10_35};
  wire [31:0]   res_hi_lo_35 = {res_hi_lo_hi_35, res_hi_lo_lo_35};
  wire [15:0]   res_hi_hi_lo_35 = {dataGroup_13_35, dataGroup_12_35};
  wire [15:0]   res_hi_hi_hi_35 = {dataGroup_15_35, dataGroup_14_35};
  wire [31:0]   res_hi_hi_35 = {res_hi_hi_hi_35, res_hi_hi_lo_35};
  wire [63:0]   res_hi_35 = {res_hi_hi_35, res_hi_lo_35};
  wire [127:0]  res_63 = {res_hi_35, res_lo_35};
  wire [255:0]  lo_lo_7 = {res_57, res_56};
  wire [255:0]  lo_hi_7 = {res_59, res_58};
  wire [511:0]  lo_7 = {lo_hi_7, lo_lo_7};
  wire [255:0]  hi_lo_7 = {res_61, res_60};
  wire [255:0]  hi_hi_7 = {res_63, res_62};
  wire [511:0]  hi_7 = {hi_hi_7, hi_lo_7};
  wire [1023:0] regroupLoadData_0_7 = {hi_7, lo_7};
  wire [511:0]  dataGroup_lo_576 = {dataGroup_lo_hi_576, dataGroup_lo_lo_576};
  wire [511:0]  dataGroup_hi_576 = {dataGroup_hi_hi_576, dataGroup_hi_lo_576};
  wire [15:0]   dataGroup_0_36 = dataGroup_lo_576[15:0];
  wire [511:0]  dataGroup_lo_577 = {dataGroup_lo_hi_577, dataGroup_lo_lo_577};
  wire [511:0]  dataGroup_hi_577 = {dataGroup_hi_hi_577, dataGroup_hi_lo_577};
  wire [15:0]   dataGroup_1_36 = dataGroup_lo_577[31:16];
  wire [511:0]  dataGroup_lo_578 = {dataGroup_lo_hi_578, dataGroup_lo_lo_578};
  wire [511:0]  dataGroup_hi_578 = {dataGroup_hi_hi_578, dataGroup_hi_lo_578};
  wire [15:0]   dataGroup_2_36 = dataGroup_lo_578[47:32];
  wire [511:0]  dataGroup_lo_579 = {dataGroup_lo_hi_579, dataGroup_lo_lo_579};
  wire [511:0]  dataGroup_hi_579 = {dataGroup_hi_hi_579, dataGroup_hi_lo_579};
  wire [15:0]   dataGroup_3_36 = dataGroup_lo_579[63:48];
  wire [511:0]  dataGroup_lo_580 = {dataGroup_lo_hi_580, dataGroup_lo_lo_580};
  wire [511:0]  dataGroup_hi_580 = {dataGroup_hi_hi_580, dataGroup_hi_lo_580};
  wire [15:0]   dataGroup_4_36 = dataGroup_lo_580[79:64];
  wire [511:0]  dataGroup_lo_581 = {dataGroup_lo_hi_581, dataGroup_lo_lo_581};
  wire [511:0]  dataGroup_hi_581 = {dataGroup_hi_hi_581, dataGroup_hi_lo_581};
  wire [15:0]   dataGroup_5_36 = dataGroup_lo_581[95:80];
  wire [511:0]  dataGroup_lo_582 = {dataGroup_lo_hi_582, dataGroup_lo_lo_582};
  wire [511:0]  dataGroup_hi_582 = {dataGroup_hi_hi_582, dataGroup_hi_lo_582};
  wire [15:0]   dataGroup_6_36 = dataGroup_lo_582[111:96];
  wire [511:0]  dataGroup_lo_583 = {dataGroup_lo_hi_583, dataGroup_lo_lo_583};
  wire [511:0]  dataGroup_hi_583 = {dataGroup_hi_hi_583, dataGroup_hi_lo_583};
  wire [15:0]   dataGroup_7_36 = dataGroup_lo_583[127:112];
  wire [31:0]   res_lo_lo_36 = {dataGroup_1_36, dataGroup_0_36};
  wire [31:0]   res_lo_hi_36 = {dataGroup_3_36, dataGroup_2_36};
  wire [63:0]   res_lo_36 = {res_lo_hi_36, res_lo_lo_36};
  wire [31:0]   res_hi_lo_36 = {dataGroup_5_36, dataGroup_4_36};
  wire [31:0]   res_hi_hi_36 = {dataGroup_7_36, dataGroup_6_36};
  wire [63:0]   res_hi_36 = {res_hi_hi_36, res_hi_lo_36};
  wire [127:0]  res_64 = {res_hi_36, res_lo_36};
  wire [255:0]  lo_lo_8 = {128'h0, res_64};
  wire [511:0]  lo_8 = {256'h0, lo_lo_8};
  wire [1023:0] regroupLoadData_1_0 = {512'h0, lo_8};
  wire [511:0]  dataGroup_lo_584 = {dataGroup_lo_hi_584, dataGroup_lo_lo_584};
  wire [511:0]  dataGroup_hi_584 = {dataGroup_hi_hi_584, dataGroup_hi_lo_584};
  wire [15:0]   dataGroup_0_37 = dataGroup_lo_584[15:0];
  wire [511:0]  dataGroup_lo_585 = {dataGroup_lo_hi_585, dataGroup_lo_lo_585};
  wire [511:0]  dataGroup_hi_585 = {dataGroup_hi_hi_585, dataGroup_hi_lo_585};
  wire [15:0]   dataGroup_1_37 = dataGroup_lo_585[47:32];
  wire [511:0]  dataGroup_lo_586 = {dataGroup_lo_hi_586, dataGroup_lo_lo_586};
  wire [511:0]  dataGroup_hi_586 = {dataGroup_hi_hi_586, dataGroup_hi_lo_586};
  wire [15:0]   dataGroup_2_37 = dataGroup_lo_586[79:64];
  wire [511:0]  dataGroup_lo_587 = {dataGroup_lo_hi_587, dataGroup_lo_lo_587};
  wire [511:0]  dataGroup_hi_587 = {dataGroup_hi_hi_587, dataGroup_hi_lo_587};
  wire [15:0]   dataGroup_3_37 = dataGroup_lo_587[111:96];
  wire [511:0]  dataGroup_lo_588 = {dataGroup_lo_hi_588, dataGroup_lo_lo_588};
  wire [511:0]  dataGroup_hi_588 = {dataGroup_hi_hi_588, dataGroup_hi_lo_588};
  wire [15:0]   dataGroup_4_37 = dataGroup_lo_588[143:128];
  wire [511:0]  dataGroup_lo_589 = {dataGroup_lo_hi_589, dataGroup_lo_lo_589};
  wire [511:0]  dataGroup_hi_589 = {dataGroup_hi_hi_589, dataGroup_hi_lo_589};
  wire [15:0]   dataGroup_5_37 = dataGroup_lo_589[175:160];
  wire [511:0]  dataGroup_lo_590 = {dataGroup_lo_hi_590, dataGroup_lo_lo_590};
  wire [511:0]  dataGroup_hi_590 = {dataGroup_hi_hi_590, dataGroup_hi_lo_590};
  wire [15:0]   dataGroup_6_37 = dataGroup_lo_590[207:192];
  wire [511:0]  dataGroup_lo_591 = {dataGroup_lo_hi_591, dataGroup_lo_lo_591};
  wire [511:0]  dataGroup_hi_591 = {dataGroup_hi_hi_591, dataGroup_hi_lo_591};
  wire [15:0]   dataGroup_7_37 = dataGroup_lo_591[239:224];
  wire [31:0]   res_lo_lo_37 = {dataGroup_1_37, dataGroup_0_37};
  wire [31:0]   res_lo_hi_37 = {dataGroup_3_37, dataGroup_2_37};
  wire [63:0]   res_lo_37 = {res_lo_hi_37, res_lo_lo_37};
  wire [31:0]   res_hi_lo_37 = {dataGroup_5_37, dataGroup_4_37};
  wire [31:0]   res_hi_hi_37 = {dataGroup_7_37, dataGroup_6_37};
  wire [63:0]   res_hi_37 = {res_hi_hi_37, res_hi_lo_37};
  wire [127:0]  res_72 = {res_hi_37, res_lo_37};
  wire [511:0]  dataGroup_lo_592 = {dataGroup_lo_hi_592, dataGroup_lo_lo_592};
  wire [511:0]  dataGroup_hi_592 = {dataGroup_hi_hi_592, dataGroup_hi_lo_592};
  wire [15:0]   dataGroup_0_38 = dataGroup_lo_592[31:16];
  wire [511:0]  dataGroup_lo_593 = {dataGroup_lo_hi_593, dataGroup_lo_lo_593};
  wire [511:0]  dataGroup_hi_593 = {dataGroup_hi_hi_593, dataGroup_hi_lo_593};
  wire [15:0]   dataGroup_1_38 = dataGroup_lo_593[63:48];
  wire [511:0]  dataGroup_lo_594 = {dataGroup_lo_hi_594, dataGroup_lo_lo_594};
  wire [511:0]  dataGroup_hi_594 = {dataGroup_hi_hi_594, dataGroup_hi_lo_594};
  wire [15:0]   dataGroup_2_38 = dataGroup_lo_594[95:80];
  wire [511:0]  dataGroup_lo_595 = {dataGroup_lo_hi_595, dataGroup_lo_lo_595};
  wire [511:0]  dataGroup_hi_595 = {dataGroup_hi_hi_595, dataGroup_hi_lo_595};
  wire [15:0]   dataGroup_3_38 = dataGroup_lo_595[127:112];
  wire [511:0]  dataGroup_lo_596 = {dataGroup_lo_hi_596, dataGroup_lo_lo_596};
  wire [511:0]  dataGroup_hi_596 = {dataGroup_hi_hi_596, dataGroup_hi_lo_596};
  wire [15:0]   dataGroup_4_38 = dataGroup_lo_596[159:144];
  wire [511:0]  dataGroup_lo_597 = {dataGroup_lo_hi_597, dataGroup_lo_lo_597};
  wire [511:0]  dataGroup_hi_597 = {dataGroup_hi_hi_597, dataGroup_hi_lo_597};
  wire [15:0]   dataGroup_5_38 = dataGroup_lo_597[191:176];
  wire [511:0]  dataGroup_lo_598 = {dataGroup_lo_hi_598, dataGroup_lo_lo_598};
  wire [511:0]  dataGroup_hi_598 = {dataGroup_hi_hi_598, dataGroup_hi_lo_598};
  wire [15:0]   dataGroup_6_38 = dataGroup_lo_598[223:208];
  wire [511:0]  dataGroup_lo_599 = {dataGroup_lo_hi_599, dataGroup_lo_lo_599};
  wire [511:0]  dataGroup_hi_599 = {dataGroup_hi_hi_599, dataGroup_hi_lo_599};
  wire [15:0]   dataGroup_7_38 = dataGroup_lo_599[255:240];
  wire [31:0]   res_lo_lo_38 = {dataGroup_1_38, dataGroup_0_38};
  wire [31:0]   res_lo_hi_38 = {dataGroup_3_38, dataGroup_2_38};
  wire [63:0]   res_lo_38 = {res_lo_hi_38, res_lo_lo_38};
  wire [31:0]   res_hi_lo_38 = {dataGroup_5_38, dataGroup_4_38};
  wire [31:0]   res_hi_hi_38 = {dataGroup_7_38, dataGroup_6_38};
  wire [63:0]   res_hi_38 = {res_hi_hi_38, res_hi_lo_38};
  wire [127:0]  res_73 = {res_hi_38, res_lo_38};
  wire [255:0]  lo_lo_9 = {res_73, res_72};
  wire [511:0]  lo_9 = {256'h0, lo_lo_9};
  wire [1023:0] regroupLoadData_1_1 = {512'h0, lo_9};
  wire [511:0]  dataGroup_lo_600 = {dataGroup_lo_hi_600, dataGroup_lo_lo_600};
  wire [511:0]  dataGroup_hi_600 = {dataGroup_hi_hi_600, dataGroup_hi_lo_600};
  wire [15:0]   dataGroup_0_39 = dataGroup_lo_600[15:0];
  wire [511:0]  dataGroup_lo_601 = {dataGroup_lo_hi_601, dataGroup_lo_lo_601};
  wire [511:0]  dataGroup_hi_601 = {dataGroup_hi_hi_601, dataGroup_hi_lo_601};
  wire [15:0]   dataGroup_1_39 = dataGroup_lo_601[63:48];
  wire [511:0]  dataGroup_lo_602 = {dataGroup_lo_hi_602, dataGroup_lo_lo_602};
  wire [511:0]  dataGroup_hi_602 = {dataGroup_hi_hi_602, dataGroup_hi_lo_602};
  wire [15:0]   dataGroup_2_39 = dataGroup_lo_602[111:96];
  wire [511:0]  dataGroup_lo_603 = {dataGroup_lo_hi_603, dataGroup_lo_lo_603};
  wire [511:0]  dataGroup_hi_603 = {dataGroup_hi_hi_603, dataGroup_hi_lo_603};
  wire [15:0]   dataGroup_3_39 = dataGroup_lo_603[159:144];
  wire [511:0]  dataGroup_lo_604 = {dataGroup_lo_hi_604, dataGroup_lo_lo_604};
  wire [511:0]  dataGroup_hi_604 = {dataGroup_hi_hi_604, dataGroup_hi_lo_604};
  wire [15:0]   dataGroup_4_39 = dataGroup_lo_604[207:192];
  wire [511:0]  dataGroup_lo_605 = {dataGroup_lo_hi_605, dataGroup_lo_lo_605};
  wire [511:0]  dataGroup_hi_605 = {dataGroup_hi_hi_605, dataGroup_hi_lo_605};
  wire [15:0]   dataGroup_5_39 = dataGroup_lo_605[255:240];
  wire [511:0]  dataGroup_lo_606 = {dataGroup_lo_hi_606, dataGroup_lo_lo_606};
  wire [511:0]  dataGroup_hi_606 = {dataGroup_hi_hi_606, dataGroup_hi_lo_606};
  wire [15:0]   dataGroup_6_39 = dataGroup_lo_606[303:288];
  wire [511:0]  dataGroup_lo_607 = {dataGroup_lo_hi_607, dataGroup_lo_lo_607};
  wire [511:0]  dataGroup_hi_607 = {dataGroup_hi_hi_607, dataGroup_hi_lo_607};
  wire [15:0]   dataGroup_7_39 = dataGroup_lo_607[351:336];
  wire [31:0]   res_lo_lo_39 = {dataGroup_1_39, dataGroup_0_39};
  wire [31:0]   res_lo_hi_39 = {dataGroup_3_39, dataGroup_2_39};
  wire [63:0]   res_lo_39 = {res_lo_hi_39, res_lo_lo_39};
  wire [31:0]   res_hi_lo_39 = {dataGroup_5_39, dataGroup_4_39};
  wire [31:0]   res_hi_hi_39 = {dataGroup_7_39, dataGroup_6_39};
  wire [63:0]   res_hi_39 = {res_hi_hi_39, res_hi_lo_39};
  wire [127:0]  res_80 = {res_hi_39, res_lo_39};
  wire [511:0]  dataGroup_lo_608 = {dataGroup_lo_hi_608, dataGroup_lo_lo_608};
  wire [511:0]  dataGroup_hi_608 = {dataGroup_hi_hi_608, dataGroup_hi_lo_608};
  wire [15:0]   dataGroup_0_40 = dataGroup_lo_608[31:16];
  wire [511:0]  dataGroup_lo_609 = {dataGroup_lo_hi_609, dataGroup_lo_lo_609};
  wire [511:0]  dataGroup_hi_609 = {dataGroup_hi_hi_609, dataGroup_hi_lo_609};
  wire [15:0]   dataGroup_1_40 = dataGroup_lo_609[79:64];
  wire [511:0]  dataGroup_lo_610 = {dataGroup_lo_hi_610, dataGroup_lo_lo_610};
  wire [511:0]  dataGroup_hi_610 = {dataGroup_hi_hi_610, dataGroup_hi_lo_610};
  wire [15:0]   dataGroup_2_40 = dataGroup_lo_610[127:112];
  wire [511:0]  dataGroup_lo_611 = {dataGroup_lo_hi_611, dataGroup_lo_lo_611};
  wire [511:0]  dataGroup_hi_611 = {dataGroup_hi_hi_611, dataGroup_hi_lo_611};
  wire [15:0]   dataGroup_3_40 = dataGroup_lo_611[175:160];
  wire [511:0]  dataGroup_lo_612 = {dataGroup_lo_hi_612, dataGroup_lo_lo_612};
  wire [511:0]  dataGroup_hi_612 = {dataGroup_hi_hi_612, dataGroup_hi_lo_612};
  wire [15:0]   dataGroup_4_40 = dataGroup_lo_612[223:208];
  wire [511:0]  dataGroup_lo_613 = {dataGroup_lo_hi_613, dataGroup_lo_lo_613};
  wire [511:0]  dataGroup_hi_613 = {dataGroup_hi_hi_613, dataGroup_hi_lo_613};
  wire [15:0]   dataGroup_5_40 = dataGroup_lo_613[271:256];
  wire [511:0]  dataGroup_lo_614 = {dataGroup_lo_hi_614, dataGroup_lo_lo_614};
  wire [511:0]  dataGroup_hi_614 = {dataGroup_hi_hi_614, dataGroup_hi_lo_614};
  wire [15:0]   dataGroup_6_40 = dataGroup_lo_614[319:304];
  wire [511:0]  dataGroup_lo_615 = {dataGroup_lo_hi_615, dataGroup_lo_lo_615};
  wire [511:0]  dataGroup_hi_615 = {dataGroup_hi_hi_615, dataGroup_hi_lo_615};
  wire [15:0]   dataGroup_7_40 = dataGroup_lo_615[367:352];
  wire [31:0]   res_lo_lo_40 = {dataGroup_1_40, dataGroup_0_40};
  wire [31:0]   res_lo_hi_40 = {dataGroup_3_40, dataGroup_2_40};
  wire [63:0]   res_lo_40 = {res_lo_hi_40, res_lo_lo_40};
  wire [31:0]   res_hi_lo_40 = {dataGroup_5_40, dataGroup_4_40};
  wire [31:0]   res_hi_hi_40 = {dataGroup_7_40, dataGroup_6_40};
  wire [63:0]   res_hi_40 = {res_hi_hi_40, res_hi_lo_40};
  wire [127:0]  res_81 = {res_hi_40, res_lo_40};
  wire [511:0]  dataGroup_lo_616 = {dataGroup_lo_hi_616, dataGroup_lo_lo_616};
  wire [511:0]  dataGroup_hi_616 = {dataGroup_hi_hi_616, dataGroup_hi_lo_616};
  wire [15:0]   dataGroup_0_41 = dataGroup_lo_616[47:32];
  wire [511:0]  dataGroup_lo_617 = {dataGroup_lo_hi_617, dataGroup_lo_lo_617};
  wire [511:0]  dataGroup_hi_617 = {dataGroup_hi_hi_617, dataGroup_hi_lo_617};
  wire [15:0]   dataGroup_1_41 = dataGroup_lo_617[95:80];
  wire [511:0]  dataGroup_lo_618 = {dataGroup_lo_hi_618, dataGroup_lo_lo_618};
  wire [511:0]  dataGroup_hi_618 = {dataGroup_hi_hi_618, dataGroup_hi_lo_618};
  wire [15:0]   dataGroup_2_41 = dataGroup_lo_618[143:128];
  wire [511:0]  dataGroup_lo_619 = {dataGroup_lo_hi_619, dataGroup_lo_lo_619};
  wire [511:0]  dataGroup_hi_619 = {dataGroup_hi_hi_619, dataGroup_hi_lo_619};
  wire [15:0]   dataGroup_3_41 = dataGroup_lo_619[191:176];
  wire [511:0]  dataGroup_lo_620 = {dataGroup_lo_hi_620, dataGroup_lo_lo_620};
  wire [511:0]  dataGroup_hi_620 = {dataGroup_hi_hi_620, dataGroup_hi_lo_620};
  wire [15:0]   dataGroup_4_41 = dataGroup_lo_620[239:224];
  wire [511:0]  dataGroup_lo_621 = {dataGroup_lo_hi_621, dataGroup_lo_lo_621};
  wire [511:0]  dataGroup_hi_621 = {dataGroup_hi_hi_621, dataGroup_hi_lo_621};
  wire [15:0]   dataGroup_5_41 = dataGroup_lo_621[287:272];
  wire [511:0]  dataGroup_lo_622 = {dataGroup_lo_hi_622, dataGroup_lo_lo_622};
  wire [511:0]  dataGroup_hi_622 = {dataGroup_hi_hi_622, dataGroup_hi_lo_622};
  wire [15:0]   dataGroup_6_41 = dataGroup_lo_622[335:320];
  wire [511:0]  dataGroup_lo_623 = {dataGroup_lo_hi_623, dataGroup_lo_lo_623};
  wire [511:0]  dataGroup_hi_623 = {dataGroup_hi_hi_623, dataGroup_hi_lo_623};
  wire [15:0]   dataGroup_7_41 = dataGroup_lo_623[383:368];
  wire [31:0]   res_lo_lo_41 = {dataGroup_1_41, dataGroup_0_41};
  wire [31:0]   res_lo_hi_41 = {dataGroup_3_41, dataGroup_2_41};
  wire [63:0]   res_lo_41 = {res_lo_hi_41, res_lo_lo_41};
  wire [31:0]   res_hi_lo_41 = {dataGroup_5_41, dataGroup_4_41};
  wire [31:0]   res_hi_hi_41 = {dataGroup_7_41, dataGroup_6_41};
  wire [63:0]   res_hi_41 = {res_hi_hi_41, res_hi_lo_41};
  wire [127:0]  res_82 = {res_hi_41, res_lo_41};
  wire [255:0]  lo_lo_10 = {res_81, res_80};
  wire [255:0]  lo_hi_10 = {128'h0, res_82};
  wire [511:0]  lo_10 = {lo_hi_10, lo_lo_10};
  wire [1023:0] regroupLoadData_1_2 = {512'h0, lo_10};
  wire [511:0]  dataGroup_lo_624 = {dataGroup_lo_hi_624, dataGroup_lo_lo_624};
  wire [511:0]  dataGroup_hi_624 = {dataGroup_hi_hi_624, dataGroup_hi_lo_624};
  wire [15:0]   dataGroup_0_42 = dataGroup_lo_624[15:0];
  wire [511:0]  dataGroup_lo_625 = {dataGroup_lo_hi_625, dataGroup_lo_lo_625};
  wire [511:0]  dataGroup_hi_625 = {dataGroup_hi_hi_625, dataGroup_hi_lo_625};
  wire [15:0]   dataGroup_1_42 = dataGroup_lo_625[79:64];
  wire [511:0]  dataGroup_lo_626 = {dataGroup_lo_hi_626, dataGroup_lo_lo_626};
  wire [511:0]  dataGroup_hi_626 = {dataGroup_hi_hi_626, dataGroup_hi_lo_626};
  wire [15:0]   dataGroup_2_42 = dataGroup_lo_626[143:128];
  wire [511:0]  dataGroup_lo_627 = {dataGroup_lo_hi_627, dataGroup_lo_lo_627};
  wire [511:0]  dataGroup_hi_627 = {dataGroup_hi_hi_627, dataGroup_hi_lo_627};
  wire [15:0]   dataGroup_3_42 = dataGroup_lo_627[207:192];
  wire [511:0]  dataGroup_lo_628 = {dataGroup_lo_hi_628, dataGroup_lo_lo_628};
  wire [511:0]  dataGroup_hi_628 = {dataGroup_hi_hi_628, dataGroup_hi_lo_628};
  wire [15:0]   dataGroup_4_42 = dataGroup_lo_628[271:256];
  wire [511:0]  dataGroup_lo_629 = {dataGroup_lo_hi_629, dataGroup_lo_lo_629};
  wire [511:0]  dataGroup_hi_629 = {dataGroup_hi_hi_629, dataGroup_hi_lo_629};
  wire [15:0]   dataGroup_5_42 = dataGroup_lo_629[335:320];
  wire [511:0]  dataGroup_lo_630 = {dataGroup_lo_hi_630, dataGroup_lo_lo_630};
  wire [511:0]  dataGroup_hi_630 = {dataGroup_hi_hi_630, dataGroup_hi_lo_630};
  wire [15:0]   dataGroup_6_42 = dataGroup_lo_630[399:384];
  wire [511:0]  dataGroup_lo_631 = {dataGroup_lo_hi_631, dataGroup_lo_lo_631};
  wire [511:0]  dataGroup_hi_631 = {dataGroup_hi_hi_631, dataGroup_hi_lo_631};
  wire [15:0]   dataGroup_7_42 = dataGroup_lo_631[463:448];
  wire [31:0]   res_lo_lo_42 = {dataGroup_1_42, dataGroup_0_42};
  wire [31:0]   res_lo_hi_42 = {dataGroup_3_42, dataGroup_2_42};
  wire [63:0]   res_lo_42 = {res_lo_hi_42, res_lo_lo_42};
  wire [31:0]   res_hi_lo_42 = {dataGroup_5_42, dataGroup_4_42};
  wire [31:0]   res_hi_hi_42 = {dataGroup_7_42, dataGroup_6_42};
  wire [63:0]   res_hi_42 = {res_hi_hi_42, res_hi_lo_42};
  wire [127:0]  res_88 = {res_hi_42, res_lo_42};
  wire [511:0]  dataGroup_lo_632 = {dataGroup_lo_hi_632, dataGroup_lo_lo_632};
  wire [511:0]  dataGroup_hi_632 = {dataGroup_hi_hi_632, dataGroup_hi_lo_632};
  wire [15:0]   dataGroup_0_43 = dataGroup_lo_632[31:16];
  wire [511:0]  dataGroup_lo_633 = {dataGroup_lo_hi_633, dataGroup_lo_lo_633};
  wire [511:0]  dataGroup_hi_633 = {dataGroup_hi_hi_633, dataGroup_hi_lo_633};
  wire [15:0]   dataGroup_1_43 = dataGroup_lo_633[95:80];
  wire [511:0]  dataGroup_lo_634 = {dataGroup_lo_hi_634, dataGroup_lo_lo_634};
  wire [511:0]  dataGroup_hi_634 = {dataGroup_hi_hi_634, dataGroup_hi_lo_634};
  wire [15:0]   dataGroup_2_43 = dataGroup_lo_634[159:144];
  wire [511:0]  dataGroup_lo_635 = {dataGroup_lo_hi_635, dataGroup_lo_lo_635};
  wire [511:0]  dataGroup_hi_635 = {dataGroup_hi_hi_635, dataGroup_hi_lo_635};
  wire [15:0]   dataGroup_3_43 = dataGroup_lo_635[223:208];
  wire [511:0]  dataGroup_lo_636 = {dataGroup_lo_hi_636, dataGroup_lo_lo_636};
  wire [511:0]  dataGroup_hi_636 = {dataGroup_hi_hi_636, dataGroup_hi_lo_636};
  wire [15:0]   dataGroup_4_43 = dataGroup_lo_636[287:272];
  wire [511:0]  dataGroup_lo_637 = {dataGroup_lo_hi_637, dataGroup_lo_lo_637};
  wire [511:0]  dataGroup_hi_637 = {dataGroup_hi_hi_637, dataGroup_hi_lo_637};
  wire [15:0]   dataGroup_5_43 = dataGroup_lo_637[351:336];
  wire [511:0]  dataGroup_lo_638 = {dataGroup_lo_hi_638, dataGroup_lo_lo_638};
  wire [511:0]  dataGroup_hi_638 = {dataGroup_hi_hi_638, dataGroup_hi_lo_638};
  wire [15:0]   dataGroup_6_43 = dataGroup_lo_638[415:400];
  wire [511:0]  dataGroup_lo_639 = {dataGroup_lo_hi_639, dataGroup_lo_lo_639};
  wire [511:0]  dataGroup_hi_639 = {dataGroup_hi_hi_639, dataGroup_hi_lo_639};
  wire [15:0]   dataGroup_7_43 = dataGroup_lo_639[479:464];
  wire [31:0]   res_lo_lo_43 = {dataGroup_1_43, dataGroup_0_43};
  wire [31:0]   res_lo_hi_43 = {dataGroup_3_43, dataGroup_2_43};
  wire [63:0]   res_lo_43 = {res_lo_hi_43, res_lo_lo_43};
  wire [31:0]   res_hi_lo_43 = {dataGroup_5_43, dataGroup_4_43};
  wire [31:0]   res_hi_hi_43 = {dataGroup_7_43, dataGroup_6_43};
  wire [63:0]   res_hi_43 = {res_hi_hi_43, res_hi_lo_43};
  wire [127:0]  res_89 = {res_hi_43, res_lo_43};
  wire [511:0]  dataGroup_lo_640 = {dataGroup_lo_hi_640, dataGroup_lo_lo_640};
  wire [511:0]  dataGroup_hi_640 = {dataGroup_hi_hi_640, dataGroup_hi_lo_640};
  wire [15:0]   dataGroup_0_44 = dataGroup_lo_640[47:32];
  wire [511:0]  dataGroup_lo_641 = {dataGroup_lo_hi_641, dataGroup_lo_lo_641};
  wire [511:0]  dataGroup_hi_641 = {dataGroup_hi_hi_641, dataGroup_hi_lo_641};
  wire [15:0]   dataGroup_1_44 = dataGroup_lo_641[111:96];
  wire [511:0]  dataGroup_lo_642 = {dataGroup_lo_hi_642, dataGroup_lo_lo_642};
  wire [511:0]  dataGroup_hi_642 = {dataGroup_hi_hi_642, dataGroup_hi_lo_642};
  wire [15:0]   dataGroup_2_44 = dataGroup_lo_642[175:160];
  wire [511:0]  dataGroup_lo_643 = {dataGroup_lo_hi_643, dataGroup_lo_lo_643};
  wire [511:0]  dataGroup_hi_643 = {dataGroup_hi_hi_643, dataGroup_hi_lo_643};
  wire [15:0]   dataGroup_3_44 = dataGroup_lo_643[239:224];
  wire [511:0]  dataGroup_lo_644 = {dataGroup_lo_hi_644, dataGroup_lo_lo_644};
  wire [511:0]  dataGroup_hi_644 = {dataGroup_hi_hi_644, dataGroup_hi_lo_644};
  wire [15:0]   dataGroup_4_44 = dataGroup_lo_644[303:288];
  wire [511:0]  dataGroup_lo_645 = {dataGroup_lo_hi_645, dataGroup_lo_lo_645};
  wire [511:0]  dataGroup_hi_645 = {dataGroup_hi_hi_645, dataGroup_hi_lo_645};
  wire [15:0]   dataGroup_5_44 = dataGroup_lo_645[367:352];
  wire [511:0]  dataGroup_lo_646 = {dataGroup_lo_hi_646, dataGroup_lo_lo_646};
  wire [511:0]  dataGroup_hi_646 = {dataGroup_hi_hi_646, dataGroup_hi_lo_646};
  wire [15:0]   dataGroup_6_44 = dataGroup_lo_646[431:416];
  wire [511:0]  dataGroup_lo_647 = {dataGroup_lo_hi_647, dataGroup_lo_lo_647};
  wire [511:0]  dataGroup_hi_647 = {dataGroup_hi_hi_647, dataGroup_hi_lo_647};
  wire [15:0]   dataGroup_7_44 = dataGroup_lo_647[495:480];
  wire [31:0]   res_lo_lo_44 = {dataGroup_1_44, dataGroup_0_44};
  wire [31:0]   res_lo_hi_44 = {dataGroup_3_44, dataGroup_2_44};
  wire [63:0]   res_lo_44 = {res_lo_hi_44, res_lo_lo_44};
  wire [31:0]   res_hi_lo_44 = {dataGroup_5_44, dataGroup_4_44};
  wire [31:0]   res_hi_hi_44 = {dataGroup_7_44, dataGroup_6_44};
  wire [63:0]   res_hi_44 = {res_hi_hi_44, res_hi_lo_44};
  wire [127:0]  res_90 = {res_hi_44, res_lo_44};
  wire [511:0]  dataGroup_lo_648 = {dataGroup_lo_hi_648, dataGroup_lo_lo_648};
  wire [511:0]  dataGroup_hi_648 = {dataGroup_hi_hi_648, dataGroup_hi_lo_648};
  wire [15:0]   dataGroup_0_45 = dataGroup_lo_648[63:48];
  wire [511:0]  dataGroup_lo_649 = {dataGroup_lo_hi_649, dataGroup_lo_lo_649};
  wire [511:0]  dataGroup_hi_649 = {dataGroup_hi_hi_649, dataGroup_hi_lo_649};
  wire [15:0]   dataGroup_1_45 = dataGroup_lo_649[127:112];
  wire [511:0]  dataGroup_lo_650 = {dataGroup_lo_hi_650, dataGroup_lo_lo_650};
  wire [511:0]  dataGroup_hi_650 = {dataGroup_hi_hi_650, dataGroup_hi_lo_650};
  wire [15:0]   dataGroup_2_45 = dataGroup_lo_650[191:176];
  wire [511:0]  dataGroup_lo_651 = {dataGroup_lo_hi_651, dataGroup_lo_lo_651};
  wire [511:0]  dataGroup_hi_651 = {dataGroup_hi_hi_651, dataGroup_hi_lo_651};
  wire [15:0]   dataGroup_3_45 = dataGroup_lo_651[255:240];
  wire [511:0]  dataGroup_lo_652 = {dataGroup_lo_hi_652, dataGroup_lo_lo_652};
  wire [511:0]  dataGroup_hi_652 = {dataGroup_hi_hi_652, dataGroup_hi_lo_652};
  wire [15:0]   dataGroup_4_45 = dataGroup_lo_652[319:304];
  wire [511:0]  dataGroup_lo_653 = {dataGroup_lo_hi_653, dataGroup_lo_lo_653};
  wire [511:0]  dataGroup_hi_653 = {dataGroup_hi_hi_653, dataGroup_hi_lo_653};
  wire [15:0]   dataGroup_5_45 = dataGroup_lo_653[383:368];
  wire [511:0]  dataGroup_lo_654 = {dataGroup_lo_hi_654, dataGroup_lo_lo_654};
  wire [511:0]  dataGroup_hi_654 = {dataGroup_hi_hi_654, dataGroup_hi_lo_654};
  wire [15:0]   dataGroup_6_45 = dataGroup_lo_654[447:432];
  wire [511:0]  dataGroup_lo_655 = {dataGroup_lo_hi_655, dataGroup_lo_lo_655};
  wire [511:0]  dataGroup_hi_655 = {dataGroup_hi_hi_655, dataGroup_hi_lo_655};
  wire [15:0]   dataGroup_7_45 = dataGroup_lo_655[511:496];
  wire [31:0]   res_lo_lo_45 = {dataGroup_1_45, dataGroup_0_45};
  wire [31:0]   res_lo_hi_45 = {dataGroup_3_45, dataGroup_2_45};
  wire [63:0]   res_lo_45 = {res_lo_hi_45, res_lo_lo_45};
  wire [31:0]   res_hi_lo_45 = {dataGroup_5_45, dataGroup_4_45};
  wire [31:0]   res_hi_hi_45 = {dataGroup_7_45, dataGroup_6_45};
  wire [63:0]   res_hi_45 = {res_hi_hi_45, res_hi_lo_45};
  wire [127:0]  res_91 = {res_hi_45, res_lo_45};
  wire [255:0]  lo_lo_11 = {res_89, res_88};
  wire [255:0]  lo_hi_11 = {res_91, res_90};
  wire [511:0]  lo_11 = {lo_hi_11, lo_lo_11};
  wire [1023:0] regroupLoadData_1_3 = {512'h0, lo_11};
  wire [511:0]  dataGroup_lo_656 = {dataGroup_lo_hi_656, dataGroup_lo_lo_656};
  wire [511:0]  dataGroup_hi_656 = {dataGroup_hi_hi_656, dataGroup_hi_lo_656};
  wire [15:0]   dataGroup_0_46 = dataGroup_lo_656[15:0];
  wire [511:0]  dataGroup_lo_657 = {dataGroup_lo_hi_657, dataGroup_lo_lo_657};
  wire [511:0]  dataGroup_hi_657 = {dataGroup_hi_hi_657, dataGroup_hi_lo_657};
  wire [15:0]   dataGroup_1_46 = dataGroup_lo_657[95:80];
  wire [511:0]  dataGroup_lo_658 = {dataGroup_lo_hi_658, dataGroup_lo_lo_658};
  wire [511:0]  dataGroup_hi_658 = {dataGroup_hi_hi_658, dataGroup_hi_lo_658};
  wire [15:0]   dataGroup_2_46 = dataGroup_lo_658[175:160];
  wire [511:0]  dataGroup_lo_659 = {dataGroup_lo_hi_659, dataGroup_lo_lo_659};
  wire [511:0]  dataGroup_hi_659 = {dataGroup_hi_hi_659, dataGroup_hi_lo_659};
  wire [15:0]   dataGroup_3_46 = dataGroup_lo_659[255:240];
  wire [511:0]  dataGroup_lo_660 = {dataGroup_lo_hi_660, dataGroup_lo_lo_660};
  wire [511:0]  dataGroup_hi_660 = {dataGroup_hi_hi_660, dataGroup_hi_lo_660};
  wire [15:0]   dataGroup_4_46 = dataGroup_lo_660[335:320];
  wire [511:0]  dataGroup_lo_661 = {dataGroup_lo_hi_661, dataGroup_lo_lo_661};
  wire [511:0]  dataGroup_hi_661 = {dataGroup_hi_hi_661, dataGroup_hi_lo_661};
  wire [15:0]   dataGroup_5_46 = dataGroup_lo_661[415:400];
  wire [511:0]  dataGroup_lo_662 = {dataGroup_lo_hi_662, dataGroup_lo_lo_662};
  wire [511:0]  dataGroup_hi_662 = {dataGroup_hi_hi_662, dataGroup_hi_lo_662};
  wire [15:0]   dataGroup_6_46 = dataGroup_lo_662[495:480];
  wire [511:0]  dataGroup_lo_663 = {dataGroup_lo_hi_663, dataGroup_lo_lo_663};
  wire [511:0]  dataGroup_hi_663 = {dataGroup_hi_hi_663, dataGroup_hi_lo_663};
  wire [15:0]   dataGroup_7_46 = dataGroup_hi_663[63:48];
  wire [31:0]   res_lo_lo_46 = {dataGroup_1_46, dataGroup_0_46};
  wire [31:0]   res_lo_hi_46 = {dataGroup_3_46, dataGroup_2_46};
  wire [63:0]   res_lo_46 = {res_lo_hi_46, res_lo_lo_46};
  wire [31:0]   res_hi_lo_46 = {dataGroup_5_46, dataGroup_4_46};
  wire [31:0]   res_hi_hi_46 = {dataGroup_7_46, dataGroup_6_46};
  wire [63:0]   res_hi_46 = {res_hi_hi_46, res_hi_lo_46};
  wire [127:0]  res_96 = {res_hi_46, res_lo_46};
  wire [511:0]  dataGroup_lo_664 = {dataGroup_lo_hi_664, dataGroup_lo_lo_664};
  wire [511:0]  dataGroup_hi_664 = {dataGroup_hi_hi_664, dataGroup_hi_lo_664};
  wire [15:0]   dataGroup_0_47 = dataGroup_lo_664[31:16];
  wire [511:0]  dataGroup_lo_665 = {dataGroup_lo_hi_665, dataGroup_lo_lo_665};
  wire [511:0]  dataGroup_hi_665 = {dataGroup_hi_hi_665, dataGroup_hi_lo_665};
  wire [15:0]   dataGroup_1_47 = dataGroup_lo_665[111:96];
  wire [511:0]  dataGroup_lo_666 = {dataGroup_lo_hi_666, dataGroup_lo_lo_666};
  wire [511:0]  dataGroup_hi_666 = {dataGroup_hi_hi_666, dataGroup_hi_lo_666};
  wire [15:0]   dataGroup_2_47 = dataGroup_lo_666[191:176];
  wire [511:0]  dataGroup_lo_667 = {dataGroup_lo_hi_667, dataGroup_lo_lo_667};
  wire [511:0]  dataGroup_hi_667 = {dataGroup_hi_hi_667, dataGroup_hi_lo_667};
  wire [15:0]   dataGroup_3_47 = dataGroup_lo_667[271:256];
  wire [511:0]  dataGroup_lo_668 = {dataGroup_lo_hi_668, dataGroup_lo_lo_668};
  wire [511:0]  dataGroup_hi_668 = {dataGroup_hi_hi_668, dataGroup_hi_lo_668};
  wire [15:0]   dataGroup_4_47 = dataGroup_lo_668[351:336];
  wire [511:0]  dataGroup_lo_669 = {dataGroup_lo_hi_669, dataGroup_lo_lo_669};
  wire [511:0]  dataGroup_hi_669 = {dataGroup_hi_hi_669, dataGroup_hi_lo_669};
  wire [15:0]   dataGroup_5_47 = dataGroup_lo_669[431:416];
  wire [511:0]  dataGroup_lo_670 = {dataGroup_lo_hi_670, dataGroup_lo_lo_670};
  wire [511:0]  dataGroup_hi_670 = {dataGroup_hi_hi_670, dataGroup_hi_lo_670};
  wire [15:0]   dataGroup_6_47 = dataGroup_lo_670[511:496];
  wire [511:0]  dataGroup_lo_671 = {dataGroup_lo_hi_671, dataGroup_lo_lo_671};
  wire [511:0]  dataGroup_hi_671 = {dataGroup_hi_hi_671, dataGroup_hi_lo_671};
  wire [15:0]   dataGroup_7_47 = dataGroup_hi_671[79:64];
  wire [31:0]   res_lo_lo_47 = {dataGroup_1_47, dataGroup_0_47};
  wire [31:0]   res_lo_hi_47 = {dataGroup_3_47, dataGroup_2_47};
  wire [63:0]   res_lo_47 = {res_lo_hi_47, res_lo_lo_47};
  wire [31:0]   res_hi_lo_47 = {dataGroup_5_47, dataGroup_4_47};
  wire [31:0]   res_hi_hi_47 = {dataGroup_7_47, dataGroup_6_47};
  wire [63:0]   res_hi_47 = {res_hi_hi_47, res_hi_lo_47};
  wire [127:0]  res_97 = {res_hi_47, res_lo_47};
  wire [511:0]  dataGroup_lo_672 = {dataGroup_lo_hi_672, dataGroup_lo_lo_672};
  wire [511:0]  dataGroup_hi_672 = {dataGroup_hi_hi_672, dataGroup_hi_lo_672};
  wire [15:0]   dataGroup_0_48 = dataGroup_lo_672[47:32];
  wire [511:0]  dataGroup_lo_673 = {dataGroup_lo_hi_673, dataGroup_lo_lo_673};
  wire [511:0]  dataGroup_hi_673 = {dataGroup_hi_hi_673, dataGroup_hi_lo_673};
  wire [15:0]   dataGroup_1_48 = dataGroup_lo_673[127:112];
  wire [511:0]  dataGroup_lo_674 = {dataGroup_lo_hi_674, dataGroup_lo_lo_674};
  wire [511:0]  dataGroup_hi_674 = {dataGroup_hi_hi_674, dataGroup_hi_lo_674};
  wire [15:0]   dataGroup_2_48 = dataGroup_lo_674[207:192];
  wire [511:0]  dataGroup_lo_675 = {dataGroup_lo_hi_675, dataGroup_lo_lo_675};
  wire [511:0]  dataGroup_hi_675 = {dataGroup_hi_hi_675, dataGroup_hi_lo_675};
  wire [15:0]   dataGroup_3_48 = dataGroup_lo_675[287:272];
  wire [511:0]  dataGroup_lo_676 = {dataGroup_lo_hi_676, dataGroup_lo_lo_676};
  wire [511:0]  dataGroup_hi_676 = {dataGroup_hi_hi_676, dataGroup_hi_lo_676};
  wire [15:0]   dataGroup_4_48 = dataGroup_lo_676[367:352];
  wire [511:0]  dataGroup_lo_677 = {dataGroup_lo_hi_677, dataGroup_lo_lo_677};
  wire [511:0]  dataGroup_hi_677 = {dataGroup_hi_hi_677, dataGroup_hi_lo_677};
  wire [15:0]   dataGroup_5_48 = dataGroup_lo_677[447:432];
  wire [511:0]  dataGroup_lo_678 = {dataGroup_lo_hi_678, dataGroup_lo_lo_678};
  wire [511:0]  dataGroup_hi_678 = {dataGroup_hi_hi_678, dataGroup_hi_lo_678};
  wire [15:0]   dataGroup_6_48 = dataGroup_hi_678[15:0];
  wire [511:0]  dataGroup_lo_679 = {dataGroup_lo_hi_679, dataGroup_lo_lo_679};
  wire [511:0]  dataGroup_hi_679 = {dataGroup_hi_hi_679, dataGroup_hi_lo_679};
  wire [15:0]   dataGroup_7_48 = dataGroup_hi_679[95:80];
  wire [31:0]   res_lo_lo_48 = {dataGroup_1_48, dataGroup_0_48};
  wire [31:0]   res_lo_hi_48 = {dataGroup_3_48, dataGroup_2_48};
  wire [63:0]   res_lo_48 = {res_lo_hi_48, res_lo_lo_48};
  wire [31:0]   res_hi_lo_48 = {dataGroup_5_48, dataGroup_4_48};
  wire [31:0]   res_hi_hi_48 = {dataGroup_7_48, dataGroup_6_48};
  wire [63:0]   res_hi_48 = {res_hi_hi_48, res_hi_lo_48};
  wire [127:0]  res_98 = {res_hi_48, res_lo_48};
  wire [511:0]  dataGroup_lo_680 = {dataGroup_lo_hi_680, dataGroup_lo_lo_680};
  wire [511:0]  dataGroup_hi_680 = {dataGroup_hi_hi_680, dataGroup_hi_lo_680};
  wire [15:0]   dataGroup_0_49 = dataGroup_lo_680[63:48];
  wire [511:0]  dataGroup_lo_681 = {dataGroup_lo_hi_681, dataGroup_lo_lo_681};
  wire [511:0]  dataGroup_hi_681 = {dataGroup_hi_hi_681, dataGroup_hi_lo_681};
  wire [15:0]   dataGroup_1_49 = dataGroup_lo_681[143:128];
  wire [511:0]  dataGroup_lo_682 = {dataGroup_lo_hi_682, dataGroup_lo_lo_682};
  wire [511:0]  dataGroup_hi_682 = {dataGroup_hi_hi_682, dataGroup_hi_lo_682};
  wire [15:0]   dataGroup_2_49 = dataGroup_lo_682[223:208];
  wire [511:0]  dataGroup_lo_683 = {dataGroup_lo_hi_683, dataGroup_lo_lo_683};
  wire [511:0]  dataGroup_hi_683 = {dataGroup_hi_hi_683, dataGroup_hi_lo_683};
  wire [15:0]   dataGroup_3_49 = dataGroup_lo_683[303:288];
  wire [511:0]  dataGroup_lo_684 = {dataGroup_lo_hi_684, dataGroup_lo_lo_684};
  wire [511:0]  dataGroup_hi_684 = {dataGroup_hi_hi_684, dataGroup_hi_lo_684};
  wire [15:0]   dataGroup_4_49 = dataGroup_lo_684[383:368];
  wire [511:0]  dataGroup_lo_685 = {dataGroup_lo_hi_685, dataGroup_lo_lo_685};
  wire [511:0]  dataGroup_hi_685 = {dataGroup_hi_hi_685, dataGroup_hi_lo_685};
  wire [15:0]   dataGroup_5_49 = dataGroup_lo_685[463:448];
  wire [511:0]  dataGroup_lo_686 = {dataGroup_lo_hi_686, dataGroup_lo_lo_686};
  wire [511:0]  dataGroup_hi_686 = {dataGroup_hi_hi_686, dataGroup_hi_lo_686};
  wire [15:0]   dataGroup_6_49 = dataGroup_hi_686[31:16];
  wire [511:0]  dataGroup_lo_687 = {dataGroup_lo_hi_687, dataGroup_lo_lo_687};
  wire [511:0]  dataGroup_hi_687 = {dataGroup_hi_hi_687, dataGroup_hi_lo_687};
  wire [15:0]   dataGroup_7_49 = dataGroup_hi_687[111:96];
  wire [31:0]   res_lo_lo_49 = {dataGroup_1_49, dataGroup_0_49};
  wire [31:0]   res_lo_hi_49 = {dataGroup_3_49, dataGroup_2_49};
  wire [63:0]   res_lo_49 = {res_lo_hi_49, res_lo_lo_49};
  wire [31:0]   res_hi_lo_49 = {dataGroup_5_49, dataGroup_4_49};
  wire [31:0]   res_hi_hi_49 = {dataGroup_7_49, dataGroup_6_49};
  wire [63:0]   res_hi_49 = {res_hi_hi_49, res_hi_lo_49};
  wire [127:0]  res_99 = {res_hi_49, res_lo_49};
  wire [511:0]  dataGroup_lo_688 = {dataGroup_lo_hi_688, dataGroup_lo_lo_688};
  wire [511:0]  dataGroup_hi_688 = {dataGroup_hi_hi_688, dataGroup_hi_lo_688};
  wire [15:0]   dataGroup_0_50 = dataGroup_lo_688[79:64];
  wire [511:0]  dataGroup_lo_689 = {dataGroup_lo_hi_689, dataGroup_lo_lo_689};
  wire [511:0]  dataGroup_hi_689 = {dataGroup_hi_hi_689, dataGroup_hi_lo_689};
  wire [15:0]   dataGroup_1_50 = dataGroup_lo_689[159:144];
  wire [511:0]  dataGroup_lo_690 = {dataGroup_lo_hi_690, dataGroup_lo_lo_690};
  wire [511:0]  dataGroup_hi_690 = {dataGroup_hi_hi_690, dataGroup_hi_lo_690};
  wire [15:0]   dataGroup_2_50 = dataGroup_lo_690[239:224];
  wire [511:0]  dataGroup_lo_691 = {dataGroup_lo_hi_691, dataGroup_lo_lo_691};
  wire [511:0]  dataGroup_hi_691 = {dataGroup_hi_hi_691, dataGroup_hi_lo_691};
  wire [15:0]   dataGroup_3_50 = dataGroup_lo_691[319:304];
  wire [511:0]  dataGroup_lo_692 = {dataGroup_lo_hi_692, dataGroup_lo_lo_692};
  wire [511:0]  dataGroup_hi_692 = {dataGroup_hi_hi_692, dataGroup_hi_lo_692};
  wire [15:0]   dataGroup_4_50 = dataGroup_lo_692[399:384];
  wire [511:0]  dataGroup_lo_693 = {dataGroup_lo_hi_693, dataGroup_lo_lo_693};
  wire [511:0]  dataGroup_hi_693 = {dataGroup_hi_hi_693, dataGroup_hi_lo_693};
  wire [15:0]   dataGroup_5_50 = dataGroup_lo_693[479:464];
  wire [511:0]  dataGroup_lo_694 = {dataGroup_lo_hi_694, dataGroup_lo_lo_694};
  wire [511:0]  dataGroup_hi_694 = {dataGroup_hi_hi_694, dataGroup_hi_lo_694};
  wire [15:0]   dataGroup_6_50 = dataGroup_hi_694[47:32];
  wire [511:0]  dataGroup_lo_695 = {dataGroup_lo_hi_695, dataGroup_lo_lo_695};
  wire [511:0]  dataGroup_hi_695 = {dataGroup_hi_hi_695, dataGroup_hi_lo_695};
  wire [15:0]   dataGroup_7_50 = dataGroup_hi_695[127:112];
  wire [31:0]   res_lo_lo_50 = {dataGroup_1_50, dataGroup_0_50};
  wire [31:0]   res_lo_hi_50 = {dataGroup_3_50, dataGroup_2_50};
  wire [63:0]   res_lo_50 = {res_lo_hi_50, res_lo_lo_50};
  wire [31:0]   res_hi_lo_50 = {dataGroup_5_50, dataGroup_4_50};
  wire [31:0]   res_hi_hi_50 = {dataGroup_7_50, dataGroup_6_50};
  wire [63:0]   res_hi_50 = {res_hi_hi_50, res_hi_lo_50};
  wire [127:0]  res_100 = {res_hi_50, res_lo_50};
  wire [255:0]  lo_lo_12 = {res_97, res_96};
  wire [255:0]  lo_hi_12 = {res_99, res_98};
  wire [511:0]  lo_12 = {lo_hi_12, lo_lo_12};
  wire [255:0]  hi_lo_12 = {128'h0, res_100};
  wire [511:0]  hi_12 = {256'h0, hi_lo_12};
  wire [1023:0] regroupLoadData_1_4 = {hi_12, lo_12};
  wire [511:0]  dataGroup_lo_696 = {dataGroup_lo_hi_696, dataGroup_lo_lo_696};
  wire [511:0]  dataGroup_hi_696 = {dataGroup_hi_hi_696, dataGroup_hi_lo_696};
  wire [15:0]   dataGroup_0_51 = dataGroup_lo_696[15:0];
  wire [511:0]  dataGroup_lo_697 = {dataGroup_lo_hi_697, dataGroup_lo_lo_697};
  wire [511:0]  dataGroup_hi_697 = {dataGroup_hi_hi_697, dataGroup_hi_lo_697};
  wire [15:0]   dataGroup_1_51 = dataGroup_lo_697[111:96];
  wire [511:0]  dataGroup_lo_698 = {dataGroup_lo_hi_698, dataGroup_lo_lo_698};
  wire [511:0]  dataGroup_hi_698 = {dataGroup_hi_hi_698, dataGroup_hi_lo_698};
  wire [15:0]   dataGroup_2_51 = dataGroup_lo_698[207:192];
  wire [511:0]  dataGroup_lo_699 = {dataGroup_lo_hi_699, dataGroup_lo_lo_699};
  wire [511:0]  dataGroup_hi_699 = {dataGroup_hi_hi_699, dataGroup_hi_lo_699};
  wire [15:0]   dataGroup_3_51 = dataGroup_lo_699[303:288];
  wire [511:0]  dataGroup_lo_700 = {dataGroup_lo_hi_700, dataGroup_lo_lo_700};
  wire [511:0]  dataGroup_hi_700 = {dataGroup_hi_hi_700, dataGroup_hi_lo_700};
  wire [15:0]   dataGroup_4_51 = dataGroup_lo_700[399:384];
  wire [511:0]  dataGroup_lo_701 = {dataGroup_lo_hi_701, dataGroup_lo_lo_701};
  wire [511:0]  dataGroup_hi_701 = {dataGroup_hi_hi_701, dataGroup_hi_lo_701};
  wire [15:0]   dataGroup_5_51 = dataGroup_lo_701[495:480];
  wire [511:0]  dataGroup_lo_702 = {dataGroup_lo_hi_702, dataGroup_lo_lo_702};
  wire [511:0]  dataGroup_hi_702 = {dataGroup_hi_hi_702, dataGroup_hi_lo_702};
  wire [15:0]   dataGroup_6_51 = dataGroup_hi_702[79:64];
  wire [511:0]  dataGroup_lo_703 = {dataGroup_lo_hi_703, dataGroup_lo_lo_703};
  wire [511:0]  dataGroup_hi_703 = {dataGroup_hi_hi_703, dataGroup_hi_lo_703};
  wire [15:0]   dataGroup_7_51 = dataGroup_hi_703[175:160];
  wire [31:0]   res_lo_lo_51 = {dataGroup_1_51, dataGroup_0_51};
  wire [31:0]   res_lo_hi_51 = {dataGroup_3_51, dataGroup_2_51};
  wire [63:0]   res_lo_51 = {res_lo_hi_51, res_lo_lo_51};
  wire [31:0]   res_hi_lo_51 = {dataGroup_5_51, dataGroup_4_51};
  wire [31:0]   res_hi_hi_51 = {dataGroup_7_51, dataGroup_6_51};
  wire [63:0]   res_hi_51 = {res_hi_hi_51, res_hi_lo_51};
  wire [127:0]  res_104 = {res_hi_51, res_lo_51};
  wire [511:0]  dataGroup_lo_704 = {dataGroup_lo_hi_704, dataGroup_lo_lo_704};
  wire [511:0]  dataGroup_hi_704 = {dataGroup_hi_hi_704, dataGroup_hi_lo_704};
  wire [15:0]   dataGroup_0_52 = dataGroup_lo_704[31:16];
  wire [511:0]  dataGroup_lo_705 = {dataGroup_lo_hi_705, dataGroup_lo_lo_705};
  wire [511:0]  dataGroup_hi_705 = {dataGroup_hi_hi_705, dataGroup_hi_lo_705};
  wire [15:0]   dataGroup_1_52 = dataGroup_lo_705[127:112];
  wire [511:0]  dataGroup_lo_706 = {dataGroup_lo_hi_706, dataGroup_lo_lo_706};
  wire [511:0]  dataGroup_hi_706 = {dataGroup_hi_hi_706, dataGroup_hi_lo_706};
  wire [15:0]   dataGroup_2_52 = dataGroup_lo_706[223:208];
  wire [511:0]  dataGroup_lo_707 = {dataGroup_lo_hi_707, dataGroup_lo_lo_707};
  wire [511:0]  dataGroup_hi_707 = {dataGroup_hi_hi_707, dataGroup_hi_lo_707};
  wire [15:0]   dataGroup_3_52 = dataGroup_lo_707[319:304];
  wire [511:0]  dataGroup_lo_708 = {dataGroup_lo_hi_708, dataGroup_lo_lo_708};
  wire [511:0]  dataGroup_hi_708 = {dataGroup_hi_hi_708, dataGroup_hi_lo_708};
  wire [15:0]   dataGroup_4_52 = dataGroup_lo_708[415:400];
  wire [511:0]  dataGroup_lo_709 = {dataGroup_lo_hi_709, dataGroup_lo_lo_709};
  wire [511:0]  dataGroup_hi_709 = {dataGroup_hi_hi_709, dataGroup_hi_lo_709};
  wire [15:0]   dataGroup_5_52 = dataGroup_lo_709[511:496];
  wire [511:0]  dataGroup_lo_710 = {dataGroup_lo_hi_710, dataGroup_lo_lo_710};
  wire [511:0]  dataGroup_hi_710 = {dataGroup_hi_hi_710, dataGroup_hi_lo_710};
  wire [15:0]   dataGroup_6_52 = dataGroup_hi_710[95:80];
  wire [511:0]  dataGroup_lo_711 = {dataGroup_lo_hi_711, dataGroup_lo_lo_711};
  wire [511:0]  dataGroup_hi_711 = {dataGroup_hi_hi_711, dataGroup_hi_lo_711};
  wire [15:0]   dataGroup_7_52 = dataGroup_hi_711[191:176];
  wire [31:0]   res_lo_lo_52 = {dataGroup_1_52, dataGroup_0_52};
  wire [31:0]   res_lo_hi_52 = {dataGroup_3_52, dataGroup_2_52};
  wire [63:0]   res_lo_52 = {res_lo_hi_52, res_lo_lo_52};
  wire [31:0]   res_hi_lo_52 = {dataGroup_5_52, dataGroup_4_52};
  wire [31:0]   res_hi_hi_52 = {dataGroup_7_52, dataGroup_6_52};
  wire [63:0]   res_hi_52 = {res_hi_hi_52, res_hi_lo_52};
  wire [127:0]  res_105 = {res_hi_52, res_lo_52};
  wire [511:0]  dataGroup_lo_712 = {dataGroup_lo_hi_712, dataGroup_lo_lo_712};
  wire [511:0]  dataGroup_hi_712 = {dataGroup_hi_hi_712, dataGroup_hi_lo_712};
  wire [15:0]   dataGroup_0_53 = dataGroup_lo_712[47:32];
  wire [511:0]  dataGroup_lo_713 = {dataGroup_lo_hi_713, dataGroup_lo_lo_713};
  wire [511:0]  dataGroup_hi_713 = {dataGroup_hi_hi_713, dataGroup_hi_lo_713};
  wire [15:0]   dataGroup_1_53 = dataGroup_lo_713[143:128];
  wire [511:0]  dataGroup_lo_714 = {dataGroup_lo_hi_714, dataGroup_lo_lo_714};
  wire [511:0]  dataGroup_hi_714 = {dataGroup_hi_hi_714, dataGroup_hi_lo_714};
  wire [15:0]   dataGroup_2_53 = dataGroup_lo_714[239:224];
  wire [511:0]  dataGroup_lo_715 = {dataGroup_lo_hi_715, dataGroup_lo_lo_715};
  wire [511:0]  dataGroup_hi_715 = {dataGroup_hi_hi_715, dataGroup_hi_lo_715};
  wire [15:0]   dataGroup_3_53 = dataGroup_lo_715[335:320];
  wire [511:0]  dataGroup_lo_716 = {dataGroup_lo_hi_716, dataGroup_lo_lo_716};
  wire [511:0]  dataGroup_hi_716 = {dataGroup_hi_hi_716, dataGroup_hi_lo_716};
  wire [15:0]   dataGroup_4_53 = dataGroup_lo_716[431:416];
  wire [511:0]  dataGroup_lo_717 = {dataGroup_lo_hi_717, dataGroup_lo_lo_717};
  wire [511:0]  dataGroup_hi_717 = {dataGroup_hi_hi_717, dataGroup_hi_lo_717};
  wire [15:0]   dataGroup_5_53 = dataGroup_hi_717[15:0];
  wire [511:0]  dataGroup_lo_718 = {dataGroup_lo_hi_718, dataGroup_lo_lo_718};
  wire [511:0]  dataGroup_hi_718 = {dataGroup_hi_hi_718, dataGroup_hi_lo_718};
  wire [15:0]   dataGroup_6_53 = dataGroup_hi_718[111:96];
  wire [511:0]  dataGroup_lo_719 = {dataGroup_lo_hi_719, dataGroup_lo_lo_719};
  wire [511:0]  dataGroup_hi_719 = {dataGroup_hi_hi_719, dataGroup_hi_lo_719};
  wire [15:0]   dataGroup_7_53 = dataGroup_hi_719[207:192];
  wire [31:0]   res_lo_lo_53 = {dataGroup_1_53, dataGroup_0_53};
  wire [31:0]   res_lo_hi_53 = {dataGroup_3_53, dataGroup_2_53};
  wire [63:0]   res_lo_53 = {res_lo_hi_53, res_lo_lo_53};
  wire [31:0]   res_hi_lo_53 = {dataGroup_5_53, dataGroup_4_53};
  wire [31:0]   res_hi_hi_53 = {dataGroup_7_53, dataGroup_6_53};
  wire [63:0]   res_hi_53 = {res_hi_hi_53, res_hi_lo_53};
  wire [127:0]  res_106 = {res_hi_53, res_lo_53};
  wire [511:0]  dataGroup_lo_720 = {dataGroup_lo_hi_720, dataGroup_lo_lo_720};
  wire [511:0]  dataGroup_hi_720 = {dataGroup_hi_hi_720, dataGroup_hi_lo_720};
  wire [15:0]   dataGroup_0_54 = dataGroup_lo_720[63:48];
  wire [511:0]  dataGroup_lo_721 = {dataGroup_lo_hi_721, dataGroup_lo_lo_721};
  wire [511:0]  dataGroup_hi_721 = {dataGroup_hi_hi_721, dataGroup_hi_lo_721};
  wire [15:0]   dataGroup_1_54 = dataGroup_lo_721[159:144];
  wire [511:0]  dataGroup_lo_722 = {dataGroup_lo_hi_722, dataGroup_lo_lo_722};
  wire [511:0]  dataGroup_hi_722 = {dataGroup_hi_hi_722, dataGroup_hi_lo_722};
  wire [15:0]   dataGroup_2_54 = dataGroup_lo_722[255:240];
  wire [511:0]  dataGroup_lo_723 = {dataGroup_lo_hi_723, dataGroup_lo_lo_723};
  wire [511:0]  dataGroup_hi_723 = {dataGroup_hi_hi_723, dataGroup_hi_lo_723};
  wire [15:0]   dataGroup_3_54 = dataGroup_lo_723[351:336];
  wire [511:0]  dataGroup_lo_724 = {dataGroup_lo_hi_724, dataGroup_lo_lo_724};
  wire [511:0]  dataGroup_hi_724 = {dataGroup_hi_hi_724, dataGroup_hi_lo_724};
  wire [15:0]   dataGroup_4_54 = dataGroup_lo_724[447:432];
  wire [511:0]  dataGroup_lo_725 = {dataGroup_lo_hi_725, dataGroup_lo_lo_725};
  wire [511:0]  dataGroup_hi_725 = {dataGroup_hi_hi_725, dataGroup_hi_lo_725};
  wire [15:0]   dataGroup_5_54 = dataGroup_hi_725[31:16];
  wire [511:0]  dataGroup_lo_726 = {dataGroup_lo_hi_726, dataGroup_lo_lo_726};
  wire [511:0]  dataGroup_hi_726 = {dataGroup_hi_hi_726, dataGroup_hi_lo_726};
  wire [15:0]   dataGroup_6_54 = dataGroup_hi_726[127:112];
  wire [511:0]  dataGroup_lo_727 = {dataGroup_lo_hi_727, dataGroup_lo_lo_727};
  wire [511:0]  dataGroup_hi_727 = {dataGroup_hi_hi_727, dataGroup_hi_lo_727};
  wire [15:0]   dataGroup_7_54 = dataGroup_hi_727[223:208];
  wire [31:0]   res_lo_lo_54 = {dataGroup_1_54, dataGroup_0_54};
  wire [31:0]   res_lo_hi_54 = {dataGroup_3_54, dataGroup_2_54};
  wire [63:0]   res_lo_54 = {res_lo_hi_54, res_lo_lo_54};
  wire [31:0]   res_hi_lo_54 = {dataGroup_5_54, dataGroup_4_54};
  wire [31:0]   res_hi_hi_54 = {dataGroup_7_54, dataGroup_6_54};
  wire [63:0]   res_hi_54 = {res_hi_hi_54, res_hi_lo_54};
  wire [127:0]  res_107 = {res_hi_54, res_lo_54};
  wire [511:0]  dataGroup_lo_728 = {dataGroup_lo_hi_728, dataGroup_lo_lo_728};
  wire [511:0]  dataGroup_hi_728 = {dataGroup_hi_hi_728, dataGroup_hi_lo_728};
  wire [15:0]   dataGroup_0_55 = dataGroup_lo_728[79:64];
  wire [511:0]  dataGroup_lo_729 = {dataGroup_lo_hi_729, dataGroup_lo_lo_729};
  wire [511:0]  dataGroup_hi_729 = {dataGroup_hi_hi_729, dataGroup_hi_lo_729};
  wire [15:0]   dataGroup_1_55 = dataGroup_lo_729[175:160];
  wire [511:0]  dataGroup_lo_730 = {dataGroup_lo_hi_730, dataGroup_lo_lo_730};
  wire [511:0]  dataGroup_hi_730 = {dataGroup_hi_hi_730, dataGroup_hi_lo_730};
  wire [15:0]   dataGroup_2_55 = dataGroup_lo_730[271:256];
  wire [511:0]  dataGroup_lo_731 = {dataGroup_lo_hi_731, dataGroup_lo_lo_731};
  wire [511:0]  dataGroup_hi_731 = {dataGroup_hi_hi_731, dataGroup_hi_lo_731};
  wire [15:0]   dataGroup_3_55 = dataGroup_lo_731[367:352];
  wire [511:0]  dataGroup_lo_732 = {dataGroup_lo_hi_732, dataGroup_lo_lo_732};
  wire [511:0]  dataGroup_hi_732 = {dataGroup_hi_hi_732, dataGroup_hi_lo_732};
  wire [15:0]   dataGroup_4_55 = dataGroup_lo_732[463:448];
  wire [511:0]  dataGroup_lo_733 = {dataGroup_lo_hi_733, dataGroup_lo_lo_733};
  wire [511:0]  dataGroup_hi_733 = {dataGroup_hi_hi_733, dataGroup_hi_lo_733};
  wire [15:0]   dataGroup_5_55 = dataGroup_hi_733[47:32];
  wire [511:0]  dataGroup_lo_734 = {dataGroup_lo_hi_734, dataGroup_lo_lo_734};
  wire [511:0]  dataGroup_hi_734 = {dataGroup_hi_hi_734, dataGroup_hi_lo_734};
  wire [15:0]   dataGroup_6_55 = dataGroup_hi_734[143:128];
  wire [511:0]  dataGroup_lo_735 = {dataGroup_lo_hi_735, dataGroup_lo_lo_735};
  wire [511:0]  dataGroup_hi_735 = {dataGroup_hi_hi_735, dataGroup_hi_lo_735};
  wire [15:0]   dataGroup_7_55 = dataGroup_hi_735[239:224];
  wire [31:0]   res_lo_lo_55 = {dataGroup_1_55, dataGroup_0_55};
  wire [31:0]   res_lo_hi_55 = {dataGroup_3_55, dataGroup_2_55};
  wire [63:0]   res_lo_55 = {res_lo_hi_55, res_lo_lo_55};
  wire [31:0]   res_hi_lo_55 = {dataGroup_5_55, dataGroup_4_55};
  wire [31:0]   res_hi_hi_55 = {dataGroup_7_55, dataGroup_6_55};
  wire [63:0]   res_hi_55 = {res_hi_hi_55, res_hi_lo_55};
  wire [127:0]  res_108 = {res_hi_55, res_lo_55};
  wire [511:0]  dataGroup_lo_736 = {dataGroup_lo_hi_736, dataGroup_lo_lo_736};
  wire [511:0]  dataGroup_hi_736 = {dataGroup_hi_hi_736, dataGroup_hi_lo_736};
  wire [15:0]   dataGroup_0_56 = dataGroup_lo_736[95:80];
  wire [511:0]  dataGroup_lo_737 = {dataGroup_lo_hi_737, dataGroup_lo_lo_737};
  wire [511:0]  dataGroup_hi_737 = {dataGroup_hi_hi_737, dataGroup_hi_lo_737};
  wire [15:0]   dataGroup_1_56 = dataGroup_lo_737[191:176];
  wire [511:0]  dataGroup_lo_738 = {dataGroup_lo_hi_738, dataGroup_lo_lo_738};
  wire [511:0]  dataGroup_hi_738 = {dataGroup_hi_hi_738, dataGroup_hi_lo_738};
  wire [15:0]   dataGroup_2_56 = dataGroup_lo_738[287:272];
  wire [511:0]  dataGroup_lo_739 = {dataGroup_lo_hi_739, dataGroup_lo_lo_739};
  wire [511:0]  dataGroup_hi_739 = {dataGroup_hi_hi_739, dataGroup_hi_lo_739};
  wire [15:0]   dataGroup_3_56 = dataGroup_lo_739[383:368];
  wire [511:0]  dataGroup_lo_740 = {dataGroup_lo_hi_740, dataGroup_lo_lo_740};
  wire [511:0]  dataGroup_hi_740 = {dataGroup_hi_hi_740, dataGroup_hi_lo_740};
  wire [15:0]   dataGroup_4_56 = dataGroup_lo_740[479:464];
  wire [511:0]  dataGroup_lo_741 = {dataGroup_lo_hi_741, dataGroup_lo_lo_741};
  wire [511:0]  dataGroup_hi_741 = {dataGroup_hi_hi_741, dataGroup_hi_lo_741};
  wire [15:0]   dataGroup_5_56 = dataGroup_hi_741[63:48];
  wire [511:0]  dataGroup_lo_742 = {dataGroup_lo_hi_742, dataGroup_lo_lo_742};
  wire [511:0]  dataGroup_hi_742 = {dataGroup_hi_hi_742, dataGroup_hi_lo_742};
  wire [15:0]   dataGroup_6_56 = dataGroup_hi_742[159:144];
  wire [511:0]  dataGroup_lo_743 = {dataGroup_lo_hi_743, dataGroup_lo_lo_743};
  wire [511:0]  dataGroup_hi_743 = {dataGroup_hi_hi_743, dataGroup_hi_lo_743};
  wire [15:0]   dataGroup_7_56 = dataGroup_hi_743[255:240];
  wire [31:0]   res_lo_lo_56 = {dataGroup_1_56, dataGroup_0_56};
  wire [31:0]   res_lo_hi_56 = {dataGroup_3_56, dataGroup_2_56};
  wire [63:0]   res_lo_56 = {res_lo_hi_56, res_lo_lo_56};
  wire [31:0]   res_hi_lo_56 = {dataGroup_5_56, dataGroup_4_56};
  wire [31:0]   res_hi_hi_56 = {dataGroup_7_56, dataGroup_6_56};
  wire [63:0]   res_hi_56 = {res_hi_hi_56, res_hi_lo_56};
  wire [127:0]  res_109 = {res_hi_56, res_lo_56};
  wire [255:0]  lo_lo_13 = {res_105, res_104};
  wire [255:0]  lo_hi_13 = {res_107, res_106};
  wire [511:0]  lo_13 = {lo_hi_13, lo_lo_13};
  wire [255:0]  hi_lo_13 = {res_109, res_108};
  wire [511:0]  hi_13 = {256'h0, hi_lo_13};
  wire [1023:0] regroupLoadData_1_5 = {hi_13, lo_13};
  wire [511:0]  dataGroup_lo_744 = {dataGroup_lo_hi_744, dataGroup_lo_lo_744};
  wire [511:0]  dataGroup_hi_744 = {dataGroup_hi_hi_744, dataGroup_hi_lo_744};
  wire [15:0]   dataGroup_0_57 = dataGroup_lo_744[15:0];
  wire [511:0]  dataGroup_lo_745 = {dataGroup_lo_hi_745, dataGroup_lo_lo_745};
  wire [511:0]  dataGroup_hi_745 = {dataGroup_hi_hi_745, dataGroup_hi_lo_745};
  wire [15:0]   dataGroup_1_57 = dataGroup_lo_745[127:112];
  wire [511:0]  dataGroup_lo_746 = {dataGroup_lo_hi_746, dataGroup_lo_lo_746};
  wire [511:0]  dataGroup_hi_746 = {dataGroup_hi_hi_746, dataGroup_hi_lo_746};
  wire [15:0]   dataGroup_2_57 = dataGroup_lo_746[239:224];
  wire [511:0]  dataGroup_lo_747 = {dataGroup_lo_hi_747, dataGroup_lo_lo_747};
  wire [511:0]  dataGroup_hi_747 = {dataGroup_hi_hi_747, dataGroup_hi_lo_747};
  wire [15:0]   dataGroup_3_57 = dataGroup_lo_747[351:336];
  wire [511:0]  dataGroup_lo_748 = {dataGroup_lo_hi_748, dataGroup_lo_lo_748};
  wire [511:0]  dataGroup_hi_748 = {dataGroup_hi_hi_748, dataGroup_hi_lo_748};
  wire [15:0]   dataGroup_4_57 = dataGroup_lo_748[463:448];
  wire [511:0]  dataGroup_lo_749 = {dataGroup_lo_hi_749, dataGroup_lo_lo_749};
  wire [511:0]  dataGroup_hi_749 = {dataGroup_hi_hi_749, dataGroup_hi_lo_749};
  wire [15:0]   dataGroup_5_57 = dataGroup_hi_749[63:48];
  wire [511:0]  dataGroup_lo_750 = {dataGroup_lo_hi_750, dataGroup_lo_lo_750};
  wire [511:0]  dataGroup_hi_750 = {dataGroup_hi_hi_750, dataGroup_hi_lo_750};
  wire [15:0]   dataGroup_6_57 = dataGroup_hi_750[175:160];
  wire [511:0]  dataGroup_lo_751 = {dataGroup_lo_hi_751, dataGroup_lo_lo_751};
  wire [511:0]  dataGroup_hi_751 = {dataGroup_hi_hi_751, dataGroup_hi_lo_751};
  wire [15:0]   dataGroup_7_57 = dataGroup_hi_751[287:272];
  wire [31:0]   res_lo_lo_57 = {dataGroup_1_57, dataGroup_0_57};
  wire [31:0]   res_lo_hi_57 = {dataGroup_3_57, dataGroup_2_57};
  wire [63:0]   res_lo_57 = {res_lo_hi_57, res_lo_lo_57};
  wire [31:0]   res_hi_lo_57 = {dataGroup_5_57, dataGroup_4_57};
  wire [31:0]   res_hi_hi_57 = {dataGroup_7_57, dataGroup_6_57};
  wire [63:0]   res_hi_57 = {res_hi_hi_57, res_hi_lo_57};
  wire [127:0]  res_112 = {res_hi_57, res_lo_57};
  wire [511:0]  dataGroup_lo_752 = {dataGroup_lo_hi_752, dataGroup_lo_lo_752};
  wire [511:0]  dataGroup_hi_752 = {dataGroup_hi_hi_752, dataGroup_hi_lo_752};
  wire [15:0]   dataGroup_0_58 = dataGroup_lo_752[31:16];
  wire [511:0]  dataGroup_lo_753 = {dataGroup_lo_hi_753, dataGroup_lo_lo_753};
  wire [511:0]  dataGroup_hi_753 = {dataGroup_hi_hi_753, dataGroup_hi_lo_753};
  wire [15:0]   dataGroup_1_58 = dataGroup_lo_753[143:128];
  wire [511:0]  dataGroup_lo_754 = {dataGroup_lo_hi_754, dataGroup_lo_lo_754};
  wire [511:0]  dataGroup_hi_754 = {dataGroup_hi_hi_754, dataGroup_hi_lo_754};
  wire [15:0]   dataGroup_2_58 = dataGroup_lo_754[255:240];
  wire [511:0]  dataGroup_lo_755 = {dataGroup_lo_hi_755, dataGroup_lo_lo_755};
  wire [511:0]  dataGroup_hi_755 = {dataGroup_hi_hi_755, dataGroup_hi_lo_755};
  wire [15:0]   dataGroup_3_58 = dataGroup_lo_755[367:352];
  wire [511:0]  dataGroup_lo_756 = {dataGroup_lo_hi_756, dataGroup_lo_lo_756};
  wire [511:0]  dataGroup_hi_756 = {dataGroup_hi_hi_756, dataGroup_hi_lo_756};
  wire [15:0]   dataGroup_4_58 = dataGroup_lo_756[479:464];
  wire [511:0]  dataGroup_lo_757 = {dataGroup_lo_hi_757, dataGroup_lo_lo_757};
  wire [511:0]  dataGroup_hi_757 = {dataGroup_hi_hi_757, dataGroup_hi_lo_757};
  wire [15:0]   dataGroup_5_58 = dataGroup_hi_757[79:64];
  wire [511:0]  dataGroup_lo_758 = {dataGroup_lo_hi_758, dataGroup_lo_lo_758};
  wire [511:0]  dataGroup_hi_758 = {dataGroup_hi_hi_758, dataGroup_hi_lo_758};
  wire [15:0]   dataGroup_6_58 = dataGroup_hi_758[191:176];
  wire [511:0]  dataGroup_lo_759 = {dataGroup_lo_hi_759, dataGroup_lo_lo_759};
  wire [511:0]  dataGroup_hi_759 = {dataGroup_hi_hi_759, dataGroup_hi_lo_759};
  wire [15:0]   dataGroup_7_58 = dataGroup_hi_759[303:288];
  wire [31:0]   res_lo_lo_58 = {dataGroup_1_58, dataGroup_0_58};
  wire [31:0]   res_lo_hi_58 = {dataGroup_3_58, dataGroup_2_58};
  wire [63:0]   res_lo_58 = {res_lo_hi_58, res_lo_lo_58};
  wire [31:0]   res_hi_lo_58 = {dataGroup_5_58, dataGroup_4_58};
  wire [31:0]   res_hi_hi_58 = {dataGroup_7_58, dataGroup_6_58};
  wire [63:0]   res_hi_58 = {res_hi_hi_58, res_hi_lo_58};
  wire [127:0]  res_113 = {res_hi_58, res_lo_58};
  wire [511:0]  dataGroup_lo_760 = {dataGroup_lo_hi_760, dataGroup_lo_lo_760};
  wire [511:0]  dataGroup_hi_760 = {dataGroup_hi_hi_760, dataGroup_hi_lo_760};
  wire [15:0]   dataGroup_0_59 = dataGroup_lo_760[47:32];
  wire [511:0]  dataGroup_lo_761 = {dataGroup_lo_hi_761, dataGroup_lo_lo_761};
  wire [511:0]  dataGroup_hi_761 = {dataGroup_hi_hi_761, dataGroup_hi_lo_761};
  wire [15:0]   dataGroup_1_59 = dataGroup_lo_761[159:144];
  wire [511:0]  dataGroup_lo_762 = {dataGroup_lo_hi_762, dataGroup_lo_lo_762};
  wire [511:0]  dataGroup_hi_762 = {dataGroup_hi_hi_762, dataGroup_hi_lo_762};
  wire [15:0]   dataGroup_2_59 = dataGroup_lo_762[271:256];
  wire [511:0]  dataGroup_lo_763 = {dataGroup_lo_hi_763, dataGroup_lo_lo_763};
  wire [511:0]  dataGroup_hi_763 = {dataGroup_hi_hi_763, dataGroup_hi_lo_763};
  wire [15:0]   dataGroup_3_59 = dataGroup_lo_763[383:368];
  wire [511:0]  dataGroup_lo_764 = {dataGroup_lo_hi_764, dataGroup_lo_lo_764};
  wire [511:0]  dataGroup_hi_764 = {dataGroup_hi_hi_764, dataGroup_hi_lo_764};
  wire [15:0]   dataGroup_4_59 = dataGroup_lo_764[495:480];
  wire [511:0]  dataGroup_lo_765 = {dataGroup_lo_hi_765, dataGroup_lo_lo_765};
  wire [511:0]  dataGroup_hi_765 = {dataGroup_hi_hi_765, dataGroup_hi_lo_765};
  wire [15:0]   dataGroup_5_59 = dataGroup_hi_765[95:80];
  wire [511:0]  dataGroup_lo_766 = {dataGroup_lo_hi_766, dataGroup_lo_lo_766};
  wire [511:0]  dataGroup_hi_766 = {dataGroup_hi_hi_766, dataGroup_hi_lo_766};
  wire [15:0]   dataGroup_6_59 = dataGroup_hi_766[207:192];
  wire [511:0]  dataGroup_lo_767 = {dataGroup_lo_hi_767, dataGroup_lo_lo_767};
  wire [511:0]  dataGroup_hi_767 = {dataGroup_hi_hi_767, dataGroup_hi_lo_767};
  wire [15:0]   dataGroup_7_59 = dataGroup_hi_767[319:304];
  wire [31:0]   res_lo_lo_59 = {dataGroup_1_59, dataGroup_0_59};
  wire [31:0]   res_lo_hi_59 = {dataGroup_3_59, dataGroup_2_59};
  wire [63:0]   res_lo_59 = {res_lo_hi_59, res_lo_lo_59};
  wire [31:0]   res_hi_lo_59 = {dataGroup_5_59, dataGroup_4_59};
  wire [31:0]   res_hi_hi_59 = {dataGroup_7_59, dataGroup_6_59};
  wire [63:0]   res_hi_59 = {res_hi_hi_59, res_hi_lo_59};
  wire [127:0]  res_114 = {res_hi_59, res_lo_59};
  wire [511:0]  dataGroup_lo_768 = {dataGroup_lo_hi_768, dataGroup_lo_lo_768};
  wire [511:0]  dataGroup_hi_768 = {dataGroup_hi_hi_768, dataGroup_hi_lo_768};
  wire [15:0]   dataGroup_0_60 = dataGroup_lo_768[63:48];
  wire [511:0]  dataGroup_lo_769 = {dataGroup_lo_hi_769, dataGroup_lo_lo_769};
  wire [511:0]  dataGroup_hi_769 = {dataGroup_hi_hi_769, dataGroup_hi_lo_769};
  wire [15:0]   dataGroup_1_60 = dataGroup_lo_769[175:160];
  wire [511:0]  dataGroup_lo_770 = {dataGroup_lo_hi_770, dataGroup_lo_lo_770};
  wire [511:0]  dataGroup_hi_770 = {dataGroup_hi_hi_770, dataGroup_hi_lo_770};
  wire [15:0]   dataGroup_2_60 = dataGroup_lo_770[287:272];
  wire [511:0]  dataGroup_lo_771 = {dataGroup_lo_hi_771, dataGroup_lo_lo_771};
  wire [511:0]  dataGroup_hi_771 = {dataGroup_hi_hi_771, dataGroup_hi_lo_771};
  wire [15:0]   dataGroup_3_60 = dataGroup_lo_771[399:384];
  wire [511:0]  dataGroup_lo_772 = {dataGroup_lo_hi_772, dataGroup_lo_lo_772};
  wire [511:0]  dataGroup_hi_772 = {dataGroup_hi_hi_772, dataGroup_hi_lo_772};
  wire [15:0]   dataGroup_4_60 = dataGroup_lo_772[511:496];
  wire [511:0]  dataGroup_lo_773 = {dataGroup_lo_hi_773, dataGroup_lo_lo_773};
  wire [511:0]  dataGroup_hi_773 = {dataGroup_hi_hi_773, dataGroup_hi_lo_773};
  wire [15:0]   dataGroup_5_60 = dataGroup_hi_773[111:96];
  wire [511:0]  dataGroup_lo_774 = {dataGroup_lo_hi_774, dataGroup_lo_lo_774};
  wire [511:0]  dataGroup_hi_774 = {dataGroup_hi_hi_774, dataGroup_hi_lo_774};
  wire [15:0]   dataGroup_6_60 = dataGroup_hi_774[223:208];
  wire [511:0]  dataGroup_lo_775 = {dataGroup_lo_hi_775, dataGroup_lo_lo_775};
  wire [511:0]  dataGroup_hi_775 = {dataGroup_hi_hi_775, dataGroup_hi_lo_775};
  wire [15:0]   dataGroup_7_60 = dataGroup_hi_775[335:320];
  wire [31:0]   res_lo_lo_60 = {dataGroup_1_60, dataGroup_0_60};
  wire [31:0]   res_lo_hi_60 = {dataGroup_3_60, dataGroup_2_60};
  wire [63:0]   res_lo_60 = {res_lo_hi_60, res_lo_lo_60};
  wire [31:0]   res_hi_lo_60 = {dataGroup_5_60, dataGroup_4_60};
  wire [31:0]   res_hi_hi_60 = {dataGroup_7_60, dataGroup_6_60};
  wire [63:0]   res_hi_60 = {res_hi_hi_60, res_hi_lo_60};
  wire [127:0]  res_115 = {res_hi_60, res_lo_60};
  wire [511:0]  dataGroup_lo_776 = {dataGroup_lo_hi_776, dataGroup_lo_lo_776};
  wire [511:0]  dataGroup_hi_776 = {dataGroup_hi_hi_776, dataGroup_hi_lo_776};
  wire [15:0]   dataGroup_0_61 = dataGroup_lo_776[79:64];
  wire [511:0]  dataGroup_lo_777 = {dataGroup_lo_hi_777, dataGroup_lo_lo_777};
  wire [511:0]  dataGroup_hi_777 = {dataGroup_hi_hi_777, dataGroup_hi_lo_777};
  wire [15:0]   dataGroup_1_61 = dataGroup_lo_777[191:176];
  wire [511:0]  dataGroup_lo_778 = {dataGroup_lo_hi_778, dataGroup_lo_lo_778};
  wire [511:0]  dataGroup_hi_778 = {dataGroup_hi_hi_778, dataGroup_hi_lo_778};
  wire [15:0]   dataGroup_2_61 = dataGroup_lo_778[303:288];
  wire [511:0]  dataGroup_lo_779 = {dataGroup_lo_hi_779, dataGroup_lo_lo_779};
  wire [511:0]  dataGroup_hi_779 = {dataGroup_hi_hi_779, dataGroup_hi_lo_779};
  wire [15:0]   dataGroup_3_61 = dataGroup_lo_779[415:400];
  wire [511:0]  dataGroup_lo_780 = {dataGroup_lo_hi_780, dataGroup_lo_lo_780};
  wire [511:0]  dataGroup_hi_780 = {dataGroup_hi_hi_780, dataGroup_hi_lo_780};
  wire [15:0]   dataGroup_4_61 = dataGroup_hi_780[15:0];
  wire [511:0]  dataGroup_lo_781 = {dataGroup_lo_hi_781, dataGroup_lo_lo_781};
  wire [511:0]  dataGroup_hi_781 = {dataGroup_hi_hi_781, dataGroup_hi_lo_781};
  wire [15:0]   dataGroup_5_61 = dataGroup_hi_781[127:112];
  wire [511:0]  dataGroup_lo_782 = {dataGroup_lo_hi_782, dataGroup_lo_lo_782};
  wire [511:0]  dataGroup_hi_782 = {dataGroup_hi_hi_782, dataGroup_hi_lo_782};
  wire [15:0]   dataGroup_6_61 = dataGroup_hi_782[239:224];
  wire [511:0]  dataGroup_lo_783 = {dataGroup_lo_hi_783, dataGroup_lo_lo_783};
  wire [511:0]  dataGroup_hi_783 = {dataGroup_hi_hi_783, dataGroup_hi_lo_783};
  wire [15:0]   dataGroup_7_61 = dataGroup_hi_783[351:336];
  wire [31:0]   res_lo_lo_61 = {dataGroup_1_61, dataGroup_0_61};
  wire [31:0]   res_lo_hi_61 = {dataGroup_3_61, dataGroup_2_61};
  wire [63:0]   res_lo_61 = {res_lo_hi_61, res_lo_lo_61};
  wire [31:0]   res_hi_lo_61 = {dataGroup_5_61, dataGroup_4_61};
  wire [31:0]   res_hi_hi_61 = {dataGroup_7_61, dataGroup_6_61};
  wire [63:0]   res_hi_61 = {res_hi_hi_61, res_hi_lo_61};
  wire [127:0]  res_116 = {res_hi_61, res_lo_61};
  wire [511:0]  dataGroup_lo_784 = {dataGroup_lo_hi_784, dataGroup_lo_lo_784};
  wire [511:0]  dataGroup_hi_784 = {dataGroup_hi_hi_784, dataGroup_hi_lo_784};
  wire [15:0]   dataGroup_0_62 = dataGroup_lo_784[95:80];
  wire [511:0]  dataGroup_lo_785 = {dataGroup_lo_hi_785, dataGroup_lo_lo_785};
  wire [511:0]  dataGroup_hi_785 = {dataGroup_hi_hi_785, dataGroup_hi_lo_785};
  wire [15:0]   dataGroup_1_62 = dataGroup_lo_785[207:192];
  wire [511:0]  dataGroup_lo_786 = {dataGroup_lo_hi_786, dataGroup_lo_lo_786};
  wire [511:0]  dataGroup_hi_786 = {dataGroup_hi_hi_786, dataGroup_hi_lo_786};
  wire [15:0]   dataGroup_2_62 = dataGroup_lo_786[319:304];
  wire [511:0]  dataGroup_lo_787 = {dataGroup_lo_hi_787, dataGroup_lo_lo_787};
  wire [511:0]  dataGroup_hi_787 = {dataGroup_hi_hi_787, dataGroup_hi_lo_787};
  wire [15:0]   dataGroup_3_62 = dataGroup_lo_787[431:416];
  wire [511:0]  dataGroup_lo_788 = {dataGroup_lo_hi_788, dataGroup_lo_lo_788};
  wire [511:0]  dataGroup_hi_788 = {dataGroup_hi_hi_788, dataGroup_hi_lo_788};
  wire [15:0]   dataGroup_4_62 = dataGroup_hi_788[31:16];
  wire [511:0]  dataGroup_lo_789 = {dataGroup_lo_hi_789, dataGroup_lo_lo_789};
  wire [511:0]  dataGroup_hi_789 = {dataGroup_hi_hi_789, dataGroup_hi_lo_789};
  wire [15:0]   dataGroup_5_62 = dataGroup_hi_789[143:128];
  wire [511:0]  dataGroup_lo_790 = {dataGroup_lo_hi_790, dataGroup_lo_lo_790};
  wire [511:0]  dataGroup_hi_790 = {dataGroup_hi_hi_790, dataGroup_hi_lo_790};
  wire [15:0]   dataGroup_6_62 = dataGroup_hi_790[255:240];
  wire [511:0]  dataGroup_lo_791 = {dataGroup_lo_hi_791, dataGroup_lo_lo_791};
  wire [511:0]  dataGroup_hi_791 = {dataGroup_hi_hi_791, dataGroup_hi_lo_791};
  wire [15:0]   dataGroup_7_62 = dataGroup_hi_791[367:352];
  wire [31:0]   res_lo_lo_62 = {dataGroup_1_62, dataGroup_0_62};
  wire [31:0]   res_lo_hi_62 = {dataGroup_3_62, dataGroup_2_62};
  wire [63:0]   res_lo_62 = {res_lo_hi_62, res_lo_lo_62};
  wire [31:0]   res_hi_lo_62 = {dataGroup_5_62, dataGroup_4_62};
  wire [31:0]   res_hi_hi_62 = {dataGroup_7_62, dataGroup_6_62};
  wire [63:0]   res_hi_62 = {res_hi_hi_62, res_hi_lo_62};
  wire [127:0]  res_117 = {res_hi_62, res_lo_62};
  wire [511:0]  dataGroup_lo_792 = {dataGroup_lo_hi_792, dataGroup_lo_lo_792};
  wire [511:0]  dataGroup_hi_792 = {dataGroup_hi_hi_792, dataGroup_hi_lo_792};
  wire [15:0]   dataGroup_0_63 = dataGroup_lo_792[111:96];
  wire [511:0]  dataGroup_lo_793 = {dataGroup_lo_hi_793, dataGroup_lo_lo_793};
  wire [511:0]  dataGroup_hi_793 = {dataGroup_hi_hi_793, dataGroup_hi_lo_793};
  wire [15:0]   dataGroup_1_63 = dataGroup_lo_793[223:208];
  wire [511:0]  dataGroup_lo_794 = {dataGroup_lo_hi_794, dataGroup_lo_lo_794};
  wire [511:0]  dataGroup_hi_794 = {dataGroup_hi_hi_794, dataGroup_hi_lo_794};
  wire [15:0]   dataGroup_2_63 = dataGroup_lo_794[335:320];
  wire [511:0]  dataGroup_lo_795 = {dataGroup_lo_hi_795, dataGroup_lo_lo_795};
  wire [511:0]  dataGroup_hi_795 = {dataGroup_hi_hi_795, dataGroup_hi_lo_795};
  wire [15:0]   dataGroup_3_63 = dataGroup_lo_795[447:432];
  wire [511:0]  dataGroup_lo_796 = {dataGroup_lo_hi_796, dataGroup_lo_lo_796};
  wire [511:0]  dataGroup_hi_796 = {dataGroup_hi_hi_796, dataGroup_hi_lo_796};
  wire [15:0]   dataGroup_4_63 = dataGroup_hi_796[47:32];
  wire [511:0]  dataGroup_lo_797 = {dataGroup_lo_hi_797, dataGroup_lo_lo_797};
  wire [511:0]  dataGroup_hi_797 = {dataGroup_hi_hi_797, dataGroup_hi_lo_797};
  wire [15:0]   dataGroup_5_63 = dataGroup_hi_797[159:144];
  wire [511:0]  dataGroup_lo_798 = {dataGroup_lo_hi_798, dataGroup_lo_lo_798};
  wire [511:0]  dataGroup_hi_798 = {dataGroup_hi_hi_798, dataGroup_hi_lo_798};
  wire [15:0]   dataGroup_6_63 = dataGroup_hi_798[271:256];
  wire [511:0]  dataGroup_lo_799 = {dataGroup_lo_hi_799, dataGroup_lo_lo_799};
  wire [511:0]  dataGroup_hi_799 = {dataGroup_hi_hi_799, dataGroup_hi_lo_799};
  wire [15:0]   dataGroup_7_63 = dataGroup_hi_799[383:368];
  wire [31:0]   res_lo_lo_63 = {dataGroup_1_63, dataGroup_0_63};
  wire [31:0]   res_lo_hi_63 = {dataGroup_3_63, dataGroup_2_63};
  wire [63:0]   res_lo_63 = {res_lo_hi_63, res_lo_lo_63};
  wire [31:0]   res_hi_lo_63 = {dataGroup_5_63, dataGroup_4_63};
  wire [31:0]   res_hi_hi_63 = {dataGroup_7_63, dataGroup_6_63};
  wire [63:0]   res_hi_63 = {res_hi_hi_63, res_hi_lo_63};
  wire [127:0]  res_118 = {res_hi_63, res_lo_63};
  wire [255:0]  lo_lo_14 = {res_113, res_112};
  wire [255:0]  lo_hi_14 = {res_115, res_114};
  wire [511:0]  lo_14 = {lo_hi_14, lo_lo_14};
  wire [255:0]  hi_lo_14 = {res_117, res_116};
  wire [255:0]  hi_hi_14 = {128'h0, res_118};
  wire [511:0]  hi_14 = {hi_hi_14, hi_lo_14};
  wire [1023:0] regroupLoadData_1_6 = {hi_14, lo_14};
  wire [511:0]  dataGroup_lo_800 = {dataGroup_lo_hi_800, dataGroup_lo_lo_800};
  wire [511:0]  dataGroup_hi_800 = {dataGroup_hi_hi_800, dataGroup_hi_lo_800};
  wire [15:0]   dataGroup_0_64 = dataGroup_lo_800[15:0];
  wire [511:0]  dataGroup_lo_801 = {dataGroup_lo_hi_801, dataGroup_lo_lo_801};
  wire [511:0]  dataGroup_hi_801 = {dataGroup_hi_hi_801, dataGroup_hi_lo_801};
  wire [15:0]   dataGroup_1_64 = dataGroup_lo_801[143:128];
  wire [511:0]  dataGroup_lo_802 = {dataGroup_lo_hi_802, dataGroup_lo_lo_802};
  wire [511:0]  dataGroup_hi_802 = {dataGroup_hi_hi_802, dataGroup_hi_lo_802};
  wire [15:0]   dataGroup_2_64 = dataGroup_lo_802[271:256];
  wire [511:0]  dataGroup_lo_803 = {dataGroup_lo_hi_803, dataGroup_lo_lo_803};
  wire [511:0]  dataGroup_hi_803 = {dataGroup_hi_hi_803, dataGroup_hi_lo_803};
  wire [15:0]   dataGroup_3_64 = dataGroup_lo_803[399:384];
  wire [511:0]  dataGroup_lo_804 = {dataGroup_lo_hi_804, dataGroup_lo_lo_804};
  wire [511:0]  dataGroup_hi_804 = {dataGroup_hi_hi_804, dataGroup_hi_lo_804};
  wire [15:0]   dataGroup_4_64 = dataGroup_hi_804[15:0];
  wire [511:0]  dataGroup_lo_805 = {dataGroup_lo_hi_805, dataGroup_lo_lo_805};
  wire [511:0]  dataGroup_hi_805 = {dataGroup_hi_hi_805, dataGroup_hi_lo_805};
  wire [15:0]   dataGroup_5_64 = dataGroup_hi_805[143:128];
  wire [511:0]  dataGroup_lo_806 = {dataGroup_lo_hi_806, dataGroup_lo_lo_806};
  wire [511:0]  dataGroup_hi_806 = {dataGroup_hi_hi_806, dataGroup_hi_lo_806};
  wire [15:0]   dataGroup_6_64 = dataGroup_hi_806[271:256];
  wire [511:0]  dataGroup_lo_807 = {dataGroup_lo_hi_807, dataGroup_lo_lo_807};
  wire [511:0]  dataGroup_hi_807 = {dataGroup_hi_hi_807, dataGroup_hi_lo_807};
  wire [15:0]   dataGroup_7_64 = dataGroup_hi_807[399:384];
  wire [31:0]   res_lo_lo_64 = {dataGroup_1_64, dataGroup_0_64};
  wire [31:0]   res_lo_hi_64 = {dataGroup_3_64, dataGroup_2_64};
  wire [63:0]   res_lo_64 = {res_lo_hi_64, res_lo_lo_64};
  wire [31:0]   res_hi_lo_64 = {dataGroup_5_64, dataGroup_4_64};
  wire [31:0]   res_hi_hi_64 = {dataGroup_7_64, dataGroup_6_64};
  wire [63:0]   res_hi_64 = {res_hi_hi_64, res_hi_lo_64};
  wire [127:0]  res_120 = {res_hi_64, res_lo_64};
  wire [511:0]  dataGroup_lo_808 = {dataGroup_lo_hi_808, dataGroup_lo_lo_808};
  wire [511:0]  dataGroup_hi_808 = {dataGroup_hi_hi_808, dataGroup_hi_lo_808};
  wire [15:0]   dataGroup_0_65 = dataGroup_lo_808[31:16];
  wire [511:0]  dataGroup_lo_809 = {dataGroup_lo_hi_809, dataGroup_lo_lo_809};
  wire [511:0]  dataGroup_hi_809 = {dataGroup_hi_hi_809, dataGroup_hi_lo_809};
  wire [15:0]   dataGroup_1_65 = dataGroup_lo_809[159:144];
  wire [511:0]  dataGroup_lo_810 = {dataGroup_lo_hi_810, dataGroup_lo_lo_810};
  wire [511:0]  dataGroup_hi_810 = {dataGroup_hi_hi_810, dataGroup_hi_lo_810};
  wire [15:0]   dataGroup_2_65 = dataGroup_lo_810[287:272];
  wire [511:0]  dataGroup_lo_811 = {dataGroup_lo_hi_811, dataGroup_lo_lo_811};
  wire [511:0]  dataGroup_hi_811 = {dataGroup_hi_hi_811, dataGroup_hi_lo_811};
  wire [15:0]   dataGroup_3_65 = dataGroup_lo_811[415:400];
  wire [511:0]  dataGroup_lo_812 = {dataGroup_lo_hi_812, dataGroup_lo_lo_812};
  wire [511:0]  dataGroup_hi_812 = {dataGroup_hi_hi_812, dataGroup_hi_lo_812};
  wire [15:0]   dataGroup_4_65 = dataGroup_hi_812[31:16];
  wire [511:0]  dataGroup_lo_813 = {dataGroup_lo_hi_813, dataGroup_lo_lo_813};
  wire [511:0]  dataGroup_hi_813 = {dataGroup_hi_hi_813, dataGroup_hi_lo_813};
  wire [15:0]   dataGroup_5_65 = dataGroup_hi_813[159:144];
  wire [511:0]  dataGroup_lo_814 = {dataGroup_lo_hi_814, dataGroup_lo_lo_814};
  wire [511:0]  dataGroup_hi_814 = {dataGroup_hi_hi_814, dataGroup_hi_lo_814};
  wire [15:0]   dataGroup_6_65 = dataGroup_hi_814[287:272];
  wire [511:0]  dataGroup_lo_815 = {dataGroup_lo_hi_815, dataGroup_lo_lo_815};
  wire [511:0]  dataGroup_hi_815 = {dataGroup_hi_hi_815, dataGroup_hi_lo_815};
  wire [15:0]   dataGroup_7_65 = dataGroup_hi_815[415:400];
  wire [31:0]   res_lo_lo_65 = {dataGroup_1_65, dataGroup_0_65};
  wire [31:0]   res_lo_hi_65 = {dataGroup_3_65, dataGroup_2_65};
  wire [63:0]   res_lo_65 = {res_lo_hi_65, res_lo_lo_65};
  wire [31:0]   res_hi_lo_65 = {dataGroup_5_65, dataGroup_4_65};
  wire [31:0]   res_hi_hi_65 = {dataGroup_7_65, dataGroup_6_65};
  wire [63:0]   res_hi_65 = {res_hi_hi_65, res_hi_lo_65};
  wire [127:0]  res_121 = {res_hi_65, res_lo_65};
  wire [511:0]  dataGroup_lo_816 = {dataGroup_lo_hi_816, dataGroup_lo_lo_816};
  wire [511:0]  dataGroup_hi_816 = {dataGroup_hi_hi_816, dataGroup_hi_lo_816};
  wire [15:0]   dataGroup_0_66 = dataGroup_lo_816[47:32];
  wire [511:0]  dataGroup_lo_817 = {dataGroup_lo_hi_817, dataGroup_lo_lo_817};
  wire [511:0]  dataGroup_hi_817 = {dataGroup_hi_hi_817, dataGroup_hi_lo_817};
  wire [15:0]   dataGroup_1_66 = dataGroup_lo_817[175:160];
  wire [511:0]  dataGroup_lo_818 = {dataGroup_lo_hi_818, dataGroup_lo_lo_818};
  wire [511:0]  dataGroup_hi_818 = {dataGroup_hi_hi_818, dataGroup_hi_lo_818};
  wire [15:0]   dataGroup_2_66 = dataGroup_lo_818[303:288];
  wire [511:0]  dataGroup_lo_819 = {dataGroup_lo_hi_819, dataGroup_lo_lo_819};
  wire [511:0]  dataGroup_hi_819 = {dataGroup_hi_hi_819, dataGroup_hi_lo_819};
  wire [15:0]   dataGroup_3_66 = dataGroup_lo_819[431:416];
  wire [511:0]  dataGroup_lo_820 = {dataGroup_lo_hi_820, dataGroup_lo_lo_820};
  wire [511:0]  dataGroup_hi_820 = {dataGroup_hi_hi_820, dataGroup_hi_lo_820};
  wire [15:0]   dataGroup_4_66 = dataGroup_hi_820[47:32];
  wire [511:0]  dataGroup_lo_821 = {dataGroup_lo_hi_821, dataGroup_lo_lo_821};
  wire [511:0]  dataGroup_hi_821 = {dataGroup_hi_hi_821, dataGroup_hi_lo_821};
  wire [15:0]   dataGroup_5_66 = dataGroup_hi_821[175:160];
  wire [511:0]  dataGroup_lo_822 = {dataGroup_lo_hi_822, dataGroup_lo_lo_822};
  wire [511:0]  dataGroup_hi_822 = {dataGroup_hi_hi_822, dataGroup_hi_lo_822};
  wire [15:0]   dataGroup_6_66 = dataGroup_hi_822[303:288];
  wire [511:0]  dataGroup_lo_823 = {dataGroup_lo_hi_823, dataGroup_lo_lo_823};
  wire [511:0]  dataGroup_hi_823 = {dataGroup_hi_hi_823, dataGroup_hi_lo_823};
  wire [15:0]   dataGroup_7_66 = dataGroup_hi_823[431:416];
  wire [31:0]   res_lo_lo_66 = {dataGroup_1_66, dataGroup_0_66};
  wire [31:0]   res_lo_hi_66 = {dataGroup_3_66, dataGroup_2_66};
  wire [63:0]   res_lo_66 = {res_lo_hi_66, res_lo_lo_66};
  wire [31:0]   res_hi_lo_66 = {dataGroup_5_66, dataGroup_4_66};
  wire [31:0]   res_hi_hi_66 = {dataGroup_7_66, dataGroup_6_66};
  wire [63:0]   res_hi_66 = {res_hi_hi_66, res_hi_lo_66};
  wire [127:0]  res_122 = {res_hi_66, res_lo_66};
  wire [511:0]  dataGroup_lo_824 = {dataGroup_lo_hi_824, dataGroup_lo_lo_824};
  wire [511:0]  dataGroup_hi_824 = {dataGroup_hi_hi_824, dataGroup_hi_lo_824};
  wire [15:0]   dataGroup_0_67 = dataGroup_lo_824[63:48];
  wire [511:0]  dataGroup_lo_825 = {dataGroup_lo_hi_825, dataGroup_lo_lo_825};
  wire [511:0]  dataGroup_hi_825 = {dataGroup_hi_hi_825, dataGroup_hi_lo_825};
  wire [15:0]   dataGroup_1_67 = dataGroup_lo_825[191:176];
  wire [511:0]  dataGroup_lo_826 = {dataGroup_lo_hi_826, dataGroup_lo_lo_826};
  wire [511:0]  dataGroup_hi_826 = {dataGroup_hi_hi_826, dataGroup_hi_lo_826};
  wire [15:0]   dataGroup_2_67 = dataGroup_lo_826[319:304];
  wire [511:0]  dataGroup_lo_827 = {dataGroup_lo_hi_827, dataGroup_lo_lo_827};
  wire [511:0]  dataGroup_hi_827 = {dataGroup_hi_hi_827, dataGroup_hi_lo_827};
  wire [15:0]   dataGroup_3_67 = dataGroup_lo_827[447:432];
  wire [511:0]  dataGroup_lo_828 = {dataGroup_lo_hi_828, dataGroup_lo_lo_828};
  wire [511:0]  dataGroup_hi_828 = {dataGroup_hi_hi_828, dataGroup_hi_lo_828};
  wire [15:0]   dataGroup_4_67 = dataGroup_hi_828[63:48];
  wire [511:0]  dataGroup_lo_829 = {dataGroup_lo_hi_829, dataGroup_lo_lo_829};
  wire [511:0]  dataGroup_hi_829 = {dataGroup_hi_hi_829, dataGroup_hi_lo_829};
  wire [15:0]   dataGroup_5_67 = dataGroup_hi_829[191:176];
  wire [511:0]  dataGroup_lo_830 = {dataGroup_lo_hi_830, dataGroup_lo_lo_830};
  wire [511:0]  dataGroup_hi_830 = {dataGroup_hi_hi_830, dataGroup_hi_lo_830};
  wire [15:0]   dataGroup_6_67 = dataGroup_hi_830[319:304];
  wire [511:0]  dataGroup_lo_831 = {dataGroup_lo_hi_831, dataGroup_lo_lo_831};
  wire [511:0]  dataGroup_hi_831 = {dataGroup_hi_hi_831, dataGroup_hi_lo_831};
  wire [15:0]   dataGroup_7_67 = dataGroup_hi_831[447:432];
  wire [31:0]   res_lo_lo_67 = {dataGroup_1_67, dataGroup_0_67};
  wire [31:0]   res_lo_hi_67 = {dataGroup_3_67, dataGroup_2_67};
  wire [63:0]   res_lo_67 = {res_lo_hi_67, res_lo_lo_67};
  wire [31:0]   res_hi_lo_67 = {dataGroup_5_67, dataGroup_4_67};
  wire [31:0]   res_hi_hi_67 = {dataGroup_7_67, dataGroup_6_67};
  wire [63:0]   res_hi_67 = {res_hi_hi_67, res_hi_lo_67};
  wire [127:0]  res_123 = {res_hi_67, res_lo_67};
  wire [511:0]  dataGroup_lo_832 = {dataGroup_lo_hi_832, dataGroup_lo_lo_832};
  wire [511:0]  dataGroup_hi_832 = {dataGroup_hi_hi_832, dataGroup_hi_lo_832};
  wire [15:0]   dataGroup_0_68 = dataGroup_lo_832[79:64];
  wire [511:0]  dataGroup_lo_833 = {dataGroup_lo_hi_833, dataGroup_lo_lo_833};
  wire [511:0]  dataGroup_hi_833 = {dataGroup_hi_hi_833, dataGroup_hi_lo_833};
  wire [15:0]   dataGroup_1_68 = dataGroup_lo_833[207:192];
  wire [511:0]  dataGroup_lo_834 = {dataGroup_lo_hi_834, dataGroup_lo_lo_834};
  wire [511:0]  dataGroup_hi_834 = {dataGroup_hi_hi_834, dataGroup_hi_lo_834};
  wire [15:0]   dataGroup_2_68 = dataGroup_lo_834[335:320];
  wire [511:0]  dataGroup_lo_835 = {dataGroup_lo_hi_835, dataGroup_lo_lo_835};
  wire [511:0]  dataGroup_hi_835 = {dataGroup_hi_hi_835, dataGroup_hi_lo_835};
  wire [15:0]   dataGroup_3_68 = dataGroup_lo_835[463:448];
  wire [511:0]  dataGroup_lo_836 = {dataGroup_lo_hi_836, dataGroup_lo_lo_836};
  wire [511:0]  dataGroup_hi_836 = {dataGroup_hi_hi_836, dataGroup_hi_lo_836};
  wire [15:0]   dataGroup_4_68 = dataGroup_hi_836[79:64];
  wire [511:0]  dataGroup_lo_837 = {dataGroup_lo_hi_837, dataGroup_lo_lo_837};
  wire [511:0]  dataGroup_hi_837 = {dataGroup_hi_hi_837, dataGroup_hi_lo_837};
  wire [15:0]   dataGroup_5_68 = dataGroup_hi_837[207:192];
  wire [511:0]  dataGroup_lo_838 = {dataGroup_lo_hi_838, dataGroup_lo_lo_838};
  wire [511:0]  dataGroup_hi_838 = {dataGroup_hi_hi_838, dataGroup_hi_lo_838};
  wire [15:0]   dataGroup_6_68 = dataGroup_hi_838[335:320];
  wire [511:0]  dataGroup_lo_839 = {dataGroup_lo_hi_839, dataGroup_lo_lo_839};
  wire [511:0]  dataGroup_hi_839 = {dataGroup_hi_hi_839, dataGroup_hi_lo_839};
  wire [15:0]   dataGroup_7_68 = dataGroup_hi_839[463:448];
  wire [31:0]   res_lo_lo_68 = {dataGroup_1_68, dataGroup_0_68};
  wire [31:0]   res_lo_hi_68 = {dataGroup_3_68, dataGroup_2_68};
  wire [63:0]   res_lo_68 = {res_lo_hi_68, res_lo_lo_68};
  wire [31:0]   res_hi_lo_68 = {dataGroup_5_68, dataGroup_4_68};
  wire [31:0]   res_hi_hi_68 = {dataGroup_7_68, dataGroup_6_68};
  wire [63:0]   res_hi_68 = {res_hi_hi_68, res_hi_lo_68};
  wire [127:0]  res_124 = {res_hi_68, res_lo_68};
  wire [511:0]  dataGroup_lo_840 = {dataGroup_lo_hi_840, dataGroup_lo_lo_840};
  wire [511:0]  dataGroup_hi_840 = {dataGroup_hi_hi_840, dataGroup_hi_lo_840};
  wire [15:0]   dataGroup_0_69 = dataGroup_lo_840[95:80];
  wire [511:0]  dataGroup_lo_841 = {dataGroup_lo_hi_841, dataGroup_lo_lo_841};
  wire [511:0]  dataGroup_hi_841 = {dataGroup_hi_hi_841, dataGroup_hi_lo_841};
  wire [15:0]   dataGroup_1_69 = dataGroup_lo_841[223:208];
  wire [511:0]  dataGroup_lo_842 = {dataGroup_lo_hi_842, dataGroup_lo_lo_842};
  wire [511:0]  dataGroup_hi_842 = {dataGroup_hi_hi_842, dataGroup_hi_lo_842};
  wire [15:0]   dataGroup_2_69 = dataGroup_lo_842[351:336];
  wire [511:0]  dataGroup_lo_843 = {dataGroup_lo_hi_843, dataGroup_lo_lo_843};
  wire [511:0]  dataGroup_hi_843 = {dataGroup_hi_hi_843, dataGroup_hi_lo_843};
  wire [15:0]   dataGroup_3_69 = dataGroup_lo_843[479:464];
  wire [511:0]  dataGroup_lo_844 = {dataGroup_lo_hi_844, dataGroup_lo_lo_844};
  wire [511:0]  dataGroup_hi_844 = {dataGroup_hi_hi_844, dataGroup_hi_lo_844};
  wire [15:0]   dataGroup_4_69 = dataGroup_hi_844[95:80];
  wire [511:0]  dataGroup_lo_845 = {dataGroup_lo_hi_845, dataGroup_lo_lo_845};
  wire [511:0]  dataGroup_hi_845 = {dataGroup_hi_hi_845, dataGroup_hi_lo_845};
  wire [15:0]   dataGroup_5_69 = dataGroup_hi_845[223:208];
  wire [511:0]  dataGroup_lo_846 = {dataGroup_lo_hi_846, dataGroup_lo_lo_846};
  wire [511:0]  dataGroup_hi_846 = {dataGroup_hi_hi_846, dataGroup_hi_lo_846};
  wire [15:0]   dataGroup_6_69 = dataGroup_hi_846[351:336];
  wire [511:0]  dataGroup_lo_847 = {dataGroup_lo_hi_847, dataGroup_lo_lo_847};
  wire [511:0]  dataGroup_hi_847 = {dataGroup_hi_hi_847, dataGroup_hi_lo_847};
  wire [15:0]   dataGroup_7_69 = dataGroup_hi_847[479:464];
  wire [31:0]   res_lo_lo_69 = {dataGroup_1_69, dataGroup_0_69};
  wire [31:0]   res_lo_hi_69 = {dataGroup_3_69, dataGroup_2_69};
  wire [63:0]   res_lo_69 = {res_lo_hi_69, res_lo_lo_69};
  wire [31:0]   res_hi_lo_69 = {dataGroup_5_69, dataGroup_4_69};
  wire [31:0]   res_hi_hi_69 = {dataGroup_7_69, dataGroup_6_69};
  wire [63:0]   res_hi_69 = {res_hi_hi_69, res_hi_lo_69};
  wire [127:0]  res_125 = {res_hi_69, res_lo_69};
  wire [511:0]  dataGroup_lo_848 = {dataGroup_lo_hi_848, dataGroup_lo_lo_848};
  wire [511:0]  dataGroup_hi_848 = {dataGroup_hi_hi_848, dataGroup_hi_lo_848};
  wire [15:0]   dataGroup_0_70 = dataGroup_lo_848[111:96];
  wire [511:0]  dataGroup_lo_849 = {dataGroup_lo_hi_849, dataGroup_lo_lo_849};
  wire [511:0]  dataGroup_hi_849 = {dataGroup_hi_hi_849, dataGroup_hi_lo_849};
  wire [15:0]   dataGroup_1_70 = dataGroup_lo_849[239:224];
  wire [511:0]  dataGroup_lo_850 = {dataGroup_lo_hi_850, dataGroup_lo_lo_850};
  wire [511:0]  dataGroup_hi_850 = {dataGroup_hi_hi_850, dataGroup_hi_lo_850};
  wire [15:0]   dataGroup_2_70 = dataGroup_lo_850[367:352];
  wire [511:0]  dataGroup_lo_851 = {dataGroup_lo_hi_851, dataGroup_lo_lo_851};
  wire [511:0]  dataGroup_hi_851 = {dataGroup_hi_hi_851, dataGroup_hi_lo_851};
  wire [15:0]   dataGroup_3_70 = dataGroup_lo_851[495:480];
  wire [511:0]  dataGroup_lo_852 = {dataGroup_lo_hi_852, dataGroup_lo_lo_852};
  wire [511:0]  dataGroup_hi_852 = {dataGroup_hi_hi_852, dataGroup_hi_lo_852};
  wire [15:0]   dataGroup_4_70 = dataGroup_hi_852[111:96];
  wire [511:0]  dataGroup_lo_853 = {dataGroup_lo_hi_853, dataGroup_lo_lo_853};
  wire [511:0]  dataGroup_hi_853 = {dataGroup_hi_hi_853, dataGroup_hi_lo_853};
  wire [15:0]   dataGroup_5_70 = dataGroup_hi_853[239:224];
  wire [511:0]  dataGroup_lo_854 = {dataGroup_lo_hi_854, dataGroup_lo_lo_854};
  wire [511:0]  dataGroup_hi_854 = {dataGroup_hi_hi_854, dataGroup_hi_lo_854};
  wire [15:0]   dataGroup_6_70 = dataGroup_hi_854[367:352];
  wire [511:0]  dataGroup_lo_855 = {dataGroup_lo_hi_855, dataGroup_lo_lo_855};
  wire [511:0]  dataGroup_hi_855 = {dataGroup_hi_hi_855, dataGroup_hi_lo_855};
  wire [15:0]   dataGroup_7_70 = dataGroup_hi_855[495:480];
  wire [31:0]   res_lo_lo_70 = {dataGroup_1_70, dataGroup_0_70};
  wire [31:0]   res_lo_hi_70 = {dataGroup_3_70, dataGroup_2_70};
  wire [63:0]   res_lo_70 = {res_lo_hi_70, res_lo_lo_70};
  wire [31:0]   res_hi_lo_70 = {dataGroup_5_70, dataGroup_4_70};
  wire [31:0]   res_hi_hi_70 = {dataGroup_7_70, dataGroup_6_70};
  wire [63:0]   res_hi_70 = {res_hi_hi_70, res_hi_lo_70};
  wire [127:0]  res_126 = {res_hi_70, res_lo_70};
  wire [511:0]  dataGroup_lo_856 = {dataGroup_lo_hi_856, dataGroup_lo_lo_856};
  wire [511:0]  dataGroup_hi_856 = {dataGroup_hi_hi_856, dataGroup_hi_lo_856};
  wire [15:0]   dataGroup_0_71 = dataGroup_lo_856[127:112];
  wire [511:0]  dataGroup_lo_857 = {dataGroup_lo_hi_857, dataGroup_lo_lo_857};
  wire [511:0]  dataGroup_hi_857 = {dataGroup_hi_hi_857, dataGroup_hi_lo_857};
  wire [15:0]   dataGroup_1_71 = dataGroup_lo_857[255:240];
  wire [511:0]  dataGroup_lo_858 = {dataGroup_lo_hi_858, dataGroup_lo_lo_858};
  wire [511:0]  dataGroup_hi_858 = {dataGroup_hi_hi_858, dataGroup_hi_lo_858};
  wire [15:0]   dataGroup_2_71 = dataGroup_lo_858[383:368];
  wire [511:0]  dataGroup_lo_859 = {dataGroup_lo_hi_859, dataGroup_lo_lo_859};
  wire [511:0]  dataGroup_hi_859 = {dataGroup_hi_hi_859, dataGroup_hi_lo_859};
  wire [15:0]   dataGroup_3_71 = dataGroup_lo_859[511:496];
  wire [511:0]  dataGroup_lo_860 = {dataGroup_lo_hi_860, dataGroup_lo_lo_860};
  wire [511:0]  dataGroup_hi_860 = {dataGroup_hi_hi_860, dataGroup_hi_lo_860};
  wire [15:0]   dataGroup_4_71 = dataGroup_hi_860[127:112];
  wire [511:0]  dataGroup_lo_861 = {dataGroup_lo_hi_861, dataGroup_lo_lo_861};
  wire [511:0]  dataGroup_hi_861 = {dataGroup_hi_hi_861, dataGroup_hi_lo_861};
  wire [15:0]   dataGroup_5_71 = dataGroup_hi_861[255:240];
  wire [511:0]  dataGroup_lo_862 = {dataGroup_lo_hi_862, dataGroup_lo_lo_862};
  wire [511:0]  dataGroup_hi_862 = {dataGroup_hi_hi_862, dataGroup_hi_lo_862};
  wire [15:0]   dataGroup_6_71 = dataGroup_hi_862[383:368];
  wire [511:0]  dataGroup_lo_863 = {dataGroup_lo_hi_863, dataGroup_lo_lo_863};
  wire [511:0]  dataGroup_hi_863 = {dataGroup_hi_hi_863, dataGroup_hi_lo_863};
  wire [15:0]   dataGroup_7_71 = dataGroup_hi_863[511:496];
  wire [31:0]   res_lo_lo_71 = {dataGroup_1_71, dataGroup_0_71};
  wire [31:0]   res_lo_hi_71 = {dataGroup_3_71, dataGroup_2_71};
  wire [63:0]   res_lo_71 = {res_lo_hi_71, res_lo_lo_71};
  wire [31:0]   res_hi_lo_71 = {dataGroup_5_71, dataGroup_4_71};
  wire [31:0]   res_hi_hi_71 = {dataGroup_7_71, dataGroup_6_71};
  wire [63:0]   res_hi_71 = {res_hi_hi_71, res_hi_lo_71};
  wire [127:0]  res_127 = {res_hi_71, res_lo_71};
  wire [255:0]  lo_lo_15 = {res_121, res_120};
  wire [255:0]  lo_hi_15 = {res_123, res_122};
  wire [511:0]  lo_15 = {lo_hi_15, lo_lo_15};
  wire [255:0]  hi_lo_15 = {res_125, res_124};
  wire [255:0]  hi_hi_15 = {res_127, res_126};
  wire [511:0]  hi_15 = {hi_hi_15, hi_lo_15};
  wire [1023:0] regroupLoadData_1_7 = {hi_15, lo_15};
  wire [511:0]  dataGroup_lo_864 = {dataGroup_lo_hi_864, dataGroup_lo_lo_864};
  wire [511:0]  dataGroup_hi_864 = {dataGroup_hi_hi_864, dataGroup_hi_lo_864};
  wire [31:0]   dataGroup_0_72 = dataGroup_lo_864[31:0];
  wire [511:0]  dataGroup_lo_865 = {dataGroup_lo_hi_865, dataGroup_lo_lo_865};
  wire [511:0]  dataGroup_hi_865 = {dataGroup_hi_hi_865, dataGroup_hi_lo_865};
  wire [31:0]   dataGroup_1_72 = dataGroup_lo_865[63:32];
  wire [511:0]  dataGroup_lo_866 = {dataGroup_lo_hi_866, dataGroup_lo_lo_866};
  wire [511:0]  dataGroup_hi_866 = {dataGroup_hi_hi_866, dataGroup_hi_lo_866};
  wire [31:0]   dataGroup_2_72 = dataGroup_lo_866[95:64];
  wire [511:0]  dataGroup_lo_867 = {dataGroup_lo_hi_867, dataGroup_lo_lo_867};
  wire [511:0]  dataGroup_hi_867 = {dataGroup_hi_hi_867, dataGroup_hi_lo_867};
  wire [31:0]   dataGroup_3_72 = dataGroup_lo_867[127:96];
  wire [63:0]   res_lo_72 = {dataGroup_1_72, dataGroup_0_72};
  wire [63:0]   res_hi_72 = {dataGroup_3_72, dataGroup_2_72};
  wire [127:0]  res_128 = {res_hi_72, res_lo_72};
  wire [255:0]  lo_lo_16 = {128'h0, res_128};
  wire [511:0]  lo_16 = {256'h0, lo_lo_16};
  wire [1023:0] regroupLoadData_2_0 = {512'h0, lo_16};
  wire [511:0]  dataGroup_lo_868 = {dataGroup_lo_hi_868, dataGroup_lo_lo_868};
  wire [511:0]  dataGroup_hi_868 = {dataGroup_hi_hi_868, dataGroup_hi_lo_868};
  wire [31:0]   dataGroup_0_73 = dataGroup_lo_868[31:0];
  wire [511:0]  dataGroup_lo_869 = {dataGroup_lo_hi_869, dataGroup_lo_lo_869};
  wire [511:0]  dataGroup_hi_869 = {dataGroup_hi_hi_869, dataGroup_hi_lo_869};
  wire [31:0]   dataGroup_1_73 = dataGroup_lo_869[95:64];
  wire [511:0]  dataGroup_lo_870 = {dataGroup_lo_hi_870, dataGroup_lo_lo_870};
  wire [511:0]  dataGroup_hi_870 = {dataGroup_hi_hi_870, dataGroup_hi_lo_870};
  wire [31:0]   dataGroup_2_73 = dataGroup_lo_870[159:128];
  wire [511:0]  dataGroup_lo_871 = {dataGroup_lo_hi_871, dataGroup_lo_lo_871};
  wire [511:0]  dataGroup_hi_871 = {dataGroup_hi_hi_871, dataGroup_hi_lo_871};
  wire [31:0]   dataGroup_3_73 = dataGroup_lo_871[223:192];
  wire [63:0]   res_lo_73 = {dataGroup_1_73, dataGroup_0_73};
  wire [63:0]   res_hi_73 = {dataGroup_3_73, dataGroup_2_73};
  wire [127:0]  res_136 = {res_hi_73, res_lo_73};
  wire [511:0]  dataGroup_lo_872 = {dataGroup_lo_hi_872, dataGroup_lo_lo_872};
  wire [511:0]  dataGroup_hi_872 = {dataGroup_hi_hi_872, dataGroup_hi_lo_872};
  wire [31:0]   dataGroup_0_74 = dataGroup_lo_872[63:32];
  wire [511:0]  dataGroup_lo_873 = {dataGroup_lo_hi_873, dataGroup_lo_lo_873};
  wire [511:0]  dataGroup_hi_873 = {dataGroup_hi_hi_873, dataGroup_hi_lo_873};
  wire [31:0]   dataGroup_1_74 = dataGroup_lo_873[127:96];
  wire [511:0]  dataGroup_lo_874 = {dataGroup_lo_hi_874, dataGroup_lo_lo_874};
  wire [511:0]  dataGroup_hi_874 = {dataGroup_hi_hi_874, dataGroup_hi_lo_874};
  wire [31:0]   dataGroup_2_74 = dataGroup_lo_874[191:160];
  wire [511:0]  dataGroup_lo_875 = {dataGroup_lo_hi_875, dataGroup_lo_lo_875};
  wire [511:0]  dataGroup_hi_875 = {dataGroup_hi_hi_875, dataGroup_hi_lo_875};
  wire [31:0]   dataGroup_3_74 = dataGroup_lo_875[255:224];
  wire [63:0]   res_lo_74 = {dataGroup_1_74, dataGroup_0_74};
  wire [63:0]   res_hi_74 = {dataGroup_3_74, dataGroup_2_74};
  wire [127:0]  res_137 = {res_hi_74, res_lo_74};
  wire [255:0]  lo_lo_17 = {res_137, res_136};
  wire [511:0]  lo_17 = {256'h0, lo_lo_17};
  wire [1023:0] regroupLoadData_2_1 = {512'h0, lo_17};
  wire [511:0]  dataGroup_lo_876 = {dataGroup_lo_hi_876, dataGroup_lo_lo_876};
  wire [511:0]  dataGroup_hi_876 = {dataGroup_hi_hi_876, dataGroup_hi_lo_876};
  wire [31:0]   dataGroup_0_75 = dataGroup_lo_876[31:0];
  wire [511:0]  dataGroup_lo_877 = {dataGroup_lo_hi_877, dataGroup_lo_lo_877};
  wire [511:0]  dataGroup_hi_877 = {dataGroup_hi_hi_877, dataGroup_hi_lo_877};
  wire [31:0]   dataGroup_1_75 = dataGroup_lo_877[127:96];
  wire [511:0]  dataGroup_lo_878 = {dataGroup_lo_hi_878, dataGroup_lo_lo_878};
  wire [511:0]  dataGroup_hi_878 = {dataGroup_hi_hi_878, dataGroup_hi_lo_878};
  wire [31:0]   dataGroup_2_75 = dataGroup_lo_878[223:192];
  wire [511:0]  dataGroup_lo_879 = {dataGroup_lo_hi_879, dataGroup_lo_lo_879};
  wire [511:0]  dataGroup_hi_879 = {dataGroup_hi_hi_879, dataGroup_hi_lo_879};
  wire [31:0]   dataGroup_3_75 = dataGroup_lo_879[319:288];
  wire [63:0]   res_lo_75 = {dataGroup_1_75, dataGroup_0_75};
  wire [63:0]   res_hi_75 = {dataGroup_3_75, dataGroup_2_75};
  wire [127:0]  res_144 = {res_hi_75, res_lo_75};
  wire [511:0]  dataGroup_lo_880 = {dataGroup_lo_hi_880, dataGroup_lo_lo_880};
  wire [511:0]  dataGroup_hi_880 = {dataGroup_hi_hi_880, dataGroup_hi_lo_880};
  wire [31:0]   dataGroup_0_76 = dataGroup_lo_880[63:32];
  wire [511:0]  dataGroup_lo_881 = {dataGroup_lo_hi_881, dataGroup_lo_lo_881};
  wire [511:0]  dataGroup_hi_881 = {dataGroup_hi_hi_881, dataGroup_hi_lo_881};
  wire [31:0]   dataGroup_1_76 = dataGroup_lo_881[159:128];
  wire [511:0]  dataGroup_lo_882 = {dataGroup_lo_hi_882, dataGroup_lo_lo_882};
  wire [511:0]  dataGroup_hi_882 = {dataGroup_hi_hi_882, dataGroup_hi_lo_882};
  wire [31:0]   dataGroup_2_76 = dataGroup_lo_882[255:224];
  wire [511:0]  dataGroup_lo_883 = {dataGroup_lo_hi_883, dataGroup_lo_lo_883};
  wire [511:0]  dataGroup_hi_883 = {dataGroup_hi_hi_883, dataGroup_hi_lo_883};
  wire [31:0]   dataGroup_3_76 = dataGroup_lo_883[351:320];
  wire [63:0]   res_lo_76 = {dataGroup_1_76, dataGroup_0_76};
  wire [63:0]   res_hi_76 = {dataGroup_3_76, dataGroup_2_76};
  wire [127:0]  res_145 = {res_hi_76, res_lo_76};
  wire [511:0]  dataGroup_lo_884 = {dataGroup_lo_hi_884, dataGroup_lo_lo_884};
  wire [511:0]  dataGroup_hi_884 = {dataGroup_hi_hi_884, dataGroup_hi_lo_884};
  wire [31:0]   dataGroup_0_77 = dataGroup_lo_884[95:64];
  wire [511:0]  dataGroup_lo_885 = {dataGroup_lo_hi_885, dataGroup_lo_lo_885};
  wire [511:0]  dataGroup_hi_885 = {dataGroup_hi_hi_885, dataGroup_hi_lo_885};
  wire [31:0]   dataGroup_1_77 = dataGroup_lo_885[191:160];
  wire [511:0]  dataGroup_lo_886 = {dataGroup_lo_hi_886, dataGroup_lo_lo_886};
  wire [511:0]  dataGroup_hi_886 = {dataGroup_hi_hi_886, dataGroup_hi_lo_886};
  wire [31:0]   dataGroup_2_77 = dataGroup_lo_886[287:256];
  wire [511:0]  dataGroup_lo_887 = {dataGroup_lo_hi_887, dataGroup_lo_lo_887};
  wire [511:0]  dataGroup_hi_887 = {dataGroup_hi_hi_887, dataGroup_hi_lo_887};
  wire [31:0]   dataGroup_3_77 = dataGroup_lo_887[383:352];
  wire [63:0]   res_lo_77 = {dataGroup_1_77, dataGroup_0_77};
  wire [63:0]   res_hi_77 = {dataGroup_3_77, dataGroup_2_77};
  wire [127:0]  res_146 = {res_hi_77, res_lo_77};
  wire [255:0]  lo_lo_18 = {res_145, res_144};
  wire [255:0]  lo_hi_18 = {128'h0, res_146};
  wire [511:0]  lo_18 = {lo_hi_18, lo_lo_18};
  wire [1023:0] regroupLoadData_2_2 = {512'h0, lo_18};
  wire [511:0]  dataGroup_lo_888 = {dataGroup_lo_hi_888, dataGroup_lo_lo_888};
  wire [511:0]  dataGroup_hi_888 = {dataGroup_hi_hi_888, dataGroup_hi_lo_888};
  wire [31:0]   dataGroup_0_78 = dataGroup_lo_888[31:0];
  wire [511:0]  dataGroup_lo_889 = {dataGroup_lo_hi_889, dataGroup_lo_lo_889};
  wire [511:0]  dataGroup_hi_889 = {dataGroup_hi_hi_889, dataGroup_hi_lo_889};
  wire [31:0]   dataGroup_1_78 = dataGroup_lo_889[159:128];
  wire [511:0]  dataGroup_lo_890 = {dataGroup_lo_hi_890, dataGroup_lo_lo_890};
  wire [511:0]  dataGroup_hi_890 = {dataGroup_hi_hi_890, dataGroup_hi_lo_890};
  wire [31:0]   dataGroup_2_78 = dataGroup_lo_890[287:256];
  wire [511:0]  dataGroup_lo_891 = {dataGroup_lo_hi_891, dataGroup_lo_lo_891};
  wire [511:0]  dataGroup_hi_891 = {dataGroup_hi_hi_891, dataGroup_hi_lo_891};
  wire [31:0]   dataGroup_3_78 = dataGroup_lo_891[415:384];
  wire [63:0]   res_lo_78 = {dataGroup_1_78, dataGroup_0_78};
  wire [63:0]   res_hi_78 = {dataGroup_3_78, dataGroup_2_78};
  wire [127:0]  res_152 = {res_hi_78, res_lo_78};
  wire [511:0]  dataGroup_lo_892 = {dataGroup_lo_hi_892, dataGroup_lo_lo_892};
  wire [511:0]  dataGroup_hi_892 = {dataGroup_hi_hi_892, dataGroup_hi_lo_892};
  wire [31:0]   dataGroup_0_79 = dataGroup_lo_892[63:32];
  wire [511:0]  dataGroup_lo_893 = {dataGroup_lo_hi_893, dataGroup_lo_lo_893};
  wire [511:0]  dataGroup_hi_893 = {dataGroup_hi_hi_893, dataGroup_hi_lo_893};
  wire [31:0]   dataGroup_1_79 = dataGroup_lo_893[191:160];
  wire [511:0]  dataGroup_lo_894 = {dataGroup_lo_hi_894, dataGroup_lo_lo_894};
  wire [511:0]  dataGroup_hi_894 = {dataGroup_hi_hi_894, dataGroup_hi_lo_894};
  wire [31:0]   dataGroup_2_79 = dataGroup_lo_894[319:288];
  wire [511:0]  dataGroup_lo_895 = {dataGroup_lo_hi_895, dataGroup_lo_lo_895};
  wire [511:0]  dataGroup_hi_895 = {dataGroup_hi_hi_895, dataGroup_hi_lo_895};
  wire [31:0]   dataGroup_3_79 = dataGroup_lo_895[447:416];
  wire [63:0]   res_lo_79 = {dataGroup_1_79, dataGroup_0_79};
  wire [63:0]   res_hi_79 = {dataGroup_3_79, dataGroup_2_79};
  wire [127:0]  res_153 = {res_hi_79, res_lo_79};
  wire [511:0]  dataGroup_lo_896 = {dataGroup_lo_hi_896, dataGroup_lo_lo_896};
  wire [511:0]  dataGroup_hi_896 = {dataGroup_hi_hi_896, dataGroup_hi_lo_896};
  wire [31:0]   dataGroup_0_80 = dataGroup_lo_896[95:64];
  wire [511:0]  dataGroup_lo_897 = {dataGroup_lo_hi_897, dataGroup_lo_lo_897};
  wire [511:0]  dataGroup_hi_897 = {dataGroup_hi_hi_897, dataGroup_hi_lo_897};
  wire [31:0]   dataGroup_1_80 = dataGroup_lo_897[223:192];
  wire [511:0]  dataGroup_lo_898 = {dataGroup_lo_hi_898, dataGroup_lo_lo_898};
  wire [511:0]  dataGroup_hi_898 = {dataGroup_hi_hi_898, dataGroup_hi_lo_898};
  wire [31:0]   dataGroup_2_80 = dataGroup_lo_898[351:320];
  wire [511:0]  dataGroup_lo_899 = {dataGroup_lo_hi_899, dataGroup_lo_lo_899};
  wire [511:0]  dataGroup_hi_899 = {dataGroup_hi_hi_899, dataGroup_hi_lo_899};
  wire [31:0]   dataGroup_3_80 = dataGroup_lo_899[479:448];
  wire [63:0]   res_lo_80 = {dataGroup_1_80, dataGroup_0_80};
  wire [63:0]   res_hi_80 = {dataGroup_3_80, dataGroup_2_80};
  wire [127:0]  res_154 = {res_hi_80, res_lo_80};
  wire [511:0]  dataGroup_lo_900 = {dataGroup_lo_hi_900, dataGroup_lo_lo_900};
  wire [511:0]  dataGroup_hi_900 = {dataGroup_hi_hi_900, dataGroup_hi_lo_900};
  wire [31:0]   dataGroup_0_81 = dataGroup_lo_900[127:96];
  wire [511:0]  dataGroup_lo_901 = {dataGroup_lo_hi_901, dataGroup_lo_lo_901};
  wire [511:0]  dataGroup_hi_901 = {dataGroup_hi_hi_901, dataGroup_hi_lo_901};
  wire [31:0]   dataGroup_1_81 = dataGroup_lo_901[255:224];
  wire [511:0]  dataGroup_lo_902 = {dataGroup_lo_hi_902, dataGroup_lo_lo_902};
  wire [511:0]  dataGroup_hi_902 = {dataGroup_hi_hi_902, dataGroup_hi_lo_902};
  wire [31:0]   dataGroup_2_81 = dataGroup_lo_902[383:352];
  wire [511:0]  dataGroup_lo_903 = {dataGroup_lo_hi_903, dataGroup_lo_lo_903};
  wire [511:0]  dataGroup_hi_903 = {dataGroup_hi_hi_903, dataGroup_hi_lo_903};
  wire [31:0]   dataGroup_3_81 = dataGroup_lo_903[511:480];
  wire [63:0]   res_lo_81 = {dataGroup_1_81, dataGroup_0_81};
  wire [63:0]   res_hi_81 = {dataGroup_3_81, dataGroup_2_81};
  wire [127:0]  res_155 = {res_hi_81, res_lo_81};
  wire [255:0]  lo_lo_19 = {res_153, res_152};
  wire [255:0]  lo_hi_19 = {res_155, res_154};
  wire [511:0]  lo_19 = {lo_hi_19, lo_lo_19};
  wire [1023:0] regroupLoadData_2_3 = {512'h0, lo_19};
  wire [511:0]  dataGroup_lo_904 = {dataGroup_lo_hi_904, dataGroup_lo_lo_904};
  wire [511:0]  dataGroup_hi_904 = {dataGroup_hi_hi_904, dataGroup_hi_lo_904};
  wire [31:0]   dataGroup_0_82 = dataGroup_lo_904[31:0];
  wire [511:0]  dataGroup_lo_905 = {dataGroup_lo_hi_905, dataGroup_lo_lo_905};
  wire [511:0]  dataGroup_hi_905 = {dataGroup_hi_hi_905, dataGroup_hi_lo_905};
  wire [31:0]   dataGroup_1_82 = dataGroup_lo_905[191:160];
  wire [511:0]  dataGroup_lo_906 = {dataGroup_lo_hi_906, dataGroup_lo_lo_906};
  wire [511:0]  dataGroup_hi_906 = {dataGroup_hi_hi_906, dataGroup_hi_lo_906};
  wire [31:0]   dataGroup_2_82 = dataGroup_lo_906[351:320];
  wire [511:0]  dataGroup_lo_907 = {dataGroup_lo_hi_907, dataGroup_lo_lo_907};
  wire [511:0]  dataGroup_hi_907 = {dataGroup_hi_hi_907, dataGroup_hi_lo_907};
  wire [31:0]   dataGroup_3_82 = dataGroup_lo_907[511:480];
  wire [63:0]   res_lo_82 = {dataGroup_1_82, dataGroup_0_82};
  wire [63:0]   res_hi_82 = {dataGroup_3_82, dataGroup_2_82};
  wire [127:0]  res_160 = {res_hi_82, res_lo_82};
  wire [511:0]  dataGroup_lo_908 = {dataGroup_lo_hi_908, dataGroup_lo_lo_908};
  wire [511:0]  dataGroup_hi_908 = {dataGroup_hi_hi_908, dataGroup_hi_lo_908};
  wire [31:0]   dataGroup_0_83 = dataGroup_lo_908[63:32];
  wire [511:0]  dataGroup_lo_909 = {dataGroup_lo_hi_909, dataGroup_lo_lo_909};
  wire [511:0]  dataGroup_hi_909 = {dataGroup_hi_hi_909, dataGroup_hi_lo_909};
  wire [31:0]   dataGroup_1_83 = dataGroup_lo_909[223:192];
  wire [511:0]  dataGroup_lo_910 = {dataGroup_lo_hi_910, dataGroup_lo_lo_910};
  wire [511:0]  dataGroup_hi_910 = {dataGroup_hi_hi_910, dataGroup_hi_lo_910};
  wire [31:0]   dataGroup_2_83 = dataGroup_lo_910[383:352];
  wire [511:0]  dataGroup_lo_911 = {dataGroup_lo_hi_911, dataGroup_lo_lo_911};
  wire [511:0]  dataGroup_hi_911 = {dataGroup_hi_hi_911, dataGroup_hi_lo_911};
  wire [31:0]   dataGroup_3_83 = dataGroup_hi_911[31:0];
  wire [63:0]   res_lo_83 = {dataGroup_1_83, dataGroup_0_83};
  wire [63:0]   res_hi_83 = {dataGroup_3_83, dataGroup_2_83};
  wire [127:0]  res_161 = {res_hi_83, res_lo_83};
  wire [511:0]  dataGroup_lo_912 = {dataGroup_lo_hi_912, dataGroup_lo_lo_912};
  wire [511:0]  dataGroup_hi_912 = {dataGroup_hi_hi_912, dataGroup_hi_lo_912};
  wire [31:0]   dataGroup_0_84 = dataGroup_lo_912[95:64];
  wire [511:0]  dataGroup_lo_913 = {dataGroup_lo_hi_913, dataGroup_lo_lo_913};
  wire [511:0]  dataGroup_hi_913 = {dataGroup_hi_hi_913, dataGroup_hi_lo_913};
  wire [31:0]   dataGroup_1_84 = dataGroup_lo_913[255:224];
  wire [511:0]  dataGroup_lo_914 = {dataGroup_lo_hi_914, dataGroup_lo_lo_914};
  wire [511:0]  dataGroup_hi_914 = {dataGroup_hi_hi_914, dataGroup_hi_lo_914};
  wire [31:0]   dataGroup_2_84 = dataGroup_lo_914[415:384];
  wire [511:0]  dataGroup_lo_915 = {dataGroup_lo_hi_915, dataGroup_lo_lo_915};
  wire [511:0]  dataGroup_hi_915 = {dataGroup_hi_hi_915, dataGroup_hi_lo_915};
  wire [31:0]   dataGroup_3_84 = dataGroup_hi_915[63:32];
  wire [63:0]   res_lo_84 = {dataGroup_1_84, dataGroup_0_84};
  wire [63:0]   res_hi_84 = {dataGroup_3_84, dataGroup_2_84};
  wire [127:0]  res_162 = {res_hi_84, res_lo_84};
  wire [511:0]  dataGroup_lo_916 = {dataGroup_lo_hi_916, dataGroup_lo_lo_916};
  wire [511:0]  dataGroup_hi_916 = {dataGroup_hi_hi_916, dataGroup_hi_lo_916};
  wire [31:0]   dataGroup_0_85 = dataGroup_lo_916[127:96];
  wire [511:0]  dataGroup_lo_917 = {dataGroup_lo_hi_917, dataGroup_lo_lo_917};
  wire [511:0]  dataGroup_hi_917 = {dataGroup_hi_hi_917, dataGroup_hi_lo_917};
  wire [31:0]   dataGroup_1_85 = dataGroup_lo_917[287:256];
  wire [511:0]  dataGroup_lo_918 = {dataGroup_lo_hi_918, dataGroup_lo_lo_918};
  wire [511:0]  dataGroup_hi_918 = {dataGroup_hi_hi_918, dataGroup_hi_lo_918};
  wire [31:0]   dataGroup_2_85 = dataGroup_lo_918[447:416];
  wire [511:0]  dataGroup_lo_919 = {dataGroup_lo_hi_919, dataGroup_lo_lo_919};
  wire [511:0]  dataGroup_hi_919 = {dataGroup_hi_hi_919, dataGroup_hi_lo_919};
  wire [31:0]   dataGroup_3_85 = dataGroup_hi_919[95:64];
  wire [63:0]   res_lo_85 = {dataGroup_1_85, dataGroup_0_85};
  wire [63:0]   res_hi_85 = {dataGroup_3_85, dataGroup_2_85};
  wire [127:0]  res_163 = {res_hi_85, res_lo_85};
  wire [511:0]  dataGroup_lo_920 = {dataGroup_lo_hi_920, dataGroup_lo_lo_920};
  wire [511:0]  dataGroup_hi_920 = {dataGroup_hi_hi_920, dataGroup_hi_lo_920};
  wire [31:0]   dataGroup_0_86 = dataGroup_lo_920[159:128];
  wire [511:0]  dataGroup_lo_921 = {dataGroup_lo_hi_921, dataGroup_lo_lo_921};
  wire [511:0]  dataGroup_hi_921 = {dataGroup_hi_hi_921, dataGroup_hi_lo_921};
  wire [31:0]   dataGroup_1_86 = dataGroup_lo_921[319:288];
  wire [511:0]  dataGroup_lo_922 = {dataGroup_lo_hi_922, dataGroup_lo_lo_922};
  wire [511:0]  dataGroup_hi_922 = {dataGroup_hi_hi_922, dataGroup_hi_lo_922};
  wire [31:0]   dataGroup_2_86 = dataGroup_lo_922[479:448];
  wire [511:0]  dataGroup_lo_923 = {dataGroup_lo_hi_923, dataGroup_lo_lo_923};
  wire [511:0]  dataGroup_hi_923 = {dataGroup_hi_hi_923, dataGroup_hi_lo_923};
  wire [31:0]   dataGroup_3_86 = dataGroup_hi_923[127:96];
  wire [63:0]   res_lo_86 = {dataGroup_1_86, dataGroup_0_86};
  wire [63:0]   res_hi_86 = {dataGroup_3_86, dataGroup_2_86};
  wire [127:0]  res_164 = {res_hi_86, res_lo_86};
  wire [255:0]  lo_lo_20 = {res_161, res_160};
  wire [255:0]  lo_hi_20 = {res_163, res_162};
  wire [511:0]  lo_20 = {lo_hi_20, lo_lo_20};
  wire [255:0]  hi_lo_20 = {128'h0, res_164};
  wire [511:0]  hi_20 = {256'h0, hi_lo_20};
  wire [1023:0] regroupLoadData_2_4 = {hi_20, lo_20};
  wire [511:0]  dataGroup_lo_924 = {dataGroup_lo_hi_924, dataGroup_lo_lo_924};
  wire [511:0]  dataGroup_hi_924 = {dataGroup_hi_hi_924, dataGroup_hi_lo_924};
  wire [31:0]   dataGroup_0_87 = dataGroup_lo_924[31:0];
  wire [511:0]  dataGroup_lo_925 = {dataGroup_lo_hi_925, dataGroup_lo_lo_925};
  wire [511:0]  dataGroup_hi_925 = {dataGroup_hi_hi_925, dataGroup_hi_lo_925};
  wire [31:0]   dataGroup_1_87 = dataGroup_lo_925[223:192];
  wire [511:0]  dataGroup_lo_926 = {dataGroup_lo_hi_926, dataGroup_lo_lo_926};
  wire [511:0]  dataGroup_hi_926 = {dataGroup_hi_hi_926, dataGroup_hi_lo_926};
  wire [31:0]   dataGroup_2_87 = dataGroup_lo_926[415:384];
  wire [511:0]  dataGroup_lo_927 = {dataGroup_lo_hi_927, dataGroup_lo_lo_927};
  wire [511:0]  dataGroup_hi_927 = {dataGroup_hi_hi_927, dataGroup_hi_lo_927};
  wire [31:0]   dataGroup_3_87 = dataGroup_hi_927[95:64];
  wire [63:0]   res_lo_87 = {dataGroup_1_87, dataGroup_0_87};
  wire [63:0]   res_hi_87 = {dataGroup_3_87, dataGroup_2_87};
  wire [127:0]  res_168 = {res_hi_87, res_lo_87};
  wire [511:0]  dataGroup_lo_928 = {dataGroup_lo_hi_928, dataGroup_lo_lo_928};
  wire [511:0]  dataGroup_hi_928 = {dataGroup_hi_hi_928, dataGroup_hi_lo_928};
  wire [31:0]   dataGroup_0_88 = dataGroup_lo_928[63:32];
  wire [511:0]  dataGroup_lo_929 = {dataGroup_lo_hi_929, dataGroup_lo_lo_929};
  wire [511:0]  dataGroup_hi_929 = {dataGroup_hi_hi_929, dataGroup_hi_lo_929};
  wire [31:0]   dataGroup_1_88 = dataGroup_lo_929[255:224];
  wire [511:0]  dataGroup_lo_930 = {dataGroup_lo_hi_930, dataGroup_lo_lo_930};
  wire [511:0]  dataGroup_hi_930 = {dataGroup_hi_hi_930, dataGroup_hi_lo_930};
  wire [31:0]   dataGroup_2_88 = dataGroup_lo_930[447:416];
  wire [511:0]  dataGroup_lo_931 = {dataGroup_lo_hi_931, dataGroup_lo_lo_931};
  wire [511:0]  dataGroup_hi_931 = {dataGroup_hi_hi_931, dataGroup_hi_lo_931};
  wire [31:0]   dataGroup_3_88 = dataGroup_hi_931[127:96];
  wire [63:0]   res_lo_88 = {dataGroup_1_88, dataGroup_0_88};
  wire [63:0]   res_hi_88 = {dataGroup_3_88, dataGroup_2_88};
  wire [127:0]  res_169 = {res_hi_88, res_lo_88};
  wire [511:0]  dataGroup_lo_932 = {dataGroup_lo_hi_932, dataGroup_lo_lo_932};
  wire [511:0]  dataGroup_hi_932 = {dataGroup_hi_hi_932, dataGroup_hi_lo_932};
  wire [31:0]   dataGroup_0_89 = dataGroup_lo_932[95:64];
  wire [511:0]  dataGroup_lo_933 = {dataGroup_lo_hi_933, dataGroup_lo_lo_933};
  wire [511:0]  dataGroup_hi_933 = {dataGroup_hi_hi_933, dataGroup_hi_lo_933};
  wire [31:0]   dataGroup_1_89 = dataGroup_lo_933[287:256];
  wire [511:0]  dataGroup_lo_934 = {dataGroup_lo_hi_934, dataGroup_lo_lo_934};
  wire [511:0]  dataGroup_hi_934 = {dataGroup_hi_hi_934, dataGroup_hi_lo_934};
  wire [31:0]   dataGroup_2_89 = dataGroup_lo_934[479:448];
  wire [511:0]  dataGroup_lo_935 = {dataGroup_lo_hi_935, dataGroup_lo_lo_935};
  wire [511:0]  dataGroup_hi_935 = {dataGroup_hi_hi_935, dataGroup_hi_lo_935};
  wire [31:0]   dataGroup_3_89 = dataGroup_hi_935[159:128];
  wire [63:0]   res_lo_89 = {dataGroup_1_89, dataGroup_0_89};
  wire [63:0]   res_hi_89 = {dataGroup_3_89, dataGroup_2_89};
  wire [127:0]  res_170 = {res_hi_89, res_lo_89};
  wire [511:0]  dataGroup_lo_936 = {dataGroup_lo_hi_936, dataGroup_lo_lo_936};
  wire [511:0]  dataGroup_hi_936 = {dataGroup_hi_hi_936, dataGroup_hi_lo_936};
  wire [31:0]   dataGroup_0_90 = dataGroup_lo_936[127:96];
  wire [511:0]  dataGroup_lo_937 = {dataGroup_lo_hi_937, dataGroup_lo_lo_937};
  wire [511:0]  dataGroup_hi_937 = {dataGroup_hi_hi_937, dataGroup_hi_lo_937};
  wire [31:0]   dataGroup_1_90 = dataGroup_lo_937[319:288];
  wire [511:0]  dataGroup_lo_938 = {dataGroup_lo_hi_938, dataGroup_lo_lo_938};
  wire [511:0]  dataGroup_hi_938 = {dataGroup_hi_hi_938, dataGroup_hi_lo_938};
  wire [31:0]   dataGroup_2_90 = dataGroup_lo_938[511:480];
  wire [511:0]  dataGroup_lo_939 = {dataGroup_lo_hi_939, dataGroup_lo_lo_939};
  wire [511:0]  dataGroup_hi_939 = {dataGroup_hi_hi_939, dataGroup_hi_lo_939};
  wire [31:0]   dataGroup_3_90 = dataGroup_hi_939[191:160];
  wire [63:0]   res_lo_90 = {dataGroup_1_90, dataGroup_0_90};
  wire [63:0]   res_hi_90 = {dataGroup_3_90, dataGroup_2_90};
  wire [127:0]  res_171 = {res_hi_90, res_lo_90};
  wire [511:0]  dataGroup_lo_940 = {dataGroup_lo_hi_940, dataGroup_lo_lo_940};
  wire [511:0]  dataGroup_hi_940 = {dataGroup_hi_hi_940, dataGroup_hi_lo_940};
  wire [31:0]   dataGroup_0_91 = dataGroup_lo_940[159:128];
  wire [511:0]  dataGroup_lo_941 = {dataGroup_lo_hi_941, dataGroup_lo_lo_941};
  wire [511:0]  dataGroup_hi_941 = {dataGroup_hi_hi_941, dataGroup_hi_lo_941};
  wire [31:0]   dataGroup_1_91 = dataGroup_lo_941[351:320];
  wire [511:0]  dataGroup_lo_942 = {dataGroup_lo_hi_942, dataGroup_lo_lo_942};
  wire [511:0]  dataGroup_hi_942 = {dataGroup_hi_hi_942, dataGroup_hi_lo_942};
  wire [31:0]   dataGroup_2_91 = dataGroup_hi_942[31:0];
  wire [511:0]  dataGroup_lo_943 = {dataGroup_lo_hi_943, dataGroup_lo_lo_943};
  wire [511:0]  dataGroup_hi_943 = {dataGroup_hi_hi_943, dataGroup_hi_lo_943};
  wire [31:0]   dataGroup_3_91 = dataGroup_hi_943[223:192];
  wire [63:0]   res_lo_91 = {dataGroup_1_91, dataGroup_0_91};
  wire [63:0]   res_hi_91 = {dataGroup_3_91, dataGroup_2_91};
  wire [127:0]  res_172 = {res_hi_91, res_lo_91};
  wire [511:0]  dataGroup_lo_944 = {dataGroup_lo_hi_944, dataGroup_lo_lo_944};
  wire [511:0]  dataGroup_hi_944 = {dataGroup_hi_hi_944, dataGroup_hi_lo_944};
  wire [31:0]   dataGroup_0_92 = dataGroup_lo_944[191:160];
  wire [511:0]  dataGroup_lo_945 = {dataGroup_lo_hi_945, dataGroup_lo_lo_945};
  wire [511:0]  dataGroup_hi_945 = {dataGroup_hi_hi_945, dataGroup_hi_lo_945};
  wire [31:0]   dataGroup_1_92 = dataGroup_lo_945[383:352];
  wire [511:0]  dataGroup_lo_946 = {dataGroup_lo_hi_946, dataGroup_lo_lo_946};
  wire [511:0]  dataGroup_hi_946 = {dataGroup_hi_hi_946, dataGroup_hi_lo_946};
  wire [31:0]   dataGroup_2_92 = dataGroup_hi_946[63:32];
  wire [511:0]  dataGroup_lo_947 = {dataGroup_lo_hi_947, dataGroup_lo_lo_947};
  wire [511:0]  dataGroup_hi_947 = {dataGroup_hi_hi_947, dataGroup_hi_lo_947};
  wire [31:0]   dataGroup_3_92 = dataGroup_hi_947[255:224];
  wire [63:0]   res_lo_92 = {dataGroup_1_92, dataGroup_0_92};
  wire [63:0]   res_hi_92 = {dataGroup_3_92, dataGroup_2_92};
  wire [127:0]  res_173 = {res_hi_92, res_lo_92};
  wire [255:0]  lo_lo_21 = {res_169, res_168};
  wire [255:0]  lo_hi_21 = {res_171, res_170};
  wire [511:0]  lo_21 = {lo_hi_21, lo_lo_21};
  wire [255:0]  hi_lo_21 = {res_173, res_172};
  wire [511:0]  hi_21 = {256'h0, hi_lo_21};
  wire [1023:0] regroupLoadData_2_5 = {hi_21, lo_21};
  wire [511:0]  dataGroup_lo_948 = {dataGroup_lo_hi_948, dataGroup_lo_lo_948};
  wire [511:0]  dataGroup_hi_948 = {dataGroup_hi_hi_948, dataGroup_hi_lo_948};
  wire [31:0]   dataGroup_0_93 = dataGroup_lo_948[31:0];
  wire [511:0]  dataGroup_lo_949 = {dataGroup_lo_hi_949, dataGroup_lo_lo_949};
  wire [511:0]  dataGroup_hi_949 = {dataGroup_hi_hi_949, dataGroup_hi_lo_949};
  wire [31:0]   dataGroup_1_93 = dataGroup_lo_949[255:224];
  wire [511:0]  dataGroup_lo_950 = {dataGroup_lo_hi_950, dataGroup_lo_lo_950};
  wire [511:0]  dataGroup_hi_950 = {dataGroup_hi_hi_950, dataGroup_hi_lo_950};
  wire [31:0]   dataGroup_2_93 = dataGroup_lo_950[479:448];
  wire [511:0]  dataGroup_lo_951 = {dataGroup_lo_hi_951, dataGroup_lo_lo_951};
  wire [511:0]  dataGroup_hi_951 = {dataGroup_hi_hi_951, dataGroup_hi_lo_951};
  wire [31:0]   dataGroup_3_93 = dataGroup_hi_951[191:160];
  wire [63:0]   res_lo_93 = {dataGroup_1_93, dataGroup_0_93};
  wire [63:0]   res_hi_93 = {dataGroup_3_93, dataGroup_2_93};
  wire [127:0]  res_176 = {res_hi_93, res_lo_93};
  wire [511:0]  dataGroup_lo_952 = {dataGroup_lo_hi_952, dataGroup_lo_lo_952};
  wire [511:0]  dataGroup_hi_952 = {dataGroup_hi_hi_952, dataGroup_hi_lo_952};
  wire [31:0]   dataGroup_0_94 = dataGroup_lo_952[63:32];
  wire [511:0]  dataGroup_lo_953 = {dataGroup_lo_hi_953, dataGroup_lo_lo_953};
  wire [511:0]  dataGroup_hi_953 = {dataGroup_hi_hi_953, dataGroup_hi_lo_953};
  wire [31:0]   dataGroup_1_94 = dataGroup_lo_953[287:256];
  wire [511:0]  dataGroup_lo_954 = {dataGroup_lo_hi_954, dataGroup_lo_lo_954};
  wire [511:0]  dataGroup_hi_954 = {dataGroup_hi_hi_954, dataGroup_hi_lo_954};
  wire [31:0]   dataGroup_2_94 = dataGroup_lo_954[511:480];
  wire [511:0]  dataGroup_lo_955 = {dataGroup_lo_hi_955, dataGroup_lo_lo_955};
  wire [511:0]  dataGroup_hi_955 = {dataGroup_hi_hi_955, dataGroup_hi_lo_955};
  wire [31:0]   dataGroup_3_94 = dataGroup_hi_955[223:192];
  wire [63:0]   res_lo_94 = {dataGroup_1_94, dataGroup_0_94};
  wire [63:0]   res_hi_94 = {dataGroup_3_94, dataGroup_2_94};
  wire [127:0]  res_177 = {res_hi_94, res_lo_94};
  wire [511:0]  dataGroup_lo_956 = {dataGroup_lo_hi_956, dataGroup_lo_lo_956};
  wire [511:0]  dataGroup_hi_956 = {dataGroup_hi_hi_956, dataGroup_hi_lo_956};
  wire [31:0]   dataGroup_0_95 = dataGroup_lo_956[95:64];
  wire [511:0]  dataGroup_lo_957 = {dataGroup_lo_hi_957, dataGroup_lo_lo_957};
  wire [511:0]  dataGroup_hi_957 = {dataGroup_hi_hi_957, dataGroup_hi_lo_957};
  wire [31:0]   dataGroup_1_95 = dataGroup_lo_957[319:288];
  wire [511:0]  dataGroup_lo_958 = {dataGroup_lo_hi_958, dataGroup_lo_lo_958};
  wire [511:0]  dataGroup_hi_958 = {dataGroup_hi_hi_958, dataGroup_hi_lo_958};
  wire [31:0]   dataGroup_2_95 = dataGroup_hi_958[31:0];
  wire [511:0]  dataGroup_lo_959 = {dataGroup_lo_hi_959, dataGroup_lo_lo_959};
  wire [511:0]  dataGroup_hi_959 = {dataGroup_hi_hi_959, dataGroup_hi_lo_959};
  wire [31:0]   dataGroup_3_95 = dataGroup_hi_959[255:224];
  wire [63:0]   res_lo_95 = {dataGroup_1_95, dataGroup_0_95};
  wire [63:0]   res_hi_95 = {dataGroup_3_95, dataGroup_2_95};
  wire [127:0]  res_178 = {res_hi_95, res_lo_95};
  wire [511:0]  dataGroup_lo_960 = {dataGroup_lo_hi_960, dataGroup_lo_lo_960};
  wire [511:0]  dataGroup_hi_960 = {dataGroup_hi_hi_960, dataGroup_hi_lo_960};
  wire [31:0]   dataGroup_0_96 = dataGroup_lo_960[127:96];
  wire [511:0]  dataGroup_lo_961 = {dataGroup_lo_hi_961, dataGroup_lo_lo_961};
  wire [511:0]  dataGroup_hi_961 = {dataGroup_hi_hi_961, dataGroup_hi_lo_961};
  wire [31:0]   dataGroup_1_96 = dataGroup_lo_961[351:320];
  wire [511:0]  dataGroup_lo_962 = {dataGroup_lo_hi_962, dataGroup_lo_lo_962};
  wire [511:0]  dataGroup_hi_962 = {dataGroup_hi_hi_962, dataGroup_hi_lo_962};
  wire [31:0]   dataGroup_2_96 = dataGroup_hi_962[63:32];
  wire [511:0]  dataGroup_lo_963 = {dataGroup_lo_hi_963, dataGroup_lo_lo_963};
  wire [511:0]  dataGroup_hi_963 = {dataGroup_hi_hi_963, dataGroup_hi_lo_963};
  wire [31:0]   dataGroup_3_96 = dataGroup_hi_963[287:256];
  wire [63:0]   res_lo_96 = {dataGroup_1_96, dataGroup_0_96};
  wire [63:0]   res_hi_96 = {dataGroup_3_96, dataGroup_2_96};
  wire [127:0]  res_179 = {res_hi_96, res_lo_96};
  wire [511:0]  dataGroup_lo_964 = {dataGroup_lo_hi_964, dataGroup_lo_lo_964};
  wire [511:0]  dataGroup_hi_964 = {dataGroup_hi_hi_964, dataGroup_hi_lo_964};
  wire [31:0]   dataGroup_0_97 = dataGroup_lo_964[159:128];
  wire [511:0]  dataGroup_lo_965 = {dataGroup_lo_hi_965, dataGroup_lo_lo_965};
  wire [511:0]  dataGroup_hi_965 = {dataGroup_hi_hi_965, dataGroup_hi_lo_965};
  wire [31:0]   dataGroup_1_97 = dataGroup_lo_965[383:352];
  wire [511:0]  dataGroup_lo_966 = {dataGroup_lo_hi_966, dataGroup_lo_lo_966};
  wire [511:0]  dataGroup_hi_966 = {dataGroup_hi_hi_966, dataGroup_hi_lo_966};
  wire [31:0]   dataGroup_2_97 = dataGroup_hi_966[95:64];
  wire [511:0]  dataGroup_lo_967 = {dataGroup_lo_hi_967, dataGroup_lo_lo_967};
  wire [511:0]  dataGroup_hi_967 = {dataGroup_hi_hi_967, dataGroup_hi_lo_967};
  wire [31:0]   dataGroup_3_97 = dataGroup_hi_967[319:288];
  wire [63:0]   res_lo_97 = {dataGroup_1_97, dataGroup_0_97};
  wire [63:0]   res_hi_97 = {dataGroup_3_97, dataGroup_2_97};
  wire [127:0]  res_180 = {res_hi_97, res_lo_97};
  wire [511:0]  dataGroup_lo_968 = {dataGroup_lo_hi_968, dataGroup_lo_lo_968};
  wire [511:0]  dataGroup_hi_968 = {dataGroup_hi_hi_968, dataGroup_hi_lo_968};
  wire [31:0]   dataGroup_0_98 = dataGroup_lo_968[191:160];
  wire [511:0]  dataGroup_lo_969 = {dataGroup_lo_hi_969, dataGroup_lo_lo_969};
  wire [511:0]  dataGroup_hi_969 = {dataGroup_hi_hi_969, dataGroup_hi_lo_969};
  wire [31:0]   dataGroup_1_98 = dataGroup_lo_969[415:384];
  wire [511:0]  dataGroup_lo_970 = {dataGroup_lo_hi_970, dataGroup_lo_lo_970};
  wire [511:0]  dataGroup_hi_970 = {dataGroup_hi_hi_970, dataGroup_hi_lo_970};
  wire [31:0]   dataGroup_2_98 = dataGroup_hi_970[127:96];
  wire [511:0]  dataGroup_lo_971 = {dataGroup_lo_hi_971, dataGroup_lo_lo_971};
  wire [511:0]  dataGroup_hi_971 = {dataGroup_hi_hi_971, dataGroup_hi_lo_971};
  wire [31:0]   dataGroup_3_98 = dataGroup_hi_971[351:320];
  wire [63:0]   res_lo_98 = {dataGroup_1_98, dataGroup_0_98};
  wire [63:0]   res_hi_98 = {dataGroup_3_98, dataGroup_2_98};
  wire [127:0]  res_181 = {res_hi_98, res_lo_98};
  wire [511:0]  dataGroup_lo_972 = {dataGroup_lo_hi_972, dataGroup_lo_lo_972};
  wire [511:0]  dataGroup_hi_972 = {dataGroup_hi_hi_972, dataGroup_hi_lo_972};
  wire [31:0]   dataGroup_0_99 = dataGroup_lo_972[223:192];
  wire [511:0]  dataGroup_lo_973 = {dataGroup_lo_hi_973, dataGroup_lo_lo_973};
  wire [511:0]  dataGroup_hi_973 = {dataGroup_hi_hi_973, dataGroup_hi_lo_973};
  wire [31:0]   dataGroup_1_99 = dataGroup_lo_973[447:416];
  wire [511:0]  dataGroup_lo_974 = {dataGroup_lo_hi_974, dataGroup_lo_lo_974};
  wire [511:0]  dataGroup_hi_974 = {dataGroup_hi_hi_974, dataGroup_hi_lo_974};
  wire [31:0]   dataGroup_2_99 = dataGroup_hi_974[159:128];
  wire [511:0]  dataGroup_lo_975 = {dataGroup_lo_hi_975, dataGroup_lo_lo_975};
  wire [511:0]  dataGroup_hi_975 = {dataGroup_hi_hi_975, dataGroup_hi_lo_975};
  wire [31:0]   dataGroup_3_99 = dataGroup_hi_975[383:352];
  wire [63:0]   res_lo_99 = {dataGroup_1_99, dataGroup_0_99};
  wire [63:0]   res_hi_99 = {dataGroup_3_99, dataGroup_2_99};
  wire [127:0]  res_182 = {res_hi_99, res_lo_99};
  wire [255:0]  lo_lo_22 = {res_177, res_176};
  wire [255:0]  lo_hi_22 = {res_179, res_178};
  wire [511:0]  lo_22 = {lo_hi_22, lo_lo_22};
  wire [255:0]  hi_lo_22 = {res_181, res_180};
  wire [255:0]  hi_hi_22 = {128'h0, res_182};
  wire [511:0]  hi_22 = {hi_hi_22, hi_lo_22};
  wire [1023:0] regroupLoadData_2_6 = {hi_22, lo_22};
  wire [511:0]  dataGroup_lo_976 = {dataGroup_lo_hi_976, dataGroup_lo_lo_976};
  wire [511:0]  dataGroup_hi_976 = {dataGroup_hi_hi_976, dataGroup_hi_lo_976};
  wire [31:0]   dataGroup_0_100 = dataGroup_lo_976[31:0];
  wire [511:0]  dataGroup_lo_977 = {dataGroup_lo_hi_977, dataGroup_lo_lo_977};
  wire [511:0]  dataGroup_hi_977 = {dataGroup_hi_hi_977, dataGroup_hi_lo_977};
  wire [31:0]   dataGroup_1_100 = dataGroup_lo_977[287:256];
  wire [511:0]  dataGroup_lo_978 = {dataGroup_lo_hi_978, dataGroup_lo_lo_978};
  wire [511:0]  dataGroup_hi_978 = {dataGroup_hi_hi_978, dataGroup_hi_lo_978};
  wire [31:0]   dataGroup_2_100 = dataGroup_hi_978[31:0];
  wire [511:0]  dataGroup_lo_979 = {dataGroup_lo_hi_979, dataGroup_lo_lo_979};
  wire [511:0]  dataGroup_hi_979 = {dataGroup_hi_hi_979, dataGroup_hi_lo_979};
  wire [31:0]   dataGroup_3_100 = dataGroup_hi_979[287:256];
  wire [63:0]   res_lo_100 = {dataGroup_1_100, dataGroup_0_100};
  wire [63:0]   res_hi_100 = {dataGroup_3_100, dataGroup_2_100};
  wire [127:0]  res_184 = {res_hi_100, res_lo_100};
  wire [511:0]  dataGroup_lo_980 = {dataGroup_lo_hi_980, dataGroup_lo_lo_980};
  wire [511:0]  dataGroup_hi_980 = {dataGroup_hi_hi_980, dataGroup_hi_lo_980};
  wire [31:0]   dataGroup_0_101 = dataGroup_lo_980[63:32];
  wire [511:0]  dataGroup_lo_981 = {dataGroup_lo_hi_981, dataGroup_lo_lo_981};
  wire [511:0]  dataGroup_hi_981 = {dataGroup_hi_hi_981, dataGroup_hi_lo_981};
  wire [31:0]   dataGroup_1_101 = dataGroup_lo_981[319:288];
  wire [511:0]  dataGroup_lo_982 = {dataGroup_lo_hi_982, dataGroup_lo_lo_982};
  wire [511:0]  dataGroup_hi_982 = {dataGroup_hi_hi_982, dataGroup_hi_lo_982};
  wire [31:0]   dataGroup_2_101 = dataGroup_hi_982[63:32];
  wire [511:0]  dataGroup_lo_983 = {dataGroup_lo_hi_983, dataGroup_lo_lo_983};
  wire [511:0]  dataGroup_hi_983 = {dataGroup_hi_hi_983, dataGroup_hi_lo_983};
  wire [31:0]   dataGroup_3_101 = dataGroup_hi_983[319:288];
  wire [63:0]   res_lo_101 = {dataGroup_1_101, dataGroup_0_101};
  wire [63:0]   res_hi_101 = {dataGroup_3_101, dataGroup_2_101};
  wire [127:0]  res_185 = {res_hi_101, res_lo_101};
  wire [511:0]  dataGroup_lo_984 = {dataGroup_lo_hi_984, dataGroup_lo_lo_984};
  wire [511:0]  dataGroup_hi_984 = {dataGroup_hi_hi_984, dataGroup_hi_lo_984};
  wire [31:0]   dataGroup_0_102 = dataGroup_lo_984[95:64];
  wire [511:0]  dataGroup_lo_985 = {dataGroup_lo_hi_985, dataGroup_lo_lo_985};
  wire [511:0]  dataGroup_hi_985 = {dataGroup_hi_hi_985, dataGroup_hi_lo_985};
  wire [31:0]   dataGroup_1_102 = dataGroup_lo_985[351:320];
  wire [511:0]  dataGroup_lo_986 = {dataGroup_lo_hi_986, dataGroup_lo_lo_986};
  wire [511:0]  dataGroup_hi_986 = {dataGroup_hi_hi_986, dataGroup_hi_lo_986};
  wire [31:0]   dataGroup_2_102 = dataGroup_hi_986[95:64];
  wire [511:0]  dataGroup_lo_987 = {dataGroup_lo_hi_987, dataGroup_lo_lo_987};
  wire [511:0]  dataGroup_hi_987 = {dataGroup_hi_hi_987, dataGroup_hi_lo_987};
  wire [31:0]   dataGroup_3_102 = dataGroup_hi_987[351:320];
  wire [63:0]   res_lo_102 = {dataGroup_1_102, dataGroup_0_102};
  wire [63:0]   res_hi_102 = {dataGroup_3_102, dataGroup_2_102};
  wire [127:0]  res_186 = {res_hi_102, res_lo_102};
  wire [511:0]  dataGroup_lo_988 = {dataGroup_lo_hi_988, dataGroup_lo_lo_988};
  wire [511:0]  dataGroup_hi_988 = {dataGroup_hi_hi_988, dataGroup_hi_lo_988};
  wire [31:0]   dataGroup_0_103 = dataGroup_lo_988[127:96];
  wire [511:0]  dataGroup_lo_989 = {dataGroup_lo_hi_989, dataGroup_lo_lo_989};
  wire [511:0]  dataGroup_hi_989 = {dataGroup_hi_hi_989, dataGroup_hi_lo_989};
  wire [31:0]   dataGroup_1_103 = dataGroup_lo_989[383:352];
  wire [511:0]  dataGroup_lo_990 = {dataGroup_lo_hi_990, dataGroup_lo_lo_990};
  wire [511:0]  dataGroup_hi_990 = {dataGroup_hi_hi_990, dataGroup_hi_lo_990};
  wire [31:0]   dataGroup_2_103 = dataGroup_hi_990[127:96];
  wire [511:0]  dataGroup_lo_991 = {dataGroup_lo_hi_991, dataGroup_lo_lo_991};
  wire [511:0]  dataGroup_hi_991 = {dataGroup_hi_hi_991, dataGroup_hi_lo_991};
  wire [31:0]   dataGroup_3_103 = dataGroup_hi_991[383:352];
  wire [63:0]   res_lo_103 = {dataGroup_1_103, dataGroup_0_103};
  wire [63:0]   res_hi_103 = {dataGroup_3_103, dataGroup_2_103};
  wire [127:0]  res_187 = {res_hi_103, res_lo_103};
  wire [511:0]  dataGroup_lo_992 = {dataGroup_lo_hi_992, dataGroup_lo_lo_992};
  wire [511:0]  dataGroup_hi_992 = {dataGroup_hi_hi_992, dataGroup_hi_lo_992};
  wire [31:0]   dataGroup_0_104 = dataGroup_lo_992[159:128];
  wire [511:0]  dataGroup_lo_993 = {dataGroup_lo_hi_993, dataGroup_lo_lo_993};
  wire [511:0]  dataGroup_hi_993 = {dataGroup_hi_hi_993, dataGroup_hi_lo_993};
  wire [31:0]   dataGroup_1_104 = dataGroup_lo_993[415:384];
  wire [511:0]  dataGroup_lo_994 = {dataGroup_lo_hi_994, dataGroup_lo_lo_994};
  wire [511:0]  dataGroup_hi_994 = {dataGroup_hi_hi_994, dataGroup_hi_lo_994};
  wire [31:0]   dataGroup_2_104 = dataGroup_hi_994[159:128];
  wire [511:0]  dataGroup_lo_995 = {dataGroup_lo_hi_995, dataGroup_lo_lo_995};
  wire [511:0]  dataGroup_hi_995 = {dataGroup_hi_hi_995, dataGroup_hi_lo_995};
  wire [31:0]   dataGroup_3_104 = dataGroup_hi_995[415:384];
  wire [63:0]   res_lo_104 = {dataGroup_1_104, dataGroup_0_104};
  wire [63:0]   res_hi_104 = {dataGroup_3_104, dataGroup_2_104};
  wire [127:0]  res_188 = {res_hi_104, res_lo_104};
  wire [511:0]  dataGroup_lo_996 = {dataGroup_lo_hi_996, dataGroup_lo_lo_996};
  wire [511:0]  dataGroup_hi_996 = {dataGroup_hi_hi_996, dataGroup_hi_lo_996};
  wire [31:0]   dataGroup_0_105 = dataGroup_lo_996[191:160];
  wire [511:0]  dataGroup_lo_997 = {dataGroup_lo_hi_997, dataGroup_lo_lo_997};
  wire [511:0]  dataGroup_hi_997 = {dataGroup_hi_hi_997, dataGroup_hi_lo_997};
  wire [31:0]   dataGroup_1_105 = dataGroup_lo_997[447:416];
  wire [511:0]  dataGroup_lo_998 = {dataGroup_lo_hi_998, dataGroup_lo_lo_998};
  wire [511:0]  dataGroup_hi_998 = {dataGroup_hi_hi_998, dataGroup_hi_lo_998};
  wire [31:0]   dataGroup_2_105 = dataGroup_hi_998[191:160];
  wire [511:0]  dataGroup_lo_999 = {dataGroup_lo_hi_999, dataGroup_lo_lo_999};
  wire [511:0]  dataGroup_hi_999 = {dataGroup_hi_hi_999, dataGroup_hi_lo_999};
  wire [31:0]   dataGroup_3_105 = dataGroup_hi_999[447:416];
  wire [63:0]   res_lo_105 = {dataGroup_1_105, dataGroup_0_105};
  wire [63:0]   res_hi_105 = {dataGroup_3_105, dataGroup_2_105};
  wire [127:0]  res_189 = {res_hi_105, res_lo_105};
  wire [511:0]  dataGroup_lo_1000 = {dataGroup_lo_hi_1000, dataGroup_lo_lo_1000};
  wire [511:0]  dataGroup_hi_1000 = {dataGroup_hi_hi_1000, dataGroup_hi_lo_1000};
  wire [31:0]   dataGroup_0_106 = dataGroup_lo_1000[223:192];
  wire [511:0]  dataGroup_lo_1001 = {dataGroup_lo_hi_1001, dataGroup_lo_lo_1001};
  wire [511:0]  dataGroup_hi_1001 = {dataGroup_hi_hi_1001, dataGroup_hi_lo_1001};
  wire [31:0]   dataGroup_1_106 = dataGroup_lo_1001[479:448];
  wire [511:0]  dataGroup_lo_1002 = {dataGroup_lo_hi_1002, dataGroup_lo_lo_1002};
  wire [511:0]  dataGroup_hi_1002 = {dataGroup_hi_hi_1002, dataGroup_hi_lo_1002};
  wire [31:0]   dataGroup_2_106 = dataGroup_hi_1002[223:192];
  wire [511:0]  dataGroup_lo_1003 = {dataGroup_lo_hi_1003, dataGroup_lo_lo_1003};
  wire [511:0]  dataGroup_hi_1003 = {dataGroup_hi_hi_1003, dataGroup_hi_lo_1003};
  wire [31:0]   dataGroup_3_106 = dataGroup_hi_1003[479:448];
  wire [63:0]   res_lo_106 = {dataGroup_1_106, dataGroup_0_106};
  wire [63:0]   res_hi_106 = {dataGroup_3_106, dataGroup_2_106};
  wire [127:0]  res_190 = {res_hi_106, res_lo_106};
  wire [511:0]  dataGroup_lo_1004 = {dataGroup_lo_hi_1004, dataGroup_lo_lo_1004};
  wire [511:0]  dataGroup_hi_1004 = {dataGroup_hi_hi_1004, dataGroup_hi_lo_1004};
  wire [31:0]   dataGroup_0_107 = dataGroup_lo_1004[255:224];
  wire [511:0]  dataGroup_lo_1005 = {dataGroup_lo_hi_1005, dataGroup_lo_lo_1005};
  wire [511:0]  dataGroup_hi_1005 = {dataGroup_hi_hi_1005, dataGroup_hi_lo_1005};
  wire [31:0]   dataGroup_1_107 = dataGroup_lo_1005[511:480];
  wire [511:0]  dataGroup_lo_1006 = {dataGroup_lo_hi_1006, dataGroup_lo_lo_1006};
  wire [511:0]  dataGroup_hi_1006 = {dataGroup_hi_hi_1006, dataGroup_hi_lo_1006};
  wire [31:0]   dataGroup_2_107 = dataGroup_hi_1006[255:224];
  wire [511:0]  dataGroup_lo_1007 = {dataGroup_lo_hi_1007, dataGroup_lo_lo_1007};
  wire [511:0]  dataGroup_hi_1007 = {dataGroup_hi_hi_1007, dataGroup_hi_lo_1007};
  wire [31:0]   dataGroup_3_107 = dataGroup_hi_1007[511:480];
  wire [63:0]   res_lo_107 = {dataGroup_1_107, dataGroup_0_107};
  wire [63:0]   res_hi_107 = {dataGroup_3_107, dataGroup_2_107};
  wire [127:0]  res_191 = {res_hi_107, res_lo_107};
  wire [255:0]  lo_lo_23 = {res_185, res_184};
  wire [255:0]  lo_hi_23 = {res_187, res_186};
  wire [511:0]  lo_23 = {lo_hi_23, lo_lo_23};
  wire [255:0]  hi_lo_23 = {res_189, res_188};
  wire [255:0]  hi_hi_23 = {res_191, res_190};
  wire [511:0]  hi_23 = {hi_hi_23, hi_lo_23};
  wire [1023:0] regroupLoadData_2_7 = {hi_23, lo_23};
  wire          vrfWritePort_0_valid_0 = accessState_0 & writeReadyReg;
  wire [3:0]    vrfWritePort_0_bits_mask_0 = maskForGroup[3:0];
  wire [3:0]    vrfWritePort_1_bits_mask_0 = maskForGroup[7:4];
  wire [3:0]    vrfWritePort_2_bits_mask_0 = maskForGroup[11:8];
  wire [3:0]    vrfWritePort_3_bits_mask_0 = maskForGroup[15:12];
  wire [7:0]    _vrfWritePort_3_bits_data_T = 8'h1 << accessPtr;
  wire [31:0]   vrfWritePort_0_bits_data_0 =
    (_vrfWritePort_3_bits_data_T[0] ? accessData_0[31:0] : 32'h0) | (_vrfWritePort_3_bits_data_T[1] ? accessData_1[31:0] : 32'h0) | (_vrfWritePort_3_bits_data_T[2] ? accessData_2[31:0] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[3] ? accessData_3[31:0] : 32'h0) | (_vrfWritePort_3_bits_data_T[4] ? accessData_4[31:0] : 32'h0) | (_vrfWritePort_3_bits_data_T[5] ? accessData_5[31:0] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[6] ? accessData_6[31:0] : 32'h0) | (_vrfWritePort_3_bits_data_T[7] ? accessData_7[31:0] : 32'h0);
  wire [3:0]    vrfWritePort_0_bits_offset_0 = dataGroup[3:0];
  wire [3:0]    vrfWritePort_1_bits_offset_0 = dataGroup[3:0];
  wire [3:0]    vrfWritePort_2_bits_offset_0 = dataGroup[3:0];
  wire [3:0]    vrfWritePort_3_bits_offset_0 = dataGroup[3:0];
  wire [4:0]    _GEN_7 = {2'h0, accessPtr} * {1'h0, segmentInstructionIndexInterval} + {2'h0, dataGroup[6:4]};
  wire [4:0]    vrfWritePort_0_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_7;
  assign accessStateUpdate_0 = ~(vrfWritePort_0_ready_0 & vrfWritePort_0_valid_0) & accessState_0;
  wire          vrfWritePort_1_valid_0 = accessState_1 & writeReadyReg;
  wire [31:0]   vrfWritePort_1_bits_data_0 =
    (_vrfWritePort_3_bits_data_T[0] ? accessData_0[63:32] : 32'h0) | (_vrfWritePort_3_bits_data_T[1] ? accessData_1[63:32] : 32'h0) | (_vrfWritePort_3_bits_data_T[2] ? accessData_2[63:32] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[3] ? accessData_3[63:32] : 32'h0) | (_vrfWritePort_3_bits_data_T[4] ? accessData_4[63:32] : 32'h0) | (_vrfWritePort_3_bits_data_T[5] ? accessData_5[63:32] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[6] ? accessData_6[63:32] : 32'h0) | (_vrfWritePort_3_bits_data_T[7] ? accessData_7[63:32] : 32'h0);
  wire [4:0]    vrfWritePort_1_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_7;
  assign accessStateUpdate_1 = ~(vrfWritePort_1_ready_0 & vrfWritePort_1_valid_0) & accessState_1;
  wire          vrfWritePort_2_valid_0 = accessState_2 & writeReadyReg;
  wire [31:0]   vrfWritePort_2_bits_data_0 =
    (_vrfWritePort_3_bits_data_T[0] ? accessData_0[95:64] : 32'h0) | (_vrfWritePort_3_bits_data_T[1] ? accessData_1[95:64] : 32'h0) | (_vrfWritePort_3_bits_data_T[2] ? accessData_2[95:64] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[3] ? accessData_3[95:64] : 32'h0) | (_vrfWritePort_3_bits_data_T[4] ? accessData_4[95:64] : 32'h0) | (_vrfWritePort_3_bits_data_T[5] ? accessData_5[95:64] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[6] ? accessData_6[95:64] : 32'h0) | (_vrfWritePort_3_bits_data_T[7] ? accessData_7[95:64] : 32'h0);
  wire [4:0]    vrfWritePort_2_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_7;
  assign accessStateUpdate_2 = ~(vrfWritePort_2_ready_0 & vrfWritePort_2_valid_0) & accessState_2;
  wire          vrfWritePort_3_valid_0 = accessState_3 & writeReadyReg;
  wire [31:0]   vrfWritePort_3_bits_data_0 =
    (_vrfWritePort_3_bits_data_T[0] ? accessData_0[127:96] : 32'h0) | (_vrfWritePort_3_bits_data_T[1] ? accessData_1[127:96] : 32'h0) | (_vrfWritePort_3_bits_data_T[2] ? accessData_2[127:96] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[3] ? accessData_3[127:96] : 32'h0) | (_vrfWritePort_3_bits_data_T[4] ? accessData_4[127:96] : 32'h0) | (_vrfWritePort_3_bits_data_T[5] ? accessData_5[127:96] : 32'h0)
    | (_vrfWritePort_3_bits_data_T[6] ? accessData_6[127:96] : 32'h0) | (_vrfWritePort_3_bits_data_T[7] ? accessData_7[127:96] : 32'h0);
  wire [4:0]    vrfWritePort_3_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_7;
  assign accessStateUpdate_3 = ~(vrfWritePort_3_ready_0 & vrfWritePort_3_valid_0) & accessState_3;
  reg           sendStateReg_0;
  reg           sendStateReg_1;
  reg           sendStateReg_2;
  reg           sendStateReg_3;
  wire          lastCacheRequest = lastRequest & _lastCacheRequest_T;
  reg           lastCacheRequestReg;
  reg           lastCacheLineAckReg;
  wire          bufferClear = ~(memResponse_valid_0 | alignedDequeue_valid | bufferFull | ~writeStageReady);
  wire          _status_idle_output = lastCacheRequestReg & lastCacheLineAckReg & bufferClear & ~sendRequest;
  reg           idleNext;
  always @(posedge clock) begin
    if (reset) begin
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 12'h0;
      csrInterfaceReg_vStart <= 12'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      requestFireNext <= 1'h0;
      dataEEW <= 2'h0;
      maskReg <= 16'h0;
      needAmend <= 1'h0;
      lastMaskAmendReg <= 15'h0;
      maskGroupCounter <= 7'h0;
      maskCounterInGroup <= 2'h0;
      maskForGroup <= 16'h0;
      isLastMaskGroup <= 1'h0;
      accessData_0 <= 128'h0;
      accessData_1 <= 128'h0;
      accessData_2 <= 128'h0;
      accessData_3 <= 128'h0;
      accessData_4 <= 128'h0;
      accessData_5 <= 128'h0;
      accessData_6 <= 128'h0;
      accessData_7 <= 128'h0;
      accessPtr <= 3'h0;
      accessState_0 <= 1'h0;
      accessState_1 <= 1'h0;
      accessState_2 <= 1'h0;
      accessState_3 <= 1'h0;
      dataGroup <= 7'h0;
      dataBuffer_0 <= 128'h0;
      dataBuffer_1 <= 128'h0;
      dataBuffer_2 <= 128'h0;
      dataBuffer_3 <= 128'h0;
      dataBuffer_4 <= 128'h0;
      dataBuffer_5 <= 128'h0;
      dataBuffer_6 <= 128'h0;
      dataBuffer_7 <= 128'h0;
      bufferBaseCacheLineIndex <= 8'h0;
      cacheLineIndexInBuffer <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      lastWriteVrfIndexReg <= 15'h0;
      lastCacheNeedPush <= 1'h0;
      cacheLineNumberReg <= 15'h0;
      sendRequest <= 1'h0;
      writeReadyReg <= 1'h0;
      unalignedCacheLine_valid <= 1'h0;
      unalignedCacheLine_bits_data <= 128'h0;
      unalignedCacheLine_bits_index <= 8'h0;
      bufferFull <= 1'h0;
      waitForFirstDataGroup <= 1'h0;
      sendStateReg_0 <= 1'h0;
      sendStateReg_1 <= 1'h0;
      sendStateReg_2 <= 1'h0;
      sendStateReg_3 <= 1'h0;
      lastCacheRequestReg <= 1'h1;
      lastCacheLineAckReg <= 1'h1;
      idleNext <= 1'h1;
    end
    else begin
      automatic logic _GEN_8 = bufferDequeueFire | accessStateCheck & ~lastPtr;
      if (lsuRequest_valid) begin
        lsuRequestReg_instructionInformation_nf <= nfCorrection;
        lsuRequestReg_instructionInformation_mew <= ~invalidInstruction & lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataEEW <= lsuRequest_bits_instructionInformation_eew;
        needAmend <= |(csrInterface_vl[3:0]);
        lastMaskAmendReg <= lastMaskAmend;
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
        lastWriteVrfIndexReg <= lastWriteVrfIndex;
        lastCacheNeedPush <= lastCacheLineIndex == lastWriteVrfIndex;
        cacheLineNumberReg <= lastCacheLineIndex;
      end
      requestFireNext <= lsuRequest_valid;
      if (_maskSelect_valid_output | lsuRequest_valid) begin
        maskReg <= maskAmend;
        isLastMaskGroup <= lsuRequest_valid ? csrInterface_vl[11:4] == 8'h0 : {1'h0, _maskSelect_bits_output} == csrInterfaceReg_vl[11:4];
      end
      if (bufferDequeueFire & isLastDataGroup)
        maskGroupCounter <= nextMaskGroup;
      else if (lsuRequest_valid)
        maskGroupCounter <= 7'h0;
      if (lsuRequest_valid | bufferDequeueFire) begin
        maskCounterInGroup <= isLastDataGroup | lsuRequest_valid ? 2'h0 : nextMaskCount;
        waitForFirstDataGroup <= lsuRequest_valid;
      end
      if (bufferDequeueFire) begin
        automatic logic [7:0]    _GEN_9;
        automatic logic [1023:0] _GEN_10;
        _GEN_9 = 8'h1 << lsuRequestReg_instructionInformation_nf;
        _GEN_10 =
          (dataEEWOH[0]
             ? (_GEN_9[0] ? regroupLoadData_0_0 : 1024'h0) | (_GEN_9[1] ? regroupLoadData_0_1 : 1024'h0) | (_GEN_9[2] ? regroupLoadData_0_2 : 1024'h0) | (_GEN_9[3] ? regroupLoadData_0_3 : 1024'h0)
               | (_GEN_9[4] ? regroupLoadData_0_4 : 1024'h0) | (_GEN_9[5] ? regroupLoadData_0_5 : 1024'h0) | (_GEN_9[6] ? regroupLoadData_0_6 : 1024'h0) | (_GEN_9[7] ? regroupLoadData_0_7 : 1024'h0)
             : 1024'h0)
          | (dataEEWOH[1]
               ? (_GEN_9[0] ? regroupLoadData_1_0 : 1024'h0) | (_GEN_9[1] ? regroupLoadData_1_1 : 1024'h0) | (_GEN_9[2] ? regroupLoadData_1_2 : 1024'h0) | (_GEN_9[3] ? regroupLoadData_1_3 : 1024'h0)
                 | (_GEN_9[4] ? regroupLoadData_1_4 : 1024'h0) | (_GEN_9[5] ? regroupLoadData_1_5 : 1024'h0) | (_GEN_9[6] ? regroupLoadData_1_6 : 1024'h0) | (_GEN_9[7] ? regroupLoadData_1_7 : 1024'h0)
               : 1024'h0)
          | (dataEEWOH[2]
               ? (_GEN_9[0] ? regroupLoadData_2_0 : 1024'h0) | (_GEN_9[1] ? regroupLoadData_2_1 : 1024'h0) | (_GEN_9[2] ? regroupLoadData_2_2 : 1024'h0) | (_GEN_9[3] ? regroupLoadData_2_3 : 1024'h0)
                 | (_GEN_9[4] ? regroupLoadData_2_4 : 1024'h0) | (_GEN_9[5] ? regroupLoadData_2_5 : 1024'h0) | (_GEN_9[6] ? regroupLoadData_2_6 : 1024'h0) | (_GEN_9[7] ? regroupLoadData_2_7 : 1024'h0)
               : 1024'h0);
        maskForGroup <= maskForGroupWire;
        accessData_0 <= _GEN_10[127:0];
        accessData_1 <= _GEN_10[255:128];
        accessData_2 <= _GEN_10[383:256];
        accessData_3 <= _GEN_10[511:384];
        accessData_4 <= _GEN_10[639:512];
        accessData_5 <= _GEN_10[767:640];
        accessData_6 <= _GEN_10[895:768];
        accessData_7 <= _GEN_10[1023:896];
        dataGroup <= waitForFirstDataGroup ? 7'h0 : dataGroup + 7'h1;
        sendStateReg_0 <= initSendState_0;
        sendStateReg_1 <= initSendState_1;
        sendStateReg_2 <= initSendState_2;
        sendStateReg_3 <= initSendState_3;
      end
      if (_GEN_8)
        accessPtr <= bufferDequeueFire ? lsuRequestReg_instructionInformation_nf : accessPtr - 3'h1;
      accessState_0 <= _GEN_8 ? (bufferDequeueFire ? initSendState_0 : sendStateReg_0) : accessStateUpdate_0;
      accessState_1 <= _GEN_8 ? (bufferDequeueFire ? initSendState_1 : sendStateReg_1) : accessStateUpdate_1;
      accessState_2 <= _GEN_8 ? (bufferDequeueFire ? initSendState_2 : sendStateReg_2) : accessStateUpdate_2;
      accessState_3 <= _GEN_8 ? (bufferDequeueFire ? initSendState_3 : sendStateReg_3) : accessStateUpdate_3;
      if (bufferEnqueueSelect[0])
        dataBuffer_0 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[1])
        dataBuffer_1 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[2])
        dataBuffer_2 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[3])
        dataBuffer_3 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[4])
        dataBuffer_4 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[5])
        dataBuffer_5 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[6])
        dataBuffer_6 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[7])
        dataBuffer_7 <= alignedDequeue_bits_data;
      if (_bufferTailFire_T & cacheLineIndexInBuffer == 3'h0)
        bufferBaseCacheLineIndex <= alignedDequeue_bits_index;
      if (_bufferTailFire_T | bufferDequeueFire)
        cacheLineIndexInBuffer <= bufferDequeueFire ? 3'h0 : cacheLineIndexInBuffer + 3'h1;
      if (validInstruction | _lastCacheRequest_T & lastRequest)
        sendRequest <= lsuRequest_valid & (|csrInterface_vl);
      writeReadyReg <= ~lsuRequest_valid;
      if (unalignedEnqueueFire ^ _bufferTailFire_T | lsuRequest_valid)
        unalignedCacheLine_valid <= unalignedEnqueueFire;
      if (unalignedEnqueueFire) begin
        unalignedCacheLine_bits_data <= memResponse_bits_data_0;
        unalignedCacheLine_bits_index <= nextIndex;
      end
      if (bufferTailFire | bufferDequeueFire)
        bufferFull <= ~bufferDequeueFire;
      if (lastCacheRequest | validInstruction)
        lastCacheRequestReg <= lastCacheRequest;
      if (anyLastCacheLineAck | validInstruction)
        lastCacheLineAckReg <= anyLastCacheLineAck;
      idleNext <= _status_idle_output;
    end
    invalidInstructionNext <= invalidInstruction & lsuRequest_valid;
    if (_lastCacheRequest_T | lsuRequest_valid)
      cacheLineIndex <= lsuRequest_valid ? 8'h0 : nextCacheLineIndex;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:76];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h4D; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        lsuRequestReg_instructionInformation_nf = _RANDOM[7'h0][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[7'h0][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[7'h0][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[7'h0][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[7'h0][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[7'h0][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[7'h0][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[7'h0][19];
        lsuRequestReg_rs1Data = {_RANDOM[7'h0][31:20], _RANDOM[7'h1][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[7'h1][31:20], _RANDOM[7'h2][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[7'h2][22:20];
        csrInterfaceReg_vl = {_RANDOM[7'h2][31:23], _RANDOM[7'h3][2:0]};
        csrInterfaceReg_vStart = _RANDOM[7'h3][14:3];
        csrInterfaceReg_vlmul = _RANDOM[7'h3][17:15];
        csrInterfaceReg_vSew = _RANDOM[7'h3][19:18];
        csrInterfaceReg_vxrm = _RANDOM[7'h3][21:20];
        csrInterfaceReg_vta = _RANDOM[7'h3][22];
        csrInterfaceReg_vma = _RANDOM[7'h3][23];
        requestFireNext = _RANDOM[7'h3][24];
        dataEEW = _RANDOM[7'h3][26:25];
        maskReg = {_RANDOM[7'h3][31:27], _RANDOM[7'h4][10:0]};
        needAmend = _RANDOM[7'h4][11];
        lastMaskAmendReg = _RANDOM[7'h4][26:12];
        maskGroupCounter = {_RANDOM[7'h4][31:27], _RANDOM[7'h5][1:0]};
        maskCounterInGroup = _RANDOM[7'h5][3:2];
        maskForGroup = _RANDOM[7'h5][19:4];
        isLastMaskGroup = _RANDOM[7'h5][20];
        accessData_0 = {_RANDOM[7'h5][31:21], _RANDOM[7'h6], _RANDOM[7'h7], _RANDOM[7'h8], _RANDOM[7'h9][20:0]};
        accessData_1 = {_RANDOM[7'h9][31:21], _RANDOM[7'hA], _RANDOM[7'hB], _RANDOM[7'hC], _RANDOM[7'hD][20:0]};
        accessData_2 = {_RANDOM[7'hD][31:21], _RANDOM[7'hE], _RANDOM[7'hF], _RANDOM[7'h10], _RANDOM[7'h11][20:0]};
        accessData_3 = {_RANDOM[7'h11][31:21], _RANDOM[7'h12], _RANDOM[7'h13], _RANDOM[7'h14], _RANDOM[7'h15][20:0]};
        accessData_4 = {_RANDOM[7'h15][31:21], _RANDOM[7'h16], _RANDOM[7'h17], _RANDOM[7'h18], _RANDOM[7'h19][20:0]};
        accessData_5 = {_RANDOM[7'h19][31:21], _RANDOM[7'h1A], _RANDOM[7'h1B], _RANDOM[7'h1C], _RANDOM[7'h1D][20:0]};
        accessData_6 = {_RANDOM[7'h1D][31:21], _RANDOM[7'h1E], _RANDOM[7'h1F], _RANDOM[7'h20], _RANDOM[7'h21][20:0]};
        accessData_7 = {_RANDOM[7'h21][31:21], _RANDOM[7'h22], _RANDOM[7'h23], _RANDOM[7'h24], _RANDOM[7'h25][20:0]};
        accessPtr = _RANDOM[7'h25][23:21];
        accessState_0 = _RANDOM[7'h25][24];
        accessState_1 = _RANDOM[7'h25][25];
        accessState_2 = _RANDOM[7'h25][26];
        accessState_3 = _RANDOM[7'h25][27];
        dataGroup = {_RANDOM[7'h25][31:28], _RANDOM[7'h26][2:0]};
        dataBuffer_0 = {_RANDOM[7'h26][31:3], _RANDOM[7'h27], _RANDOM[7'h28], _RANDOM[7'h29], _RANDOM[7'h2A][2:0]};
        dataBuffer_1 = {_RANDOM[7'h2A][31:3], _RANDOM[7'h2B], _RANDOM[7'h2C], _RANDOM[7'h2D], _RANDOM[7'h2E][2:0]};
        dataBuffer_2 = {_RANDOM[7'h2E][31:3], _RANDOM[7'h2F], _RANDOM[7'h30], _RANDOM[7'h31], _RANDOM[7'h32][2:0]};
        dataBuffer_3 = {_RANDOM[7'h32][31:3], _RANDOM[7'h33], _RANDOM[7'h34], _RANDOM[7'h35], _RANDOM[7'h36][2:0]};
        dataBuffer_4 = {_RANDOM[7'h36][31:3], _RANDOM[7'h37], _RANDOM[7'h38], _RANDOM[7'h39], _RANDOM[7'h3A][2:0]};
        dataBuffer_5 = {_RANDOM[7'h3A][31:3], _RANDOM[7'h3B], _RANDOM[7'h3C], _RANDOM[7'h3D], _RANDOM[7'h3E][2:0]};
        dataBuffer_6 = {_RANDOM[7'h3E][31:3], _RANDOM[7'h3F], _RANDOM[7'h40], _RANDOM[7'h41], _RANDOM[7'h42][2:0]};
        dataBuffer_7 = {_RANDOM[7'h42][31:3], _RANDOM[7'h43], _RANDOM[7'h44], _RANDOM[7'h45], _RANDOM[7'h46][2:0]};
        bufferBaseCacheLineIndex = _RANDOM[7'h46][10:3];
        cacheLineIndexInBuffer = _RANDOM[7'h46][13:11];
        invalidInstructionNext = _RANDOM[7'h46][14];
        segmentInstructionIndexInterval = _RANDOM[7'h46][18:15];
        lastWriteVrfIndexReg = {_RANDOM[7'h46][31:19], _RANDOM[7'h47][1:0]};
        lastCacheNeedPush = _RANDOM[7'h47][2];
        cacheLineNumberReg = _RANDOM[7'h47][17:3];
        cacheLineIndex = _RANDOM[7'h47][25:18];
        sendRequest = _RANDOM[7'h47][26];
        writeReadyReg = _RANDOM[7'h47][27];
        unalignedCacheLine_valid = _RANDOM[7'h47][28];
        unalignedCacheLine_bits_data = {_RANDOM[7'h47][31:29], _RANDOM[7'h48], _RANDOM[7'h49], _RANDOM[7'h4A], _RANDOM[7'h4B][28:0]};
        unalignedCacheLine_bits_index = {_RANDOM[7'h4B][31:29], _RANDOM[7'h4C][4:0]};
        bufferFull = _RANDOM[7'h4C][5];
        waitForFirstDataGroup = _RANDOM[7'h4C][6];
        sendStateReg_0 = _RANDOM[7'h4C][7];
        sendStateReg_1 = _RANDOM[7'h4C][8];
        sendStateReg_2 = _RANDOM[7'h4C][9];
        sendStateReg_3 = _RANDOM[7'h4C][10];
        lastCacheRequestReg = _RANDOM[7'h4C][11];
        lastCacheLineAckReg = _RANDOM[7'h4C][12];
        idleNext = _RANDOM[7'h4C][13];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign maskSelect_valid = _maskSelect_valid_output;
  assign maskSelect_bits = _maskSelect_bits_output;
  assign memRequest_valid = memRequest_valid_0;
  assign memRequest_bits_src = memRequest_bits_src_0;
  assign memRequest_bits_address = memRequest_bits_address_0;
  assign memResponse_ready = memResponse_ready_0;
  assign status_idle = _status_idle_output;
  assign status_last = ~idleNext & _status_idle_output | invalidInstructionNext;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_changeMaskGroup = _maskSelect_valid_output & ~lsuRequest_valid;
  assign status_startAddress = requestAddress;
  assign status_endAddress = {lsuRequestReg_rs1Data[31:4] + {13'h0, cacheLineNumberReg}, 4'h0};
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_offset = vrfWritePort_0_bits_offset_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_offset = vrfWritePort_1_bits_offset_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_offset = vrfWritePort_2_bits_offset_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_offset = vrfWritePort_3_bits_offset_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
endmodule

