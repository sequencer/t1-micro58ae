
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module LoadUnit(
  input          clock,
                 reset,
                 lsuRequest_valid,
  input  [2:0]   lsuRequest_bits_instructionInformation_nf,
  input          lsuRequest_bits_instructionInformation_mew,
  input  [1:0]   lsuRequest_bits_instructionInformation_mop,
  input  [4:0]   lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]   lsuRequest_bits_instructionInformation_eew,
  input  [4:0]   lsuRequest_bits_instructionInformation_vs3,
  input          lsuRequest_bits_instructionInformation_isStore,
                 lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  lsuRequest_bits_rs1Data,
                 lsuRequest_bits_rs2Data,
  input  [2:0]   lsuRequest_bits_instructionIndex,
  input  [11:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
  input  [31:0]  maskInput,
  output         maskSelect_valid,
  output [5:0]   maskSelect_bits,
  input          addressConflict,
                 memRequest_ready,
  output         memRequest_valid,
  output [6:0]   memRequest_bits_src,
  output [31:0]  memRequest_bits_address,
  output         memResponse_ready,
  input          memResponse_valid,
  input  [255:0] memResponse_bits_data,
  input  [6:0]   memResponse_bits_index,
  output         status_idle,
                 status_last,
  output [2:0]   status_instructionIndex,
  output         status_changeMaskGroup,
  output [31:0]  status_startAddress,
                 status_endAddress,
  input          vrfWritePort_0_ready,
  output         vrfWritePort_0_valid,
  output [4:0]   vrfWritePort_0_bits_vd,
  output [2:0]   vrfWritePort_0_bits_offset,
  output [3:0]   vrfWritePort_0_bits_mask,
  output [31:0]  vrfWritePort_0_bits_data,
  output [2:0]   vrfWritePort_0_bits_instructionIndex,
  input          vrfWritePort_1_ready,
  output         vrfWritePort_1_valid,
  output [4:0]   vrfWritePort_1_bits_vd,
  output [2:0]   vrfWritePort_1_bits_offset,
  output [3:0]   vrfWritePort_1_bits_mask,
  output [31:0]  vrfWritePort_1_bits_data,
  output [2:0]   vrfWritePort_1_bits_instructionIndex,
  input          vrfWritePort_2_ready,
  output         vrfWritePort_2_valid,
  output [4:0]   vrfWritePort_2_bits_vd,
  output [2:0]   vrfWritePort_2_bits_offset,
  output [3:0]   vrfWritePort_2_bits_mask,
  output [31:0]  vrfWritePort_2_bits_data,
  output [2:0]   vrfWritePort_2_bits_instructionIndex,
  input          vrfWritePort_3_ready,
  output         vrfWritePort_3_valid,
  output [4:0]   vrfWritePort_3_bits_vd,
  output [2:0]   vrfWritePort_3_bits_offset,
  output [3:0]   vrfWritePort_3_bits_mask,
  output [31:0]  vrfWritePort_3_bits_data,
  output [2:0]   vrfWritePort_3_bits_instructionIndex,
  input          vrfWritePort_4_ready,
  output         vrfWritePort_4_valid,
  output [4:0]   vrfWritePort_4_bits_vd,
  output [2:0]   vrfWritePort_4_bits_offset,
  output [3:0]   vrfWritePort_4_bits_mask,
  output [31:0]  vrfWritePort_4_bits_data,
  output [2:0]   vrfWritePort_4_bits_instructionIndex,
  input          vrfWritePort_5_ready,
  output         vrfWritePort_5_valid,
  output [4:0]   vrfWritePort_5_bits_vd,
  output [2:0]   vrfWritePort_5_bits_offset,
  output [3:0]   vrfWritePort_5_bits_mask,
  output [31:0]  vrfWritePort_5_bits_data,
  output [2:0]   vrfWritePort_5_bits_instructionIndex,
  input          vrfWritePort_6_ready,
  output         vrfWritePort_6_valid,
  output [4:0]   vrfWritePort_6_bits_vd,
  output [2:0]   vrfWritePort_6_bits_offset,
  output [3:0]   vrfWritePort_6_bits_mask,
  output [31:0]  vrfWritePort_6_bits_data,
  output [2:0]   vrfWritePort_6_bits_instructionIndex,
  input          vrfWritePort_7_ready,
  output         vrfWritePort_7_valid,
  output [4:0]   vrfWritePort_7_bits_vd,
  output [2:0]   vrfWritePort_7_bits_offset,
  output [3:0]   vrfWritePort_7_bits_mask,
  output [31:0]  vrfWritePort_7_bits_data,
  output [2:0]   vrfWritePort_7_bits_instructionIndex
);

  wire          memRequest_ready_0 = memRequest_ready;
  wire          memResponse_valid_0 = memResponse_valid;
  wire [255:0]  memResponse_bits_data_0 = memResponse_bits_data;
  wire [6:0]    memResponse_bits_index_0 = memResponse_bits_index;
  wire          vrfWritePort_0_ready_0 = vrfWritePort_0_ready;
  wire          vrfWritePort_1_ready_0 = vrfWritePort_1_ready;
  wire          vrfWritePort_2_ready_0 = vrfWritePort_2_ready;
  wire          vrfWritePort_3_ready_0 = vrfWritePort_3_ready;
  wire          vrfWritePort_4_ready_0 = vrfWritePort_4_ready;
  wire          vrfWritePort_5_ready_0 = vrfWritePort_5_ready;
  wire          vrfWritePort_6_ready_0 = vrfWritePort_6_ready;
  wire          vrfWritePort_7_ready_0 = vrfWritePort_7_ready;
  wire [1023:0] hi = 1024'h0;
  wire [1023:0] hi_1 = 1024'h0;
  wire [1023:0] hi_2 = 1024'h0;
  wire [1023:0] hi_3 = 1024'h0;
  wire [1023:0] hi_8 = 1024'h0;
  wire [1023:0] hi_9 = 1024'h0;
  wire [1023:0] hi_10 = 1024'h0;
  wire [1023:0] hi_11 = 1024'h0;
  wire [1023:0] hi_16 = 1024'h0;
  wire [1023:0] hi_17 = 1024'h0;
  wire [1023:0] hi_18 = 1024'h0;
  wire [1023:0] hi_19 = 1024'h0;
  wire [511:0]  lo_hi = 512'h0;
  wire [511:0]  hi_lo = 512'h0;
  wire [511:0]  hi_hi = 512'h0;
  wire [511:0]  lo_hi_1 = 512'h0;
  wire [511:0]  hi_lo_1 = 512'h0;
  wire [511:0]  hi_hi_1 = 512'h0;
  wire [511:0]  hi_lo_2 = 512'h0;
  wire [511:0]  hi_hi_2 = 512'h0;
  wire [511:0]  hi_lo_3 = 512'h0;
  wire [511:0]  hi_hi_3 = 512'h0;
  wire [511:0]  hi_hi_4 = 512'h0;
  wire [511:0]  hi_hi_5 = 512'h0;
  wire [511:0]  lo_hi_8 = 512'h0;
  wire [511:0]  hi_lo_8 = 512'h0;
  wire [511:0]  hi_hi_8 = 512'h0;
  wire [511:0]  lo_hi_9 = 512'h0;
  wire [511:0]  hi_lo_9 = 512'h0;
  wire [511:0]  hi_hi_9 = 512'h0;
  wire [511:0]  hi_lo_10 = 512'h0;
  wire [511:0]  hi_hi_10 = 512'h0;
  wire [511:0]  hi_lo_11 = 512'h0;
  wire [511:0]  hi_hi_11 = 512'h0;
  wire [511:0]  hi_hi_12 = 512'h0;
  wire [511:0]  hi_hi_13 = 512'h0;
  wire [511:0]  lo_hi_16 = 512'h0;
  wire [511:0]  hi_lo_16 = 512'h0;
  wire [511:0]  hi_hi_16 = 512'h0;
  wire [511:0]  lo_hi_17 = 512'h0;
  wire [511:0]  hi_lo_17 = 512'h0;
  wire [511:0]  hi_hi_17 = 512'h0;
  wire [511:0]  hi_lo_18 = 512'h0;
  wire [511:0]  hi_hi_18 = 512'h0;
  wire [511:0]  hi_lo_19 = 512'h0;
  wire [511:0]  hi_hi_19 = 512'h0;
  wire [511:0]  hi_hi_20 = 512'h0;
  wire [511:0]  hi_hi_21 = 512'h0;
  wire [255:0]  res_1 = 256'h0;
  wire [255:0]  res_2 = 256'h0;
  wire [255:0]  res_3 = 256'h0;
  wire [255:0]  res_4 = 256'h0;
  wire [255:0]  res_5 = 256'h0;
  wire [255:0]  res_6 = 256'h0;
  wire [255:0]  res_7 = 256'h0;
  wire [255:0]  res_10 = 256'h0;
  wire [255:0]  res_11 = 256'h0;
  wire [255:0]  res_12 = 256'h0;
  wire [255:0]  res_13 = 256'h0;
  wire [255:0]  res_14 = 256'h0;
  wire [255:0]  res_15 = 256'h0;
  wire [255:0]  res_19 = 256'h0;
  wire [255:0]  res_20 = 256'h0;
  wire [255:0]  res_21 = 256'h0;
  wire [255:0]  res_22 = 256'h0;
  wire [255:0]  res_23 = 256'h0;
  wire [255:0]  res_28 = 256'h0;
  wire [255:0]  res_29 = 256'h0;
  wire [255:0]  res_30 = 256'h0;
  wire [255:0]  res_31 = 256'h0;
  wire [255:0]  res_37 = 256'h0;
  wire [255:0]  res_38 = 256'h0;
  wire [255:0]  res_39 = 256'h0;
  wire [255:0]  res_46 = 256'h0;
  wire [255:0]  res_47 = 256'h0;
  wire [255:0]  res_55 = 256'h0;
  wire [255:0]  res_65 = 256'h0;
  wire [255:0]  res_66 = 256'h0;
  wire [255:0]  res_67 = 256'h0;
  wire [255:0]  res_68 = 256'h0;
  wire [255:0]  res_69 = 256'h0;
  wire [255:0]  res_70 = 256'h0;
  wire [255:0]  res_71 = 256'h0;
  wire [255:0]  res_74 = 256'h0;
  wire [255:0]  res_75 = 256'h0;
  wire [255:0]  res_76 = 256'h0;
  wire [255:0]  res_77 = 256'h0;
  wire [255:0]  res_78 = 256'h0;
  wire [255:0]  res_79 = 256'h0;
  wire [255:0]  res_83 = 256'h0;
  wire [255:0]  res_84 = 256'h0;
  wire [255:0]  res_85 = 256'h0;
  wire [255:0]  res_86 = 256'h0;
  wire [255:0]  res_87 = 256'h0;
  wire [255:0]  res_92 = 256'h0;
  wire [255:0]  res_93 = 256'h0;
  wire [255:0]  res_94 = 256'h0;
  wire [255:0]  res_95 = 256'h0;
  wire [255:0]  res_101 = 256'h0;
  wire [255:0]  res_102 = 256'h0;
  wire [255:0]  res_103 = 256'h0;
  wire [255:0]  res_110 = 256'h0;
  wire [255:0]  res_111 = 256'h0;
  wire [255:0]  res_119 = 256'h0;
  wire [255:0]  res_129 = 256'h0;
  wire [255:0]  res_130 = 256'h0;
  wire [255:0]  res_131 = 256'h0;
  wire [255:0]  res_132 = 256'h0;
  wire [255:0]  res_133 = 256'h0;
  wire [255:0]  res_134 = 256'h0;
  wire [255:0]  res_135 = 256'h0;
  wire [255:0]  res_138 = 256'h0;
  wire [255:0]  res_139 = 256'h0;
  wire [255:0]  res_140 = 256'h0;
  wire [255:0]  res_141 = 256'h0;
  wire [255:0]  res_142 = 256'h0;
  wire [255:0]  res_143 = 256'h0;
  wire [255:0]  res_147 = 256'h0;
  wire [255:0]  res_148 = 256'h0;
  wire [255:0]  res_149 = 256'h0;
  wire [255:0]  res_150 = 256'h0;
  wire [255:0]  res_151 = 256'h0;
  wire [255:0]  res_156 = 256'h0;
  wire [255:0]  res_157 = 256'h0;
  wire [255:0]  res_158 = 256'h0;
  wire [255:0]  res_159 = 256'h0;
  wire [255:0]  res_165 = 256'h0;
  wire [255:0]  res_166 = 256'h0;
  wire [255:0]  res_167 = 256'h0;
  wire [255:0]  res_174 = 256'h0;
  wire [255:0]  res_175 = 256'h0;
  wire [255:0]  res_183 = 256'h0;
  wire          vrfWritePort_0_bits_last = 1'h0;
  wire          vrfWritePort_1_bits_last = 1'h0;
  wire          vrfWritePort_2_bits_last = 1'h0;
  wire          vrfWritePort_3_bits_last = 1'h0;
  wire          vrfWritePort_4_bits_last = 1'h0;
  wire          vrfWritePort_5_bits_last = 1'h0;
  wire          vrfWritePort_6_bits_last = 1'h0;
  wire          vrfWritePort_7_bits_last = 1'h0;
  wire [31:0]   requestAddress;
  wire          unalignedEnqueueReady;
  reg  [2:0]    lsuRequestReg_instructionInformation_nf;
  reg           lsuRequestReg_instructionInformation_mew;
  reg  [1:0]    lsuRequestReg_instructionInformation_mop;
  reg  [4:0]    lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]    lsuRequestReg_instructionInformation_eew;
  reg  [4:0]    lsuRequestReg_instructionInformation_vs3;
  reg           lsuRequestReg_instructionInformation_isStore;
  reg           lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]   lsuRequestReg_rs1Data;
  reg  [31:0]   lsuRequestReg_rs2Data;
  reg  [2:0]    lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_0_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_1_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_2_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_3_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_4_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_5_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_6_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]    vrfWritePort_7_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [11:0]   csrInterfaceReg_vl;
  reg  [11:0]   csrInterfaceReg_vStart;
  reg  [2:0]    csrInterfaceReg_vlmul;
  reg  [1:0]    csrInterfaceReg_vSew;
  reg  [1:0]    csrInterfaceReg_vxrm;
  reg           csrInterfaceReg_vta;
  reg           csrInterfaceReg_vma;
  reg           requestFireNext;
  reg  [1:0]    dataEEW;
  wire [3:0]    _dataEEWOH_T = 4'h1 << dataEEW;
  wire [2:0]    dataEEWOH = _dataEEWOH_T[2:0];
  wire          isMaskType = lsuRequest_valid ? lsuRequest_bits_instructionInformation_maskedLoadStore : lsuRequestReg_instructionInformation_maskedLoadStore;
  wire [31:0]   maskAmend = isMaskType ? maskInput : 32'hFFFFFFFF;
  reg  [31:0]   maskReg;
  wire [31:0]   _lastMaskAmend_T_1 = 32'h1 << csrInterface_vl[4:0];
  wire [29:0]   _GEN = _lastMaskAmend_T_1[30:1] | _lastMaskAmend_T_1[31:2];
  wire [28:0]   _GEN_0 = _GEN[28:0] | {_lastMaskAmend_T_1[31], _GEN[29:2]};
  wire [26:0]   _GEN_1 = _GEN_0[26:0] | {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:4]};
  wire [22:0]   _GEN_2 = _GEN_1[22:0] | {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:27], _GEN_1[26:8]};
  wire [30:0]   lastMaskAmend = {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:27], _GEN_1[26:23], _GEN_2[22:15], _GEN_2[14:0] | {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:27], _GEN_1[26:23], _GEN_2[22:16]}};
  reg           needAmend;
  reg  [30:0]   lastMaskAmendReg;
  wire [1:0]    countEndForGroup = {1'h0, dataEEWOH[1]} | {2{dataEEWOH[2]}};
  reg  [5:0]    maskGroupCounter;
  wire [5:0]    nextMaskGroup = maskGroupCounter + 6'h1;
  reg  [1:0]    maskCounterInGroup;
  wire [1:0]    nextMaskCount = maskCounterInGroup + 2'h1;
  wire          isLastDataGroup = maskCounterInGroup == countEndForGroup;
  wire [5:0]    _maskSelect_bits_output = lsuRequest_valid ? 6'h0 : nextMaskGroup;
  reg  [31:0]   maskForGroup;
  reg           isLastMaskGroup;
  wire [31:0]   maskWire = maskReg & (needAmend & isLastMaskGroup ? {1'h0, lastMaskAmendReg} : 32'hFFFFFFFF);
  wire [3:0]    maskForGroupWire_lo_lo_lo_lo = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]    maskForGroupWire_lo_lo_lo_hi = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo = {maskForGroupWire_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo};
  wire [3:0]    maskForGroupWire_lo_lo_hi_lo = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi_hi = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi = {maskForGroupWire_lo_lo_hi_hi, maskForGroupWire_lo_lo_hi_lo};
  wire [15:0]   maskForGroupWire_lo_lo = {maskForGroupWire_lo_lo_hi, maskForGroupWire_lo_lo_lo};
  wire [3:0]    maskForGroupWire_lo_hi_lo_lo = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]    maskForGroupWire_lo_hi_lo_hi = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo = {maskForGroupWire_lo_hi_lo_hi, maskForGroupWire_lo_hi_lo_lo};
  wire [3:0]    maskForGroupWire_lo_hi_hi_lo = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi_hi = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi = {maskForGroupWire_lo_hi_hi_hi, maskForGroupWire_lo_hi_hi_lo};
  wire [15:0]   maskForGroupWire_lo_hi = {maskForGroupWire_lo_hi_hi, maskForGroupWire_lo_hi_lo};
  wire [31:0]   maskForGroupWire_lo = {maskForGroupWire_lo_hi, maskForGroupWire_lo_lo};
  wire [3:0]    maskForGroupWire_hi_lo_lo_lo = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]    maskForGroupWire_hi_lo_lo_hi = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo = {maskForGroupWire_hi_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo};
  wire [3:0]    maskForGroupWire_hi_lo_hi_lo = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi_hi = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi = {maskForGroupWire_hi_lo_hi_hi, maskForGroupWire_hi_lo_hi_lo};
  wire [15:0]   maskForGroupWire_hi_lo = {maskForGroupWire_hi_lo_hi, maskForGroupWire_hi_lo_lo};
  wire [3:0]    maskForGroupWire_hi_hi_lo_lo = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]    maskForGroupWire_hi_hi_lo_hi = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo = {maskForGroupWire_hi_hi_lo_hi, maskForGroupWire_hi_hi_lo_lo};
  wire [3:0]    maskForGroupWire_hi_hi_hi_lo = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi_hi = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_lo};
  wire [15:0]   maskForGroupWire_hi_hi = {maskForGroupWire_hi_hi_hi, maskForGroupWire_hi_hi_lo};
  wire [31:0]   maskForGroupWire_hi = {maskForGroupWire_hi_hi, maskForGroupWire_hi_lo};
  wire [3:0]    maskForGroupWire_lo_lo_lo_lo_1 = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]    maskForGroupWire_lo_lo_lo_hi_1 = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_lo_hi_lo_1 = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]    maskForGroupWire_lo_lo_hi_hi_1 = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_1 = {maskForGroupWire_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_hi_lo_1};
  wire [15:0]   maskForGroupWire_lo_lo_1 = {maskForGroupWire_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_hi_lo_lo_1 = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]    maskForGroupWire_lo_hi_lo_hi_1 = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_1 = {maskForGroupWire_lo_hi_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_lo_hi_hi_lo_1 = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]    maskForGroupWire_lo_hi_hi_hi_1 = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_lo_1};
  wire [15:0]   maskForGroupWire_lo_hi_1 = {maskForGroupWire_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_1};
  wire [31:0]   maskForGroupWire_lo_1 = {maskForGroupWire_lo_hi_1, maskForGroupWire_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_lo_lo_lo_1 = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]    maskForGroupWire_hi_lo_lo_hi_1 = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_1 = {maskForGroupWire_hi_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_lo_hi_lo_1 = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]    maskForGroupWire_hi_lo_hi_hi_1 = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_1 = {maskForGroupWire_hi_lo_hi_hi_1, maskForGroupWire_hi_lo_hi_lo_1};
  wire [15:0]   maskForGroupWire_hi_lo_1 = {maskForGroupWire_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_hi_lo_lo_1 = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]    maskForGroupWire_hi_hi_lo_hi_1 = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_1 = {maskForGroupWire_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_1};
  wire [3:0]    maskForGroupWire_hi_hi_hi_lo_1 = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]    maskForGroupWire_hi_hi_hi_hi_1 = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_lo_1};
  wire [15:0]   maskForGroupWire_hi_hi_1 = {maskForGroupWire_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_1};
  wire [31:0]   maskForGroupWire_hi_1 = {maskForGroupWire_hi_hi_1, maskForGroupWire_hi_lo_1};
  wire [3:0]    _maskForGroupWire_T_133 = 4'h1 << maskCounterInGroup;
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_2 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_2 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_2 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_2 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_2 = {maskForGroupWire_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_hi_lo_2};
  wire [31:0]   maskForGroupWire_lo_lo_2 = {maskForGroupWire_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_2 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_2 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_2 = {maskForGroupWire_lo_hi_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_2 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_2 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_lo_2};
  wire [31:0]   maskForGroupWire_lo_hi_2 = {maskForGroupWire_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_2};
  wire [63:0]   maskForGroupWire_lo_2 = {maskForGroupWire_lo_hi_2, maskForGroupWire_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_2 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_2 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_2 = {maskForGroupWire_hi_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_2 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_2 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_2 = {maskForGroupWire_hi_lo_hi_hi_2, maskForGroupWire_hi_lo_hi_lo_2};
  wire [31:0]   maskForGroupWire_hi_lo_2 = {maskForGroupWire_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_2 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_2 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_2 = {maskForGroupWire_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_2};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_2 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_2 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_lo_2};
  wire [31:0]   maskForGroupWire_hi_hi_2 = {maskForGroupWire_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_2};
  wire [63:0]   maskForGroupWire_hi_2 = {maskForGroupWire_hi_hi_2, maskForGroupWire_hi_lo_2};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_3 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_3 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_3 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_3 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_3 = {maskForGroupWire_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_hi_lo_3};
  wire [31:0]   maskForGroupWire_lo_lo_3 = {maskForGroupWire_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_3 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_3 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_3 = {maskForGroupWire_lo_hi_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_3 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_3 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_lo_3};
  wire [31:0]   maskForGroupWire_lo_hi_3 = {maskForGroupWire_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_3};
  wire [63:0]   maskForGroupWire_lo_3 = {maskForGroupWire_lo_hi_3, maskForGroupWire_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_3 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_3 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_3 = {maskForGroupWire_hi_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_3 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_3 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_3 = {maskForGroupWire_hi_lo_hi_hi_3, maskForGroupWire_hi_lo_hi_lo_3};
  wire [31:0]   maskForGroupWire_hi_lo_3 = {maskForGroupWire_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_3 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_3 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_3 = {maskForGroupWire_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_3};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_3 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_3 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_lo_3};
  wire [31:0]   maskForGroupWire_hi_hi_3 = {maskForGroupWire_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_3};
  wire [63:0]   maskForGroupWire_hi_3 = {maskForGroupWire_hi_hi_3, maskForGroupWire_hi_lo_3};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_4 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_4 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_4 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_4 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_4 = {maskForGroupWire_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_hi_lo_4};
  wire [31:0]   maskForGroupWire_lo_lo_4 = {maskForGroupWire_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_4 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_4 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_4 = {maskForGroupWire_lo_hi_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_4 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_4 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_lo_4};
  wire [31:0]   maskForGroupWire_lo_hi_4 = {maskForGroupWire_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_4};
  wire [63:0]   maskForGroupWire_lo_4 = {maskForGroupWire_lo_hi_4, maskForGroupWire_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_4 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_4 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_4 = {maskForGroupWire_hi_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_4 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_4 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_4 = {maskForGroupWire_hi_lo_hi_hi_4, maskForGroupWire_hi_lo_hi_lo_4};
  wire [31:0]   maskForGroupWire_hi_lo_4 = {maskForGroupWire_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_4 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_4 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_4 = {maskForGroupWire_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_4};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_4 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_4 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_lo_4};
  wire [31:0]   maskForGroupWire_hi_hi_4 = {maskForGroupWire_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_4};
  wire [63:0]   maskForGroupWire_hi_4 = {maskForGroupWire_hi_hi_4, maskForGroupWire_hi_lo_4};
  wire [7:0]    maskForGroupWire_lo_lo_lo_lo_5 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]    maskForGroupWire_lo_lo_lo_hi_5 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]   maskForGroupWire_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_lo_hi_lo_5 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]    maskForGroupWire_lo_lo_hi_hi_5 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]   maskForGroupWire_lo_lo_hi_5 = {maskForGroupWire_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_hi_lo_5};
  wire [31:0]   maskForGroupWire_lo_lo_5 = {maskForGroupWire_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_hi_lo_lo_5 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]    maskForGroupWire_lo_hi_lo_hi_5 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]   maskForGroupWire_lo_hi_lo_5 = {maskForGroupWire_lo_hi_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_lo_hi_hi_lo_5 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]    maskForGroupWire_lo_hi_hi_hi_5 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]   maskForGroupWire_lo_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_lo_5};
  wire [31:0]   maskForGroupWire_lo_hi_5 = {maskForGroupWire_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_5};
  wire [63:0]   maskForGroupWire_lo_5 = {maskForGroupWire_lo_hi_5, maskForGroupWire_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_lo_lo_lo_5 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]    maskForGroupWire_hi_lo_lo_hi_5 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]   maskForGroupWire_hi_lo_lo_5 = {maskForGroupWire_hi_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_lo_hi_lo_5 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]    maskForGroupWire_hi_lo_hi_hi_5 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]   maskForGroupWire_hi_lo_hi_5 = {maskForGroupWire_hi_lo_hi_hi_5, maskForGroupWire_hi_lo_hi_lo_5};
  wire [31:0]   maskForGroupWire_hi_lo_5 = {maskForGroupWire_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_hi_lo_lo_5 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]    maskForGroupWire_hi_hi_lo_hi_5 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]   maskForGroupWire_hi_hi_lo_5 = {maskForGroupWire_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_5};
  wire [7:0]    maskForGroupWire_hi_hi_hi_lo_5 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]    maskForGroupWire_hi_hi_hi_hi_5 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]   maskForGroupWire_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_lo_5};
  wire [31:0]   maskForGroupWire_hi_hi_5 = {maskForGroupWire_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_5};
  wire [63:0]   maskForGroupWire_hi_5 = {maskForGroupWire_hi_hi_5, maskForGroupWire_hi_lo_5};
  wire [31:0]   maskForGroupWire =
    (dataEEWOH[0] ? maskWire : 32'h0) | (dataEEWOH[1] ? (maskCounterInGroup[0] ? maskForGroupWire_hi : maskForGroupWire_lo_1) : 32'h0)
    | (dataEEWOH[2]
         ? (_maskForGroupWire_T_133[0] ? maskForGroupWire_lo_2[31:0] : 32'h0) | (_maskForGroupWire_T_133[1] ? maskForGroupWire_lo_3[63:32] : 32'h0) | (_maskForGroupWire_T_133[2] ? maskForGroupWire_hi_4[31:0] : 32'h0)
           | (_maskForGroupWire_T_133[3] ? maskForGroupWire_hi_5[63:32] : 32'h0)
         : 32'h0);
  wire [1:0]    initSendState_lo = maskForGroupWire[1:0];
  wire [1:0]    initSendState_hi = maskForGroupWire[3:2];
  wire          initSendState_0 = |{initSendState_hi, initSendState_lo};
  wire [1:0]    initSendState_lo_1 = maskForGroupWire[5:4];
  wire [1:0]    initSendState_hi_1 = maskForGroupWire[7:6];
  wire          initSendState_1 = |{initSendState_hi_1, initSendState_lo_1};
  wire [1:0]    initSendState_lo_2 = maskForGroupWire[9:8];
  wire [1:0]    initSendState_hi_2 = maskForGroupWire[11:10];
  wire          initSendState_2 = |{initSendState_hi_2, initSendState_lo_2};
  wire [1:0]    initSendState_lo_3 = maskForGroupWire[13:12];
  wire [1:0]    initSendState_hi_3 = maskForGroupWire[15:14];
  wire          initSendState_3 = |{initSendState_hi_3, initSendState_lo_3};
  wire [1:0]    initSendState_lo_4 = maskForGroupWire[17:16];
  wire [1:0]    initSendState_hi_4 = maskForGroupWire[19:18];
  wire          initSendState_4 = |{initSendState_hi_4, initSendState_lo_4};
  wire [1:0]    initSendState_lo_5 = maskForGroupWire[21:20];
  wire [1:0]    initSendState_hi_5 = maskForGroupWire[23:22];
  wire          initSendState_5 = |{initSendState_hi_5, initSendState_lo_5};
  wire [1:0]    initSendState_lo_6 = maskForGroupWire[25:24];
  wire [1:0]    initSendState_hi_6 = maskForGroupWire[27:26];
  wire          initSendState_6 = |{initSendState_hi_6, initSendState_lo_6};
  wire [1:0]    initSendState_lo_7 = maskForGroupWire[29:28];
  wire [1:0]    initSendState_hi_7 = maskForGroupWire[31:30];
  wire          initSendState_7 = |{initSendState_hi_7, initSendState_lo_7};
  reg  [255:0]  accessData_0;
  reg  [255:0]  accessData_1;
  reg  [255:0]  accessData_2;
  reg  [255:0]  accessData_3;
  reg  [255:0]  accessData_4;
  reg  [255:0]  accessData_5;
  reg  [255:0]  accessData_6;
  reg  [255:0]  accessData_7;
  reg  [2:0]    accessPtr;
  reg           accessState_0;
  reg           accessState_1;
  reg           accessState_2;
  reg           accessState_3;
  reg           accessState_4;
  reg           accessState_5;
  reg           accessState_6;
  reg           accessState_7;
  wire          accessStateUpdate_0;
  wire          accessStateUpdate_1;
  wire [1:0]    accessStateCheck_lo_lo = {accessStateUpdate_1, accessStateUpdate_0};
  wire          accessStateUpdate_2;
  wire          accessStateUpdate_3;
  wire [1:0]    accessStateCheck_lo_hi = {accessStateUpdate_3, accessStateUpdate_2};
  wire [3:0]    accessStateCheck_lo = {accessStateCheck_lo_hi, accessStateCheck_lo_lo};
  wire          accessStateUpdate_4;
  wire          accessStateUpdate_5;
  wire [1:0]    accessStateCheck_hi_lo = {accessStateUpdate_5, accessStateUpdate_4};
  wire          accessStateUpdate_6;
  wire          accessStateUpdate_7;
  wire [1:0]    accessStateCheck_hi_hi = {accessStateUpdate_7, accessStateUpdate_6};
  wire [3:0]    accessStateCheck_hi = {accessStateCheck_hi_hi, accessStateCheck_hi_lo};
  wire          accessStateCheck = {accessStateCheck_hi, accessStateCheck_lo} == 8'h0;
  reg  [5:0]    dataGroup;
  reg  [255:0]  dataBuffer_0;
  reg  [255:0]  dataBuffer_1;
  reg  [255:0]  dataBuffer_2;
  reg  [255:0]  dataBuffer_3;
  reg  [255:0]  dataBuffer_4;
  reg  [255:0]  dataBuffer_5;
  reg  [255:0]  dataBuffer_6;
  reg  [255:0]  dataBuffer_7;
  reg  [6:0]    bufferBaseCacheLineIndex;
  reg  [2:0]    cacheLineIndexInBuffer;
  wire [4:0]    initOffset = lsuRequestReg_rs1Data[4:0];
  wire          invalidInstruction = csrInterface_vl == 12'h0;
  reg           invalidInstructionNext;
  wire          wholeType = lsuRequest_bits_instructionInformation_lumop[3];
  wire [2:0]    nfCorrection = wholeType ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [3:0]    segmentInstructionIndexInterval;
  wire [18:0]   bytePerInstruction = {3'h0, {12'h0, {1'h0, nfCorrection} + 4'h1} * {4'h0, csrInterface_vl}} << lsuRequest_bits_instructionInformation_eew;
  wire [18:0]   accessMemSize = bytePerInstruction + {14'h0, lsuRequest_bits_rs1Data[4:0]};
  wire [13:0]   lastCacheLineIndex = accessMemSize[18:5] - {13'h0, accessMemSize[4:0] == 5'h0};
  wire [13:0]   lastWriteVrfIndex = bytePerInstruction[18:5] - {13'h0, bytePerInstruction[4:0] == 5'h0};
  reg  [13:0]   lastWriteVrfIndexReg;
  reg           lastCacheNeedPush;
  reg  [13:0]   cacheLineNumberReg;
  wire          memRequest_valid_0;
  wire          _lastCacheRequest_T = memRequest_ready_0 & memRequest_valid_0;
  reg  [6:0]    cacheLineIndex;
  wire [6:0]    memRequest_bits_src_0 = cacheLineIndex;
  wire [6:0]    nextCacheLineIndex = cacheLineIndex + 7'h1;
  wire          validInstruction = ~invalidInstruction & lsuRequest_valid;
  wire          lastRequest = cacheLineNumberReg == {7'h0, cacheLineIndex};
  reg           sendRequest;
  assign requestAddress = {lsuRequestReg_rs1Data[31:5] + {20'h0, cacheLineIndex}, 5'h0};
  wire [31:0]   memRequest_bits_address_0 = requestAddress;
  reg           writeReadyReg;
  assign memRequest_valid_0 = sendRequest & ~addressConflict;
  wire          memResponse_ready_0;
  wire          unalignedEnqueueFire = memResponse_ready_0 & memResponse_valid_0;
  wire          anyLastCacheLineAck = unalignedEnqueueFire & {7'h0, memResponse_bits_index_0} == cacheLineNumberReg;
  wire          alignedDequeueValid;
  wire [255:0]  alignedDequeue_bits_data_lo_72;
  reg           unalignedCacheLine_valid;
  reg  [255:0]  unalignedCacheLine_bits_data;
  reg  [6:0]    unalignedCacheLine_bits_index;
  wire [6:0]    alignedDequeue_bits_index = unalignedCacheLine_bits_index;
  wire          alignedDequeue_ready;
  assign unalignedEnqueueReady = alignedDequeue_ready | ~unalignedCacheLine_valid;
  assign memResponse_ready_0 = unalignedEnqueueReady;
  wire [6:0]    nextIndex = unalignedCacheLine_valid ? unalignedCacheLine_bits_index + 7'h1 : 7'h0;
  assign alignedDequeueValid = unalignedCacheLine_valid & (memResponse_valid_0 | {7'h0, unalignedCacheLine_bits_index} == cacheLineNumberReg & lastCacheNeedPush);
  wire          alignedDequeue_valid = alignedDequeueValid;
  wire          _bufferTailFire_T = alignedDequeue_ready & alignedDequeue_valid;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo = {unalignedCacheLine_bits_data[8], unalignedCacheLine_bits_data[0]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi = {unalignedCacheLine_bits_data[24], unalignedCacheLine_bits_data[16]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo = {alignedDequeue_bits_data_lo_lo_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo = {unalignedCacheLine_bits_data[40], unalignedCacheLine_bits_data[32]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi = {unalignedCacheLine_bits_data[56], unalignedCacheLine_bits_data[48]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi = {alignedDequeue_bits_data_lo_lo_lo_hi_hi, alignedDequeue_bits_data_lo_lo_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo = {alignedDequeue_bits_data_lo_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo = {unalignedCacheLine_bits_data[72], unalignedCacheLine_bits_data[64]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi = {unalignedCacheLine_bits_data[88], unalignedCacheLine_bits_data[80]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo = {alignedDequeue_bits_data_lo_lo_hi_lo_hi, alignedDequeue_bits_data_lo_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo = {unalignedCacheLine_bits_data[104], unalignedCacheLine_bits_data[96]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi = {unalignedCacheLine_bits_data[120], unalignedCacheLine_bits_data[112]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi = {alignedDequeue_bits_data_lo_lo_hi_hi_hi, alignedDequeue_bits_data_lo_lo_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi = {alignedDequeue_bits_data_lo_lo_hi_hi, alignedDequeue_bits_data_lo_lo_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_lo_lo = {alignedDequeue_bits_data_lo_lo_hi, alignedDequeue_bits_data_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo = {unalignedCacheLine_bits_data[136], unalignedCacheLine_bits_data[128]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi = {unalignedCacheLine_bits_data[152], unalignedCacheLine_bits_data[144]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo = {alignedDequeue_bits_data_lo_hi_lo_lo_hi, alignedDequeue_bits_data_lo_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo = {unalignedCacheLine_bits_data[168], unalignedCacheLine_bits_data[160]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi = {unalignedCacheLine_bits_data[184], unalignedCacheLine_bits_data[176]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi = {alignedDequeue_bits_data_lo_hi_lo_hi_hi, alignedDequeue_bits_data_lo_hi_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo = {alignedDequeue_bits_data_lo_hi_lo_hi, alignedDequeue_bits_data_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo = {unalignedCacheLine_bits_data[200], unalignedCacheLine_bits_data[192]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi = {unalignedCacheLine_bits_data[216], unalignedCacheLine_bits_data[208]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo = {alignedDequeue_bits_data_lo_hi_hi_lo_hi, alignedDequeue_bits_data_lo_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo = {unalignedCacheLine_bits_data[232], unalignedCacheLine_bits_data[224]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi = {unalignedCacheLine_bits_data[248], unalignedCacheLine_bits_data[240]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi = {alignedDequeue_bits_data_lo_hi_hi_hi_hi, alignedDequeue_bits_data_lo_hi_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi = {alignedDequeue_bits_data_lo_hi_hi_hi, alignedDequeue_bits_data_lo_hi_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_lo_hi = {alignedDequeue_bits_data_lo_hi_hi, alignedDequeue_bits_data_lo_hi_lo};
  wire [31:0]   alignedDequeue_bits_data_lo = {alignedDequeue_bits_data_lo_hi, alignedDequeue_bits_data_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo = {memResponse_bits_data_0[8], memResponse_bits_data_0[0]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi = {memResponse_bits_data_0[24], memResponse_bits_data_0[16]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo = {alignedDequeue_bits_data_hi_lo_lo_lo_hi, alignedDequeue_bits_data_hi_lo_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo = {memResponse_bits_data_0[40], memResponse_bits_data_0[32]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi = {memResponse_bits_data_0[56], memResponse_bits_data_0[48]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi = {alignedDequeue_bits_data_hi_lo_lo_hi_hi, alignedDequeue_bits_data_hi_lo_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo = {alignedDequeue_bits_data_hi_lo_lo_hi, alignedDequeue_bits_data_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo = {memResponse_bits_data_0[72], memResponse_bits_data_0[64]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi = {memResponse_bits_data_0[88], memResponse_bits_data_0[80]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo = {alignedDequeue_bits_data_hi_lo_hi_lo_hi, alignedDequeue_bits_data_hi_lo_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo = {memResponse_bits_data_0[104], memResponse_bits_data_0[96]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi = {memResponse_bits_data_0[120], memResponse_bits_data_0[112]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi = {alignedDequeue_bits_data_hi_lo_hi_hi_hi, alignedDequeue_bits_data_hi_lo_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi = {alignedDequeue_bits_data_hi_lo_hi_hi, alignedDequeue_bits_data_hi_lo_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_hi_lo = {alignedDequeue_bits_data_hi_lo_hi, alignedDequeue_bits_data_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo = {memResponse_bits_data_0[136], memResponse_bits_data_0[128]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi = {memResponse_bits_data_0[152], memResponse_bits_data_0[144]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo = {alignedDequeue_bits_data_hi_hi_lo_lo_hi, alignedDequeue_bits_data_hi_hi_lo_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo = {memResponse_bits_data_0[168], memResponse_bits_data_0[160]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi = {memResponse_bits_data_0[184], memResponse_bits_data_0[176]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi = {alignedDequeue_bits_data_hi_hi_lo_hi_hi, alignedDequeue_bits_data_hi_hi_lo_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo = {alignedDequeue_bits_data_hi_hi_lo_hi, alignedDequeue_bits_data_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo = {memResponse_bits_data_0[200], memResponse_bits_data_0[192]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi = {memResponse_bits_data_0[216], memResponse_bits_data_0[208]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo = {alignedDequeue_bits_data_hi_hi_hi_lo_hi, alignedDequeue_bits_data_hi_hi_hi_lo_lo};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo = {memResponse_bits_data_0[232], memResponse_bits_data_0[224]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi = {memResponse_bits_data_0[248], memResponse_bits_data_0[240]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi = {alignedDequeue_bits_data_hi_hi_hi_hi_hi, alignedDequeue_bits_data_hi_hi_hi_hi_lo};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi = {alignedDequeue_bits_data_hi_hi_hi_hi, alignedDequeue_bits_data_hi_hi_hi_lo};
  wire [15:0]   alignedDequeue_bits_data_hi_hi = {alignedDequeue_bits_data_hi_hi_hi, alignedDequeue_bits_data_hi_hi_lo};
  wire [31:0]   alignedDequeue_bits_data_hi = {alignedDequeue_bits_data_hi_hi, alignedDequeue_bits_data_hi_lo};
  wire [63:0]   _GEN_3 = {59'h0, initOffset};
  wire [63:0]   _alignedDequeue_bits_data_T_514 = {alignedDequeue_bits_data_hi, alignedDequeue_bits_data_lo} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_1 = {unalignedCacheLine_bits_data[9], unalignedCacheLine_bits_data[1]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_1 = {unalignedCacheLine_bits_data[25], unalignedCacheLine_bits_data[17]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_1 = {unalignedCacheLine_bits_data[41], unalignedCacheLine_bits_data[33]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_1 = {unalignedCacheLine_bits_data[57], unalignedCacheLine_bits_data[49]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_1 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_1, alignedDequeue_bits_data_lo_lo_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_1 = {unalignedCacheLine_bits_data[73], unalignedCacheLine_bits_data[65]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_1 = {unalignedCacheLine_bits_data[89], unalignedCacheLine_bits_data[81]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_1 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_1, alignedDequeue_bits_data_lo_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_1 = {unalignedCacheLine_bits_data[105], unalignedCacheLine_bits_data[97]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_1 = {unalignedCacheLine_bits_data[121], unalignedCacheLine_bits_data[113]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_1 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_1, alignedDequeue_bits_data_lo_lo_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_1 = {alignedDequeue_bits_data_lo_lo_hi_hi_1, alignedDequeue_bits_data_lo_lo_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_1 = {alignedDequeue_bits_data_lo_lo_hi_1, alignedDequeue_bits_data_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_1 = {unalignedCacheLine_bits_data[137], unalignedCacheLine_bits_data[129]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_1 = {unalignedCacheLine_bits_data[153], unalignedCacheLine_bits_data[145]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_1 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_1, alignedDequeue_bits_data_lo_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_1 = {unalignedCacheLine_bits_data[169], unalignedCacheLine_bits_data[161]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_1 = {unalignedCacheLine_bits_data[185], unalignedCacheLine_bits_data[177]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_1 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_1, alignedDequeue_bits_data_lo_hi_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_1 = {alignedDequeue_bits_data_lo_hi_lo_hi_1, alignedDequeue_bits_data_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_1 = {unalignedCacheLine_bits_data[201], unalignedCacheLine_bits_data[193]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_1 = {unalignedCacheLine_bits_data[217], unalignedCacheLine_bits_data[209]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_1 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_1, alignedDequeue_bits_data_lo_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_1 = {unalignedCacheLine_bits_data[233], unalignedCacheLine_bits_data[225]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_1 = {unalignedCacheLine_bits_data[249], unalignedCacheLine_bits_data[241]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_1, alignedDequeue_bits_data_lo_hi_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_hi_1, alignedDequeue_bits_data_lo_hi_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_1 = {alignedDequeue_bits_data_lo_hi_hi_1, alignedDequeue_bits_data_lo_hi_lo_1};
  wire [31:0]   alignedDequeue_bits_data_lo_1 = {alignedDequeue_bits_data_lo_hi_1, alignedDequeue_bits_data_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_1 = {memResponse_bits_data_0[9], memResponse_bits_data_0[1]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_1 = {memResponse_bits_data_0[25], memResponse_bits_data_0[17]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_1 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_1 = {memResponse_bits_data_0[41], memResponse_bits_data_0[33]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_1 = {memResponse_bits_data_0[57], memResponse_bits_data_0[49]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_1 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_1, alignedDequeue_bits_data_hi_lo_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_1 = {alignedDequeue_bits_data_hi_lo_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_1 = {memResponse_bits_data_0[73], memResponse_bits_data_0[65]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_1 = {memResponse_bits_data_0[89], memResponse_bits_data_0[81]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_1 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_1, alignedDequeue_bits_data_hi_lo_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_1 = {memResponse_bits_data_0[105], memResponse_bits_data_0[97]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_1 = {memResponse_bits_data_0[121], memResponse_bits_data_0[113]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_1 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_1, alignedDequeue_bits_data_hi_lo_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_1 = {alignedDequeue_bits_data_hi_lo_hi_hi_1, alignedDequeue_bits_data_hi_lo_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_1 = {alignedDequeue_bits_data_hi_lo_hi_1, alignedDequeue_bits_data_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_1 = {memResponse_bits_data_0[137], memResponse_bits_data_0[129]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_1 = {memResponse_bits_data_0[153], memResponse_bits_data_0[145]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_1 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_1, alignedDequeue_bits_data_hi_hi_lo_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_1 = {memResponse_bits_data_0[169], memResponse_bits_data_0[161]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_1 = {memResponse_bits_data_0[185], memResponse_bits_data_0[177]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_1 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_1, alignedDequeue_bits_data_hi_hi_lo_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_1 = {alignedDequeue_bits_data_hi_hi_lo_hi_1, alignedDequeue_bits_data_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_1 = {memResponse_bits_data_0[201], memResponse_bits_data_0[193]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_1 = {memResponse_bits_data_0[217], memResponse_bits_data_0[209]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_1 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_1, alignedDequeue_bits_data_hi_hi_hi_lo_lo_1};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_1 = {memResponse_bits_data_0[233], memResponse_bits_data_0[225]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_1 = {memResponse_bits_data_0[249], memResponse_bits_data_0[241]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_hi_hi_lo_1};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_hi_lo_1};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_1 = {alignedDequeue_bits_data_hi_hi_hi_1, alignedDequeue_bits_data_hi_hi_lo_1};
  wire [31:0]   alignedDequeue_bits_data_hi_1 = {alignedDequeue_bits_data_hi_hi_1, alignedDequeue_bits_data_hi_lo_1};
  wire [63:0]   _alignedDequeue_bits_data_T_580 = {alignedDequeue_bits_data_hi_1, alignedDequeue_bits_data_lo_1} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_2 = {unalignedCacheLine_bits_data[10], unalignedCacheLine_bits_data[2]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_2 = {unalignedCacheLine_bits_data[26], unalignedCacheLine_bits_data[18]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_2 = {unalignedCacheLine_bits_data[42], unalignedCacheLine_bits_data[34]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_2 = {unalignedCacheLine_bits_data[58], unalignedCacheLine_bits_data[50]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_2 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_2, alignedDequeue_bits_data_lo_lo_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_2 = {unalignedCacheLine_bits_data[74], unalignedCacheLine_bits_data[66]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_2 = {unalignedCacheLine_bits_data[90], unalignedCacheLine_bits_data[82]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_2 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_2, alignedDequeue_bits_data_lo_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_2 = {unalignedCacheLine_bits_data[106], unalignedCacheLine_bits_data[98]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_2 = {unalignedCacheLine_bits_data[122], unalignedCacheLine_bits_data[114]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_2 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_2, alignedDequeue_bits_data_lo_lo_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_2 = {alignedDequeue_bits_data_lo_lo_hi_hi_2, alignedDequeue_bits_data_lo_lo_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_2 = {alignedDequeue_bits_data_lo_lo_hi_2, alignedDequeue_bits_data_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_2 = {unalignedCacheLine_bits_data[138], unalignedCacheLine_bits_data[130]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_2 = {unalignedCacheLine_bits_data[154], unalignedCacheLine_bits_data[146]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_2 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_2, alignedDequeue_bits_data_lo_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_2 = {unalignedCacheLine_bits_data[170], unalignedCacheLine_bits_data[162]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_2 = {unalignedCacheLine_bits_data[186], unalignedCacheLine_bits_data[178]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_2 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_2, alignedDequeue_bits_data_lo_hi_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_2 = {alignedDequeue_bits_data_lo_hi_lo_hi_2, alignedDequeue_bits_data_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_2 = {unalignedCacheLine_bits_data[202], unalignedCacheLine_bits_data[194]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_2 = {unalignedCacheLine_bits_data[218], unalignedCacheLine_bits_data[210]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_2 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_2, alignedDequeue_bits_data_lo_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_2 = {unalignedCacheLine_bits_data[234], unalignedCacheLine_bits_data[226]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_2 = {unalignedCacheLine_bits_data[250], unalignedCacheLine_bits_data[242]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_2, alignedDequeue_bits_data_lo_hi_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_hi_2, alignedDequeue_bits_data_lo_hi_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_2 = {alignedDequeue_bits_data_lo_hi_hi_2, alignedDequeue_bits_data_lo_hi_lo_2};
  wire [31:0]   alignedDequeue_bits_data_lo_2 = {alignedDequeue_bits_data_lo_hi_2, alignedDequeue_bits_data_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_2 = {memResponse_bits_data_0[10], memResponse_bits_data_0[2]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_2 = {memResponse_bits_data_0[26], memResponse_bits_data_0[18]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_2 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_2 = {memResponse_bits_data_0[42], memResponse_bits_data_0[34]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_2 = {memResponse_bits_data_0[58], memResponse_bits_data_0[50]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_2 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_2, alignedDequeue_bits_data_hi_lo_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_2 = {alignedDequeue_bits_data_hi_lo_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_2 = {memResponse_bits_data_0[74], memResponse_bits_data_0[66]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_2 = {memResponse_bits_data_0[90], memResponse_bits_data_0[82]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_2 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_2, alignedDequeue_bits_data_hi_lo_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_2 = {memResponse_bits_data_0[106], memResponse_bits_data_0[98]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_2 = {memResponse_bits_data_0[122], memResponse_bits_data_0[114]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_2 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_2, alignedDequeue_bits_data_hi_lo_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_2 = {alignedDequeue_bits_data_hi_lo_hi_hi_2, alignedDequeue_bits_data_hi_lo_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_2 = {alignedDequeue_bits_data_hi_lo_hi_2, alignedDequeue_bits_data_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_2 = {memResponse_bits_data_0[138], memResponse_bits_data_0[130]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_2 = {memResponse_bits_data_0[154], memResponse_bits_data_0[146]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_2 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_2, alignedDequeue_bits_data_hi_hi_lo_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_2 = {memResponse_bits_data_0[170], memResponse_bits_data_0[162]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_2 = {memResponse_bits_data_0[186], memResponse_bits_data_0[178]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_2 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_2, alignedDequeue_bits_data_hi_hi_lo_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_2 = {alignedDequeue_bits_data_hi_hi_lo_hi_2, alignedDequeue_bits_data_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_2 = {memResponse_bits_data_0[202], memResponse_bits_data_0[194]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_2 = {memResponse_bits_data_0[218], memResponse_bits_data_0[210]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_2 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_2, alignedDequeue_bits_data_hi_hi_hi_lo_lo_2};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_2 = {memResponse_bits_data_0[234], memResponse_bits_data_0[226]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_2 = {memResponse_bits_data_0[250], memResponse_bits_data_0[242]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_hi_hi_lo_2};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_hi_lo_2};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_2 = {alignedDequeue_bits_data_hi_hi_hi_2, alignedDequeue_bits_data_hi_hi_lo_2};
  wire [31:0]   alignedDequeue_bits_data_hi_2 = {alignedDequeue_bits_data_hi_hi_2, alignedDequeue_bits_data_hi_lo_2};
  wire [63:0]   _alignedDequeue_bits_data_T_646 = {alignedDequeue_bits_data_hi_2, alignedDequeue_bits_data_lo_2} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_3 = {unalignedCacheLine_bits_data[11], unalignedCacheLine_bits_data[3]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_3 = {unalignedCacheLine_bits_data[27], unalignedCacheLine_bits_data[19]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_3 = {unalignedCacheLine_bits_data[43], unalignedCacheLine_bits_data[35]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_3 = {unalignedCacheLine_bits_data[59], unalignedCacheLine_bits_data[51]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_3 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_3, alignedDequeue_bits_data_lo_lo_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_3 = {unalignedCacheLine_bits_data[75], unalignedCacheLine_bits_data[67]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_3 = {unalignedCacheLine_bits_data[91], unalignedCacheLine_bits_data[83]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_3 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_3, alignedDequeue_bits_data_lo_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_3 = {unalignedCacheLine_bits_data[107], unalignedCacheLine_bits_data[99]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_3 = {unalignedCacheLine_bits_data[123], unalignedCacheLine_bits_data[115]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_3 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_3, alignedDequeue_bits_data_lo_lo_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_3 = {alignedDequeue_bits_data_lo_lo_hi_hi_3, alignedDequeue_bits_data_lo_lo_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_3 = {alignedDequeue_bits_data_lo_lo_hi_3, alignedDequeue_bits_data_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_3 = {unalignedCacheLine_bits_data[139], unalignedCacheLine_bits_data[131]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_3 = {unalignedCacheLine_bits_data[155], unalignedCacheLine_bits_data[147]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_3 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_3, alignedDequeue_bits_data_lo_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_3 = {unalignedCacheLine_bits_data[171], unalignedCacheLine_bits_data[163]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_3 = {unalignedCacheLine_bits_data[187], unalignedCacheLine_bits_data[179]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_3 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_3, alignedDequeue_bits_data_lo_hi_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_3 = {alignedDequeue_bits_data_lo_hi_lo_hi_3, alignedDequeue_bits_data_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_3 = {unalignedCacheLine_bits_data[203], unalignedCacheLine_bits_data[195]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_3 = {unalignedCacheLine_bits_data[219], unalignedCacheLine_bits_data[211]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_3 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_3, alignedDequeue_bits_data_lo_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_3 = {unalignedCacheLine_bits_data[235], unalignedCacheLine_bits_data[227]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_3 = {unalignedCacheLine_bits_data[251], unalignedCacheLine_bits_data[243]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_3, alignedDequeue_bits_data_lo_hi_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_hi_3, alignedDequeue_bits_data_lo_hi_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_3 = {alignedDequeue_bits_data_lo_hi_hi_3, alignedDequeue_bits_data_lo_hi_lo_3};
  wire [31:0]   alignedDequeue_bits_data_lo_3 = {alignedDequeue_bits_data_lo_hi_3, alignedDequeue_bits_data_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_3 = {memResponse_bits_data_0[11], memResponse_bits_data_0[3]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_3 = {memResponse_bits_data_0[27], memResponse_bits_data_0[19]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_3 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_3 = {memResponse_bits_data_0[43], memResponse_bits_data_0[35]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_3 = {memResponse_bits_data_0[59], memResponse_bits_data_0[51]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_3 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_3, alignedDequeue_bits_data_hi_lo_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_3 = {alignedDequeue_bits_data_hi_lo_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_3 = {memResponse_bits_data_0[75], memResponse_bits_data_0[67]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_3 = {memResponse_bits_data_0[91], memResponse_bits_data_0[83]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_3 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_3, alignedDequeue_bits_data_hi_lo_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_3 = {memResponse_bits_data_0[107], memResponse_bits_data_0[99]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_3 = {memResponse_bits_data_0[123], memResponse_bits_data_0[115]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_3 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_3, alignedDequeue_bits_data_hi_lo_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_3 = {alignedDequeue_bits_data_hi_lo_hi_hi_3, alignedDequeue_bits_data_hi_lo_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_3 = {alignedDequeue_bits_data_hi_lo_hi_3, alignedDequeue_bits_data_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_3 = {memResponse_bits_data_0[139], memResponse_bits_data_0[131]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_3 = {memResponse_bits_data_0[155], memResponse_bits_data_0[147]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_3 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_3, alignedDequeue_bits_data_hi_hi_lo_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_3 = {memResponse_bits_data_0[171], memResponse_bits_data_0[163]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_3 = {memResponse_bits_data_0[187], memResponse_bits_data_0[179]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_3 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_3, alignedDequeue_bits_data_hi_hi_lo_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_3 = {alignedDequeue_bits_data_hi_hi_lo_hi_3, alignedDequeue_bits_data_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_3 = {memResponse_bits_data_0[203], memResponse_bits_data_0[195]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_3 = {memResponse_bits_data_0[219], memResponse_bits_data_0[211]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_3 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_3, alignedDequeue_bits_data_hi_hi_hi_lo_lo_3};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_3 = {memResponse_bits_data_0[235], memResponse_bits_data_0[227]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_3 = {memResponse_bits_data_0[251], memResponse_bits_data_0[243]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_hi_hi_lo_3};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_hi_lo_3};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_3 = {alignedDequeue_bits_data_hi_hi_hi_3, alignedDequeue_bits_data_hi_hi_lo_3};
  wire [31:0]   alignedDequeue_bits_data_hi_3 = {alignedDequeue_bits_data_hi_hi_3, alignedDequeue_bits_data_hi_lo_3};
  wire [63:0]   _alignedDequeue_bits_data_T_712 = {alignedDequeue_bits_data_hi_3, alignedDequeue_bits_data_lo_3} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_4 = {unalignedCacheLine_bits_data[12], unalignedCacheLine_bits_data[4]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_4 = {unalignedCacheLine_bits_data[28], unalignedCacheLine_bits_data[20]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_4 = {unalignedCacheLine_bits_data[44], unalignedCacheLine_bits_data[36]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_4 = {unalignedCacheLine_bits_data[60], unalignedCacheLine_bits_data[52]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_4 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_4, alignedDequeue_bits_data_lo_lo_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_4 = {unalignedCacheLine_bits_data[76], unalignedCacheLine_bits_data[68]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_4 = {unalignedCacheLine_bits_data[92], unalignedCacheLine_bits_data[84]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_4 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_4, alignedDequeue_bits_data_lo_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_4 = {unalignedCacheLine_bits_data[108], unalignedCacheLine_bits_data[100]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_4 = {unalignedCacheLine_bits_data[124], unalignedCacheLine_bits_data[116]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_4 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_4, alignedDequeue_bits_data_lo_lo_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_4 = {alignedDequeue_bits_data_lo_lo_hi_hi_4, alignedDequeue_bits_data_lo_lo_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_4 = {alignedDequeue_bits_data_lo_lo_hi_4, alignedDequeue_bits_data_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_4 = {unalignedCacheLine_bits_data[140], unalignedCacheLine_bits_data[132]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_4 = {unalignedCacheLine_bits_data[156], unalignedCacheLine_bits_data[148]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_4 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_4, alignedDequeue_bits_data_lo_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_4 = {unalignedCacheLine_bits_data[172], unalignedCacheLine_bits_data[164]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_4 = {unalignedCacheLine_bits_data[188], unalignedCacheLine_bits_data[180]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_4 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_4, alignedDequeue_bits_data_lo_hi_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_4 = {alignedDequeue_bits_data_lo_hi_lo_hi_4, alignedDequeue_bits_data_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_4 = {unalignedCacheLine_bits_data[204], unalignedCacheLine_bits_data[196]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_4 = {unalignedCacheLine_bits_data[220], unalignedCacheLine_bits_data[212]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_4 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_4, alignedDequeue_bits_data_lo_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_4 = {unalignedCacheLine_bits_data[236], unalignedCacheLine_bits_data[228]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_4 = {unalignedCacheLine_bits_data[252], unalignedCacheLine_bits_data[244]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_4, alignedDequeue_bits_data_lo_hi_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_hi_4, alignedDequeue_bits_data_lo_hi_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_4 = {alignedDequeue_bits_data_lo_hi_hi_4, alignedDequeue_bits_data_lo_hi_lo_4};
  wire [31:0]   alignedDequeue_bits_data_lo_4 = {alignedDequeue_bits_data_lo_hi_4, alignedDequeue_bits_data_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_4 = {memResponse_bits_data_0[12], memResponse_bits_data_0[4]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_4 = {memResponse_bits_data_0[28], memResponse_bits_data_0[20]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_4 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_4 = {memResponse_bits_data_0[44], memResponse_bits_data_0[36]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_4 = {memResponse_bits_data_0[60], memResponse_bits_data_0[52]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_4 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_4, alignedDequeue_bits_data_hi_lo_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_4 = {alignedDequeue_bits_data_hi_lo_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_4 = {memResponse_bits_data_0[76], memResponse_bits_data_0[68]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_4 = {memResponse_bits_data_0[92], memResponse_bits_data_0[84]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_4 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_4, alignedDequeue_bits_data_hi_lo_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_4 = {memResponse_bits_data_0[108], memResponse_bits_data_0[100]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_4 = {memResponse_bits_data_0[124], memResponse_bits_data_0[116]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_4 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_4, alignedDequeue_bits_data_hi_lo_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_4 = {alignedDequeue_bits_data_hi_lo_hi_hi_4, alignedDequeue_bits_data_hi_lo_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_4 = {alignedDequeue_bits_data_hi_lo_hi_4, alignedDequeue_bits_data_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_4 = {memResponse_bits_data_0[140], memResponse_bits_data_0[132]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_4 = {memResponse_bits_data_0[156], memResponse_bits_data_0[148]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_4 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_4, alignedDequeue_bits_data_hi_hi_lo_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_4 = {memResponse_bits_data_0[172], memResponse_bits_data_0[164]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_4 = {memResponse_bits_data_0[188], memResponse_bits_data_0[180]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_4 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_4, alignedDequeue_bits_data_hi_hi_lo_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_4 = {alignedDequeue_bits_data_hi_hi_lo_hi_4, alignedDequeue_bits_data_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_4 = {memResponse_bits_data_0[204], memResponse_bits_data_0[196]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_4 = {memResponse_bits_data_0[220], memResponse_bits_data_0[212]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_4 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_4, alignedDequeue_bits_data_hi_hi_hi_lo_lo_4};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_4 = {memResponse_bits_data_0[236], memResponse_bits_data_0[228]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_4 = {memResponse_bits_data_0[252], memResponse_bits_data_0[244]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_hi_hi_lo_4};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_hi_lo_4};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_4 = {alignedDequeue_bits_data_hi_hi_hi_4, alignedDequeue_bits_data_hi_hi_lo_4};
  wire [31:0]   alignedDequeue_bits_data_hi_4 = {alignedDequeue_bits_data_hi_hi_4, alignedDequeue_bits_data_hi_lo_4};
  wire [63:0]   _alignedDequeue_bits_data_T_778 = {alignedDequeue_bits_data_hi_4, alignedDequeue_bits_data_lo_4} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_5 = {unalignedCacheLine_bits_data[13], unalignedCacheLine_bits_data[5]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_5 = {unalignedCacheLine_bits_data[29], unalignedCacheLine_bits_data[21]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_5 = {unalignedCacheLine_bits_data[45], unalignedCacheLine_bits_data[37]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_5 = {unalignedCacheLine_bits_data[61], unalignedCacheLine_bits_data[53]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_5 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_5, alignedDequeue_bits_data_lo_lo_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_5 = {unalignedCacheLine_bits_data[77], unalignedCacheLine_bits_data[69]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_5 = {unalignedCacheLine_bits_data[93], unalignedCacheLine_bits_data[85]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_5 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_5, alignedDequeue_bits_data_lo_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_5 = {unalignedCacheLine_bits_data[109], unalignedCacheLine_bits_data[101]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_5 = {unalignedCacheLine_bits_data[125], unalignedCacheLine_bits_data[117]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_5 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_5, alignedDequeue_bits_data_lo_lo_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_5 = {alignedDequeue_bits_data_lo_lo_hi_hi_5, alignedDequeue_bits_data_lo_lo_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_5 = {alignedDequeue_bits_data_lo_lo_hi_5, alignedDequeue_bits_data_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_5 = {unalignedCacheLine_bits_data[141], unalignedCacheLine_bits_data[133]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_5 = {unalignedCacheLine_bits_data[157], unalignedCacheLine_bits_data[149]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_5 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_5, alignedDequeue_bits_data_lo_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_5 = {unalignedCacheLine_bits_data[173], unalignedCacheLine_bits_data[165]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_5 = {unalignedCacheLine_bits_data[189], unalignedCacheLine_bits_data[181]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_5 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_5, alignedDequeue_bits_data_lo_hi_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_5 = {alignedDequeue_bits_data_lo_hi_lo_hi_5, alignedDequeue_bits_data_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_5 = {unalignedCacheLine_bits_data[205], unalignedCacheLine_bits_data[197]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_5 = {unalignedCacheLine_bits_data[221], unalignedCacheLine_bits_data[213]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_5 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_5, alignedDequeue_bits_data_lo_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_5 = {unalignedCacheLine_bits_data[237], unalignedCacheLine_bits_data[229]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_5 = {unalignedCacheLine_bits_data[253], unalignedCacheLine_bits_data[245]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_5, alignedDequeue_bits_data_lo_hi_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_hi_5, alignedDequeue_bits_data_lo_hi_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_5 = {alignedDequeue_bits_data_lo_hi_hi_5, alignedDequeue_bits_data_lo_hi_lo_5};
  wire [31:0]   alignedDequeue_bits_data_lo_5 = {alignedDequeue_bits_data_lo_hi_5, alignedDequeue_bits_data_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_5 = {memResponse_bits_data_0[13], memResponse_bits_data_0[5]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_5 = {memResponse_bits_data_0[29], memResponse_bits_data_0[21]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_5 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_5 = {memResponse_bits_data_0[45], memResponse_bits_data_0[37]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_5 = {memResponse_bits_data_0[61], memResponse_bits_data_0[53]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_5 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_5, alignedDequeue_bits_data_hi_lo_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_5 = {alignedDequeue_bits_data_hi_lo_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_5 = {memResponse_bits_data_0[77], memResponse_bits_data_0[69]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_5 = {memResponse_bits_data_0[93], memResponse_bits_data_0[85]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_5 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_5, alignedDequeue_bits_data_hi_lo_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_5 = {memResponse_bits_data_0[109], memResponse_bits_data_0[101]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_5 = {memResponse_bits_data_0[125], memResponse_bits_data_0[117]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_5 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_5, alignedDequeue_bits_data_hi_lo_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_5 = {alignedDequeue_bits_data_hi_lo_hi_hi_5, alignedDequeue_bits_data_hi_lo_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_5 = {alignedDequeue_bits_data_hi_lo_hi_5, alignedDequeue_bits_data_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_5 = {memResponse_bits_data_0[141], memResponse_bits_data_0[133]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_5 = {memResponse_bits_data_0[157], memResponse_bits_data_0[149]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_5 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_5, alignedDequeue_bits_data_hi_hi_lo_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_5 = {memResponse_bits_data_0[173], memResponse_bits_data_0[165]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_5 = {memResponse_bits_data_0[189], memResponse_bits_data_0[181]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_5 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_5, alignedDequeue_bits_data_hi_hi_lo_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_5 = {alignedDequeue_bits_data_hi_hi_lo_hi_5, alignedDequeue_bits_data_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_5 = {memResponse_bits_data_0[205], memResponse_bits_data_0[197]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_5 = {memResponse_bits_data_0[221], memResponse_bits_data_0[213]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_5 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_5, alignedDequeue_bits_data_hi_hi_hi_lo_lo_5};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_5 = {memResponse_bits_data_0[237], memResponse_bits_data_0[229]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_5 = {memResponse_bits_data_0[253], memResponse_bits_data_0[245]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_hi_hi_lo_5};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_hi_lo_5};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_5 = {alignedDequeue_bits_data_hi_hi_hi_5, alignedDequeue_bits_data_hi_hi_lo_5};
  wire [31:0]   alignedDequeue_bits_data_hi_5 = {alignedDequeue_bits_data_hi_hi_5, alignedDequeue_bits_data_hi_lo_5};
  wire [63:0]   _alignedDequeue_bits_data_T_844 = {alignedDequeue_bits_data_hi_5, alignedDequeue_bits_data_lo_5} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_6 = {unalignedCacheLine_bits_data[14], unalignedCacheLine_bits_data[6]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_6 = {unalignedCacheLine_bits_data[30], unalignedCacheLine_bits_data[22]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_6 = {unalignedCacheLine_bits_data[46], unalignedCacheLine_bits_data[38]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_6 = {unalignedCacheLine_bits_data[62], unalignedCacheLine_bits_data[54]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_6 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_6, alignedDequeue_bits_data_lo_lo_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_6 = {unalignedCacheLine_bits_data[78], unalignedCacheLine_bits_data[70]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_6 = {unalignedCacheLine_bits_data[94], unalignedCacheLine_bits_data[86]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_6 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_6, alignedDequeue_bits_data_lo_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_6 = {unalignedCacheLine_bits_data[110], unalignedCacheLine_bits_data[102]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_6 = {unalignedCacheLine_bits_data[126], unalignedCacheLine_bits_data[118]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_6 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_6, alignedDequeue_bits_data_lo_lo_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_6 = {alignedDequeue_bits_data_lo_lo_hi_hi_6, alignedDequeue_bits_data_lo_lo_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_6 = {alignedDequeue_bits_data_lo_lo_hi_6, alignedDequeue_bits_data_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_6 = {unalignedCacheLine_bits_data[142], unalignedCacheLine_bits_data[134]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_6 = {unalignedCacheLine_bits_data[158], unalignedCacheLine_bits_data[150]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_6 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_6, alignedDequeue_bits_data_lo_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_6 = {unalignedCacheLine_bits_data[174], unalignedCacheLine_bits_data[166]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_6 = {unalignedCacheLine_bits_data[190], unalignedCacheLine_bits_data[182]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_6 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_6, alignedDequeue_bits_data_lo_hi_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_6 = {alignedDequeue_bits_data_lo_hi_lo_hi_6, alignedDequeue_bits_data_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_6 = {unalignedCacheLine_bits_data[206], unalignedCacheLine_bits_data[198]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_6 = {unalignedCacheLine_bits_data[222], unalignedCacheLine_bits_data[214]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_6 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_6, alignedDequeue_bits_data_lo_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_6 = {unalignedCacheLine_bits_data[238], unalignedCacheLine_bits_data[230]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_6 = {unalignedCacheLine_bits_data[254], unalignedCacheLine_bits_data[246]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_6, alignedDequeue_bits_data_lo_hi_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_hi_6, alignedDequeue_bits_data_lo_hi_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_6 = {alignedDequeue_bits_data_lo_hi_hi_6, alignedDequeue_bits_data_lo_hi_lo_6};
  wire [31:0]   alignedDequeue_bits_data_lo_6 = {alignedDequeue_bits_data_lo_hi_6, alignedDequeue_bits_data_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_6 = {memResponse_bits_data_0[14], memResponse_bits_data_0[6]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_6 = {memResponse_bits_data_0[30], memResponse_bits_data_0[22]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_6 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_6 = {memResponse_bits_data_0[46], memResponse_bits_data_0[38]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_6 = {memResponse_bits_data_0[62], memResponse_bits_data_0[54]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_6 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_6, alignedDequeue_bits_data_hi_lo_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_6 = {alignedDequeue_bits_data_hi_lo_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_6 = {memResponse_bits_data_0[78], memResponse_bits_data_0[70]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_6 = {memResponse_bits_data_0[94], memResponse_bits_data_0[86]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_6 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_6, alignedDequeue_bits_data_hi_lo_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_6 = {memResponse_bits_data_0[110], memResponse_bits_data_0[102]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_6 = {memResponse_bits_data_0[126], memResponse_bits_data_0[118]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_6 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_6, alignedDequeue_bits_data_hi_lo_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_6 = {alignedDequeue_bits_data_hi_lo_hi_hi_6, alignedDequeue_bits_data_hi_lo_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_6 = {alignedDequeue_bits_data_hi_lo_hi_6, alignedDequeue_bits_data_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_6 = {memResponse_bits_data_0[142], memResponse_bits_data_0[134]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_6 = {memResponse_bits_data_0[158], memResponse_bits_data_0[150]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_6 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_6, alignedDequeue_bits_data_hi_hi_lo_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_6 = {memResponse_bits_data_0[174], memResponse_bits_data_0[166]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_6 = {memResponse_bits_data_0[190], memResponse_bits_data_0[182]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_6 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_6, alignedDequeue_bits_data_hi_hi_lo_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_6 = {alignedDequeue_bits_data_hi_hi_lo_hi_6, alignedDequeue_bits_data_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_6 = {memResponse_bits_data_0[206], memResponse_bits_data_0[198]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_6 = {memResponse_bits_data_0[222], memResponse_bits_data_0[214]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_6 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_6, alignedDequeue_bits_data_hi_hi_hi_lo_lo_6};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_6 = {memResponse_bits_data_0[238], memResponse_bits_data_0[230]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_6 = {memResponse_bits_data_0[254], memResponse_bits_data_0[246]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_hi_hi_lo_6};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_hi_lo_6};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_6 = {alignedDequeue_bits_data_hi_hi_hi_6, alignedDequeue_bits_data_hi_hi_lo_6};
  wire [31:0]   alignedDequeue_bits_data_hi_6 = {alignedDequeue_bits_data_hi_hi_6, alignedDequeue_bits_data_hi_lo_6};
  wire [63:0]   _alignedDequeue_bits_data_T_910 = {alignedDequeue_bits_data_hi_6, alignedDequeue_bits_data_lo_6} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_lo_7 = {unalignedCacheLine_bits_data[15], unalignedCacheLine_bits_data[7]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_lo_hi_7 = {unalignedCacheLine_bits_data[31], unalignedCacheLine_bits_data[23]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_lo_7 = {unalignedCacheLine_bits_data[47], unalignedCacheLine_bits_data[39]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_lo_hi_hi_7 = {unalignedCacheLine_bits_data[63], unalignedCacheLine_bits_data[55]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_lo_hi_7 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_7, alignedDequeue_bits_data_lo_lo_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_lo_7 = {unalignedCacheLine_bits_data[79], unalignedCacheLine_bits_data[71]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_lo_hi_7 = {unalignedCacheLine_bits_data[95], unalignedCacheLine_bits_data[87]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_lo_7 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_7, alignedDequeue_bits_data_lo_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_lo_7 = {unalignedCacheLine_bits_data[111], unalignedCacheLine_bits_data[103]};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_hi_hi_hi_7 = {unalignedCacheLine_bits_data[127], unalignedCacheLine_bits_data[119]};
  wire [3:0]    alignedDequeue_bits_data_lo_lo_hi_hi_7 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_7, alignedDequeue_bits_data_lo_lo_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_lo_hi_7 = {alignedDequeue_bits_data_lo_lo_hi_hi_7, alignedDequeue_bits_data_lo_lo_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_7 = {alignedDequeue_bits_data_lo_lo_hi_7, alignedDequeue_bits_data_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_lo_7 = {unalignedCacheLine_bits_data[143], unalignedCacheLine_bits_data[135]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_lo_hi_7 = {unalignedCacheLine_bits_data[159], unalignedCacheLine_bits_data[151]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_lo_7 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_7, alignedDequeue_bits_data_lo_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_lo_7 = {unalignedCacheLine_bits_data[175], unalignedCacheLine_bits_data[167]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_lo_hi_hi_7 = {unalignedCacheLine_bits_data[191], unalignedCacheLine_bits_data[183]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_lo_hi_7 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_7, alignedDequeue_bits_data_lo_hi_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_lo_7 = {alignedDequeue_bits_data_lo_hi_lo_hi_7, alignedDequeue_bits_data_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_lo_7 = {unalignedCacheLine_bits_data[207], unalignedCacheLine_bits_data[199]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_lo_hi_7 = {unalignedCacheLine_bits_data[223], unalignedCacheLine_bits_data[215]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_lo_7 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_7, alignedDequeue_bits_data_lo_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_lo_7 = {unalignedCacheLine_bits_data[239], unalignedCacheLine_bits_data[231]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_hi_hi_hi_7 = {unalignedCacheLine_bits_data[255], unalignedCacheLine_bits_data[247]};
  wire [3:0]    alignedDequeue_bits_data_lo_hi_hi_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_7, alignedDequeue_bits_data_lo_hi_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_lo_hi_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_hi_7, alignedDequeue_bits_data_lo_hi_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_7 = {alignedDequeue_bits_data_lo_hi_hi_7, alignedDequeue_bits_data_lo_hi_lo_7};
  wire [31:0]   alignedDequeue_bits_data_lo_7 = {alignedDequeue_bits_data_lo_hi_7, alignedDequeue_bits_data_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_lo_7 = {memResponse_bits_data_0[15], memResponse_bits_data_0[7]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_lo_hi_7 = {memResponse_bits_data_0[31], memResponse_bits_data_0[23]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_lo_7 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_lo_7 = {memResponse_bits_data_0[47], memResponse_bits_data_0[39]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_lo_hi_hi_7 = {memResponse_bits_data_0[63], memResponse_bits_data_0[55]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_lo_hi_7 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_7, alignedDequeue_bits_data_hi_lo_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_lo_7 = {alignedDequeue_bits_data_hi_lo_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_lo_7 = {memResponse_bits_data_0[79], memResponse_bits_data_0[71]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_lo_hi_7 = {memResponse_bits_data_0[95], memResponse_bits_data_0[87]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_lo_7 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_7, alignedDequeue_bits_data_hi_lo_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_lo_7 = {memResponse_bits_data_0[111], memResponse_bits_data_0[103]};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_hi_hi_hi_7 = {memResponse_bits_data_0[127], memResponse_bits_data_0[119]};
  wire [3:0]    alignedDequeue_bits_data_hi_lo_hi_hi_7 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_7, alignedDequeue_bits_data_hi_lo_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_lo_hi_7 = {alignedDequeue_bits_data_hi_lo_hi_hi_7, alignedDequeue_bits_data_hi_lo_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_7 = {alignedDequeue_bits_data_hi_lo_hi_7, alignedDequeue_bits_data_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_lo_7 = {memResponse_bits_data_0[143], memResponse_bits_data_0[135]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_lo_hi_7 = {memResponse_bits_data_0[159], memResponse_bits_data_0[151]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_lo_7 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_7, alignedDequeue_bits_data_hi_hi_lo_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_lo_7 = {memResponse_bits_data_0[175], memResponse_bits_data_0[167]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_lo_hi_hi_7 = {memResponse_bits_data_0[191], memResponse_bits_data_0[183]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_lo_hi_7 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_7, alignedDequeue_bits_data_hi_hi_lo_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_lo_7 = {alignedDequeue_bits_data_hi_hi_lo_hi_7, alignedDequeue_bits_data_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_lo_7 = {memResponse_bits_data_0[207], memResponse_bits_data_0[199]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_lo_hi_7 = {memResponse_bits_data_0[223], memResponse_bits_data_0[215]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_lo_7 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_7, alignedDequeue_bits_data_hi_hi_hi_lo_lo_7};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_lo_7 = {memResponse_bits_data_0[239], memResponse_bits_data_0[231]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_hi_hi_hi_7 = {memResponse_bits_data_0[255], memResponse_bits_data_0[247]};
  wire [3:0]    alignedDequeue_bits_data_hi_hi_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_hi_hi_lo_7};
  wire [7:0]    alignedDequeue_bits_data_hi_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_hi_lo_7};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_7 = {alignedDequeue_bits_data_hi_hi_hi_7, alignedDequeue_bits_data_hi_hi_lo_7};
  wire [31:0]   alignedDequeue_bits_data_hi_7 = {alignedDequeue_bits_data_hi_hi_7, alignedDequeue_bits_data_hi_lo_7};
  wire [63:0]   _alignedDequeue_bits_data_T_976 = {alignedDequeue_bits_data_hi_7, alignedDequeue_bits_data_lo_7} >> _GEN_3;
  wire [1:0]    alignedDequeue_bits_data_lo_lo_8 = {_alignedDequeue_bits_data_T_580[0], _alignedDequeue_bits_data_T_514[0]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_8 = {_alignedDequeue_bits_data_T_712[0], _alignedDequeue_bits_data_T_646[0]};
  wire [3:0]    alignedDequeue_bits_data_lo_8 = {alignedDequeue_bits_data_lo_hi_8, alignedDequeue_bits_data_lo_lo_8};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_8 = {_alignedDequeue_bits_data_T_844[0], _alignedDequeue_bits_data_T_778[0]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_8 = {_alignedDequeue_bits_data_T_976[0], _alignedDequeue_bits_data_T_910[0]};
  wire [3:0]    alignedDequeue_bits_data_hi_8 = {alignedDequeue_bits_data_hi_hi_8, alignedDequeue_bits_data_hi_lo_8};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_9 = {_alignedDequeue_bits_data_T_580[1], _alignedDequeue_bits_data_T_514[1]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_9 = {_alignedDequeue_bits_data_T_712[1], _alignedDequeue_bits_data_T_646[1]};
  wire [3:0]    alignedDequeue_bits_data_lo_9 = {alignedDequeue_bits_data_lo_hi_9, alignedDequeue_bits_data_lo_lo_9};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_9 = {_alignedDequeue_bits_data_T_844[1], _alignedDequeue_bits_data_T_778[1]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_9 = {_alignedDequeue_bits_data_T_976[1], _alignedDequeue_bits_data_T_910[1]};
  wire [3:0]    alignedDequeue_bits_data_hi_9 = {alignedDequeue_bits_data_hi_hi_9, alignedDequeue_bits_data_hi_lo_9};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_10 = {_alignedDequeue_bits_data_T_580[2], _alignedDequeue_bits_data_T_514[2]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_10 = {_alignedDequeue_bits_data_T_712[2], _alignedDequeue_bits_data_T_646[2]};
  wire [3:0]    alignedDequeue_bits_data_lo_10 = {alignedDequeue_bits_data_lo_hi_10, alignedDequeue_bits_data_lo_lo_10};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_10 = {_alignedDequeue_bits_data_T_844[2], _alignedDequeue_bits_data_T_778[2]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_10 = {_alignedDequeue_bits_data_T_976[2], _alignedDequeue_bits_data_T_910[2]};
  wire [3:0]    alignedDequeue_bits_data_hi_10 = {alignedDequeue_bits_data_hi_hi_10, alignedDequeue_bits_data_hi_lo_10};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_11 = {_alignedDequeue_bits_data_T_580[3], _alignedDequeue_bits_data_T_514[3]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_11 = {_alignedDequeue_bits_data_T_712[3], _alignedDequeue_bits_data_T_646[3]};
  wire [3:0]    alignedDequeue_bits_data_lo_11 = {alignedDequeue_bits_data_lo_hi_11, alignedDequeue_bits_data_lo_lo_11};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_11 = {_alignedDequeue_bits_data_T_844[3], _alignedDequeue_bits_data_T_778[3]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_11 = {_alignedDequeue_bits_data_T_976[3], _alignedDequeue_bits_data_T_910[3]};
  wire [3:0]    alignedDequeue_bits_data_hi_11 = {alignedDequeue_bits_data_hi_hi_11, alignedDequeue_bits_data_hi_lo_11};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_12 = {_alignedDequeue_bits_data_T_580[4], _alignedDequeue_bits_data_T_514[4]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_12 = {_alignedDequeue_bits_data_T_712[4], _alignedDequeue_bits_data_T_646[4]};
  wire [3:0]    alignedDequeue_bits_data_lo_12 = {alignedDequeue_bits_data_lo_hi_12, alignedDequeue_bits_data_lo_lo_12};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_12 = {_alignedDequeue_bits_data_T_844[4], _alignedDequeue_bits_data_T_778[4]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_12 = {_alignedDequeue_bits_data_T_976[4], _alignedDequeue_bits_data_T_910[4]};
  wire [3:0]    alignedDequeue_bits_data_hi_12 = {alignedDequeue_bits_data_hi_hi_12, alignedDequeue_bits_data_hi_lo_12};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_13 = {_alignedDequeue_bits_data_T_580[5], _alignedDequeue_bits_data_T_514[5]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_13 = {_alignedDequeue_bits_data_T_712[5], _alignedDequeue_bits_data_T_646[5]};
  wire [3:0]    alignedDequeue_bits_data_lo_13 = {alignedDequeue_bits_data_lo_hi_13, alignedDequeue_bits_data_lo_lo_13};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_13 = {_alignedDequeue_bits_data_T_844[5], _alignedDequeue_bits_data_T_778[5]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_13 = {_alignedDequeue_bits_data_T_976[5], _alignedDequeue_bits_data_T_910[5]};
  wire [3:0]    alignedDequeue_bits_data_hi_13 = {alignedDequeue_bits_data_hi_hi_13, alignedDequeue_bits_data_hi_lo_13};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_14 = {_alignedDequeue_bits_data_T_580[6], _alignedDequeue_bits_data_T_514[6]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_14 = {_alignedDequeue_bits_data_T_712[6], _alignedDequeue_bits_data_T_646[6]};
  wire [3:0]    alignedDequeue_bits_data_lo_14 = {alignedDequeue_bits_data_lo_hi_14, alignedDequeue_bits_data_lo_lo_14};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_14 = {_alignedDequeue_bits_data_T_844[6], _alignedDequeue_bits_data_T_778[6]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_14 = {_alignedDequeue_bits_data_T_976[6], _alignedDequeue_bits_data_T_910[6]};
  wire [3:0]    alignedDequeue_bits_data_hi_14 = {alignedDequeue_bits_data_hi_hi_14, alignedDequeue_bits_data_hi_lo_14};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_15 = {_alignedDequeue_bits_data_T_580[7], _alignedDequeue_bits_data_T_514[7]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_15 = {_alignedDequeue_bits_data_T_712[7], _alignedDequeue_bits_data_T_646[7]};
  wire [3:0]    alignedDequeue_bits_data_lo_15 = {alignedDequeue_bits_data_lo_hi_15, alignedDequeue_bits_data_lo_lo_15};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_15 = {_alignedDequeue_bits_data_T_844[7], _alignedDequeue_bits_data_T_778[7]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_15 = {_alignedDequeue_bits_data_T_976[7], _alignedDequeue_bits_data_T_910[7]};
  wire [3:0]    alignedDequeue_bits_data_hi_15 = {alignedDequeue_bits_data_hi_hi_15, alignedDequeue_bits_data_hi_lo_15};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_16 = {_alignedDequeue_bits_data_T_580[8], _alignedDequeue_bits_data_T_514[8]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_16 = {_alignedDequeue_bits_data_T_712[8], _alignedDequeue_bits_data_T_646[8]};
  wire [3:0]    alignedDequeue_bits_data_lo_16 = {alignedDequeue_bits_data_lo_hi_16, alignedDequeue_bits_data_lo_lo_16};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_16 = {_alignedDequeue_bits_data_T_844[8], _alignedDequeue_bits_data_T_778[8]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_16 = {_alignedDequeue_bits_data_T_976[8], _alignedDequeue_bits_data_T_910[8]};
  wire [3:0]    alignedDequeue_bits_data_hi_16 = {alignedDequeue_bits_data_hi_hi_16, alignedDequeue_bits_data_hi_lo_16};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_17 = {_alignedDequeue_bits_data_T_580[9], _alignedDequeue_bits_data_T_514[9]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_17 = {_alignedDequeue_bits_data_T_712[9], _alignedDequeue_bits_data_T_646[9]};
  wire [3:0]    alignedDequeue_bits_data_lo_17 = {alignedDequeue_bits_data_lo_hi_17, alignedDequeue_bits_data_lo_lo_17};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_17 = {_alignedDequeue_bits_data_T_844[9], _alignedDequeue_bits_data_T_778[9]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_17 = {_alignedDequeue_bits_data_T_976[9], _alignedDequeue_bits_data_T_910[9]};
  wire [3:0]    alignedDequeue_bits_data_hi_17 = {alignedDequeue_bits_data_hi_hi_17, alignedDequeue_bits_data_hi_lo_17};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_18 = {_alignedDequeue_bits_data_T_580[10], _alignedDequeue_bits_data_T_514[10]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_18 = {_alignedDequeue_bits_data_T_712[10], _alignedDequeue_bits_data_T_646[10]};
  wire [3:0]    alignedDequeue_bits_data_lo_18 = {alignedDequeue_bits_data_lo_hi_18, alignedDequeue_bits_data_lo_lo_18};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_18 = {_alignedDequeue_bits_data_T_844[10], _alignedDequeue_bits_data_T_778[10]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_18 = {_alignedDequeue_bits_data_T_976[10], _alignedDequeue_bits_data_T_910[10]};
  wire [3:0]    alignedDequeue_bits_data_hi_18 = {alignedDequeue_bits_data_hi_hi_18, alignedDequeue_bits_data_hi_lo_18};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_19 = {_alignedDequeue_bits_data_T_580[11], _alignedDequeue_bits_data_T_514[11]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_19 = {_alignedDequeue_bits_data_T_712[11], _alignedDequeue_bits_data_T_646[11]};
  wire [3:0]    alignedDequeue_bits_data_lo_19 = {alignedDequeue_bits_data_lo_hi_19, alignedDequeue_bits_data_lo_lo_19};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_19 = {_alignedDequeue_bits_data_T_844[11], _alignedDequeue_bits_data_T_778[11]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_19 = {_alignedDequeue_bits_data_T_976[11], _alignedDequeue_bits_data_T_910[11]};
  wire [3:0]    alignedDequeue_bits_data_hi_19 = {alignedDequeue_bits_data_hi_hi_19, alignedDequeue_bits_data_hi_lo_19};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_20 = {_alignedDequeue_bits_data_T_580[12], _alignedDequeue_bits_data_T_514[12]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_20 = {_alignedDequeue_bits_data_T_712[12], _alignedDequeue_bits_data_T_646[12]};
  wire [3:0]    alignedDequeue_bits_data_lo_20 = {alignedDequeue_bits_data_lo_hi_20, alignedDequeue_bits_data_lo_lo_20};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_20 = {_alignedDequeue_bits_data_T_844[12], _alignedDequeue_bits_data_T_778[12]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_20 = {_alignedDequeue_bits_data_T_976[12], _alignedDequeue_bits_data_T_910[12]};
  wire [3:0]    alignedDequeue_bits_data_hi_20 = {alignedDequeue_bits_data_hi_hi_20, alignedDequeue_bits_data_hi_lo_20};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_21 = {_alignedDequeue_bits_data_T_580[13], _alignedDequeue_bits_data_T_514[13]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_21 = {_alignedDequeue_bits_data_T_712[13], _alignedDequeue_bits_data_T_646[13]};
  wire [3:0]    alignedDequeue_bits_data_lo_21 = {alignedDequeue_bits_data_lo_hi_21, alignedDequeue_bits_data_lo_lo_21};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_21 = {_alignedDequeue_bits_data_T_844[13], _alignedDequeue_bits_data_T_778[13]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_21 = {_alignedDequeue_bits_data_T_976[13], _alignedDequeue_bits_data_T_910[13]};
  wire [3:0]    alignedDequeue_bits_data_hi_21 = {alignedDequeue_bits_data_hi_hi_21, alignedDequeue_bits_data_hi_lo_21};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_22 = {_alignedDequeue_bits_data_T_580[14], _alignedDequeue_bits_data_T_514[14]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_22 = {_alignedDequeue_bits_data_T_712[14], _alignedDequeue_bits_data_T_646[14]};
  wire [3:0]    alignedDequeue_bits_data_lo_22 = {alignedDequeue_bits_data_lo_hi_22, alignedDequeue_bits_data_lo_lo_22};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_22 = {_alignedDequeue_bits_data_T_844[14], _alignedDequeue_bits_data_T_778[14]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_22 = {_alignedDequeue_bits_data_T_976[14], _alignedDequeue_bits_data_T_910[14]};
  wire [3:0]    alignedDequeue_bits_data_hi_22 = {alignedDequeue_bits_data_hi_hi_22, alignedDequeue_bits_data_hi_lo_22};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_23 = {_alignedDequeue_bits_data_T_580[15], _alignedDequeue_bits_data_T_514[15]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_23 = {_alignedDequeue_bits_data_T_712[15], _alignedDequeue_bits_data_T_646[15]};
  wire [3:0]    alignedDequeue_bits_data_lo_23 = {alignedDequeue_bits_data_lo_hi_23, alignedDequeue_bits_data_lo_lo_23};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_23 = {_alignedDequeue_bits_data_T_844[15], _alignedDequeue_bits_data_T_778[15]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_23 = {_alignedDequeue_bits_data_T_976[15], _alignedDequeue_bits_data_T_910[15]};
  wire [3:0]    alignedDequeue_bits_data_hi_23 = {alignedDequeue_bits_data_hi_hi_23, alignedDequeue_bits_data_hi_lo_23};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_24 = {_alignedDequeue_bits_data_T_580[16], _alignedDequeue_bits_data_T_514[16]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_24 = {_alignedDequeue_bits_data_T_712[16], _alignedDequeue_bits_data_T_646[16]};
  wire [3:0]    alignedDequeue_bits_data_lo_24 = {alignedDequeue_bits_data_lo_hi_24, alignedDequeue_bits_data_lo_lo_24};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_24 = {_alignedDequeue_bits_data_T_844[16], _alignedDequeue_bits_data_T_778[16]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_24 = {_alignedDequeue_bits_data_T_976[16], _alignedDequeue_bits_data_T_910[16]};
  wire [3:0]    alignedDequeue_bits_data_hi_24 = {alignedDequeue_bits_data_hi_hi_24, alignedDequeue_bits_data_hi_lo_24};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_25 = {_alignedDequeue_bits_data_T_580[17], _alignedDequeue_bits_data_T_514[17]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_25 = {_alignedDequeue_bits_data_T_712[17], _alignedDequeue_bits_data_T_646[17]};
  wire [3:0]    alignedDequeue_bits_data_lo_25 = {alignedDequeue_bits_data_lo_hi_25, alignedDequeue_bits_data_lo_lo_25};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_25 = {_alignedDequeue_bits_data_T_844[17], _alignedDequeue_bits_data_T_778[17]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_25 = {_alignedDequeue_bits_data_T_976[17], _alignedDequeue_bits_data_T_910[17]};
  wire [3:0]    alignedDequeue_bits_data_hi_25 = {alignedDequeue_bits_data_hi_hi_25, alignedDequeue_bits_data_hi_lo_25};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_26 = {_alignedDequeue_bits_data_T_580[18], _alignedDequeue_bits_data_T_514[18]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_26 = {_alignedDequeue_bits_data_T_712[18], _alignedDequeue_bits_data_T_646[18]};
  wire [3:0]    alignedDequeue_bits_data_lo_26 = {alignedDequeue_bits_data_lo_hi_26, alignedDequeue_bits_data_lo_lo_26};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_26 = {_alignedDequeue_bits_data_T_844[18], _alignedDequeue_bits_data_T_778[18]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_26 = {_alignedDequeue_bits_data_T_976[18], _alignedDequeue_bits_data_T_910[18]};
  wire [3:0]    alignedDequeue_bits_data_hi_26 = {alignedDequeue_bits_data_hi_hi_26, alignedDequeue_bits_data_hi_lo_26};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_27 = {_alignedDequeue_bits_data_T_580[19], _alignedDequeue_bits_data_T_514[19]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_27 = {_alignedDequeue_bits_data_T_712[19], _alignedDequeue_bits_data_T_646[19]};
  wire [3:0]    alignedDequeue_bits_data_lo_27 = {alignedDequeue_bits_data_lo_hi_27, alignedDequeue_bits_data_lo_lo_27};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_27 = {_alignedDequeue_bits_data_T_844[19], _alignedDequeue_bits_data_T_778[19]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_27 = {_alignedDequeue_bits_data_T_976[19], _alignedDequeue_bits_data_T_910[19]};
  wire [3:0]    alignedDequeue_bits_data_hi_27 = {alignedDequeue_bits_data_hi_hi_27, alignedDequeue_bits_data_hi_lo_27};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_28 = {_alignedDequeue_bits_data_T_580[20], _alignedDequeue_bits_data_T_514[20]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_28 = {_alignedDequeue_bits_data_T_712[20], _alignedDequeue_bits_data_T_646[20]};
  wire [3:0]    alignedDequeue_bits_data_lo_28 = {alignedDequeue_bits_data_lo_hi_28, alignedDequeue_bits_data_lo_lo_28};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_28 = {_alignedDequeue_bits_data_T_844[20], _alignedDequeue_bits_data_T_778[20]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_28 = {_alignedDequeue_bits_data_T_976[20], _alignedDequeue_bits_data_T_910[20]};
  wire [3:0]    alignedDequeue_bits_data_hi_28 = {alignedDequeue_bits_data_hi_hi_28, alignedDequeue_bits_data_hi_lo_28};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_29 = {_alignedDequeue_bits_data_T_580[21], _alignedDequeue_bits_data_T_514[21]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_29 = {_alignedDequeue_bits_data_T_712[21], _alignedDequeue_bits_data_T_646[21]};
  wire [3:0]    alignedDequeue_bits_data_lo_29 = {alignedDequeue_bits_data_lo_hi_29, alignedDequeue_bits_data_lo_lo_29};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_29 = {_alignedDequeue_bits_data_T_844[21], _alignedDequeue_bits_data_T_778[21]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_29 = {_alignedDequeue_bits_data_T_976[21], _alignedDequeue_bits_data_T_910[21]};
  wire [3:0]    alignedDequeue_bits_data_hi_29 = {alignedDequeue_bits_data_hi_hi_29, alignedDequeue_bits_data_hi_lo_29};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_30 = {_alignedDequeue_bits_data_T_580[22], _alignedDequeue_bits_data_T_514[22]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_30 = {_alignedDequeue_bits_data_T_712[22], _alignedDequeue_bits_data_T_646[22]};
  wire [3:0]    alignedDequeue_bits_data_lo_30 = {alignedDequeue_bits_data_lo_hi_30, alignedDequeue_bits_data_lo_lo_30};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_30 = {_alignedDequeue_bits_data_T_844[22], _alignedDequeue_bits_data_T_778[22]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_30 = {_alignedDequeue_bits_data_T_976[22], _alignedDequeue_bits_data_T_910[22]};
  wire [3:0]    alignedDequeue_bits_data_hi_30 = {alignedDequeue_bits_data_hi_hi_30, alignedDequeue_bits_data_hi_lo_30};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_31 = {_alignedDequeue_bits_data_T_580[23], _alignedDequeue_bits_data_T_514[23]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_31 = {_alignedDequeue_bits_data_T_712[23], _alignedDequeue_bits_data_T_646[23]};
  wire [3:0]    alignedDequeue_bits_data_lo_31 = {alignedDequeue_bits_data_lo_hi_31, alignedDequeue_bits_data_lo_lo_31};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_31 = {_alignedDequeue_bits_data_T_844[23], _alignedDequeue_bits_data_T_778[23]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_31 = {_alignedDequeue_bits_data_T_976[23], _alignedDequeue_bits_data_T_910[23]};
  wire [3:0]    alignedDequeue_bits_data_hi_31 = {alignedDequeue_bits_data_hi_hi_31, alignedDequeue_bits_data_hi_lo_31};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_32 = {_alignedDequeue_bits_data_T_580[24], _alignedDequeue_bits_data_T_514[24]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_32 = {_alignedDequeue_bits_data_T_712[24], _alignedDequeue_bits_data_T_646[24]};
  wire [3:0]    alignedDequeue_bits_data_lo_32 = {alignedDequeue_bits_data_lo_hi_32, alignedDequeue_bits_data_lo_lo_32};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_32 = {_alignedDequeue_bits_data_T_844[24], _alignedDequeue_bits_data_T_778[24]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_32 = {_alignedDequeue_bits_data_T_976[24], _alignedDequeue_bits_data_T_910[24]};
  wire [3:0]    alignedDequeue_bits_data_hi_32 = {alignedDequeue_bits_data_hi_hi_32, alignedDequeue_bits_data_hi_lo_32};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_33 = {_alignedDequeue_bits_data_T_580[25], _alignedDequeue_bits_data_T_514[25]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_33 = {_alignedDequeue_bits_data_T_712[25], _alignedDequeue_bits_data_T_646[25]};
  wire [3:0]    alignedDequeue_bits_data_lo_33 = {alignedDequeue_bits_data_lo_hi_33, alignedDequeue_bits_data_lo_lo_33};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_33 = {_alignedDequeue_bits_data_T_844[25], _alignedDequeue_bits_data_T_778[25]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_33 = {_alignedDequeue_bits_data_T_976[25], _alignedDequeue_bits_data_T_910[25]};
  wire [3:0]    alignedDequeue_bits_data_hi_33 = {alignedDequeue_bits_data_hi_hi_33, alignedDequeue_bits_data_hi_lo_33};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_34 = {_alignedDequeue_bits_data_T_580[26], _alignedDequeue_bits_data_T_514[26]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_34 = {_alignedDequeue_bits_data_T_712[26], _alignedDequeue_bits_data_T_646[26]};
  wire [3:0]    alignedDequeue_bits_data_lo_34 = {alignedDequeue_bits_data_lo_hi_34, alignedDequeue_bits_data_lo_lo_34};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_34 = {_alignedDequeue_bits_data_T_844[26], _alignedDequeue_bits_data_T_778[26]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_34 = {_alignedDequeue_bits_data_T_976[26], _alignedDequeue_bits_data_T_910[26]};
  wire [3:0]    alignedDequeue_bits_data_hi_34 = {alignedDequeue_bits_data_hi_hi_34, alignedDequeue_bits_data_hi_lo_34};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_35 = {_alignedDequeue_bits_data_T_580[27], _alignedDequeue_bits_data_T_514[27]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_35 = {_alignedDequeue_bits_data_T_712[27], _alignedDequeue_bits_data_T_646[27]};
  wire [3:0]    alignedDequeue_bits_data_lo_35 = {alignedDequeue_bits_data_lo_hi_35, alignedDequeue_bits_data_lo_lo_35};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_35 = {_alignedDequeue_bits_data_T_844[27], _alignedDequeue_bits_data_T_778[27]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_35 = {_alignedDequeue_bits_data_T_976[27], _alignedDequeue_bits_data_T_910[27]};
  wire [3:0]    alignedDequeue_bits_data_hi_35 = {alignedDequeue_bits_data_hi_hi_35, alignedDequeue_bits_data_hi_lo_35};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_36 = {_alignedDequeue_bits_data_T_580[28], _alignedDequeue_bits_data_T_514[28]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_36 = {_alignedDequeue_bits_data_T_712[28], _alignedDequeue_bits_data_T_646[28]};
  wire [3:0]    alignedDequeue_bits_data_lo_36 = {alignedDequeue_bits_data_lo_hi_36, alignedDequeue_bits_data_lo_lo_36};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_36 = {_alignedDequeue_bits_data_T_844[28], _alignedDequeue_bits_data_T_778[28]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_36 = {_alignedDequeue_bits_data_T_976[28], _alignedDequeue_bits_data_T_910[28]};
  wire [3:0]    alignedDequeue_bits_data_hi_36 = {alignedDequeue_bits_data_hi_hi_36, alignedDequeue_bits_data_hi_lo_36};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_37 = {_alignedDequeue_bits_data_T_580[29], _alignedDequeue_bits_data_T_514[29]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_37 = {_alignedDequeue_bits_data_T_712[29], _alignedDequeue_bits_data_T_646[29]};
  wire [3:0]    alignedDequeue_bits_data_lo_37 = {alignedDequeue_bits_data_lo_hi_37, alignedDequeue_bits_data_lo_lo_37};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_37 = {_alignedDequeue_bits_data_T_844[29], _alignedDequeue_bits_data_T_778[29]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_37 = {_alignedDequeue_bits_data_T_976[29], _alignedDequeue_bits_data_T_910[29]};
  wire [3:0]    alignedDequeue_bits_data_hi_37 = {alignedDequeue_bits_data_hi_hi_37, alignedDequeue_bits_data_hi_lo_37};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_38 = {_alignedDequeue_bits_data_T_580[30], _alignedDequeue_bits_data_T_514[30]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_38 = {_alignedDequeue_bits_data_T_712[30], _alignedDequeue_bits_data_T_646[30]};
  wire [3:0]    alignedDequeue_bits_data_lo_38 = {alignedDequeue_bits_data_lo_hi_38, alignedDequeue_bits_data_lo_lo_38};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_38 = {_alignedDequeue_bits_data_T_844[30], _alignedDequeue_bits_data_T_778[30]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_38 = {_alignedDequeue_bits_data_T_976[30], _alignedDequeue_bits_data_T_910[30]};
  wire [3:0]    alignedDequeue_bits_data_hi_38 = {alignedDequeue_bits_data_hi_hi_38, alignedDequeue_bits_data_hi_lo_38};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_39 = {_alignedDequeue_bits_data_T_580[31], _alignedDequeue_bits_data_T_514[31]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_39 = {_alignedDequeue_bits_data_T_712[31], _alignedDequeue_bits_data_T_646[31]};
  wire [3:0]    alignedDequeue_bits_data_lo_39 = {alignedDequeue_bits_data_lo_hi_39, alignedDequeue_bits_data_lo_lo_39};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_39 = {_alignedDequeue_bits_data_T_844[31], _alignedDequeue_bits_data_T_778[31]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_39 = {_alignedDequeue_bits_data_T_976[31], _alignedDequeue_bits_data_T_910[31]};
  wire [3:0]    alignedDequeue_bits_data_hi_39 = {alignedDequeue_bits_data_hi_hi_39, alignedDequeue_bits_data_hi_lo_39};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_40 = {_alignedDequeue_bits_data_T_580[32], _alignedDequeue_bits_data_T_514[32]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_40 = {_alignedDequeue_bits_data_T_712[32], _alignedDequeue_bits_data_T_646[32]};
  wire [3:0]    alignedDequeue_bits_data_lo_40 = {alignedDequeue_bits_data_lo_hi_40, alignedDequeue_bits_data_lo_lo_40};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_40 = {_alignedDequeue_bits_data_T_844[32], _alignedDequeue_bits_data_T_778[32]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_40 = {_alignedDequeue_bits_data_T_976[32], _alignedDequeue_bits_data_T_910[32]};
  wire [3:0]    alignedDequeue_bits_data_hi_40 = {alignedDequeue_bits_data_hi_hi_40, alignedDequeue_bits_data_hi_lo_40};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_41 = {_alignedDequeue_bits_data_T_580[33], _alignedDequeue_bits_data_T_514[33]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_41 = {_alignedDequeue_bits_data_T_712[33], _alignedDequeue_bits_data_T_646[33]};
  wire [3:0]    alignedDequeue_bits_data_lo_41 = {alignedDequeue_bits_data_lo_hi_41, alignedDequeue_bits_data_lo_lo_41};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_41 = {_alignedDequeue_bits_data_T_844[33], _alignedDequeue_bits_data_T_778[33]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_41 = {_alignedDequeue_bits_data_T_976[33], _alignedDequeue_bits_data_T_910[33]};
  wire [3:0]    alignedDequeue_bits_data_hi_41 = {alignedDequeue_bits_data_hi_hi_41, alignedDequeue_bits_data_hi_lo_41};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_42 = {_alignedDequeue_bits_data_T_580[34], _alignedDequeue_bits_data_T_514[34]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_42 = {_alignedDequeue_bits_data_T_712[34], _alignedDequeue_bits_data_T_646[34]};
  wire [3:0]    alignedDequeue_bits_data_lo_42 = {alignedDequeue_bits_data_lo_hi_42, alignedDequeue_bits_data_lo_lo_42};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_42 = {_alignedDequeue_bits_data_T_844[34], _alignedDequeue_bits_data_T_778[34]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_42 = {_alignedDequeue_bits_data_T_976[34], _alignedDequeue_bits_data_T_910[34]};
  wire [3:0]    alignedDequeue_bits_data_hi_42 = {alignedDequeue_bits_data_hi_hi_42, alignedDequeue_bits_data_hi_lo_42};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_43 = {_alignedDequeue_bits_data_T_580[35], _alignedDequeue_bits_data_T_514[35]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_43 = {_alignedDequeue_bits_data_T_712[35], _alignedDequeue_bits_data_T_646[35]};
  wire [3:0]    alignedDequeue_bits_data_lo_43 = {alignedDequeue_bits_data_lo_hi_43, alignedDequeue_bits_data_lo_lo_43};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_43 = {_alignedDequeue_bits_data_T_844[35], _alignedDequeue_bits_data_T_778[35]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_43 = {_alignedDequeue_bits_data_T_976[35], _alignedDequeue_bits_data_T_910[35]};
  wire [3:0]    alignedDequeue_bits_data_hi_43 = {alignedDequeue_bits_data_hi_hi_43, alignedDequeue_bits_data_hi_lo_43};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_44 = {_alignedDequeue_bits_data_T_580[36], _alignedDequeue_bits_data_T_514[36]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_44 = {_alignedDequeue_bits_data_T_712[36], _alignedDequeue_bits_data_T_646[36]};
  wire [3:0]    alignedDequeue_bits_data_lo_44 = {alignedDequeue_bits_data_lo_hi_44, alignedDequeue_bits_data_lo_lo_44};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_44 = {_alignedDequeue_bits_data_T_844[36], _alignedDequeue_bits_data_T_778[36]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_44 = {_alignedDequeue_bits_data_T_976[36], _alignedDequeue_bits_data_T_910[36]};
  wire [3:0]    alignedDequeue_bits_data_hi_44 = {alignedDequeue_bits_data_hi_hi_44, alignedDequeue_bits_data_hi_lo_44};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_45 = {_alignedDequeue_bits_data_T_580[37], _alignedDequeue_bits_data_T_514[37]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_45 = {_alignedDequeue_bits_data_T_712[37], _alignedDequeue_bits_data_T_646[37]};
  wire [3:0]    alignedDequeue_bits_data_lo_45 = {alignedDequeue_bits_data_lo_hi_45, alignedDequeue_bits_data_lo_lo_45};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_45 = {_alignedDequeue_bits_data_T_844[37], _alignedDequeue_bits_data_T_778[37]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_45 = {_alignedDequeue_bits_data_T_976[37], _alignedDequeue_bits_data_T_910[37]};
  wire [3:0]    alignedDequeue_bits_data_hi_45 = {alignedDequeue_bits_data_hi_hi_45, alignedDequeue_bits_data_hi_lo_45};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_46 = {_alignedDequeue_bits_data_T_580[38], _alignedDequeue_bits_data_T_514[38]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_46 = {_alignedDequeue_bits_data_T_712[38], _alignedDequeue_bits_data_T_646[38]};
  wire [3:0]    alignedDequeue_bits_data_lo_46 = {alignedDequeue_bits_data_lo_hi_46, alignedDequeue_bits_data_lo_lo_46};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_46 = {_alignedDequeue_bits_data_T_844[38], _alignedDequeue_bits_data_T_778[38]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_46 = {_alignedDequeue_bits_data_T_976[38], _alignedDequeue_bits_data_T_910[38]};
  wire [3:0]    alignedDequeue_bits_data_hi_46 = {alignedDequeue_bits_data_hi_hi_46, alignedDequeue_bits_data_hi_lo_46};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_47 = {_alignedDequeue_bits_data_T_580[39], _alignedDequeue_bits_data_T_514[39]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_47 = {_alignedDequeue_bits_data_T_712[39], _alignedDequeue_bits_data_T_646[39]};
  wire [3:0]    alignedDequeue_bits_data_lo_47 = {alignedDequeue_bits_data_lo_hi_47, alignedDequeue_bits_data_lo_lo_47};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_47 = {_alignedDequeue_bits_data_T_844[39], _alignedDequeue_bits_data_T_778[39]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_47 = {_alignedDequeue_bits_data_T_976[39], _alignedDequeue_bits_data_T_910[39]};
  wire [3:0]    alignedDequeue_bits_data_hi_47 = {alignedDequeue_bits_data_hi_hi_47, alignedDequeue_bits_data_hi_lo_47};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_48 = {_alignedDequeue_bits_data_T_580[40], _alignedDequeue_bits_data_T_514[40]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_48 = {_alignedDequeue_bits_data_T_712[40], _alignedDequeue_bits_data_T_646[40]};
  wire [3:0]    alignedDequeue_bits_data_lo_48 = {alignedDequeue_bits_data_lo_hi_48, alignedDequeue_bits_data_lo_lo_48};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_48 = {_alignedDequeue_bits_data_T_844[40], _alignedDequeue_bits_data_T_778[40]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_48 = {_alignedDequeue_bits_data_T_976[40], _alignedDequeue_bits_data_T_910[40]};
  wire [3:0]    alignedDequeue_bits_data_hi_48 = {alignedDequeue_bits_data_hi_hi_48, alignedDequeue_bits_data_hi_lo_48};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_49 = {_alignedDequeue_bits_data_T_580[41], _alignedDequeue_bits_data_T_514[41]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_49 = {_alignedDequeue_bits_data_T_712[41], _alignedDequeue_bits_data_T_646[41]};
  wire [3:0]    alignedDequeue_bits_data_lo_49 = {alignedDequeue_bits_data_lo_hi_49, alignedDequeue_bits_data_lo_lo_49};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_49 = {_alignedDequeue_bits_data_T_844[41], _alignedDequeue_bits_data_T_778[41]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_49 = {_alignedDequeue_bits_data_T_976[41], _alignedDequeue_bits_data_T_910[41]};
  wire [3:0]    alignedDequeue_bits_data_hi_49 = {alignedDequeue_bits_data_hi_hi_49, alignedDequeue_bits_data_hi_lo_49};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_50 = {_alignedDequeue_bits_data_T_580[42], _alignedDequeue_bits_data_T_514[42]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_50 = {_alignedDequeue_bits_data_T_712[42], _alignedDequeue_bits_data_T_646[42]};
  wire [3:0]    alignedDequeue_bits_data_lo_50 = {alignedDequeue_bits_data_lo_hi_50, alignedDequeue_bits_data_lo_lo_50};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_50 = {_alignedDequeue_bits_data_T_844[42], _alignedDequeue_bits_data_T_778[42]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_50 = {_alignedDequeue_bits_data_T_976[42], _alignedDequeue_bits_data_T_910[42]};
  wire [3:0]    alignedDequeue_bits_data_hi_50 = {alignedDequeue_bits_data_hi_hi_50, alignedDequeue_bits_data_hi_lo_50};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_51 = {_alignedDequeue_bits_data_T_580[43], _alignedDequeue_bits_data_T_514[43]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_51 = {_alignedDequeue_bits_data_T_712[43], _alignedDequeue_bits_data_T_646[43]};
  wire [3:0]    alignedDequeue_bits_data_lo_51 = {alignedDequeue_bits_data_lo_hi_51, alignedDequeue_bits_data_lo_lo_51};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_51 = {_alignedDequeue_bits_data_T_844[43], _alignedDequeue_bits_data_T_778[43]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_51 = {_alignedDequeue_bits_data_T_976[43], _alignedDequeue_bits_data_T_910[43]};
  wire [3:0]    alignedDequeue_bits_data_hi_51 = {alignedDequeue_bits_data_hi_hi_51, alignedDequeue_bits_data_hi_lo_51};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_52 = {_alignedDequeue_bits_data_T_580[44], _alignedDequeue_bits_data_T_514[44]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_52 = {_alignedDequeue_bits_data_T_712[44], _alignedDequeue_bits_data_T_646[44]};
  wire [3:0]    alignedDequeue_bits_data_lo_52 = {alignedDequeue_bits_data_lo_hi_52, alignedDequeue_bits_data_lo_lo_52};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_52 = {_alignedDequeue_bits_data_T_844[44], _alignedDequeue_bits_data_T_778[44]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_52 = {_alignedDequeue_bits_data_T_976[44], _alignedDequeue_bits_data_T_910[44]};
  wire [3:0]    alignedDequeue_bits_data_hi_52 = {alignedDequeue_bits_data_hi_hi_52, alignedDequeue_bits_data_hi_lo_52};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_53 = {_alignedDequeue_bits_data_T_580[45], _alignedDequeue_bits_data_T_514[45]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_53 = {_alignedDequeue_bits_data_T_712[45], _alignedDequeue_bits_data_T_646[45]};
  wire [3:0]    alignedDequeue_bits_data_lo_53 = {alignedDequeue_bits_data_lo_hi_53, alignedDequeue_bits_data_lo_lo_53};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_53 = {_alignedDequeue_bits_data_T_844[45], _alignedDequeue_bits_data_T_778[45]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_53 = {_alignedDequeue_bits_data_T_976[45], _alignedDequeue_bits_data_T_910[45]};
  wire [3:0]    alignedDequeue_bits_data_hi_53 = {alignedDequeue_bits_data_hi_hi_53, alignedDequeue_bits_data_hi_lo_53};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_54 = {_alignedDequeue_bits_data_T_580[46], _alignedDequeue_bits_data_T_514[46]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_54 = {_alignedDequeue_bits_data_T_712[46], _alignedDequeue_bits_data_T_646[46]};
  wire [3:0]    alignedDequeue_bits_data_lo_54 = {alignedDequeue_bits_data_lo_hi_54, alignedDequeue_bits_data_lo_lo_54};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_54 = {_alignedDequeue_bits_data_T_844[46], _alignedDequeue_bits_data_T_778[46]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_54 = {_alignedDequeue_bits_data_T_976[46], _alignedDequeue_bits_data_T_910[46]};
  wire [3:0]    alignedDequeue_bits_data_hi_54 = {alignedDequeue_bits_data_hi_hi_54, alignedDequeue_bits_data_hi_lo_54};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_55 = {_alignedDequeue_bits_data_T_580[47], _alignedDequeue_bits_data_T_514[47]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_55 = {_alignedDequeue_bits_data_T_712[47], _alignedDequeue_bits_data_T_646[47]};
  wire [3:0]    alignedDequeue_bits_data_lo_55 = {alignedDequeue_bits_data_lo_hi_55, alignedDequeue_bits_data_lo_lo_55};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_55 = {_alignedDequeue_bits_data_T_844[47], _alignedDequeue_bits_data_T_778[47]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_55 = {_alignedDequeue_bits_data_T_976[47], _alignedDequeue_bits_data_T_910[47]};
  wire [3:0]    alignedDequeue_bits_data_hi_55 = {alignedDequeue_bits_data_hi_hi_55, alignedDequeue_bits_data_hi_lo_55};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_56 = {_alignedDequeue_bits_data_T_580[48], _alignedDequeue_bits_data_T_514[48]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_56 = {_alignedDequeue_bits_data_T_712[48], _alignedDequeue_bits_data_T_646[48]};
  wire [3:0]    alignedDequeue_bits_data_lo_56 = {alignedDequeue_bits_data_lo_hi_56, alignedDequeue_bits_data_lo_lo_56};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_56 = {_alignedDequeue_bits_data_T_844[48], _alignedDequeue_bits_data_T_778[48]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_56 = {_alignedDequeue_bits_data_T_976[48], _alignedDequeue_bits_data_T_910[48]};
  wire [3:0]    alignedDequeue_bits_data_hi_56 = {alignedDequeue_bits_data_hi_hi_56, alignedDequeue_bits_data_hi_lo_56};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_57 = {_alignedDequeue_bits_data_T_580[49], _alignedDequeue_bits_data_T_514[49]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_57 = {_alignedDequeue_bits_data_T_712[49], _alignedDequeue_bits_data_T_646[49]};
  wire [3:0]    alignedDequeue_bits_data_lo_57 = {alignedDequeue_bits_data_lo_hi_57, alignedDequeue_bits_data_lo_lo_57};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_57 = {_alignedDequeue_bits_data_T_844[49], _alignedDequeue_bits_data_T_778[49]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_57 = {_alignedDequeue_bits_data_T_976[49], _alignedDequeue_bits_data_T_910[49]};
  wire [3:0]    alignedDequeue_bits_data_hi_57 = {alignedDequeue_bits_data_hi_hi_57, alignedDequeue_bits_data_hi_lo_57};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_58 = {_alignedDequeue_bits_data_T_580[50], _alignedDequeue_bits_data_T_514[50]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_58 = {_alignedDequeue_bits_data_T_712[50], _alignedDequeue_bits_data_T_646[50]};
  wire [3:0]    alignedDequeue_bits_data_lo_58 = {alignedDequeue_bits_data_lo_hi_58, alignedDequeue_bits_data_lo_lo_58};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_58 = {_alignedDequeue_bits_data_T_844[50], _alignedDequeue_bits_data_T_778[50]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_58 = {_alignedDequeue_bits_data_T_976[50], _alignedDequeue_bits_data_T_910[50]};
  wire [3:0]    alignedDequeue_bits_data_hi_58 = {alignedDequeue_bits_data_hi_hi_58, alignedDequeue_bits_data_hi_lo_58};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_59 = {_alignedDequeue_bits_data_T_580[51], _alignedDequeue_bits_data_T_514[51]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_59 = {_alignedDequeue_bits_data_T_712[51], _alignedDequeue_bits_data_T_646[51]};
  wire [3:0]    alignedDequeue_bits_data_lo_59 = {alignedDequeue_bits_data_lo_hi_59, alignedDequeue_bits_data_lo_lo_59};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_59 = {_alignedDequeue_bits_data_T_844[51], _alignedDequeue_bits_data_T_778[51]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_59 = {_alignedDequeue_bits_data_T_976[51], _alignedDequeue_bits_data_T_910[51]};
  wire [3:0]    alignedDequeue_bits_data_hi_59 = {alignedDequeue_bits_data_hi_hi_59, alignedDequeue_bits_data_hi_lo_59};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_60 = {_alignedDequeue_bits_data_T_580[52], _alignedDequeue_bits_data_T_514[52]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_60 = {_alignedDequeue_bits_data_T_712[52], _alignedDequeue_bits_data_T_646[52]};
  wire [3:0]    alignedDequeue_bits_data_lo_60 = {alignedDequeue_bits_data_lo_hi_60, alignedDequeue_bits_data_lo_lo_60};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_60 = {_alignedDequeue_bits_data_T_844[52], _alignedDequeue_bits_data_T_778[52]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_60 = {_alignedDequeue_bits_data_T_976[52], _alignedDequeue_bits_data_T_910[52]};
  wire [3:0]    alignedDequeue_bits_data_hi_60 = {alignedDequeue_bits_data_hi_hi_60, alignedDequeue_bits_data_hi_lo_60};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_61 = {_alignedDequeue_bits_data_T_580[53], _alignedDequeue_bits_data_T_514[53]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_61 = {_alignedDequeue_bits_data_T_712[53], _alignedDequeue_bits_data_T_646[53]};
  wire [3:0]    alignedDequeue_bits_data_lo_61 = {alignedDequeue_bits_data_lo_hi_61, alignedDequeue_bits_data_lo_lo_61};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_61 = {_alignedDequeue_bits_data_T_844[53], _alignedDequeue_bits_data_T_778[53]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_61 = {_alignedDequeue_bits_data_T_976[53], _alignedDequeue_bits_data_T_910[53]};
  wire [3:0]    alignedDequeue_bits_data_hi_61 = {alignedDequeue_bits_data_hi_hi_61, alignedDequeue_bits_data_hi_lo_61};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_62 = {_alignedDequeue_bits_data_T_580[54], _alignedDequeue_bits_data_T_514[54]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_62 = {_alignedDequeue_bits_data_T_712[54], _alignedDequeue_bits_data_T_646[54]};
  wire [3:0]    alignedDequeue_bits_data_lo_62 = {alignedDequeue_bits_data_lo_hi_62, alignedDequeue_bits_data_lo_lo_62};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_62 = {_alignedDequeue_bits_data_T_844[54], _alignedDequeue_bits_data_T_778[54]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_62 = {_alignedDequeue_bits_data_T_976[54], _alignedDequeue_bits_data_T_910[54]};
  wire [3:0]    alignedDequeue_bits_data_hi_62 = {alignedDequeue_bits_data_hi_hi_62, alignedDequeue_bits_data_hi_lo_62};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_63 = {_alignedDequeue_bits_data_T_580[55], _alignedDequeue_bits_data_T_514[55]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_63 = {_alignedDequeue_bits_data_T_712[55], _alignedDequeue_bits_data_T_646[55]};
  wire [3:0]    alignedDequeue_bits_data_lo_63 = {alignedDequeue_bits_data_lo_hi_63, alignedDequeue_bits_data_lo_lo_63};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_63 = {_alignedDequeue_bits_data_T_844[55], _alignedDequeue_bits_data_T_778[55]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_63 = {_alignedDequeue_bits_data_T_976[55], _alignedDequeue_bits_data_T_910[55]};
  wire [3:0]    alignedDequeue_bits_data_hi_63 = {alignedDequeue_bits_data_hi_hi_63, alignedDequeue_bits_data_hi_lo_63};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_64 = {_alignedDequeue_bits_data_T_580[56], _alignedDequeue_bits_data_T_514[56]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_64 = {_alignedDequeue_bits_data_T_712[56], _alignedDequeue_bits_data_T_646[56]};
  wire [3:0]    alignedDequeue_bits_data_lo_64 = {alignedDequeue_bits_data_lo_hi_64, alignedDequeue_bits_data_lo_lo_64};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_64 = {_alignedDequeue_bits_data_T_844[56], _alignedDequeue_bits_data_T_778[56]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_64 = {_alignedDequeue_bits_data_T_976[56], _alignedDequeue_bits_data_T_910[56]};
  wire [3:0]    alignedDequeue_bits_data_hi_64 = {alignedDequeue_bits_data_hi_hi_64, alignedDequeue_bits_data_hi_lo_64};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_65 = {_alignedDequeue_bits_data_T_580[57], _alignedDequeue_bits_data_T_514[57]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_65 = {_alignedDequeue_bits_data_T_712[57], _alignedDequeue_bits_data_T_646[57]};
  wire [3:0]    alignedDequeue_bits_data_lo_65 = {alignedDequeue_bits_data_lo_hi_65, alignedDequeue_bits_data_lo_lo_65};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_65 = {_alignedDequeue_bits_data_T_844[57], _alignedDequeue_bits_data_T_778[57]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_65 = {_alignedDequeue_bits_data_T_976[57], _alignedDequeue_bits_data_T_910[57]};
  wire [3:0]    alignedDequeue_bits_data_hi_65 = {alignedDequeue_bits_data_hi_hi_65, alignedDequeue_bits_data_hi_lo_65};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_66 = {_alignedDequeue_bits_data_T_580[58], _alignedDequeue_bits_data_T_514[58]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_66 = {_alignedDequeue_bits_data_T_712[58], _alignedDequeue_bits_data_T_646[58]};
  wire [3:0]    alignedDequeue_bits_data_lo_66 = {alignedDequeue_bits_data_lo_hi_66, alignedDequeue_bits_data_lo_lo_66};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_66 = {_alignedDequeue_bits_data_T_844[58], _alignedDequeue_bits_data_T_778[58]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_66 = {_alignedDequeue_bits_data_T_976[58], _alignedDequeue_bits_data_T_910[58]};
  wire [3:0]    alignedDequeue_bits_data_hi_66 = {alignedDequeue_bits_data_hi_hi_66, alignedDequeue_bits_data_hi_lo_66};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_67 = {_alignedDequeue_bits_data_T_580[59], _alignedDequeue_bits_data_T_514[59]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_67 = {_alignedDequeue_bits_data_T_712[59], _alignedDequeue_bits_data_T_646[59]};
  wire [3:0]    alignedDequeue_bits_data_lo_67 = {alignedDequeue_bits_data_lo_hi_67, alignedDequeue_bits_data_lo_lo_67};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_67 = {_alignedDequeue_bits_data_T_844[59], _alignedDequeue_bits_data_T_778[59]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_67 = {_alignedDequeue_bits_data_T_976[59], _alignedDequeue_bits_data_T_910[59]};
  wire [3:0]    alignedDequeue_bits_data_hi_67 = {alignedDequeue_bits_data_hi_hi_67, alignedDequeue_bits_data_hi_lo_67};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_68 = {_alignedDequeue_bits_data_T_580[60], _alignedDequeue_bits_data_T_514[60]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_68 = {_alignedDequeue_bits_data_T_712[60], _alignedDequeue_bits_data_T_646[60]};
  wire [3:0]    alignedDequeue_bits_data_lo_68 = {alignedDequeue_bits_data_lo_hi_68, alignedDequeue_bits_data_lo_lo_68};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_68 = {_alignedDequeue_bits_data_T_844[60], _alignedDequeue_bits_data_T_778[60]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_68 = {_alignedDequeue_bits_data_T_976[60], _alignedDequeue_bits_data_T_910[60]};
  wire [3:0]    alignedDequeue_bits_data_hi_68 = {alignedDequeue_bits_data_hi_hi_68, alignedDequeue_bits_data_hi_lo_68};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_69 = {_alignedDequeue_bits_data_T_580[61], _alignedDequeue_bits_data_T_514[61]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_69 = {_alignedDequeue_bits_data_T_712[61], _alignedDequeue_bits_data_T_646[61]};
  wire [3:0]    alignedDequeue_bits_data_lo_69 = {alignedDequeue_bits_data_lo_hi_69, alignedDequeue_bits_data_lo_lo_69};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_69 = {_alignedDequeue_bits_data_T_844[61], _alignedDequeue_bits_data_T_778[61]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_69 = {_alignedDequeue_bits_data_T_976[61], _alignedDequeue_bits_data_T_910[61]};
  wire [3:0]    alignedDequeue_bits_data_hi_69 = {alignedDequeue_bits_data_hi_hi_69, alignedDequeue_bits_data_hi_lo_69};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_70 = {_alignedDequeue_bits_data_T_580[62], _alignedDequeue_bits_data_T_514[62]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_70 = {_alignedDequeue_bits_data_T_712[62], _alignedDequeue_bits_data_T_646[62]};
  wire [3:0]    alignedDequeue_bits_data_lo_70 = {alignedDequeue_bits_data_lo_hi_70, alignedDequeue_bits_data_lo_lo_70};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_70 = {_alignedDequeue_bits_data_T_844[62], _alignedDequeue_bits_data_T_778[62]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_70 = {_alignedDequeue_bits_data_T_976[62], _alignedDequeue_bits_data_T_910[62]};
  wire [3:0]    alignedDequeue_bits_data_hi_70 = {alignedDequeue_bits_data_hi_hi_70, alignedDequeue_bits_data_hi_lo_70};
  wire [1:0]    alignedDequeue_bits_data_lo_lo_71 = {_alignedDequeue_bits_data_T_580[63], _alignedDequeue_bits_data_T_514[63]};
  wire [1:0]    alignedDequeue_bits_data_lo_hi_71 = {_alignedDequeue_bits_data_T_712[63], _alignedDequeue_bits_data_T_646[63]};
  wire [3:0]    alignedDequeue_bits_data_lo_71 = {alignedDequeue_bits_data_lo_hi_71, alignedDequeue_bits_data_lo_lo_71};
  wire [1:0]    alignedDequeue_bits_data_hi_lo_71 = {_alignedDequeue_bits_data_T_844[63], _alignedDequeue_bits_data_T_778[63]};
  wire [1:0]    alignedDequeue_bits_data_hi_hi_71 = {_alignedDequeue_bits_data_T_976[63], _alignedDequeue_bits_data_T_910[63]};
  wire [3:0]    alignedDequeue_bits_data_hi_71 = {alignedDequeue_bits_data_hi_hi_71, alignedDequeue_bits_data_hi_lo_71};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_9, alignedDequeue_bits_data_lo_9, alignedDequeue_bits_data_hi_8, alignedDequeue_bits_data_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_11, alignedDequeue_bits_data_lo_11, alignedDequeue_bits_data_hi_10, alignedDequeue_bits_data_lo_10};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_lo_lo_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_13, alignedDequeue_bits_data_lo_13, alignedDequeue_bits_data_hi_12, alignedDequeue_bits_data_lo_12};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_15, alignedDequeue_bits_data_lo_15, alignedDequeue_bits_data_hi_14, alignedDequeue_bits_data_lo_14};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_lo_lo_lo_hi_hi_8, alignedDequeue_bits_data_lo_lo_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_lo_lo_8 = {alignedDequeue_bits_data_lo_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_17, alignedDequeue_bits_data_lo_17, alignedDequeue_bits_data_hi_16, alignedDequeue_bits_data_lo_16};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_19, alignedDequeue_bits_data_lo_19, alignedDequeue_bits_data_hi_18, alignedDequeue_bits_data_lo_18};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_lo_lo_hi_lo_hi_8, alignedDequeue_bits_data_lo_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_21, alignedDequeue_bits_data_lo_21, alignedDequeue_bits_data_hi_20, alignedDequeue_bits_data_lo_20};
  wire [15:0]   alignedDequeue_bits_data_lo_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_23, alignedDequeue_bits_data_lo_23, alignedDequeue_bits_data_hi_22, alignedDequeue_bits_data_lo_22};
  wire [31:0]   alignedDequeue_bits_data_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_lo_lo_hi_hi_hi_8, alignedDequeue_bits_data_lo_lo_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_lo_hi_8 = {alignedDequeue_bits_data_lo_lo_hi_hi_8, alignedDequeue_bits_data_lo_lo_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_lo_lo_72 = {alignedDequeue_bits_data_lo_lo_hi_8, alignedDequeue_bits_data_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_25, alignedDequeue_bits_data_lo_25, alignedDequeue_bits_data_hi_24, alignedDequeue_bits_data_lo_24};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_27, alignedDequeue_bits_data_lo_27, alignedDequeue_bits_data_hi_26, alignedDequeue_bits_data_lo_26};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_lo_hi_lo_lo_hi_8, alignedDequeue_bits_data_lo_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_29, alignedDequeue_bits_data_lo_29, alignedDequeue_bits_data_hi_28, alignedDequeue_bits_data_lo_28};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_31, alignedDequeue_bits_data_lo_31, alignedDequeue_bits_data_hi_30, alignedDequeue_bits_data_lo_30};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_lo_hi_lo_hi_hi_8, alignedDequeue_bits_data_lo_hi_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_hi_lo_8 = {alignedDequeue_bits_data_lo_hi_lo_hi_8, alignedDequeue_bits_data_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_33, alignedDequeue_bits_data_lo_33, alignedDequeue_bits_data_hi_32, alignedDequeue_bits_data_lo_32};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_35, alignedDequeue_bits_data_lo_35, alignedDequeue_bits_data_hi_34, alignedDequeue_bits_data_lo_34};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_lo_hi_hi_lo_hi_8, alignedDequeue_bits_data_lo_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_37, alignedDequeue_bits_data_lo_37, alignedDequeue_bits_data_hi_36, alignedDequeue_bits_data_lo_36};
  wire [15:0]   alignedDequeue_bits_data_lo_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_39, alignedDequeue_bits_data_lo_39, alignedDequeue_bits_data_hi_38, alignedDequeue_bits_data_lo_38};
  wire [31:0]   alignedDequeue_bits_data_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_lo_hi_hi_hi_hi_8, alignedDequeue_bits_data_lo_hi_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_lo_hi_hi_8 = {alignedDequeue_bits_data_lo_hi_hi_hi_8, alignedDequeue_bits_data_lo_hi_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_lo_hi_72 = {alignedDequeue_bits_data_lo_hi_hi_8, alignedDequeue_bits_data_lo_hi_lo_8};
  assign alignedDequeue_bits_data_lo_72 = {alignedDequeue_bits_data_lo_hi_72, alignedDequeue_bits_data_lo_lo_72};
  wire [255:0]  alignedDequeue_bits_data = alignedDequeue_bits_data_lo_72;
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_41, alignedDequeue_bits_data_lo_41, alignedDequeue_bits_data_hi_40, alignedDequeue_bits_data_lo_40};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_43, alignedDequeue_bits_data_lo_43, alignedDequeue_bits_data_hi_42, alignedDequeue_bits_data_lo_42};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_lo_lo_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_45, alignedDequeue_bits_data_lo_45, alignedDequeue_bits_data_hi_44, alignedDequeue_bits_data_lo_44};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_47, alignedDequeue_bits_data_lo_47, alignedDequeue_bits_data_hi_46, alignedDequeue_bits_data_lo_46};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_lo_lo_hi_hi_8, alignedDequeue_bits_data_hi_lo_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_lo_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_49, alignedDequeue_bits_data_lo_49, alignedDequeue_bits_data_hi_48, alignedDequeue_bits_data_lo_48};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_51, alignedDequeue_bits_data_lo_51, alignedDequeue_bits_data_hi_50, alignedDequeue_bits_data_lo_50};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_lo_hi_lo_hi_8, alignedDequeue_bits_data_hi_lo_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_53, alignedDequeue_bits_data_lo_53, alignedDequeue_bits_data_hi_52, alignedDequeue_bits_data_lo_52};
  wire [15:0]   alignedDequeue_bits_data_hi_lo_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_55, alignedDequeue_bits_data_lo_55, alignedDequeue_bits_data_hi_54, alignedDequeue_bits_data_lo_54};
  wire [31:0]   alignedDequeue_bits_data_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_lo_hi_hi_hi_8, alignedDequeue_bits_data_hi_lo_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_lo_hi_hi_8, alignedDequeue_bits_data_hi_lo_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_hi_lo_72 = {alignedDequeue_bits_data_hi_lo_hi_8, alignedDequeue_bits_data_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_lo_lo_8 = {alignedDequeue_bits_data_hi_57, alignedDequeue_bits_data_lo_57, alignedDequeue_bits_data_hi_56, alignedDequeue_bits_data_lo_56};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_lo_hi_8 = {alignedDequeue_bits_data_hi_59, alignedDequeue_bits_data_lo_59, alignedDequeue_bits_data_hi_58, alignedDequeue_bits_data_lo_58};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_hi_lo_lo_hi_8, alignedDequeue_bits_data_hi_hi_lo_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_hi_lo_8 = {alignedDequeue_bits_data_hi_61, alignedDequeue_bits_data_lo_61, alignedDequeue_bits_data_hi_60, alignedDequeue_bits_data_lo_60};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_lo_hi_hi_8 = {alignedDequeue_bits_data_hi_63, alignedDequeue_bits_data_lo_63, alignedDequeue_bits_data_hi_62, alignedDequeue_bits_data_lo_62};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_hi_lo_hi_hi_8, alignedDequeue_bits_data_hi_hi_lo_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_hi_lo_hi_8, alignedDequeue_bits_data_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_lo_lo_8 = {alignedDequeue_bits_data_hi_65, alignedDequeue_bits_data_lo_65, alignedDequeue_bits_data_hi_64, alignedDequeue_bits_data_lo_64};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_lo_hi_8 = {alignedDequeue_bits_data_hi_67, alignedDequeue_bits_data_lo_67, alignedDequeue_bits_data_hi_66, alignedDequeue_bits_data_lo_66};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_hi_hi_lo_hi_8, alignedDequeue_bits_data_hi_hi_hi_lo_lo_8};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_hi_lo_8 = {alignedDequeue_bits_data_hi_69, alignedDequeue_bits_data_lo_69, alignedDequeue_bits_data_hi_68, alignedDequeue_bits_data_lo_68};
  wire [15:0]   alignedDequeue_bits_data_hi_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_71, alignedDequeue_bits_data_lo_71, alignedDequeue_bits_data_hi_70, alignedDequeue_bits_data_lo_70};
  wire [31:0]   alignedDequeue_bits_data_hi_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_hi_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_hi_hi_lo_8};
  wire [63:0]   alignedDequeue_bits_data_hi_hi_hi_8 = {alignedDequeue_bits_data_hi_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_hi_lo_8};
  wire [127:0]  alignedDequeue_bits_data_hi_hi_72 = {alignedDequeue_bits_data_hi_hi_hi_8, alignedDequeue_bits_data_hi_hi_lo_8};
  wire [255:0]  alignedDequeue_bits_data_hi_72 = {alignedDequeue_bits_data_hi_hi_72, alignedDequeue_bits_data_hi_lo_72};
  reg           bufferFull;
  wire          bufferTailFire;
  wire          bufferDequeueValid = bufferFull | bufferTailFire;
  wire          writeStageReady;
  wire          bufferDequeueReady;
  wire          bufferDequeueFire = bufferDequeueReady & bufferDequeueValid;
  assign alignedDequeue_ready = ~bufferFull;
  wire [7:0]    bufferEnqueueSelect = _bufferTailFire_T ? 8'h1 << cacheLineIndexInBuffer : 8'h0;
  wire [255:0]  dataBufferUpdate_0 = bufferEnqueueSelect[0] ? alignedDequeue_bits_data : dataBuffer_0;
  wire [255:0]  dataBufferUpdate_1 = bufferEnqueueSelect[1] ? alignedDequeue_bits_data : dataBuffer_1;
  wire [255:0]  dataBufferUpdate_2 = bufferEnqueueSelect[2] ? alignedDequeue_bits_data : dataBuffer_2;
  wire [255:0]  dataBufferUpdate_3 = bufferEnqueueSelect[3] ? alignedDequeue_bits_data : dataBuffer_3;
  wire [255:0]  dataBufferUpdate_4 = bufferEnqueueSelect[4] ? alignedDequeue_bits_data : dataBuffer_4;
  wire [255:0]  dataBufferUpdate_5 = bufferEnqueueSelect[5] ? alignedDequeue_bits_data : dataBuffer_5;
  wire [255:0]  dataBufferUpdate_6 = bufferEnqueueSelect[6] ? alignedDequeue_bits_data : dataBuffer_6;
  wire [255:0]  dataBufferUpdate_7 = bufferEnqueueSelect[7] ? alignedDequeue_bits_data : dataBuffer_7;
  wire [255:0]  dataSelect_0 = bufferFull ? dataBuffer_0 : dataBufferUpdate_0;
  wire [255:0]  dataSelect_1 = bufferFull ? dataBuffer_1 : dataBufferUpdate_1;
  wire [255:0]  dataSelect_2 = bufferFull ? dataBuffer_2 : dataBufferUpdate_2;
  wire [255:0]  dataSelect_3 = bufferFull ? dataBuffer_3 : dataBufferUpdate_3;
  wire [255:0]  dataSelect_4 = bufferFull ? dataBuffer_4 : dataBufferUpdate_4;
  wire [255:0]  dataSelect_5 = bufferFull ? dataBuffer_5 : dataBufferUpdate_5;
  wire [255:0]  dataSelect_6 = bufferFull ? dataBuffer_6 : dataBufferUpdate_6;
  wire [255:0]  dataSelect_7 = bufferFull ? dataBuffer_7 : dataBufferUpdate_7;
  wire          lastCacheLineForThisGroup = cacheLineIndexInBuffer == lsuRequestReg_instructionInformation_nf;
  wire          lastCacheLineForInst = {7'h0, alignedDequeue_bits_index} == lastWriteVrfIndexReg;
  assign bufferTailFire = _bufferTailFire_T & (lastCacheLineForThisGroup | lastCacheLineForInst);
  reg           waitForFirstDataGroup;
  wire          lastPtr = accessPtr == 3'h0;
  assign writeStageReady = lastPtr & accessStateCheck;
  assign bufferDequeueReady = writeStageReady;
  wire          _maskSelect_valid_output = bufferDequeueFire & isLastDataGroup;
  wire [511:0]  _GEN_4 = {dataSelect_1, dataSelect_0};
  wire [511:0]  dataGroup_lo_lo;
  assign dataGroup_lo_lo = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1;
  assign dataGroup_lo_lo_1 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2;
  assign dataGroup_lo_lo_2 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_3;
  assign dataGroup_lo_lo_3 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_4;
  assign dataGroup_lo_lo_4 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_5;
  assign dataGroup_lo_lo_5 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_6;
  assign dataGroup_lo_lo_6 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_7;
  assign dataGroup_lo_lo_7 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_8;
  assign dataGroup_lo_lo_8 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_9;
  assign dataGroup_lo_lo_9 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_10;
  assign dataGroup_lo_lo_10 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_11;
  assign dataGroup_lo_lo_11 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_12;
  assign dataGroup_lo_lo_12 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_13;
  assign dataGroup_lo_lo_13 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_14;
  assign dataGroup_lo_lo_14 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_15;
  assign dataGroup_lo_lo_15 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_16;
  assign dataGroup_lo_lo_16 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_17;
  assign dataGroup_lo_lo_17 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_18;
  assign dataGroup_lo_lo_18 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_19;
  assign dataGroup_lo_lo_19 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_20;
  assign dataGroup_lo_lo_20 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_21;
  assign dataGroup_lo_lo_21 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_22;
  assign dataGroup_lo_lo_22 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_23;
  assign dataGroup_lo_lo_23 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_24;
  assign dataGroup_lo_lo_24 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_25;
  assign dataGroup_lo_lo_25 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_26;
  assign dataGroup_lo_lo_26 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_27;
  assign dataGroup_lo_lo_27 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_28;
  assign dataGroup_lo_lo_28 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_29;
  assign dataGroup_lo_lo_29 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_30;
  assign dataGroup_lo_lo_30 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_31;
  assign dataGroup_lo_lo_31 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_32;
  assign dataGroup_lo_lo_32 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_33;
  assign dataGroup_lo_lo_33 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_34;
  assign dataGroup_lo_lo_34 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_35;
  assign dataGroup_lo_lo_35 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_36;
  assign dataGroup_lo_lo_36 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_37;
  assign dataGroup_lo_lo_37 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_38;
  assign dataGroup_lo_lo_38 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_39;
  assign dataGroup_lo_lo_39 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_40;
  assign dataGroup_lo_lo_40 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_41;
  assign dataGroup_lo_lo_41 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_42;
  assign dataGroup_lo_lo_42 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_43;
  assign dataGroup_lo_lo_43 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_44;
  assign dataGroup_lo_lo_44 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_45;
  assign dataGroup_lo_lo_45 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_46;
  assign dataGroup_lo_lo_46 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_47;
  assign dataGroup_lo_lo_47 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_48;
  assign dataGroup_lo_lo_48 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_49;
  assign dataGroup_lo_lo_49 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_50;
  assign dataGroup_lo_lo_50 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_51;
  assign dataGroup_lo_lo_51 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_52;
  assign dataGroup_lo_lo_52 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_53;
  assign dataGroup_lo_lo_53 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_54;
  assign dataGroup_lo_lo_54 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_55;
  assign dataGroup_lo_lo_55 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_56;
  assign dataGroup_lo_lo_56 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_57;
  assign dataGroup_lo_lo_57 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_58;
  assign dataGroup_lo_lo_58 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_59;
  assign dataGroup_lo_lo_59 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_60;
  assign dataGroup_lo_lo_60 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_61;
  assign dataGroup_lo_lo_61 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_62;
  assign dataGroup_lo_lo_62 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_63;
  assign dataGroup_lo_lo_63 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_64;
  assign dataGroup_lo_lo_64 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_65;
  assign dataGroup_lo_lo_65 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_66;
  assign dataGroup_lo_lo_66 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_67;
  assign dataGroup_lo_lo_67 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_68;
  assign dataGroup_lo_lo_68 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_69;
  assign dataGroup_lo_lo_69 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_70;
  assign dataGroup_lo_lo_70 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_71;
  assign dataGroup_lo_lo_71 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_72;
  assign dataGroup_lo_lo_72 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_73;
  assign dataGroup_lo_lo_73 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_74;
  assign dataGroup_lo_lo_74 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_75;
  assign dataGroup_lo_lo_75 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_76;
  assign dataGroup_lo_lo_76 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_77;
  assign dataGroup_lo_lo_77 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_78;
  assign dataGroup_lo_lo_78 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_79;
  assign dataGroup_lo_lo_79 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_80;
  assign dataGroup_lo_lo_80 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_81;
  assign dataGroup_lo_lo_81 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_82;
  assign dataGroup_lo_lo_82 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_83;
  assign dataGroup_lo_lo_83 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_84;
  assign dataGroup_lo_lo_84 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_85;
  assign dataGroup_lo_lo_85 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_86;
  assign dataGroup_lo_lo_86 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_87;
  assign dataGroup_lo_lo_87 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_88;
  assign dataGroup_lo_lo_88 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_89;
  assign dataGroup_lo_lo_89 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_90;
  assign dataGroup_lo_lo_90 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_91;
  assign dataGroup_lo_lo_91 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_92;
  assign dataGroup_lo_lo_92 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_93;
  assign dataGroup_lo_lo_93 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_94;
  assign dataGroup_lo_lo_94 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_95;
  assign dataGroup_lo_lo_95 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_96;
  assign dataGroup_lo_lo_96 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_97;
  assign dataGroup_lo_lo_97 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_98;
  assign dataGroup_lo_lo_98 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_99;
  assign dataGroup_lo_lo_99 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_100;
  assign dataGroup_lo_lo_100 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_101;
  assign dataGroup_lo_lo_101 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_102;
  assign dataGroup_lo_lo_102 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_103;
  assign dataGroup_lo_lo_103 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_104;
  assign dataGroup_lo_lo_104 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_105;
  assign dataGroup_lo_lo_105 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_106;
  assign dataGroup_lo_lo_106 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_107;
  assign dataGroup_lo_lo_107 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_108;
  assign dataGroup_lo_lo_108 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_109;
  assign dataGroup_lo_lo_109 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_110;
  assign dataGroup_lo_lo_110 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_111;
  assign dataGroup_lo_lo_111 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_112;
  assign dataGroup_lo_lo_112 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_113;
  assign dataGroup_lo_lo_113 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_114;
  assign dataGroup_lo_lo_114 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_115;
  assign dataGroup_lo_lo_115 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_116;
  assign dataGroup_lo_lo_116 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_117;
  assign dataGroup_lo_lo_117 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_118;
  assign dataGroup_lo_lo_118 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_119;
  assign dataGroup_lo_lo_119 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_120;
  assign dataGroup_lo_lo_120 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_121;
  assign dataGroup_lo_lo_121 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_122;
  assign dataGroup_lo_lo_122 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_123;
  assign dataGroup_lo_lo_123 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_124;
  assign dataGroup_lo_lo_124 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_125;
  assign dataGroup_lo_lo_125 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_126;
  assign dataGroup_lo_lo_126 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_127;
  assign dataGroup_lo_lo_127 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_128;
  assign dataGroup_lo_lo_128 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_129;
  assign dataGroup_lo_lo_129 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_130;
  assign dataGroup_lo_lo_130 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_131;
  assign dataGroup_lo_lo_131 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_132;
  assign dataGroup_lo_lo_132 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_133;
  assign dataGroup_lo_lo_133 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_134;
  assign dataGroup_lo_lo_134 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_135;
  assign dataGroup_lo_lo_135 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_136;
  assign dataGroup_lo_lo_136 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_137;
  assign dataGroup_lo_lo_137 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_138;
  assign dataGroup_lo_lo_138 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_139;
  assign dataGroup_lo_lo_139 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_140;
  assign dataGroup_lo_lo_140 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_141;
  assign dataGroup_lo_lo_141 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_142;
  assign dataGroup_lo_lo_142 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_143;
  assign dataGroup_lo_lo_143 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_144;
  assign dataGroup_lo_lo_144 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_145;
  assign dataGroup_lo_lo_145 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_146;
  assign dataGroup_lo_lo_146 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_147;
  assign dataGroup_lo_lo_147 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_148;
  assign dataGroup_lo_lo_148 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_149;
  assign dataGroup_lo_lo_149 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_150;
  assign dataGroup_lo_lo_150 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_151;
  assign dataGroup_lo_lo_151 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_152;
  assign dataGroup_lo_lo_152 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_153;
  assign dataGroup_lo_lo_153 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_154;
  assign dataGroup_lo_lo_154 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_155;
  assign dataGroup_lo_lo_155 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_156;
  assign dataGroup_lo_lo_156 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_157;
  assign dataGroup_lo_lo_157 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_158;
  assign dataGroup_lo_lo_158 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_159;
  assign dataGroup_lo_lo_159 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_160;
  assign dataGroup_lo_lo_160 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_161;
  assign dataGroup_lo_lo_161 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_162;
  assign dataGroup_lo_lo_162 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_163;
  assign dataGroup_lo_lo_163 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_164;
  assign dataGroup_lo_lo_164 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_165;
  assign dataGroup_lo_lo_165 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_166;
  assign dataGroup_lo_lo_166 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_167;
  assign dataGroup_lo_lo_167 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_168;
  assign dataGroup_lo_lo_168 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_169;
  assign dataGroup_lo_lo_169 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_170;
  assign dataGroup_lo_lo_170 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_171;
  assign dataGroup_lo_lo_171 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_172;
  assign dataGroup_lo_lo_172 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_173;
  assign dataGroup_lo_lo_173 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_174;
  assign dataGroup_lo_lo_174 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_175;
  assign dataGroup_lo_lo_175 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_176;
  assign dataGroup_lo_lo_176 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_177;
  assign dataGroup_lo_lo_177 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_178;
  assign dataGroup_lo_lo_178 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_179;
  assign dataGroup_lo_lo_179 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_180;
  assign dataGroup_lo_lo_180 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_181;
  assign dataGroup_lo_lo_181 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_182;
  assign dataGroup_lo_lo_182 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_183;
  assign dataGroup_lo_lo_183 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_184;
  assign dataGroup_lo_lo_184 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_185;
  assign dataGroup_lo_lo_185 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_186;
  assign dataGroup_lo_lo_186 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_187;
  assign dataGroup_lo_lo_187 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_188;
  assign dataGroup_lo_lo_188 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_189;
  assign dataGroup_lo_lo_189 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_190;
  assign dataGroup_lo_lo_190 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_191;
  assign dataGroup_lo_lo_191 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_192;
  assign dataGroup_lo_lo_192 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_193;
  assign dataGroup_lo_lo_193 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_194;
  assign dataGroup_lo_lo_194 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_195;
  assign dataGroup_lo_lo_195 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_196;
  assign dataGroup_lo_lo_196 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_197;
  assign dataGroup_lo_lo_197 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_198;
  assign dataGroup_lo_lo_198 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_199;
  assign dataGroup_lo_lo_199 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_200;
  assign dataGroup_lo_lo_200 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_201;
  assign dataGroup_lo_lo_201 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_202;
  assign dataGroup_lo_lo_202 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_203;
  assign dataGroup_lo_lo_203 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_204;
  assign dataGroup_lo_lo_204 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_205;
  assign dataGroup_lo_lo_205 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_206;
  assign dataGroup_lo_lo_206 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_207;
  assign dataGroup_lo_lo_207 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_208;
  assign dataGroup_lo_lo_208 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_209;
  assign dataGroup_lo_lo_209 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_210;
  assign dataGroup_lo_lo_210 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_211;
  assign dataGroup_lo_lo_211 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_212;
  assign dataGroup_lo_lo_212 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_213;
  assign dataGroup_lo_lo_213 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_214;
  assign dataGroup_lo_lo_214 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_215;
  assign dataGroup_lo_lo_215 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_216;
  assign dataGroup_lo_lo_216 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_217;
  assign dataGroup_lo_lo_217 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_218;
  assign dataGroup_lo_lo_218 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_219;
  assign dataGroup_lo_lo_219 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_220;
  assign dataGroup_lo_lo_220 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_221;
  assign dataGroup_lo_lo_221 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_222;
  assign dataGroup_lo_lo_222 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_223;
  assign dataGroup_lo_lo_223 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_224;
  assign dataGroup_lo_lo_224 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_225;
  assign dataGroup_lo_lo_225 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_226;
  assign dataGroup_lo_lo_226 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_227;
  assign dataGroup_lo_lo_227 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_228;
  assign dataGroup_lo_lo_228 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_229;
  assign dataGroup_lo_lo_229 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_230;
  assign dataGroup_lo_lo_230 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_231;
  assign dataGroup_lo_lo_231 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_232;
  assign dataGroup_lo_lo_232 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_233;
  assign dataGroup_lo_lo_233 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_234;
  assign dataGroup_lo_lo_234 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_235;
  assign dataGroup_lo_lo_235 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_236;
  assign dataGroup_lo_lo_236 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_237;
  assign dataGroup_lo_lo_237 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_238;
  assign dataGroup_lo_lo_238 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_239;
  assign dataGroup_lo_lo_239 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_240;
  assign dataGroup_lo_lo_240 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_241;
  assign dataGroup_lo_lo_241 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_242;
  assign dataGroup_lo_lo_242 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_243;
  assign dataGroup_lo_lo_243 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_244;
  assign dataGroup_lo_lo_244 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_245;
  assign dataGroup_lo_lo_245 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_246;
  assign dataGroup_lo_lo_246 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_247;
  assign dataGroup_lo_lo_247 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_248;
  assign dataGroup_lo_lo_248 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_249;
  assign dataGroup_lo_lo_249 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_250;
  assign dataGroup_lo_lo_250 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_251;
  assign dataGroup_lo_lo_251 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_252;
  assign dataGroup_lo_lo_252 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_253;
  assign dataGroup_lo_lo_253 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_254;
  assign dataGroup_lo_lo_254 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_255;
  assign dataGroup_lo_lo_255 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_256;
  assign dataGroup_lo_lo_256 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_257;
  assign dataGroup_lo_lo_257 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_258;
  assign dataGroup_lo_lo_258 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_259;
  assign dataGroup_lo_lo_259 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_260;
  assign dataGroup_lo_lo_260 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_261;
  assign dataGroup_lo_lo_261 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_262;
  assign dataGroup_lo_lo_262 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_263;
  assign dataGroup_lo_lo_263 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_264;
  assign dataGroup_lo_lo_264 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_265;
  assign dataGroup_lo_lo_265 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_266;
  assign dataGroup_lo_lo_266 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_267;
  assign dataGroup_lo_lo_267 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_268;
  assign dataGroup_lo_lo_268 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_269;
  assign dataGroup_lo_lo_269 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_270;
  assign dataGroup_lo_lo_270 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_271;
  assign dataGroup_lo_lo_271 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_272;
  assign dataGroup_lo_lo_272 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_273;
  assign dataGroup_lo_lo_273 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_274;
  assign dataGroup_lo_lo_274 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_275;
  assign dataGroup_lo_lo_275 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_276;
  assign dataGroup_lo_lo_276 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_277;
  assign dataGroup_lo_lo_277 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_278;
  assign dataGroup_lo_lo_278 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_279;
  assign dataGroup_lo_lo_279 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_280;
  assign dataGroup_lo_lo_280 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_281;
  assign dataGroup_lo_lo_281 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_282;
  assign dataGroup_lo_lo_282 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_283;
  assign dataGroup_lo_lo_283 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_284;
  assign dataGroup_lo_lo_284 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_285;
  assign dataGroup_lo_lo_285 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_286;
  assign dataGroup_lo_lo_286 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_287;
  assign dataGroup_lo_lo_287 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_288;
  assign dataGroup_lo_lo_288 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_289;
  assign dataGroup_lo_lo_289 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_290;
  assign dataGroup_lo_lo_290 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_291;
  assign dataGroup_lo_lo_291 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_292;
  assign dataGroup_lo_lo_292 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_293;
  assign dataGroup_lo_lo_293 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_294;
  assign dataGroup_lo_lo_294 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_295;
  assign dataGroup_lo_lo_295 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_296;
  assign dataGroup_lo_lo_296 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_297;
  assign dataGroup_lo_lo_297 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_298;
  assign dataGroup_lo_lo_298 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_299;
  assign dataGroup_lo_lo_299 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_300;
  assign dataGroup_lo_lo_300 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_301;
  assign dataGroup_lo_lo_301 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_302;
  assign dataGroup_lo_lo_302 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_303;
  assign dataGroup_lo_lo_303 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_304;
  assign dataGroup_lo_lo_304 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_305;
  assign dataGroup_lo_lo_305 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_306;
  assign dataGroup_lo_lo_306 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_307;
  assign dataGroup_lo_lo_307 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_308;
  assign dataGroup_lo_lo_308 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_309;
  assign dataGroup_lo_lo_309 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_310;
  assign dataGroup_lo_lo_310 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_311;
  assign dataGroup_lo_lo_311 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_312;
  assign dataGroup_lo_lo_312 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_313;
  assign dataGroup_lo_lo_313 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_314;
  assign dataGroup_lo_lo_314 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_315;
  assign dataGroup_lo_lo_315 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_316;
  assign dataGroup_lo_lo_316 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_317;
  assign dataGroup_lo_lo_317 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_318;
  assign dataGroup_lo_lo_318 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_319;
  assign dataGroup_lo_lo_319 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_320;
  assign dataGroup_lo_lo_320 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_321;
  assign dataGroup_lo_lo_321 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_322;
  assign dataGroup_lo_lo_322 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_323;
  assign dataGroup_lo_lo_323 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_324;
  assign dataGroup_lo_lo_324 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_325;
  assign dataGroup_lo_lo_325 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_326;
  assign dataGroup_lo_lo_326 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_327;
  assign dataGroup_lo_lo_327 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_328;
  assign dataGroup_lo_lo_328 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_329;
  assign dataGroup_lo_lo_329 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_330;
  assign dataGroup_lo_lo_330 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_331;
  assign dataGroup_lo_lo_331 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_332;
  assign dataGroup_lo_lo_332 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_333;
  assign dataGroup_lo_lo_333 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_334;
  assign dataGroup_lo_lo_334 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_335;
  assign dataGroup_lo_lo_335 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_336;
  assign dataGroup_lo_lo_336 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_337;
  assign dataGroup_lo_lo_337 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_338;
  assign dataGroup_lo_lo_338 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_339;
  assign dataGroup_lo_lo_339 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_340;
  assign dataGroup_lo_lo_340 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_341;
  assign dataGroup_lo_lo_341 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_342;
  assign dataGroup_lo_lo_342 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_343;
  assign dataGroup_lo_lo_343 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_344;
  assign dataGroup_lo_lo_344 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_345;
  assign dataGroup_lo_lo_345 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_346;
  assign dataGroup_lo_lo_346 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_347;
  assign dataGroup_lo_lo_347 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_348;
  assign dataGroup_lo_lo_348 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_349;
  assign dataGroup_lo_lo_349 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_350;
  assign dataGroup_lo_lo_350 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_351;
  assign dataGroup_lo_lo_351 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_352;
  assign dataGroup_lo_lo_352 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_353;
  assign dataGroup_lo_lo_353 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_354;
  assign dataGroup_lo_lo_354 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_355;
  assign dataGroup_lo_lo_355 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_356;
  assign dataGroup_lo_lo_356 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_357;
  assign dataGroup_lo_lo_357 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_358;
  assign dataGroup_lo_lo_358 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_359;
  assign dataGroup_lo_lo_359 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_360;
  assign dataGroup_lo_lo_360 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_361;
  assign dataGroup_lo_lo_361 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_362;
  assign dataGroup_lo_lo_362 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_363;
  assign dataGroup_lo_lo_363 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_364;
  assign dataGroup_lo_lo_364 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_365;
  assign dataGroup_lo_lo_365 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_366;
  assign dataGroup_lo_lo_366 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_367;
  assign dataGroup_lo_lo_367 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_368;
  assign dataGroup_lo_lo_368 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_369;
  assign dataGroup_lo_lo_369 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_370;
  assign dataGroup_lo_lo_370 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_371;
  assign dataGroup_lo_lo_371 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_372;
  assign dataGroup_lo_lo_372 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_373;
  assign dataGroup_lo_lo_373 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_374;
  assign dataGroup_lo_lo_374 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_375;
  assign dataGroup_lo_lo_375 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_376;
  assign dataGroup_lo_lo_376 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_377;
  assign dataGroup_lo_lo_377 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_378;
  assign dataGroup_lo_lo_378 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_379;
  assign dataGroup_lo_lo_379 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_380;
  assign dataGroup_lo_lo_380 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_381;
  assign dataGroup_lo_lo_381 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_382;
  assign dataGroup_lo_lo_382 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_383;
  assign dataGroup_lo_lo_383 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_384;
  assign dataGroup_lo_lo_384 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_385;
  assign dataGroup_lo_lo_385 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_386;
  assign dataGroup_lo_lo_386 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_387;
  assign dataGroup_lo_lo_387 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_388;
  assign dataGroup_lo_lo_388 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_389;
  assign dataGroup_lo_lo_389 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_390;
  assign dataGroup_lo_lo_390 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_391;
  assign dataGroup_lo_lo_391 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_392;
  assign dataGroup_lo_lo_392 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_393;
  assign dataGroup_lo_lo_393 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_394;
  assign dataGroup_lo_lo_394 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_395;
  assign dataGroup_lo_lo_395 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_396;
  assign dataGroup_lo_lo_396 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_397;
  assign dataGroup_lo_lo_397 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_398;
  assign dataGroup_lo_lo_398 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_399;
  assign dataGroup_lo_lo_399 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_400;
  assign dataGroup_lo_lo_400 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_401;
  assign dataGroup_lo_lo_401 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_402;
  assign dataGroup_lo_lo_402 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_403;
  assign dataGroup_lo_lo_403 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_404;
  assign dataGroup_lo_lo_404 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_405;
  assign dataGroup_lo_lo_405 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_406;
  assign dataGroup_lo_lo_406 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_407;
  assign dataGroup_lo_lo_407 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_408;
  assign dataGroup_lo_lo_408 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_409;
  assign dataGroup_lo_lo_409 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_410;
  assign dataGroup_lo_lo_410 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_411;
  assign dataGroup_lo_lo_411 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_412;
  assign dataGroup_lo_lo_412 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_413;
  assign dataGroup_lo_lo_413 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_414;
  assign dataGroup_lo_lo_414 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_415;
  assign dataGroup_lo_lo_415 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_416;
  assign dataGroup_lo_lo_416 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_417;
  assign dataGroup_lo_lo_417 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_418;
  assign dataGroup_lo_lo_418 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_419;
  assign dataGroup_lo_lo_419 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_420;
  assign dataGroup_lo_lo_420 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_421;
  assign dataGroup_lo_lo_421 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_422;
  assign dataGroup_lo_lo_422 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_423;
  assign dataGroup_lo_lo_423 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_424;
  assign dataGroup_lo_lo_424 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_425;
  assign dataGroup_lo_lo_425 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_426;
  assign dataGroup_lo_lo_426 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_427;
  assign dataGroup_lo_lo_427 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_428;
  assign dataGroup_lo_lo_428 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_429;
  assign dataGroup_lo_lo_429 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_430;
  assign dataGroup_lo_lo_430 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_431;
  assign dataGroup_lo_lo_431 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_432;
  assign dataGroup_lo_lo_432 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_433;
  assign dataGroup_lo_lo_433 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_434;
  assign dataGroup_lo_lo_434 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_435;
  assign dataGroup_lo_lo_435 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_436;
  assign dataGroup_lo_lo_436 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_437;
  assign dataGroup_lo_lo_437 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_438;
  assign dataGroup_lo_lo_438 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_439;
  assign dataGroup_lo_lo_439 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_440;
  assign dataGroup_lo_lo_440 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_441;
  assign dataGroup_lo_lo_441 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_442;
  assign dataGroup_lo_lo_442 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_443;
  assign dataGroup_lo_lo_443 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_444;
  assign dataGroup_lo_lo_444 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_445;
  assign dataGroup_lo_lo_445 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_446;
  assign dataGroup_lo_lo_446 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_447;
  assign dataGroup_lo_lo_447 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_448;
  assign dataGroup_lo_lo_448 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_449;
  assign dataGroup_lo_lo_449 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_450;
  assign dataGroup_lo_lo_450 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_451;
  assign dataGroup_lo_lo_451 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_452;
  assign dataGroup_lo_lo_452 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_453;
  assign dataGroup_lo_lo_453 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_454;
  assign dataGroup_lo_lo_454 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_455;
  assign dataGroup_lo_lo_455 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_456;
  assign dataGroup_lo_lo_456 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_457;
  assign dataGroup_lo_lo_457 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_458;
  assign dataGroup_lo_lo_458 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_459;
  assign dataGroup_lo_lo_459 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_460;
  assign dataGroup_lo_lo_460 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_461;
  assign dataGroup_lo_lo_461 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_462;
  assign dataGroup_lo_lo_462 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_463;
  assign dataGroup_lo_lo_463 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_464;
  assign dataGroup_lo_lo_464 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_465;
  assign dataGroup_lo_lo_465 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_466;
  assign dataGroup_lo_lo_466 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_467;
  assign dataGroup_lo_lo_467 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_468;
  assign dataGroup_lo_lo_468 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_469;
  assign dataGroup_lo_lo_469 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_470;
  assign dataGroup_lo_lo_470 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_471;
  assign dataGroup_lo_lo_471 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_472;
  assign dataGroup_lo_lo_472 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_473;
  assign dataGroup_lo_lo_473 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_474;
  assign dataGroup_lo_lo_474 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_475;
  assign dataGroup_lo_lo_475 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_476;
  assign dataGroup_lo_lo_476 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_477;
  assign dataGroup_lo_lo_477 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_478;
  assign dataGroup_lo_lo_478 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_479;
  assign dataGroup_lo_lo_479 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_480;
  assign dataGroup_lo_lo_480 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_481;
  assign dataGroup_lo_lo_481 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_482;
  assign dataGroup_lo_lo_482 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_483;
  assign dataGroup_lo_lo_483 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_484;
  assign dataGroup_lo_lo_484 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_485;
  assign dataGroup_lo_lo_485 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_486;
  assign dataGroup_lo_lo_486 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_487;
  assign dataGroup_lo_lo_487 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_488;
  assign dataGroup_lo_lo_488 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_489;
  assign dataGroup_lo_lo_489 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_490;
  assign dataGroup_lo_lo_490 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_491;
  assign dataGroup_lo_lo_491 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_492;
  assign dataGroup_lo_lo_492 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_493;
  assign dataGroup_lo_lo_493 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_494;
  assign dataGroup_lo_lo_494 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_495;
  assign dataGroup_lo_lo_495 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_496;
  assign dataGroup_lo_lo_496 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_497;
  assign dataGroup_lo_lo_497 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_498;
  assign dataGroup_lo_lo_498 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_499;
  assign dataGroup_lo_lo_499 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_500;
  assign dataGroup_lo_lo_500 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_501;
  assign dataGroup_lo_lo_501 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_502;
  assign dataGroup_lo_lo_502 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_503;
  assign dataGroup_lo_lo_503 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_504;
  assign dataGroup_lo_lo_504 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_505;
  assign dataGroup_lo_lo_505 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_506;
  assign dataGroup_lo_lo_506 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_507;
  assign dataGroup_lo_lo_507 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_508;
  assign dataGroup_lo_lo_508 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_509;
  assign dataGroup_lo_lo_509 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_510;
  assign dataGroup_lo_lo_510 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_511;
  assign dataGroup_lo_lo_511 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_512;
  assign dataGroup_lo_lo_512 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_513;
  assign dataGroup_lo_lo_513 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_514;
  assign dataGroup_lo_lo_514 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_515;
  assign dataGroup_lo_lo_515 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_516;
  assign dataGroup_lo_lo_516 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_517;
  assign dataGroup_lo_lo_517 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_518;
  assign dataGroup_lo_lo_518 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_519;
  assign dataGroup_lo_lo_519 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_520;
  assign dataGroup_lo_lo_520 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_521;
  assign dataGroup_lo_lo_521 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_522;
  assign dataGroup_lo_lo_522 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_523;
  assign dataGroup_lo_lo_523 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_524;
  assign dataGroup_lo_lo_524 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_525;
  assign dataGroup_lo_lo_525 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_526;
  assign dataGroup_lo_lo_526 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_527;
  assign dataGroup_lo_lo_527 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_528;
  assign dataGroup_lo_lo_528 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_529;
  assign dataGroup_lo_lo_529 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_530;
  assign dataGroup_lo_lo_530 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_531;
  assign dataGroup_lo_lo_531 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_532;
  assign dataGroup_lo_lo_532 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_533;
  assign dataGroup_lo_lo_533 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_534;
  assign dataGroup_lo_lo_534 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_535;
  assign dataGroup_lo_lo_535 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_536;
  assign dataGroup_lo_lo_536 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_537;
  assign dataGroup_lo_lo_537 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_538;
  assign dataGroup_lo_lo_538 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_539;
  assign dataGroup_lo_lo_539 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_540;
  assign dataGroup_lo_lo_540 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_541;
  assign dataGroup_lo_lo_541 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_542;
  assign dataGroup_lo_lo_542 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_543;
  assign dataGroup_lo_lo_543 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_544;
  assign dataGroup_lo_lo_544 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_545;
  assign dataGroup_lo_lo_545 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_546;
  assign dataGroup_lo_lo_546 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_547;
  assign dataGroup_lo_lo_547 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_548;
  assign dataGroup_lo_lo_548 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_549;
  assign dataGroup_lo_lo_549 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_550;
  assign dataGroup_lo_lo_550 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_551;
  assign dataGroup_lo_lo_551 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_552;
  assign dataGroup_lo_lo_552 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_553;
  assign dataGroup_lo_lo_553 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_554;
  assign dataGroup_lo_lo_554 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_555;
  assign dataGroup_lo_lo_555 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_556;
  assign dataGroup_lo_lo_556 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_557;
  assign dataGroup_lo_lo_557 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_558;
  assign dataGroup_lo_lo_558 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_559;
  assign dataGroup_lo_lo_559 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_560;
  assign dataGroup_lo_lo_560 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_561;
  assign dataGroup_lo_lo_561 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_562;
  assign dataGroup_lo_lo_562 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_563;
  assign dataGroup_lo_lo_563 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_564;
  assign dataGroup_lo_lo_564 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_565;
  assign dataGroup_lo_lo_565 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_566;
  assign dataGroup_lo_lo_566 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_567;
  assign dataGroup_lo_lo_567 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_568;
  assign dataGroup_lo_lo_568 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_569;
  assign dataGroup_lo_lo_569 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_570;
  assign dataGroup_lo_lo_570 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_571;
  assign dataGroup_lo_lo_571 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_572;
  assign dataGroup_lo_lo_572 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_573;
  assign dataGroup_lo_lo_573 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_574;
  assign dataGroup_lo_lo_574 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_575;
  assign dataGroup_lo_lo_575 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_576;
  assign dataGroup_lo_lo_576 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_577;
  assign dataGroup_lo_lo_577 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_578;
  assign dataGroup_lo_lo_578 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_579;
  assign dataGroup_lo_lo_579 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_580;
  assign dataGroup_lo_lo_580 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_581;
  assign dataGroup_lo_lo_581 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_582;
  assign dataGroup_lo_lo_582 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_583;
  assign dataGroup_lo_lo_583 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_584;
  assign dataGroup_lo_lo_584 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_585;
  assign dataGroup_lo_lo_585 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_586;
  assign dataGroup_lo_lo_586 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_587;
  assign dataGroup_lo_lo_587 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_588;
  assign dataGroup_lo_lo_588 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_589;
  assign dataGroup_lo_lo_589 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_590;
  assign dataGroup_lo_lo_590 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_591;
  assign dataGroup_lo_lo_591 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_592;
  assign dataGroup_lo_lo_592 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_593;
  assign dataGroup_lo_lo_593 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_594;
  assign dataGroup_lo_lo_594 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_595;
  assign dataGroup_lo_lo_595 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_596;
  assign dataGroup_lo_lo_596 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_597;
  assign dataGroup_lo_lo_597 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_598;
  assign dataGroup_lo_lo_598 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_599;
  assign dataGroup_lo_lo_599 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_600;
  assign dataGroup_lo_lo_600 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_601;
  assign dataGroup_lo_lo_601 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_602;
  assign dataGroup_lo_lo_602 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_603;
  assign dataGroup_lo_lo_603 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_604;
  assign dataGroup_lo_lo_604 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_605;
  assign dataGroup_lo_lo_605 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_606;
  assign dataGroup_lo_lo_606 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_607;
  assign dataGroup_lo_lo_607 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_608;
  assign dataGroup_lo_lo_608 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_609;
  assign dataGroup_lo_lo_609 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_610;
  assign dataGroup_lo_lo_610 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_611;
  assign dataGroup_lo_lo_611 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_612;
  assign dataGroup_lo_lo_612 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_613;
  assign dataGroup_lo_lo_613 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_614;
  assign dataGroup_lo_lo_614 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_615;
  assign dataGroup_lo_lo_615 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_616;
  assign dataGroup_lo_lo_616 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_617;
  assign dataGroup_lo_lo_617 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_618;
  assign dataGroup_lo_lo_618 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_619;
  assign dataGroup_lo_lo_619 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_620;
  assign dataGroup_lo_lo_620 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_621;
  assign dataGroup_lo_lo_621 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_622;
  assign dataGroup_lo_lo_622 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_623;
  assign dataGroup_lo_lo_623 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_624;
  assign dataGroup_lo_lo_624 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_625;
  assign dataGroup_lo_lo_625 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_626;
  assign dataGroup_lo_lo_626 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_627;
  assign dataGroup_lo_lo_627 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_628;
  assign dataGroup_lo_lo_628 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_629;
  assign dataGroup_lo_lo_629 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_630;
  assign dataGroup_lo_lo_630 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_631;
  assign dataGroup_lo_lo_631 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_632;
  assign dataGroup_lo_lo_632 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_633;
  assign dataGroup_lo_lo_633 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_634;
  assign dataGroup_lo_lo_634 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_635;
  assign dataGroup_lo_lo_635 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_636;
  assign dataGroup_lo_lo_636 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_637;
  assign dataGroup_lo_lo_637 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_638;
  assign dataGroup_lo_lo_638 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_639;
  assign dataGroup_lo_lo_639 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_640;
  assign dataGroup_lo_lo_640 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_641;
  assign dataGroup_lo_lo_641 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_642;
  assign dataGroup_lo_lo_642 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_643;
  assign dataGroup_lo_lo_643 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_644;
  assign dataGroup_lo_lo_644 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_645;
  assign dataGroup_lo_lo_645 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_646;
  assign dataGroup_lo_lo_646 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_647;
  assign dataGroup_lo_lo_647 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_648;
  assign dataGroup_lo_lo_648 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_649;
  assign dataGroup_lo_lo_649 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_650;
  assign dataGroup_lo_lo_650 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_651;
  assign dataGroup_lo_lo_651 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_652;
  assign dataGroup_lo_lo_652 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_653;
  assign dataGroup_lo_lo_653 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_654;
  assign dataGroup_lo_lo_654 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_655;
  assign dataGroup_lo_lo_655 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_656;
  assign dataGroup_lo_lo_656 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_657;
  assign dataGroup_lo_lo_657 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_658;
  assign dataGroup_lo_lo_658 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_659;
  assign dataGroup_lo_lo_659 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_660;
  assign dataGroup_lo_lo_660 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_661;
  assign dataGroup_lo_lo_661 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_662;
  assign dataGroup_lo_lo_662 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_663;
  assign dataGroup_lo_lo_663 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_664;
  assign dataGroup_lo_lo_664 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_665;
  assign dataGroup_lo_lo_665 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_666;
  assign dataGroup_lo_lo_666 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_667;
  assign dataGroup_lo_lo_667 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_668;
  assign dataGroup_lo_lo_668 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_669;
  assign dataGroup_lo_lo_669 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_670;
  assign dataGroup_lo_lo_670 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_671;
  assign dataGroup_lo_lo_671 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_672;
  assign dataGroup_lo_lo_672 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_673;
  assign dataGroup_lo_lo_673 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_674;
  assign dataGroup_lo_lo_674 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_675;
  assign dataGroup_lo_lo_675 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_676;
  assign dataGroup_lo_lo_676 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_677;
  assign dataGroup_lo_lo_677 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_678;
  assign dataGroup_lo_lo_678 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_679;
  assign dataGroup_lo_lo_679 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_680;
  assign dataGroup_lo_lo_680 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_681;
  assign dataGroup_lo_lo_681 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_682;
  assign dataGroup_lo_lo_682 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_683;
  assign dataGroup_lo_lo_683 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_684;
  assign dataGroup_lo_lo_684 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_685;
  assign dataGroup_lo_lo_685 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_686;
  assign dataGroup_lo_lo_686 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_687;
  assign dataGroup_lo_lo_687 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_688;
  assign dataGroup_lo_lo_688 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_689;
  assign dataGroup_lo_lo_689 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_690;
  assign dataGroup_lo_lo_690 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_691;
  assign dataGroup_lo_lo_691 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_692;
  assign dataGroup_lo_lo_692 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_693;
  assign dataGroup_lo_lo_693 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_694;
  assign dataGroup_lo_lo_694 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_695;
  assign dataGroup_lo_lo_695 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_696;
  assign dataGroup_lo_lo_696 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_697;
  assign dataGroup_lo_lo_697 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_698;
  assign dataGroup_lo_lo_698 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_699;
  assign dataGroup_lo_lo_699 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_700;
  assign dataGroup_lo_lo_700 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_701;
  assign dataGroup_lo_lo_701 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_702;
  assign dataGroup_lo_lo_702 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_703;
  assign dataGroup_lo_lo_703 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_704;
  assign dataGroup_lo_lo_704 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_705;
  assign dataGroup_lo_lo_705 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_706;
  assign dataGroup_lo_lo_706 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_707;
  assign dataGroup_lo_lo_707 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_708;
  assign dataGroup_lo_lo_708 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_709;
  assign dataGroup_lo_lo_709 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_710;
  assign dataGroup_lo_lo_710 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_711;
  assign dataGroup_lo_lo_711 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_712;
  assign dataGroup_lo_lo_712 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_713;
  assign dataGroup_lo_lo_713 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_714;
  assign dataGroup_lo_lo_714 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_715;
  assign dataGroup_lo_lo_715 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_716;
  assign dataGroup_lo_lo_716 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_717;
  assign dataGroup_lo_lo_717 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_718;
  assign dataGroup_lo_lo_718 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_719;
  assign dataGroup_lo_lo_719 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_720;
  assign dataGroup_lo_lo_720 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_721;
  assign dataGroup_lo_lo_721 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_722;
  assign dataGroup_lo_lo_722 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_723;
  assign dataGroup_lo_lo_723 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_724;
  assign dataGroup_lo_lo_724 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_725;
  assign dataGroup_lo_lo_725 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_726;
  assign dataGroup_lo_lo_726 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_727;
  assign dataGroup_lo_lo_727 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_728;
  assign dataGroup_lo_lo_728 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_729;
  assign dataGroup_lo_lo_729 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_730;
  assign dataGroup_lo_lo_730 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_731;
  assign dataGroup_lo_lo_731 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_732;
  assign dataGroup_lo_lo_732 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_733;
  assign dataGroup_lo_lo_733 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_734;
  assign dataGroup_lo_lo_734 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_735;
  assign dataGroup_lo_lo_735 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_736;
  assign dataGroup_lo_lo_736 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_737;
  assign dataGroup_lo_lo_737 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_738;
  assign dataGroup_lo_lo_738 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_739;
  assign dataGroup_lo_lo_739 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_740;
  assign dataGroup_lo_lo_740 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_741;
  assign dataGroup_lo_lo_741 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_742;
  assign dataGroup_lo_lo_742 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_743;
  assign dataGroup_lo_lo_743 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_744;
  assign dataGroup_lo_lo_744 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_745;
  assign dataGroup_lo_lo_745 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_746;
  assign dataGroup_lo_lo_746 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_747;
  assign dataGroup_lo_lo_747 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_748;
  assign dataGroup_lo_lo_748 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_749;
  assign dataGroup_lo_lo_749 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_750;
  assign dataGroup_lo_lo_750 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_751;
  assign dataGroup_lo_lo_751 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_752;
  assign dataGroup_lo_lo_752 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_753;
  assign dataGroup_lo_lo_753 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_754;
  assign dataGroup_lo_lo_754 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_755;
  assign dataGroup_lo_lo_755 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_756;
  assign dataGroup_lo_lo_756 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_757;
  assign dataGroup_lo_lo_757 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_758;
  assign dataGroup_lo_lo_758 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_759;
  assign dataGroup_lo_lo_759 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_760;
  assign dataGroup_lo_lo_760 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_761;
  assign dataGroup_lo_lo_761 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_762;
  assign dataGroup_lo_lo_762 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_763;
  assign dataGroup_lo_lo_763 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_764;
  assign dataGroup_lo_lo_764 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_765;
  assign dataGroup_lo_lo_765 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_766;
  assign dataGroup_lo_lo_766 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_767;
  assign dataGroup_lo_lo_767 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_768;
  assign dataGroup_lo_lo_768 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_769;
  assign dataGroup_lo_lo_769 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_770;
  assign dataGroup_lo_lo_770 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_771;
  assign dataGroup_lo_lo_771 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_772;
  assign dataGroup_lo_lo_772 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_773;
  assign dataGroup_lo_lo_773 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_774;
  assign dataGroup_lo_lo_774 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_775;
  assign dataGroup_lo_lo_775 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_776;
  assign dataGroup_lo_lo_776 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_777;
  assign dataGroup_lo_lo_777 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_778;
  assign dataGroup_lo_lo_778 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_779;
  assign dataGroup_lo_lo_779 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_780;
  assign dataGroup_lo_lo_780 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_781;
  assign dataGroup_lo_lo_781 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_782;
  assign dataGroup_lo_lo_782 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_783;
  assign dataGroup_lo_lo_783 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_784;
  assign dataGroup_lo_lo_784 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_785;
  assign dataGroup_lo_lo_785 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_786;
  assign dataGroup_lo_lo_786 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_787;
  assign dataGroup_lo_lo_787 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_788;
  assign dataGroup_lo_lo_788 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_789;
  assign dataGroup_lo_lo_789 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_790;
  assign dataGroup_lo_lo_790 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_791;
  assign dataGroup_lo_lo_791 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_792;
  assign dataGroup_lo_lo_792 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_793;
  assign dataGroup_lo_lo_793 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_794;
  assign dataGroup_lo_lo_794 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_795;
  assign dataGroup_lo_lo_795 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_796;
  assign dataGroup_lo_lo_796 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_797;
  assign dataGroup_lo_lo_797 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_798;
  assign dataGroup_lo_lo_798 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_799;
  assign dataGroup_lo_lo_799 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_800;
  assign dataGroup_lo_lo_800 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_801;
  assign dataGroup_lo_lo_801 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_802;
  assign dataGroup_lo_lo_802 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_803;
  assign dataGroup_lo_lo_803 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_804;
  assign dataGroup_lo_lo_804 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_805;
  assign dataGroup_lo_lo_805 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_806;
  assign dataGroup_lo_lo_806 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_807;
  assign dataGroup_lo_lo_807 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_808;
  assign dataGroup_lo_lo_808 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_809;
  assign dataGroup_lo_lo_809 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_810;
  assign dataGroup_lo_lo_810 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_811;
  assign dataGroup_lo_lo_811 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_812;
  assign dataGroup_lo_lo_812 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_813;
  assign dataGroup_lo_lo_813 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_814;
  assign dataGroup_lo_lo_814 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_815;
  assign dataGroup_lo_lo_815 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_816;
  assign dataGroup_lo_lo_816 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_817;
  assign dataGroup_lo_lo_817 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_818;
  assign dataGroup_lo_lo_818 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_819;
  assign dataGroup_lo_lo_819 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_820;
  assign dataGroup_lo_lo_820 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_821;
  assign dataGroup_lo_lo_821 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_822;
  assign dataGroup_lo_lo_822 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_823;
  assign dataGroup_lo_lo_823 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_824;
  assign dataGroup_lo_lo_824 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_825;
  assign dataGroup_lo_lo_825 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_826;
  assign dataGroup_lo_lo_826 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_827;
  assign dataGroup_lo_lo_827 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_828;
  assign dataGroup_lo_lo_828 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_829;
  assign dataGroup_lo_lo_829 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_830;
  assign dataGroup_lo_lo_830 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_831;
  assign dataGroup_lo_lo_831 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_832;
  assign dataGroup_lo_lo_832 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_833;
  assign dataGroup_lo_lo_833 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_834;
  assign dataGroup_lo_lo_834 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_835;
  assign dataGroup_lo_lo_835 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_836;
  assign dataGroup_lo_lo_836 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_837;
  assign dataGroup_lo_lo_837 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_838;
  assign dataGroup_lo_lo_838 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_839;
  assign dataGroup_lo_lo_839 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_840;
  assign dataGroup_lo_lo_840 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_841;
  assign dataGroup_lo_lo_841 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_842;
  assign dataGroup_lo_lo_842 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_843;
  assign dataGroup_lo_lo_843 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_844;
  assign dataGroup_lo_lo_844 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_845;
  assign dataGroup_lo_lo_845 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_846;
  assign dataGroup_lo_lo_846 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_847;
  assign dataGroup_lo_lo_847 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_848;
  assign dataGroup_lo_lo_848 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_849;
  assign dataGroup_lo_lo_849 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_850;
  assign dataGroup_lo_lo_850 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_851;
  assign dataGroup_lo_lo_851 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_852;
  assign dataGroup_lo_lo_852 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_853;
  assign dataGroup_lo_lo_853 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_854;
  assign dataGroup_lo_lo_854 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_855;
  assign dataGroup_lo_lo_855 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_856;
  assign dataGroup_lo_lo_856 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_857;
  assign dataGroup_lo_lo_857 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_858;
  assign dataGroup_lo_lo_858 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_859;
  assign dataGroup_lo_lo_859 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_860;
  assign dataGroup_lo_lo_860 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_861;
  assign dataGroup_lo_lo_861 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_862;
  assign dataGroup_lo_lo_862 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_863;
  assign dataGroup_lo_lo_863 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_864;
  assign dataGroup_lo_lo_864 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_865;
  assign dataGroup_lo_lo_865 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_866;
  assign dataGroup_lo_lo_866 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_867;
  assign dataGroup_lo_lo_867 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_868;
  assign dataGroup_lo_lo_868 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_869;
  assign dataGroup_lo_lo_869 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_870;
  assign dataGroup_lo_lo_870 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_871;
  assign dataGroup_lo_lo_871 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_872;
  assign dataGroup_lo_lo_872 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_873;
  assign dataGroup_lo_lo_873 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_874;
  assign dataGroup_lo_lo_874 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_875;
  assign dataGroup_lo_lo_875 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_876;
  assign dataGroup_lo_lo_876 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_877;
  assign dataGroup_lo_lo_877 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_878;
  assign dataGroup_lo_lo_878 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_879;
  assign dataGroup_lo_lo_879 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_880;
  assign dataGroup_lo_lo_880 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_881;
  assign dataGroup_lo_lo_881 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_882;
  assign dataGroup_lo_lo_882 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_883;
  assign dataGroup_lo_lo_883 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_884;
  assign dataGroup_lo_lo_884 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_885;
  assign dataGroup_lo_lo_885 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_886;
  assign dataGroup_lo_lo_886 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_887;
  assign dataGroup_lo_lo_887 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_888;
  assign dataGroup_lo_lo_888 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_889;
  assign dataGroup_lo_lo_889 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_890;
  assign dataGroup_lo_lo_890 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_891;
  assign dataGroup_lo_lo_891 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_892;
  assign dataGroup_lo_lo_892 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_893;
  assign dataGroup_lo_lo_893 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_894;
  assign dataGroup_lo_lo_894 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_895;
  assign dataGroup_lo_lo_895 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_896;
  assign dataGroup_lo_lo_896 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_897;
  assign dataGroup_lo_lo_897 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_898;
  assign dataGroup_lo_lo_898 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_899;
  assign dataGroup_lo_lo_899 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_900;
  assign dataGroup_lo_lo_900 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_901;
  assign dataGroup_lo_lo_901 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_902;
  assign dataGroup_lo_lo_902 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_903;
  assign dataGroup_lo_lo_903 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_904;
  assign dataGroup_lo_lo_904 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_905;
  assign dataGroup_lo_lo_905 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_906;
  assign dataGroup_lo_lo_906 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_907;
  assign dataGroup_lo_lo_907 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_908;
  assign dataGroup_lo_lo_908 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_909;
  assign dataGroup_lo_lo_909 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_910;
  assign dataGroup_lo_lo_910 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_911;
  assign dataGroup_lo_lo_911 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_912;
  assign dataGroup_lo_lo_912 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_913;
  assign dataGroup_lo_lo_913 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_914;
  assign dataGroup_lo_lo_914 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_915;
  assign dataGroup_lo_lo_915 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_916;
  assign dataGroup_lo_lo_916 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_917;
  assign dataGroup_lo_lo_917 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_918;
  assign dataGroup_lo_lo_918 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_919;
  assign dataGroup_lo_lo_919 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_920;
  assign dataGroup_lo_lo_920 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_921;
  assign dataGroup_lo_lo_921 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_922;
  assign dataGroup_lo_lo_922 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_923;
  assign dataGroup_lo_lo_923 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_924;
  assign dataGroup_lo_lo_924 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_925;
  assign dataGroup_lo_lo_925 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_926;
  assign dataGroup_lo_lo_926 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_927;
  assign dataGroup_lo_lo_927 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_928;
  assign dataGroup_lo_lo_928 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_929;
  assign dataGroup_lo_lo_929 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_930;
  assign dataGroup_lo_lo_930 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_931;
  assign dataGroup_lo_lo_931 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_932;
  assign dataGroup_lo_lo_932 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_933;
  assign dataGroup_lo_lo_933 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_934;
  assign dataGroup_lo_lo_934 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_935;
  assign dataGroup_lo_lo_935 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_936;
  assign dataGroup_lo_lo_936 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_937;
  assign dataGroup_lo_lo_937 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_938;
  assign dataGroup_lo_lo_938 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_939;
  assign dataGroup_lo_lo_939 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_940;
  assign dataGroup_lo_lo_940 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_941;
  assign dataGroup_lo_lo_941 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_942;
  assign dataGroup_lo_lo_942 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_943;
  assign dataGroup_lo_lo_943 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_944;
  assign dataGroup_lo_lo_944 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_945;
  assign dataGroup_lo_lo_945 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_946;
  assign dataGroup_lo_lo_946 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_947;
  assign dataGroup_lo_lo_947 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_948;
  assign dataGroup_lo_lo_948 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_949;
  assign dataGroup_lo_lo_949 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_950;
  assign dataGroup_lo_lo_950 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_951;
  assign dataGroup_lo_lo_951 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_952;
  assign dataGroup_lo_lo_952 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_953;
  assign dataGroup_lo_lo_953 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_954;
  assign dataGroup_lo_lo_954 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_955;
  assign dataGroup_lo_lo_955 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_956;
  assign dataGroup_lo_lo_956 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_957;
  assign dataGroup_lo_lo_957 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_958;
  assign dataGroup_lo_lo_958 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_959;
  assign dataGroup_lo_lo_959 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_960;
  assign dataGroup_lo_lo_960 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_961;
  assign dataGroup_lo_lo_961 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_962;
  assign dataGroup_lo_lo_962 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_963;
  assign dataGroup_lo_lo_963 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_964;
  assign dataGroup_lo_lo_964 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_965;
  assign dataGroup_lo_lo_965 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_966;
  assign dataGroup_lo_lo_966 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_967;
  assign dataGroup_lo_lo_967 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_968;
  assign dataGroup_lo_lo_968 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_969;
  assign dataGroup_lo_lo_969 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_970;
  assign dataGroup_lo_lo_970 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_971;
  assign dataGroup_lo_lo_971 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_972;
  assign dataGroup_lo_lo_972 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_973;
  assign dataGroup_lo_lo_973 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_974;
  assign dataGroup_lo_lo_974 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_975;
  assign dataGroup_lo_lo_975 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_976;
  assign dataGroup_lo_lo_976 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_977;
  assign dataGroup_lo_lo_977 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_978;
  assign dataGroup_lo_lo_978 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_979;
  assign dataGroup_lo_lo_979 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_980;
  assign dataGroup_lo_lo_980 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_981;
  assign dataGroup_lo_lo_981 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_982;
  assign dataGroup_lo_lo_982 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_983;
  assign dataGroup_lo_lo_983 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_984;
  assign dataGroup_lo_lo_984 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_985;
  assign dataGroup_lo_lo_985 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_986;
  assign dataGroup_lo_lo_986 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_987;
  assign dataGroup_lo_lo_987 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_988;
  assign dataGroup_lo_lo_988 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_989;
  assign dataGroup_lo_lo_989 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_990;
  assign dataGroup_lo_lo_990 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_991;
  assign dataGroup_lo_lo_991 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_992;
  assign dataGroup_lo_lo_992 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_993;
  assign dataGroup_lo_lo_993 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_994;
  assign dataGroup_lo_lo_994 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_995;
  assign dataGroup_lo_lo_995 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_996;
  assign dataGroup_lo_lo_996 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_997;
  assign dataGroup_lo_lo_997 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_998;
  assign dataGroup_lo_lo_998 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_999;
  assign dataGroup_lo_lo_999 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1000;
  assign dataGroup_lo_lo_1000 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1001;
  assign dataGroup_lo_lo_1001 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1002;
  assign dataGroup_lo_lo_1002 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1003;
  assign dataGroup_lo_lo_1003 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1004;
  assign dataGroup_lo_lo_1004 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1005;
  assign dataGroup_lo_lo_1005 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1006;
  assign dataGroup_lo_lo_1006 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1007;
  assign dataGroup_lo_lo_1007 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1008;
  assign dataGroup_lo_lo_1008 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1009;
  assign dataGroup_lo_lo_1009 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1010;
  assign dataGroup_lo_lo_1010 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1011;
  assign dataGroup_lo_lo_1011 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1012;
  assign dataGroup_lo_lo_1012 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1013;
  assign dataGroup_lo_lo_1013 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1014;
  assign dataGroup_lo_lo_1014 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1015;
  assign dataGroup_lo_lo_1015 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1016;
  assign dataGroup_lo_lo_1016 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1017;
  assign dataGroup_lo_lo_1017 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1018;
  assign dataGroup_lo_lo_1018 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1019;
  assign dataGroup_lo_lo_1019 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1020;
  assign dataGroup_lo_lo_1020 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1021;
  assign dataGroup_lo_lo_1021 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1022;
  assign dataGroup_lo_lo_1022 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1023;
  assign dataGroup_lo_lo_1023 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1024;
  assign dataGroup_lo_lo_1024 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1025;
  assign dataGroup_lo_lo_1025 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1026;
  assign dataGroup_lo_lo_1026 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1027;
  assign dataGroup_lo_lo_1027 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1028;
  assign dataGroup_lo_lo_1028 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1029;
  assign dataGroup_lo_lo_1029 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1030;
  assign dataGroup_lo_lo_1030 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1031;
  assign dataGroup_lo_lo_1031 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1032;
  assign dataGroup_lo_lo_1032 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1033;
  assign dataGroup_lo_lo_1033 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1034;
  assign dataGroup_lo_lo_1034 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1035;
  assign dataGroup_lo_lo_1035 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1036;
  assign dataGroup_lo_lo_1036 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1037;
  assign dataGroup_lo_lo_1037 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1038;
  assign dataGroup_lo_lo_1038 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1039;
  assign dataGroup_lo_lo_1039 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1040;
  assign dataGroup_lo_lo_1040 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1041;
  assign dataGroup_lo_lo_1041 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1042;
  assign dataGroup_lo_lo_1042 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1043;
  assign dataGroup_lo_lo_1043 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1044;
  assign dataGroup_lo_lo_1044 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1045;
  assign dataGroup_lo_lo_1045 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1046;
  assign dataGroup_lo_lo_1046 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1047;
  assign dataGroup_lo_lo_1047 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1048;
  assign dataGroup_lo_lo_1048 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1049;
  assign dataGroup_lo_lo_1049 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1050;
  assign dataGroup_lo_lo_1050 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1051;
  assign dataGroup_lo_lo_1051 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1052;
  assign dataGroup_lo_lo_1052 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1053;
  assign dataGroup_lo_lo_1053 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1054;
  assign dataGroup_lo_lo_1054 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1055;
  assign dataGroup_lo_lo_1055 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1056;
  assign dataGroup_lo_lo_1056 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1057;
  assign dataGroup_lo_lo_1057 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1058;
  assign dataGroup_lo_lo_1058 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1059;
  assign dataGroup_lo_lo_1059 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1060;
  assign dataGroup_lo_lo_1060 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1061;
  assign dataGroup_lo_lo_1061 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1062;
  assign dataGroup_lo_lo_1062 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1063;
  assign dataGroup_lo_lo_1063 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1064;
  assign dataGroup_lo_lo_1064 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1065;
  assign dataGroup_lo_lo_1065 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1066;
  assign dataGroup_lo_lo_1066 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1067;
  assign dataGroup_lo_lo_1067 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1068;
  assign dataGroup_lo_lo_1068 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1069;
  assign dataGroup_lo_lo_1069 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1070;
  assign dataGroup_lo_lo_1070 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1071;
  assign dataGroup_lo_lo_1071 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1072;
  assign dataGroup_lo_lo_1072 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1073;
  assign dataGroup_lo_lo_1073 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1074;
  assign dataGroup_lo_lo_1074 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1075;
  assign dataGroup_lo_lo_1075 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1076;
  assign dataGroup_lo_lo_1076 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1077;
  assign dataGroup_lo_lo_1077 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1078;
  assign dataGroup_lo_lo_1078 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1079;
  assign dataGroup_lo_lo_1079 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1080;
  assign dataGroup_lo_lo_1080 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1081;
  assign dataGroup_lo_lo_1081 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1082;
  assign dataGroup_lo_lo_1082 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1083;
  assign dataGroup_lo_lo_1083 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1084;
  assign dataGroup_lo_lo_1084 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1085;
  assign dataGroup_lo_lo_1085 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1086;
  assign dataGroup_lo_lo_1086 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1087;
  assign dataGroup_lo_lo_1087 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1088;
  assign dataGroup_lo_lo_1088 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1089;
  assign dataGroup_lo_lo_1089 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1090;
  assign dataGroup_lo_lo_1090 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1091;
  assign dataGroup_lo_lo_1091 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1092;
  assign dataGroup_lo_lo_1092 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1093;
  assign dataGroup_lo_lo_1093 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1094;
  assign dataGroup_lo_lo_1094 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1095;
  assign dataGroup_lo_lo_1095 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1096;
  assign dataGroup_lo_lo_1096 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1097;
  assign dataGroup_lo_lo_1097 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1098;
  assign dataGroup_lo_lo_1098 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1099;
  assign dataGroup_lo_lo_1099 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1100;
  assign dataGroup_lo_lo_1100 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1101;
  assign dataGroup_lo_lo_1101 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1102;
  assign dataGroup_lo_lo_1102 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1103;
  assign dataGroup_lo_lo_1103 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1104;
  assign dataGroup_lo_lo_1104 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1105;
  assign dataGroup_lo_lo_1105 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1106;
  assign dataGroup_lo_lo_1106 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1107;
  assign dataGroup_lo_lo_1107 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1108;
  assign dataGroup_lo_lo_1108 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1109;
  assign dataGroup_lo_lo_1109 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1110;
  assign dataGroup_lo_lo_1110 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1111;
  assign dataGroup_lo_lo_1111 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1112;
  assign dataGroup_lo_lo_1112 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1113;
  assign dataGroup_lo_lo_1113 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1114;
  assign dataGroup_lo_lo_1114 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1115;
  assign dataGroup_lo_lo_1115 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1116;
  assign dataGroup_lo_lo_1116 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1117;
  assign dataGroup_lo_lo_1117 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1118;
  assign dataGroup_lo_lo_1118 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1119;
  assign dataGroup_lo_lo_1119 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1120;
  assign dataGroup_lo_lo_1120 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1121;
  assign dataGroup_lo_lo_1121 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1122;
  assign dataGroup_lo_lo_1122 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1123;
  assign dataGroup_lo_lo_1123 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1124;
  assign dataGroup_lo_lo_1124 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1125;
  assign dataGroup_lo_lo_1125 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1126;
  assign dataGroup_lo_lo_1126 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1127;
  assign dataGroup_lo_lo_1127 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1128;
  assign dataGroup_lo_lo_1128 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1129;
  assign dataGroup_lo_lo_1129 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1130;
  assign dataGroup_lo_lo_1130 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1131;
  assign dataGroup_lo_lo_1131 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1132;
  assign dataGroup_lo_lo_1132 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1133;
  assign dataGroup_lo_lo_1133 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1134;
  assign dataGroup_lo_lo_1134 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1135;
  assign dataGroup_lo_lo_1135 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1136;
  assign dataGroup_lo_lo_1136 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1137;
  assign dataGroup_lo_lo_1137 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1138;
  assign dataGroup_lo_lo_1138 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1139;
  assign dataGroup_lo_lo_1139 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1140;
  assign dataGroup_lo_lo_1140 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1141;
  assign dataGroup_lo_lo_1141 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1142;
  assign dataGroup_lo_lo_1142 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1143;
  assign dataGroup_lo_lo_1143 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1144;
  assign dataGroup_lo_lo_1144 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1145;
  assign dataGroup_lo_lo_1145 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1146;
  assign dataGroup_lo_lo_1146 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1147;
  assign dataGroup_lo_lo_1147 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1148;
  assign dataGroup_lo_lo_1148 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1149;
  assign dataGroup_lo_lo_1149 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1150;
  assign dataGroup_lo_lo_1150 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1151;
  assign dataGroup_lo_lo_1151 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1152;
  assign dataGroup_lo_lo_1152 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1153;
  assign dataGroup_lo_lo_1153 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1154;
  assign dataGroup_lo_lo_1154 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1155;
  assign dataGroup_lo_lo_1155 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1156;
  assign dataGroup_lo_lo_1156 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1157;
  assign dataGroup_lo_lo_1157 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1158;
  assign dataGroup_lo_lo_1158 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1159;
  assign dataGroup_lo_lo_1159 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1160;
  assign dataGroup_lo_lo_1160 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1161;
  assign dataGroup_lo_lo_1161 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1162;
  assign dataGroup_lo_lo_1162 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1163;
  assign dataGroup_lo_lo_1163 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1164;
  assign dataGroup_lo_lo_1164 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1165;
  assign dataGroup_lo_lo_1165 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1166;
  assign dataGroup_lo_lo_1166 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1167;
  assign dataGroup_lo_lo_1167 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1168;
  assign dataGroup_lo_lo_1168 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1169;
  assign dataGroup_lo_lo_1169 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1170;
  assign dataGroup_lo_lo_1170 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1171;
  assign dataGroup_lo_lo_1171 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1172;
  assign dataGroup_lo_lo_1172 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1173;
  assign dataGroup_lo_lo_1173 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1174;
  assign dataGroup_lo_lo_1174 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1175;
  assign dataGroup_lo_lo_1175 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1176;
  assign dataGroup_lo_lo_1176 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1177;
  assign dataGroup_lo_lo_1177 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1178;
  assign dataGroup_lo_lo_1178 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1179;
  assign dataGroup_lo_lo_1179 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1180;
  assign dataGroup_lo_lo_1180 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1181;
  assign dataGroup_lo_lo_1181 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1182;
  assign dataGroup_lo_lo_1182 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1183;
  assign dataGroup_lo_lo_1183 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1184;
  assign dataGroup_lo_lo_1184 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1185;
  assign dataGroup_lo_lo_1185 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1186;
  assign dataGroup_lo_lo_1186 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1187;
  assign dataGroup_lo_lo_1187 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1188;
  assign dataGroup_lo_lo_1188 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1189;
  assign dataGroup_lo_lo_1189 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1190;
  assign dataGroup_lo_lo_1190 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1191;
  assign dataGroup_lo_lo_1191 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1192;
  assign dataGroup_lo_lo_1192 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1193;
  assign dataGroup_lo_lo_1193 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1194;
  assign dataGroup_lo_lo_1194 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1195;
  assign dataGroup_lo_lo_1195 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1196;
  assign dataGroup_lo_lo_1196 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1197;
  assign dataGroup_lo_lo_1197 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1198;
  assign dataGroup_lo_lo_1198 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1199;
  assign dataGroup_lo_lo_1199 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1200;
  assign dataGroup_lo_lo_1200 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1201;
  assign dataGroup_lo_lo_1201 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1202;
  assign dataGroup_lo_lo_1202 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1203;
  assign dataGroup_lo_lo_1203 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1204;
  assign dataGroup_lo_lo_1204 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1205;
  assign dataGroup_lo_lo_1205 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1206;
  assign dataGroup_lo_lo_1206 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1207;
  assign dataGroup_lo_lo_1207 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1208;
  assign dataGroup_lo_lo_1208 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1209;
  assign dataGroup_lo_lo_1209 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1210;
  assign dataGroup_lo_lo_1210 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1211;
  assign dataGroup_lo_lo_1211 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1212;
  assign dataGroup_lo_lo_1212 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1213;
  assign dataGroup_lo_lo_1213 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1214;
  assign dataGroup_lo_lo_1214 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1215;
  assign dataGroup_lo_lo_1215 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1216;
  assign dataGroup_lo_lo_1216 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1217;
  assign dataGroup_lo_lo_1217 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1218;
  assign dataGroup_lo_lo_1218 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1219;
  assign dataGroup_lo_lo_1219 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1220;
  assign dataGroup_lo_lo_1220 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1221;
  assign dataGroup_lo_lo_1221 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1222;
  assign dataGroup_lo_lo_1222 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1223;
  assign dataGroup_lo_lo_1223 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1224;
  assign dataGroup_lo_lo_1224 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1225;
  assign dataGroup_lo_lo_1225 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1226;
  assign dataGroup_lo_lo_1226 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1227;
  assign dataGroup_lo_lo_1227 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1228;
  assign dataGroup_lo_lo_1228 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1229;
  assign dataGroup_lo_lo_1229 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1230;
  assign dataGroup_lo_lo_1230 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1231;
  assign dataGroup_lo_lo_1231 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1232;
  assign dataGroup_lo_lo_1232 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1233;
  assign dataGroup_lo_lo_1233 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1234;
  assign dataGroup_lo_lo_1234 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1235;
  assign dataGroup_lo_lo_1235 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1236;
  assign dataGroup_lo_lo_1236 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1237;
  assign dataGroup_lo_lo_1237 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1238;
  assign dataGroup_lo_lo_1238 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1239;
  assign dataGroup_lo_lo_1239 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1240;
  assign dataGroup_lo_lo_1240 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1241;
  assign dataGroup_lo_lo_1241 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1242;
  assign dataGroup_lo_lo_1242 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1243;
  assign dataGroup_lo_lo_1243 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1244;
  assign dataGroup_lo_lo_1244 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1245;
  assign dataGroup_lo_lo_1245 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1246;
  assign dataGroup_lo_lo_1246 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1247;
  assign dataGroup_lo_lo_1247 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1248;
  assign dataGroup_lo_lo_1248 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1249;
  assign dataGroup_lo_lo_1249 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1250;
  assign dataGroup_lo_lo_1250 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1251;
  assign dataGroup_lo_lo_1251 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1252;
  assign dataGroup_lo_lo_1252 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1253;
  assign dataGroup_lo_lo_1253 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1254;
  assign dataGroup_lo_lo_1254 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1255;
  assign dataGroup_lo_lo_1255 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1256;
  assign dataGroup_lo_lo_1256 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1257;
  assign dataGroup_lo_lo_1257 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1258;
  assign dataGroup_lo_lo_1258 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1259;
  assign dataGroup_lo_lo_1259 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1260;
  assign dataGroup_lo_lo_1260 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1261;
  assign dataGroup_lo_lo_1261 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1262;
  assign dataGroup_lo_lo_1262 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1263;
  assign dataGroup_lo_lo_1263 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1264;
  assign dataGroup_lo_lo_1264 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1265;
  assign dataGroup_lo_lo_1265 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1266;
  assign dataGroup_lo_lo_1266 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1267;
  assign dataGroup_lo_lo_1267 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1268;
  assign dataGroup_lo_lo_1268 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1269;
  assign dataGroup_lo_lo_1269 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1270;
  assign dataGroup_lo_lo_1270 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1271;
  assign dataGroup_lo_lo_1271 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1272;
  assign dataGroup_lo_lo_1272 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1273;
  assign dataGroup_lo_lo_1273 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1274;
  assign dataGroup_lo_lo_1274 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1275;
  assign dataGroup_lo_lo_1275 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1276;
  assign dataGroup_lo_lo_1276 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1277;
  assign dataGroup_lo_lo_1277 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1278;
  assign dataGroup_lo_lo_1278 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1279;
  assign dataGroup_lo_lo_1279 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1280;
  assign dataGroup_lo_lo_1280 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1281;
  assign dataGroup_lo_lo_1281 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1282;
  assign dataGroup_lo_lo_1282 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1283;
  assign dataGroup_lo_lo_1283 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1284;
  assign dataGroup_lo_lo_1284 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1285;
  assign dataGroup_lo_lo_1285 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1286;
  assign dataGroup_lo_lo_1286 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1287;
  assign dataGroup_lo_lo_1287 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1288;
  assign dataGroup_lo_lo_1288 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1289;
  assign dataGroup_lo_lo_1289 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1290;
  assign dataGroup_lo_lo_1290 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1291;
  assign dataGroup_lo_lo_1291 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1292;
  assign dataGroup_lo_lo_1292 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1293;
  assign dataGroup_lo_lo_1293 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1294;
  assign dataGroup_lo_lo_1294 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1295;
  assign dataGroup_lo_lo_1295 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1296;
  assign dataGroup_lo_lo_1296 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1297;
  assign dataGroup_lo_lo_1297 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1298;
  assign dataGroup_lo_lo_1298 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1299;
  assign dataGroup_lo_lo_1299 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1300;
  assign dataGroup_lo_lo_1300 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1301;
  assign dataGroup_lo_lo_1301 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1302;
  assign dataGroup_lo_lo_1302 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1303;
  assign dataGroup_lo_lo_1303 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1304;
  assign dataGroup_lo_lo_1304 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1305;
  assign dataGroup_lo_lo_1305 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1306;
  assign dataGroup_lo_lo_1306 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1307;
  assign dataGroup_lo_lo_1307 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1308;
  assign dataGroup_lo_lo_1308 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1309;
  assign dataGroup_lo_lo_1309 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1310;
  assign dataGroup_lo_lo_1310 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1311;
  assign dataGroup_lo_lo_1311 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1312;
  assign dataGroup_lo_lo_1312 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1313;
  assign dataGroup_lo_lo_1313 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1314;
  assign dataGroup_lo_lo_1314 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1315;
  assign dataGroup_lo_lo_1315 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1316;
  assign dataGroup_lo_lo_1316 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1317;
  assign dataGroup_lo_lo_1317 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1318;
  assign dataGroup_lo_lo_1318 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1319;
  assign dataGroup_lo_lo_1319 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1320;
  assign dataGroup_lo_lo_1320 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1321;
  assign dataGroup_lo_lo_1321 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1322;
  assign dataGroup_lo_lo_1322 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1323;
  assign dataGroup_lo_lo_1323 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1324;
  assign dataGroup_lo_lo_1324 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1325;
  assign dataGroup_lo_lo_1325 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1326;
  assign dataGroup_lo_lo_1326 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1327;
  assign dataGroup_lo_lo_1327 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1328;
  assign dataGroup_lo_lo_1328 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1329;
  assign dataGroup_lo_lo_1329 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1330;
  assign dataGroup_lo_lo_1330 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1331;
  assign dataGroup_lo_lo_1331 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1332;
  assign dataGroup_lo_lo_1332 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1333;
  assign dataGroup_lo_lo_1333 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1334;
  assign dataGroup_lo_lo_1334 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1335;
  assign dataGroup_lo_lo_1335 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1336;
  assign dataGroup_lo_lo_1336 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1337;
  assign dataGroup_lo_lo_1337 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1338;
  assign dataGroup_lo_lo_1338 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1339;
  assign dataGroup_lo_lo_1339 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1340;
  assign dataGroup_lo_lo_1340 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1341;
  assign dataGroup_lo_lo_1341 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1342;
  assign dataGroup_lo_lo_1342 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1343;
  assign dataGroup_lo_lo_1343 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1344;
  assign dataGroup_lo_lo_1344 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1345;
  assign dataGroup_lo_lo_1345 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1346;
  assign dataGroup_lo_lo_1346 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1347;
  assign dataGroup_lo_lo_1347 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1348;
  assign dataGroup_lo_lo_1348 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1349;
  assign dataGroup_lo_lo_1349 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1350;
  assign dataGroup_lo_lo_1350 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1351;
  assign dataGroup_lo_lo_1351 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1352;
  assign dataGroup_lo_lo_1352 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1353;
  assign dataGroup_lo_lo_1353 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1354;
  assign dataGroup_lo_lo_1354 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1355;
  assign dataGroup_lo_lo_1355 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1356;
  assign dataGroup_lo_lo_1356 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1357;
  assign dataGroup_lo_lo_1357 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1358;
  assign dataGroup_lo_lo_1358 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1359;
  assign dataGroup_lo_lo_1359 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1360;
  assign dataGroup_lo_lo_1360 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1361;
  assign dataGroup_lo_lo_1361 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1362;
  assign dataGroup_lo_lo_1362 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1363;
  assign dataGroup_lo_lo_1363 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1364;
  assign dataGroup_lo_lo_1364 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1365;
  assign dataGroup_lo_lo_1365 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1366;
  assign dataGroup_lo_lo_1366 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1367;
  assign dataGroup_lo_lo_1367 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1368;
  assign dataGroup_lo_lo_1368 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1369;
  assign dataGroup_lo_lo_1369 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1370;
  assign dataGroup_lo_lo_1370 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1371;
  assign dataGroup_lo_lo_1371 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1372;
  assign dataGroup_lo_lo_1372 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1373;
  assign dataGroup_lo_lo_1373 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1374;
  assign dataGroup_lo_lo_1374 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1375;
  assign dataGroup_lo_lo_1375 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1376;
  assign dataGroup_lo_lo_1376 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1377;
  assign dataGroup_lo_lo_1377 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1378;
  assign dataGroup_lo_lo_1378 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1379;
  assign dataGroup_lo_lo_1379 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1380;
  assign dataGroup_lo_lo_1380 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1381;
  assign dataGroup_lo_lo_1381 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1382;
  assign dataGroup_lo_lo_1382 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1383;
  assign dataGroup_lo_lo_1383 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1384;
  assign dataGroup_lo_lo_1384 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1385;
  assign dataGroup_lo_lo_1385 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1386;
  assign dataGroup_lo_lo_1386 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1387;
  assign dataGroup_lo_lo_1387 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1388;
  assign dataGroup_lo_lo_1388 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1389;
  assign dataGroup_lo_lo_1389 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1390;
  assign dataGroup_lo_lo_1390 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1391;
  assign dataGroup_lo_lo_1391 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1392;
  assign dataGroup_lo_lo_1392 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1393;
  assign dataGroup_lo_lo_1393 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1394;
  assign dataGroup_lo_lo_1394 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1395;
  assign dataGroup_lo_lo_1395 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1396;
  assign dataGroup_lo_lo_1396 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1397;
  assign dataGroup_lo_lo_1397 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1398;
  assign dataGroup_lo_lo_1398 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1399;
  assign dataGroup_lo_lo_1399 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1400;
  assign dataGroup_lo_lo_1400 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1401;
  assign dataGroup_lo_lo_1401 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1402;
  assign dataGroup_lo_lo_1402 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1403;
  assign dataGroup_lo_lo_1403 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1404;
  assign dataGroup_lo_lo_1404 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1405;
  assign dataGroup_lo_lo_1405 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1406;
  assign dataGroup_lo_lo_1406 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1407;
  assign dataGroup_lo_lo_1407 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1408;
  assign dataGroup_lo_lo_1408 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1409;
  assign dataGroup_lo_lo_1409 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1410;
  assign dataGroup_lo_lo_1410 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1411;
  assign dataGroup_lo_lo_1411 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1412;
  assign dataGroup_lo_lo_1412 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1413;
  assign dataGroup_lo_lo_1413 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1414;
  assign dataGroup_lo_lo_1414 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1415;
  assign dataGroup_lo_lo_1415 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1416;
  assign dataGroup_lo_lo_1416 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1417;
  assign dataGroup_lo_lo_1417 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1418;
  assign dataGroup_lo_lo_1418 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1419;
  assign dataGroup_lo_lo_1419 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1420;
  assign dataGroup_lo_lo_1420 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1421;
  assign dataGroup_lo_lo_1421 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1422;
  assign dataGroup_lo_lo_1422 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1423;
  assign dataGroup_lo_lo_1423 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1424;
  assign dataGroup_lo_lo_1424 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1425;
  assign dataGroup_lo_lo_1425 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1426;
  assign dataGroup_lo_lo_1426 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1427;
  assign dataGroup_lo_lo_1427 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1428;
  assign dataGroup_lo_lo_1428 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1429;
  assign dataGroup_lo_lo_1429 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1430;
  assign dataGroup_lo_lo_1430 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1431;
  assign dataGroup_lo_lo_1431 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1432;
  assign dataGroup_lo_lo_1432 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1433;
  assign dataGroup_lo_lo_1433 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1434;
  assign dataGroup_lo_lo_1434 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1435;
  assign dataGroup_lo_lo_1435 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1436;
  assign dataGroup_lo_lo_1436 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1437;
  assign dataGroup_lo_lo_1437 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1438;
  assign dataGroup_lo_lo_1438 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1439;
  assign dataGroup_lo_lo_1439 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1440;
  assign dataGroup_lo_lo_1440 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1441;
  assign dataGroup_lo_lo_1441 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1442;
  assign dataGroup_lo_lo_1442 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1443;
  assign dataGroup_lo_lo_1443 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1444;
  assign dataGroup_lo_lo_1444 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1445;
  assign dataGroup_lo_lo_1445 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1446;
  assign dataGroup_lo_lo_1446 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1447;
  assign dataGroup_lo_lo_1447 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1448;
  assign dataGroup_lo_lo_1448 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1449;
  assign dataGroup_lo_lo_1449 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1450;
  assign dataGroup_lo_lo_1450 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1451;
  assign dataGroup_lo_lo_1451 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1452;
  assign dataGroup_lo_lo_1452 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1453;
  assign dataGroup_lo_lo_1453 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1454;
  assign dataGroup_lo_lo_1454 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1455;
  assign dataGroup_lo_lo_1455 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1456;
  assign dataGroup_lo_lo_1456 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1457;
  assign dataGroup_lo_lo_1457 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1458;
  assign dataGroup_lo_lo_1458 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1459;
  assign dataGroup_lo_lo_1459 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1460;
  assign dataGroup_lo_lo_1460 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1461;
  assign dataGroup_lo_lo_1461 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1462;
  assign dataGroup_lo_lo_1462 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1463;
  assign dataGroup_lo_lo_1463 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1464;
  assign dataGroup_lo_lo_1464 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1465;
  assign dataGroup_lo_lo_1465 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1466;
  assign dataGroup_lo_lo_1466 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1467;
  assign dataGroup_lo_lo_1467 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1468;
  assign dataGroup_lo_lo_1468 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1469;
  assign dataGroup_lo_lo_1469 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1470;
  assign dataGroup_lo_lo_1470 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1471;
  assign dataGroup_lo_lo_1471 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1472;
  assign dataGroup_lo_lo_1472 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1473;
  assign dataGroup_lo_lo_1473 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1474;
  assign dataGroup_lo_lo_1474 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1475;
  assign dataGroup_lo_lo_1475 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1476;
  assign dataGroup_lo_lo_1476 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1477;
  assign dataGroup_lo_lo_1477 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1478;
  assign dataGroup_lo_lo_1478 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1479;
  assign dataGroup_lo_lo_1479 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1480;
  assign dataGroup_lo_lo_1480 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1481;
  assign dataGroup_lo_lo_1481 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1482;
  assign dataGroup_lo_lo_1482 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1483;
  assign dataGroup_lo_lo_1483 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1484;
  assign dataGroup_lo_lo_1484 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1485;
  assign dataGroup_lo_lo_1485 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1486;
  assign dataGroup_lo_lo_1486 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1487;
  assign dataGroup_lo_lo_1487 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1488;
  assign dataGroup_lo_lo_1488 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1489;
  assign dataGroup_lo_lo_1489 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1490;
  assign dataGroup_lo_lo_1490 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1491;
  assign dataGroup_lo_lo_1491 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1492;
  assign dataGroup_lo_lo_1492 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1493;
  assign dataGroup_lo_lo_1493 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1494;
  assign dataGroup_lo_lo_1494 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1495;
  assign dataGroup_lo_lo_1495 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1496;
  assign dataGroup_lo_lo_1496 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1497;
  assign dataGroup_lo_lo_1497 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1498;
  assign dataGroup_lo_lo_1498 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1499;
  assign dataGroup_lo_lo_1499 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1500;
  assign dataGroup_lo_lo_1500 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1501;
  assign dataGroup_lo_lo_1501 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1502;
  assign dataGroup_lo_lo_1502 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1503;
  assign dataGroup_lo_lo_1503 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1504;
  assign dataGroup_lo_lo_1504 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1505;
  assign dataGroup_lo_lo_1505 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1506;
  assign dataGroup_lo_lo_1506 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1507;
  assign dataGroup_lo_lo_1507 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1508;
  assign dataGroup_lo_lo_1508 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1509;
  assign dataGroup_lo_lo_1509 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1510;
  assign dataGroup_lo_lo_1510 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1511;
  assign dataGroup_lo_lo_1511 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1512;
  assign dataGroup_lo_lo_1512 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1513;
  assign dataGroup_lo_lo_1513 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1514;
  assign dataGroup_lo_lo_1514 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1515;
  assign dataGroup_lo_lo_1515 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1516;
  assign dataGroup_lo_lo_1516 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1517;
  assign dataGroup_lo_lo_1517 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1518;
  assign dataGroup_lo_lo_1518 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1519;
  assign dataGroup_lo_lo_1519 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1520;
  assign dataGroup_lo_lo_1520 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1521;
  assign dataGroup_lo_lo_1521 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1522;
  assign dataGroup_lo_lo_1522 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1523;
  assign dataGroup_lo_lo_1523 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1524;
  assign dataGroup_lo_lo_1524 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1525;
  assign dataGroup_lo_lo_1525 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1526;
  assign dataGroup_lo_lo_1526 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1527;
  assign dataGroup_lo_lo_1527 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1528;
  assign dataGroup_lo_lo_1528 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1529;
  assign dataGroup_lo_lo_1529 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1530;
  assign dataGroup_lo_lo_1530 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1531;
  assign dataGroup_lo_lo_1531 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1532;
  assign dataGroup_lo_lo_1532 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1533;
  assign dataGroup_lo_lo_1533 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1534;
  assign dataGroup_lo_lo_1534 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1535;
  assign dataGroup_lo_lo_1535 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1536;
  assign dataGroup_lo_lo_1536 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1537;
  assign dataGroup_lo_lo_1537 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1538;
  assign dataGroup_lo_lo_1538 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1539;
  assign dataGroup_lo_lo_1539 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1540;
  assign dataGroup_lo_lo_1540 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1541;
  assign dataGroup_lo_lo_1541 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1542;
  assign dataGroup_lo_lo_1542 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1543;
  assign dataGroup_lo_lo_1543 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1544;
  assign dataGroup_lo_lo_1544 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1545;
  assign dataGroup_lo_lo_1545 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1546;
  assign dataGroup_lo_lo_1546 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1547;
  assign dataGroup_lo_lo_1547 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1548;
  assign dataGroup_lo_lo_1548 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1549;
  assign dataGroup_lo_lo_1549 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1550;
  assign dataGroup_lo_lo_1550 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1551;
  assign dataGroup_lo_lo_1551 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1552;
  assign dataGroup_lo_lo_1552 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1553;
  assign dataGroup_lo_lo_1553 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1554;
  assign dataGroup_lo_lo_1554 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1555;
  assign dataGroup_lo_lo_1555 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1556;
  assign dataGroup_lo_lo_1556 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1557;
  assign dataGroup_lo_lo_1557 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1558;
  assign dataGroup_lo_lo_1558 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1559;
  assign dataGroup_lo_lo_1559 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1560;
  assign dataGroup_lo_lo_1560 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1561;
  assign dataGroup_lo_lo_1561 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1562;
  assign dataGroup_lo_lo_1562 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1563;
  assign dataGroup_lo_lo_1563 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1564;
  assign dataGroup_lo_lo_1564 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1565;
  assign dataGroup_lo_lo_1565 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1566;
  assign dataGroup_lo_lo_1566 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1567;
  assign dataGroup_lo_lo_1567 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1568;
  assign dataGroup_lo_lo_1568 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1569;
  assign dataGroup_lo_lo_1569 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1570;
  assign dataGroup_lo_lo_1570 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1571;
  assign dataGroup_lo_lo_1571 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1572;
  assign dataGroup_lo_lo_1572 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1573;
  assign dataGroup_lo_lo_1573 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1574;
  assign dataGroup_lo_lo_1574 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1575;
  assign dataGroup_lo_lo_1575 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1576;
  assign dataGroup_lo_lo_1576 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1577;
  assign dataGroup_lo_lo_1577 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1578;
  assign dataGroup_lo_lo_1578 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1579;
  assign dataGroup_lo_lo_1579 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1580;
  assign dataGroup_lo_lo_1580 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1581;
  assign dataGroup_lo_lo_1581 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1582;
  assign dataGroup_lo_lo_1582 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1583;
  assign dataGroup_lo_lo_1583 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1584;
  assign dataGroup_lo_lo_1584 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1585;
  assign dataGroup_lo_lo_1585 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1586;
  assign dataGroup_lo_lo_1586 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1587;
  assign dataGroup_lo_lo_1587 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1588;
  assign dataGroup_lo_lo_1588 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1589;
  assign dataGroup_lo_lo_1589 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1590;
  assign dataGroup_lo_lo_1590 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1591;
  assign dataGroup_lo_lo_1591 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1592;
  assign dataGroup_lo_lo_1592 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1593;
  assign dataGroup_lo_lo_1593 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1594;
  assign dataGroup_lo_lo_1594 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1595;
  assign dataGroup_lo_lo_1595 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1596;
  assign dataGroup_lo_lo_1596 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1597;
  assign dataGroup_lo_lo_1597 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1598;
  assign dataGroup_lo_lo_1598 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1599;
  assign dataGroup_lo_lo_1599 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1600;
  assign dataGroup_lo_lo_1600 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1601;
  assign dataGroup_lo_lo_1601 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1602;
  assign dataGroup_lo_lo_1602 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1603;
  assign dataGroup_lo_lo_1603 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1604;
  assign dataGroup_lo_lo_1604 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1605;
  assign dataGroup_lo_lo_1605 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1606;
  assign dataGroup_lo_lo_1606 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1607;
  assign dataGroup_lo_lo_1607 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1608;
  assign dataGroup_lo_lo_1608 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1609;
  assign dataGroup_lo_lo_1609 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1610;
  assign dataGroup_lo_lo_1610 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1611;
  assign dataGroup_lo_lo_1611 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1612;
  assign dataGroup_lo_lo_1612 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1613;
  assign dataGroup_lo_lo_1613 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1614;
  assign dataGroup_lo_lo_1614 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1615;
  assign dataGroup_lo_lo_1615 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1616;
  assign dataGroup_lo_lo_1616 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1617;
  assign dataGroup_lo_lo_1617 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1618;
  assign dataGroup_lo_lo_1618 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1619;
  assign dataGroup_lo_lo_1619 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1620;
  assign dataGroup_lo_lo_1620 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1621;
  assign dataGroup_lo_lo_1621 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1622;
  assign dataGroup_lo_lo_1622 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1623;
  assign dataGroup_lo_lo_1623 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1624;
  assign dataGroup_lo_lo_1624 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1625;
  assign dataGroup_lo_lo_1625 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1626;
  assign dataGroup_lo_lo_1626 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1627;
  assign dataGroup_lo_lo_1627 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1628;
  assign dataGroup_lo_lo_1628 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1629;
  assign dataGroup_lo_lo_1629 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1630;
  assign dataGroup_lo_lo_1630 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1631;
  assign dataGroup_lo_lo_1631 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1632;
  assign dataGroup_lo_lo_1632 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1633;
  assign dataGroup_lo_lo_1633 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1634;
  assign dataGroup_lo_lo_1634 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1635;
  assign dataGroup_lo_lo_1635 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1636;
  assign dataGroup_lo_lo_1636 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1637;
  assign dataGroup_lo_lo_1637 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1638;
  assign dataGroup_lo_lo_1638 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1639;
  assign dataGroup_lo_lo_1639 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1640;
  assign dataGroup_lo_lo_1640 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1641;
  assign dataGroup_lo_lo_1641 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1642;
  assign dataGroup_lo_lo_1642 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1643;
  assign dataGroup_lo_lo_1643 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1644;
  assign dataGroup_lo_lo_1644 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1645;
  assign dataGroup_lo_lo_1645 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1646;
  assign dataGroup_lo_lo_1646 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1647;
  assign dataGroup_lo_lo_1647 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1648;
  assign dataGroup_lo_lo_1648 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1649;
  assign dataGroup_lo_lo_1649 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1650;
  assign dataGroup_lo_lo_1650 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1651;
  assign dataGroup_lo_lo_1651 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1652;
  assign dataGroup_lo_lo_1652 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1653;
  assign dataGroup_lo_lo_1653 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1654;
  assign dataGroup_lo_lo_1654 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1655;
  assign dataGroup_lo_lo_1655 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1656;
  assign dataGroup_lo_lo_1656 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1657;
  assign dataGroup_lo_lo_1657 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1658;
  assign dataGroup_lo_lo_1658 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1659;
  assign dataGroup_lo_lo_1659 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1660;
  assign dataGroup_lo_lo_1660 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1661;
  assign dataGroup_lo_lo_1661 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1662;
  assign dataGroup_lo_lo_1662 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1663;
  assign dataGroup_lo_lo_1663 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1664;
  assign dataGroup_lo_lo_1664 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1665;
  assign dataGroup_lo_lo_1665 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1666;
  assign dataGroup_lo_lo_1666 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1667;
  assign dataGroup_lo_lo_1667 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1668;
  assign dataGroup_lo_lo_1668 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1669;
  assign dataGroup_lo_lo_1669 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1670;
  assign dataGroup_lo_lo_1670 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1671;
  assign dataGroup_lo_lo_1671 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1672;
  assign dataGroup_lo_lo_1672 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1673;
  assign dataGroup_lo_lo_1673 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1674;
  assign dataGroup_lo_lo_1674 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1675;
  assign dataGroup_lo_lo_1675 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1676;
  assign dataGroup_lo_lo_1676 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1677;
  assign dataGroup_lo_lo_1677 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1678;
  assign dataGroup_lo_lo_1678 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1679;
  assign dataGroup_lo_lo_1679 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1680;
  assign dataGroup_lo_lo_1680 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1681;
  assign dataGroup_lo_lo_1681 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1682;
  assign dataGroup_lo_lo_1682 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1683;
  assign dataGroup_lo_lo_1683 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1684;
  assign dataGroup_lo_lo_1684 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1685;
  assign dataGroup_lo_lo_1685 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1686;
  assign dataGroup_lo_lo_1686 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1687;
  assign dataGroup_lo_lo_1687 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1688;
  assign dataGroup_lo_lo_1688 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1689;
  assign dataGroup_lo_lo_1689 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1690;
  assign dataGroup_lo_lo_1690 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1691;
  assign dataGroup_lo_lo_1691 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1692;
  assign dataGroup_lo_lo_1692 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1693;
  assign dataGroup_lo_lo_1693 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1694;
  assign dataGroup_lo_lo_1694 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1695;
  assign dataGroup_lo_lo_1695 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1696;
  assign dataGroup_lo_lo_1696 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1697;
  assign dataGroup_lo_lo_1697 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1698;
  assign dataGroup_lo_lo_1698 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1699;
  assign dataGroup_lo_lo_1699 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1700;
  assign dataGroup_lo_lo_1700 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1701;
  assign dataGroup_lo_lo_1701 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1702;
  assign dataGroup_lo_lo_1702 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1703;
  assign dataGroup_lo_lo_1703 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1704;
  assign dataGroup_lo_lo_1704 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1705;
  assign dataGroup_lo_lo_1705 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1706;
  assign dataGroup_lo_lo_1706 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1707;
  assign dataGroup_lo_lo_1707 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1708;
  assign dataGroup_lo_lo_1708 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1709;
  assign dataGroup_lo_lo_1709 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1710;
  assign dataGroup_lo_lo_1710 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1711;
  assign dataGroup_lo_lo_1711 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1712;
  assign dataGroup_lo_lo_1712 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1713;
  assign dataGroup_lo_lo_1713 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1714;
  assign dataGroup_lo_lo_1714 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1715;
  assign dataGroup_lo_lo_1715 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1716;
  assign dataGroup_lo_lo_1716 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1717;
  assign dataGroup_lo_lo_1717 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1718;
  assign dataGroup_lo_lo_1718 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1719;
  assign dataGroup_lo_lo_1719 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1720;
  assign dataGroup_lo_lo_1720 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1721;
  assign dataGroup_lo_lo_1721 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1722;
  assign dataGroup_lo_lo_1722 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1723;
  assign dataGroup_lo_lo_1723 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1724;
  assign dataGroup_lo_lo_1724 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1725;
  assign dataGroup_lo_lo_1725 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1726;
  assign dataGroup_lo_lo_1726 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1727;
  assign dataGroup_lo_lo_1727 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1728;
  assign dataGroup_lo_lo_1728 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1729;
  assign dataGroup_lo_lo_1729 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1730;
  assign dataGroup_lo_lo_1730 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1731;
  assign dataGroup_lo_lo_1731 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1732;
  assign dataGroup_lo_lo_1732 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1733;
  assign dataGroup_lo_lo_1733 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1734;
  assign dataGroup_lo_lo_1734 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1735;
  assign dataGroup_lo_lo_1735 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1736;
  assign dataGroup_lo_lo_1736 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1737;
  assign dataGroup_lo_lo_1737 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1738;
  assign dataGroup_lo_lo_1738 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1739;
  assign dataGroup_lo_lo_1739 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1740;
  assign dataGroup_lo_lo_1740 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1741;
  assign dataGroup_lo_lo_1741 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1742;
  assign dataGroup_lo_lo_1742 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1743;
  assign dataGroup_lo_lo_1743 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1744;
  assign dataGroup_lo_lo_1744 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1745;
  assign dataGroup_lo_lo_1745 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1746;
  assign dataGroup_lo_lo_1746 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1747;
  assign dataGroup_lo_lo_1747 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1748;
  assign dataGroup_lo_lo_1748 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1749;
  assign dataGroup_lo_lo_1749 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1750;
  assign dataGroup_lo_lo_1750 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1751;
  assign dataGroup_lo_lo_1751 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1752;
  assign dataGroup_lo_lo_1752 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1753;
  assign dataGroup_lo_lo_1753 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1754;
  assign dataGroup_lo_lo_1754 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1755;
  assign dataGroup_lo_lo_1755 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1756;
  assign dataGroup_lo_lo_1756 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1757;
  assign dataGroup_lo_lo_1757 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1758;
  assign dataGroup_lo_lo_1758 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1759;
  assign dataGroup_lo_lo_1759 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1760;
  assign dataGroup_lo_lo_1760 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1761;
  assign dataGroup_lo_lo_1761 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1762;
  assign dataGroup_lo_lo_1762 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1763;
  assign dataGroup_lo_lo_1763 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1764;
  assign dataGroup_lo_lo_1764 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1765;
  assign dataGroup_lo_lo_1765 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1766;
  assign dataGroup_lo_lo_1766 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1767;
  assign dataGroup_lo_lo_1767 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1768;
  assign dataGroup_lo_lo_1768 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1769;
  assign dataGroup_lo_lo_1769 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1770;
  assign dataGroup_lo_lo_1770 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1771;
  assign dataGroup_lo_lo_1771 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1772;
  assign dataGroup_lo_lo_1772 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1773;
  assign dataGroup_lo_lo_1773 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1774;
  assign dataGroup_lo_lo_1774 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1775;
  assign dataGroup_lo_lo_1775 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1776;
  assign dataGroup_lo_lo_1776 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1777;
  assign dataGroup_lo_lo_1777 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1778;
  assign dataGroup_lo_lo_1778 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1779;
  assign dataGroup_lo_lo_1779 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1780;
  assign dataGroup_lo_lo_1780 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1781;
  assign dataGroup_lo_lo_1781 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1782;
  assign dataGroup_lo_lo_1782 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1783;
  assign dataGroup_lo_lo_1783 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1784;
  assign dataGroup_lo_lo_1784 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1785;
  assign dataGroup_lo_lo_1785 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1786;
  assign dataGroup_lo_lo_1786 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1787;
  assign dataGroup_lo_lo_1787 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1788;
  assign dataGroup_lo_lo_1788 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1789;
  assign dataGroup_lo_lo_1789 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1790;
  assign dataGroup_lo_lo_1790 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1791;
  assign dataGroup_lo_lo_1791 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1792;
  assign dataGroup_lo_lo_1792 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1793;
  assign dataGroup_lo_lo_1793 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1794;
  assign dataGroup_lo_lo_1794 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1795;
  assign dataGroup_lo_lo_1795 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1796;
  assign dataGroup_lo_lo_1796 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1797;
  assign dataGroup_lo_lo_1797 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1798;
  assign dataGroup_lo_lo_1798 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1799;
  assign dataGroup_lo_lo_1799 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1800;
  assign dataGroup_lo_lo_1800 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1801;
  assign dataGroup_lo_lo_1801 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1802;
  assign dataGroup_lo_lo_1802 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1803;
  assign dataGroup_lo_lo_1803 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1804;
  assign dataGroup_lo_lo_1804 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1805;
  assign dataGroup_lo_lo_1805 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1806;
  assign dataGroup_lo_lo_1806 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1807;
  assign dataGroup_lo_lo_1807 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1808;
  assign dataGroup_lo_lo_1808 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1809;
  assign dataGroup_lo_lo_1809 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1810;
  assign dataGroup_lo_lo_1810 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1811;
  assign dataGroup_lo_lo_1811 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1812;
  assign dataGroup_lo_lo_1812 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1813;
  assign dataGroup_lo_lo_1813 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1814;
  assign dataGroup_lo_lo_1814 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1815;
  assign dataGroup_lo_lo_1815 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1816;
  assign dataGroup_lo_lo_1816 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1817;
  assign dataGroup_lo_lo_1817 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1818;
  assign dataGroup_lo_lo_1818 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1819;
  assign dataGroup_lo_lo_1819 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1820;
  assign dataGroup_lo_lo_1820 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1821;
  assign dataGroup_lo_lo_1821 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1822;
  assign dataGroup_lo_lo_1822 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1823;
  assign dataGroup_lo_lo_1823 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1824;
  assign dataGroup_lo_lo_1824 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1825;
  assign dataGroup_lo_lo_1825 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1826;
  assign dataGroup_lo_lo_1826 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1827;
  assign dataGroup_lo_lo_1827 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1828;
  assign dataGroup_lo_lo_1828 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1829;
  assign dataGroup_lo_lo_1829 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1830;
  assign dataGroup_lo_lo_1830 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1831;
  assign dataGroup_lo_lo_1831 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1832;
  assign dataGroup_lo_lo_1832 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1833;
  assign dataGroup_lo_lo_1833 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1834;
  assign dataGroup_lo_lo_1834 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1835;
  assign dataGroup_lo_lo_1835 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1836;
  assign dataGroup_lo_lo_1836 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1837;
  assign dataGroup_lo_lo_1837 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1838;
  assign dataGroup_lo_lo_1838 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1839;
  assign dataGroup_lo_lo_1839 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1840;
  assign dataGroup_lo_lo_1840 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1841;
  assign dataGroup_lo_lo_1841 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1842;
  assign dataGroup_lo_lo_1842 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1843;
  assign dataGroup_lo_lo_1843 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1844;
  assign dataGroup_lo_lo_1844 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1845;
  assign dataGroup_lo_lo_1845 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1846;
  assign dataGroup_lo_lo_1846 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1847;
  assign dataGroup_lo_lo_1847 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1848;
  assign dataGroup_lo_lo_1848 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1849;
  assign dataGroup_lo_lo_1849 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1850;
  assign dataGroup_lo_lo_1850 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1851;
  assign dataGroup_lo_lo_1851 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1852;
  assign dataGroup_lo_lo_1852 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1853;
  assign dataGroup_lo_lo_1853 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1854;
  assign dataGroup_lo_lo_1854 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1855;
  assign dataGroup_lo_lo_1855 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1856;
  assign dataGroup_lo_lo_1856 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1857;
  assign dataGroup_lo_lo_1857 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1858;
  assign dataGroup_lo_lo_1858 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1859;
  assign dataGroup_lo_lo_1859 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1860;
  assign dataGroup_lo_lo_1860 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1861;
  assign dataGroup_lo_lo_1861 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1862;
  assign dataGroup_lo_lo_1862 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1863;
  assign dataGroup_lo_lo_1863 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1864;
  assign dataGroup_lo_lo_1864 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1865;
  assign dataGroup_lo_lo_1865 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1866;
  assign dataGroup_lo_lo_1866 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1867;
  assign dataGroup_lo_lo_1867 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1868;
  assign dataGroup_lo_lo_1868 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1869;
  assign dataGroup_lo_lo_1869 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1870;
  assign dataGroup_lo_lo_1870 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1871;
  assign dataGroup_lo_lo_1871 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1872;
  assign dataGroup_lo_lo_1872 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1873;
  assign dataGroup_lo_lo_1873 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1874;
  assign dataGroup_lo_lo_1874 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1875;
  assign dataGroup_lo_lo_1875 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1876;
  assign dataGroup_lo_lo_1876 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1877;
  assign dataGroup_lo_lo_1877 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1878;
  assign dataGroup_lo_lo_1878 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1879;
  assign dataGroup_lo_lo_1879 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1880;
  assign dataGroup_lo_lo_1880 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1881;
  assign dataGroup_lo_lo_1881 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1882;
  assign dataGroup_lo_lo_1882 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1883;
  assign dataGroup_lo_lo_1883 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1884;
  assign dataGroup_lo_lo_1884 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1885;
  assign dataGroup_lo_lo_1885 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1886;
  assign dataGroup_lo_lo_1886 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1887;
  assign dataGroup_lo_lo_1887 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1888;
  assign dataGroup_lo_lo_1888 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1889;
  assign dataGroup_lo_lo_1889 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1890;
  assign dataGroup_lo_lo_1890 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1891;
  assign dataGroup_lo_lo_1891 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1892;
  assign dataGroup_lo_lo_1892 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1893;
  assign dataGroup_lo_lo_1893 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1894;
  assign dataGroup_lo_lo_1894 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1895;
  assign dataGroup_lo_lo_1895 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1896;
  assign dataGroup_lo_lo_1896 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1897;
  assign dataGroup_lo_lo_1897 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1898;
  assign dataGroup_lo_lo_1898 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1899;
  assign dataGroup_lo_lo_1899 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1900;
  assign dataGroup_lo_lo_1900 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1901;
  assign dataGroup_lo_lo_1901 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1902;
  assign dataGroup_lo_lo_1902 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1903;
  assign dataGroup_lo_lo_1903 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1904;
  assign dataGroup_lo_lo_1904 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1905;
  assign dataGroup_lo_lo_1905 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1906;
  assign dataGroup_lo_lo_1906 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1907;
  assign dataGroup_lo_lo_1907 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1908;
  assign dataGroup_lo_lo_1908 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1909;
  assign dataGroup_lo_lo_1909 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1910;
  assign dataGroup_lo_lo_1910 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1911;
  assign dataGroup_lo_lo_1911 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1912;
  assign dataGroup_lo_lo_1912 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1913;
  assign dataGroup_lo_lo_1913 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1914;
  assign dataGroup_lo_lo_1914 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1915;
  assign dataGroup_lo_lo_1915 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1916;
  assign dataGroup_lo_lo_1916 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1917;
  assign dataGroup_lo_lo_1917 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1918;
  assign dataGroup_lo_lo_1918 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1919;
  assign dataGroup_lo_lo_1919 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1920;
  assign dataGroup_lo_lo_1920 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1921;
  assign dataGroup_lo_lo_1921 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1922;
  assign dataGroup_lo_lo_1922 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1923;
  assign dataGroup_lo_lo_1923 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1924;
  assign dataGroup_lo_lo_1924 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1925;
  assign dataGroup_lo_lo_1925 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1926;
  assign dataGroup_lo_lo_1926 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1927;
  assign dataGroup_lo_lo_1927 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1928;
  assign dataGroup_lo_lo_1928 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1929;
  assign dataGroup_lo_lo_1929 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1930;
  assign dataGroup_lo_lo_1930 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1931;
  assign dataGroup_lo_lo_1931 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1932;
  assign dataGroup_lo_lo_1932 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1933;
  assign dataGroup_lo_lo_1933 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1934;
  assign dataGroup_lo_lo_1934 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1935;
  assign dataGroup_lo_lo_1935 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1936;
  assign dataGroup_lo_lo_1936 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1937;
  assign dataGroup_lo_lo_1937 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1938;
  assign dataGroup_lo_lo_1938 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1939;
  assign dataGroup_lo_lo_1939 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1940;
  assign dataGroup_lo_lo_1940 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1941;
  assign dataGroup_lo_lo_1941 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1942;
  assign dataGroup_lo_lo_1942 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1943;
  assign dataGroup_lo_lo_1943 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1944;
  assign dataGroup_lo_lo_1944 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1945;
  assign dataGroup_lo_lo_1945 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1946;
  assign dataGroup_lo_lo_1946 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1947;
  assign dataGroup_lo_lo_1947 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1948;
  assign dataGroup_lo_lo_1948 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1949;
  assign dataGroup_lo_lo_1949 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1950;
  assign dataGroup_lo_lo_1950 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1951;
  assign dataGroup_lo_lo_1951 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1952;
  assign dataGroup_lo_lo_1952 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1953;
  assign dataGroup_lo_lo_1953 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1954;
  assign dataGroup_lo_lo_1954 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1955;
  assign dataGroup_lo_lo_1955 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1956;
  assign dataGroup_lo_lo_1956 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1957;
  assign dataGroup_lo_lo_1957 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1958;
  assign dataGroup_lo_lo_1958 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1959;
  assign dataGroup_lo_lo_1959 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1960;
  assign dataGroup_lo_lo_1960 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1961;
  assign dataGroup_lo_lo_1961 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1962;
  assign dataGroup_lo_lo_1962 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1963;
  assign dataGroup_lo_lo_1963 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1964;
  assign dataGroup_lo_lo_1964 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1965;
  assign dataGroup_lo_lo_1965 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1966;
  assign dataGroup_lo_lo_1966 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1967;
  assign dataGroup_lo_lo_1967 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1968;
  assign dataGroup_lo_lo_1968 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1969;
  assign dataGroup_lo_lo_1969 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1970;
  assign dataGroup_lo_lo_1970 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1971;
  assign dataGroup_lo_lo_1971 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1972;
  assign dataGroup_lo_lo_1972 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1973;
  assign dataGroup_lo_lo_1973 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1974;
  assign dataGroup_lo_lo_1974 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1975;
  assign dataGroup_lo_lo_1975 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1976;
  assign dataGroup_lo_lo_1976 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1977;
  assign dataGroup_lo_lo_1977 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1978;
  assign dataGroup_lo_lo_1978 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1979;
  assign dataGroup_lo_lo_1979 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1980;
  assign dataGroup_lo_lo_1980 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1981;
  assign dataGroup_lo_lo_1981 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1982;
  assign dataGroup_lo_lo_1982 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1983;
  assign dataGroup_lo_lo_1983 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1984;
  assign dataGroup_lo_lo_1984 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1985;
  assign dataGroup_lo_lo_1985 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1986;
  assign dataGroup_lo_lo_1986 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1987;
  assign dataGroup_lo_lo_1987 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1988;
  assign dataGroup_lo_lo_1988 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1989;
  assign dataGroup_lo_lo_1989 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1990;
  assign dataGroup_lo_lo_1990 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1991;
  assign dataGroup_lo_lo_1991 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1992;
  assign dataGroup_lo_lo_1992 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1993;
  assign dataGroup_lo_lo_1993 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1994;
  assign dataGroup_lo_lo_1994 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1995;
  assign dataGroup_lo_lo_1995 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1996;
  assign dataGroup_lo_lo_1996 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1997;
  assign dataGroup_lo_lo_1997 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1998;
  assign dataGroup_lo_lo_1998 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_1999;
  assign dataGroup_lo_lo_1999 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2000;
  assign dataGroup_lo_lo_2000 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2001;
  assign dataGroup_lo_lo_2001 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2002;
  assign dataGroup_lo_lo_2002 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2003;
  assign dataGroup_lo_lo_2003 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2004;
  assign dataGroup_lo_lo_2004 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2005;
  assign dataGroup_lo_lo_2005 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2006;
  assign dataGroup_lo_lo_2006 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2007;
  assign dataGroup_lo_lo_2007 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2008;
  assign dataGroup_lo_lo_2008 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2009;
  assign dataGroup_lo_lo_2009 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2010;
  assign dataGroup_lo_lo_2010 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2011;
  assign dataGroup_lo_lo_2011 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2012;
  assign dataGroup_lo_lo_2012 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2013;
  assign dataGroup_lo_lo_2013 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2014;
  assign dataGroup_lo_lo_2014 = _GEN_4;
  wire [511:0]  dataGroup_lo_lo_2015;
  assign dataGroup_lo_lo_2015 = _GEN_4;
  wire [511:0]  _GEN_5 = {dataSelect_3, dataSelect_2};
  wire [511:0]  dataGroup_lo_hi;
  assign dataGroup_lo_hi = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1;
  assign dataGroup_lo_hi_1 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2;
  assign dataGroup_lo_hi_2 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_3;
  assign dataGroup_lo_hi_3 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_4;
  assign dataGroup_lo_hi_4 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_5;
  assign dataGroup_lo_hi_5 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_6;
  assign dataGroup_lo_hi_6 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_7;
  assign dataGroup_lo_hi_7 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_8;
  assign dataGroup_lo_hi_8 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_9;
  assign dataGroup_lo_hi_9 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_10;
  assign dataGroup_lo_hi_10 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_11;
  assign dataGroup_lo_hi_11 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_12;
  assign dataGroup_lo_hi_12 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_13;
  assign dataGroup_lo_hi_13 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_14;
  assign dataGroup_lo_hi_14 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_15;
  assign dataGroup_lo_hi_15 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_16;
  assign dataGroup_lo_hi_16 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_17;
  assign dataGroup_lo_hi_17 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_18;
  assign dataGroup_lo_hi_18 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_19;
  assign dataGroup_lo_hi_19 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_20;
  assign dataGroup_lo_hi_20 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_21;
  assign dataGroup_lo_hi_21 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_22;
  assign dataGroup_lo_hi_22 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_23;
  assign dataGroup_lo_hi_23 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_24;
  assign dataGroup_lo_hi_24 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_25;
  assign dataGroup_lo_hi_25 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_26;
  assign dataGroup_lo_hi_26 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_27;
  assign dataGroup_lo_hi_27 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_28;
  assign dataGroup_lo_hi_28 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_29;
  assign dataGroup_lo_hi_29 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_30;
  assign dataGroup_lo_hi_30 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_31;
  assign dataGroup_lo_hi_31 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_32;
  assign dataGroup_lo_hi_32 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_33;
  assign dataGroup_lo_hi_33 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_34;
  assign dataGroup_lo_hi_34 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_35;
  assign dataGroup_lo_hi_35 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_36;
  assign dataGroup_lo_hi_36 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_37;
  assign dataGroup_lo_hi_37 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_38;
  assign dataGroup_lo_hi_38 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_39;
  assign dataGroup_lo_hi_39 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_40;
  assign dataGroup_lo_hi_40 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_41;
  assign dataGroup_lo_hi_41 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_42;
  assign dataGroup_lo_hi_42 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_43;
  assign dataGroup_lo_hi_43 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_44;
  assign dataGroup_lo_hi_44 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_45;
  assign dataGroup_lo_hi_45 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_46;
  assign dataGroup_lo_hi_46 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_47;
  assign dataGroup_lo_hi_47 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_48;
  assign dataGroup_lo_hi_48 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_49;
  assign dataGroup_lo_hi_49 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_50;
  assign dataGroup_lo_hi_50 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_51;
  assign dataGroup_lo_hi_51 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_52;
  assign dataGroup_lo_hi_52 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_53;
  assign dataGroup_lo_hi_53 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_54;
  assign dataGroup_lo_hi_54 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_55;
  assign dataGroup_lo_hi_55 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_56;
  assign dataGroup_lo_hi_56 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_57;
  assign dataGroup_lo_hi_57 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_58;
  assign dataGroup_lo_hi_58 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_59;
  assign dataGroup_lo_hi_59 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_60;
  assign dataGroup_lo_hi_60 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_61;
  assign dataGroup_lo_hi_61 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_62;
  assign dataGroup_lo_hi_62 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_63;
  assign dataGroup_lo_hi_63 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_64;
  assign dataGroup_lo_hi_64 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_65;
  assign dataGroup_lo_hi_65 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_66;
  assign dataGroup_lo_hi_66 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_67;
  assign dataGroup_lo_hi_67 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_68;
  assign dataGroup_lo_hi_68 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_69;
  assign dataGroup_lo_hi_69 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_70;
  assign dataGroup_lo_hi_70 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_71;
  assign dataGroup_lo_hi_71 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_72;
  assign dataGroup_lo_hi_72 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_73;
  assign dataGroup_lo_hi_73 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_74;
  assign dataGroup_lo_hi_74 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_75;
  assign dataGroup_lo_hi_75 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_76;
  assign dataGroup_lo_hi_76 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_77;
  assign dataGroup_lo_hi_77 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_78;
  assign dataGroup_lo_hi_78 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_79;
  assign dataGroup_lo_hi_79 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_80;
  assign dataGroup_lo_hi_80 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_81;
  assign dataGroup_lo_hi_81 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_82;
  assign dataGroup_lo_hi_82 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_83;
  assign dataGroup_lo_hi_83 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_84;
  assign dataGroup_lo_hi_84 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_85;
  assign dataGroup_lo_hi_85 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_86;
  assign dataGroup_lo_hi_86 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_87;
  assign dataGroup_lo_hi_87 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_88;
  assign dataGroup_lo_hi_88 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_89;
  assign dataGroup_lo_hi_89 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_90;
  assign dataGroup_lo_hi_90 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_91;
  assign dataGroup_lo_hi_91 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_92;
  assign dataGroup_lo_hi_92 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_93;
  assign dataGroup_lo_hi_93 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_94;
  assign dataGroup_lo_hi_94 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_95;
  assign dataGroup_lo_hi_95 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_96;
  assign dataGroup_lo_hi_96 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_97;
  assign dataGroup_lo_hi_97 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_98;
  assign dataGroup_lo_hi_98 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_99;
  assign dataGroup_lo_hi_99 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_100;
  assign dataGroup_lo_hi_100 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_101;
  assign dataGroup_lo_hi_101 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_102;
  assign dataGroup_lo_hi_102 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_103;
  assign dataGroup_lo_hi_103 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_104;
  assign dataGroup_lo_hi_104 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_105;
  assign dataGroup_lo_hi_105 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_106;
  assign dataGroup_lo_hi_106 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_107;
  assign dataGroup_lo_hi_107 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_108;
  assign dataGroup_lo_hi_108 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_109;
  assign dataGroup_lo_hi_109 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_110;
  assign dataGroup_lo_hi_110 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_111;
  assign dataGroup_lo_hi_111 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_112;
  assign dataGroup_lo_hi_112 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_113;
  assign dataGroup_lo_hi_113 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_114;
  assign dataGroup_lo_hi_114 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_115;
  assign dataGroup_lo_hi_115 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_116;
  assign dataGroup_lo_hi_116 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_117;
  assign dataGroup_lo_hi_117 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_118;
  assign dataGroup_lo_hi_118 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_119;
  assign dataGroup_lo_hi_119 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_120;
  assign dataGroup_lo_hi_120 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_121;
  assign dataGroup_lo_hi_121 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_122;
  assign dataGroup_lo_hi_122 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_123;
  assign dataGroup_lo_hi_123 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_124;
  assign dataGroup_lo_hi_124 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_125;
  assign dataGroup_lo_hi_125 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_126;
  assign dataGroup_lo_hi_126 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_127;
  assign dataGroup_lo_hi_127 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_128;
  assign dataGroup_lo_hi_128 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_129;
  assign dataGroup_lo_hi_129 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_130;
  assign dataGroup_lo_hi_130 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_131;
  assign dataGroup_lo_hi_131 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_132;
  assign dataGroup_lo_hi_132 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_133;
  assign dataGroup_lo_hi_133 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_134;
  assign dataGroup_lo_hi_134 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_135;
  assign dataGroup_lo_hi_135 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_136;
  assign dataGroup_lo_hi_136 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_137;
  assign dataGroup_lo_hi_137 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_138;
  assign dataGroup_lo_hi_138 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_139;
  assign dataGroup_lo_hi_139 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_140;
  assign dataGroup_lo_hi_140 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_141;
  assign dataGroup_lo_hi_141 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_142;
  assign dataGroup_lo_hi_142 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_143;
  assign dataGroup_lo_hi_143 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_144;
  assign dataGroup_lo_hi_144 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_145;
  assign dataGroup_lo_hi_145 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_146;
  assign dataGroup_lo_hi_146 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_147;
  assign dataGroup_lo_hi_147 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_148;
  assign dataGroup_lo_hi_148 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_149;
  assign dataGroup_lo_hi_149 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_150;
  assign dataGroup_lo_hi_150 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_151;
  assign dataGroup_lo_hi_151 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_152;
  assign dataGroup_lo_hi_152 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_153;
  assign dataGroup_lo_hi_153 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_154;
  assign dataGroup_lo_hi_154 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_155;
  assign dataGroup_lo_hi_155 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_156;
  assign dataGroup_lo_hi_156 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_157;
  assign dataGroup_lo_hi_157 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_158;
  assign dataGroup_lo_hi_158 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_159;
  assign dataGroup_lo_hi_159 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_160;
  assign dataGroup_lo_hi_160 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_161;
  assign dataGroup_lo_hi_161 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_162;
  assign dataGroup_lo_hi_162 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_163;
  assign dataGroup_lo_hi_163 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_164;
  assign dataGroup_lo_hi_164 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_165;
  assign dataGroup_lo_hi_165 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_166;
  assign dataGroup_lo_hi_166 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_167;
  assign dataGroup_lo_hi_167 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_168;
  assign dataGroup_lo_hi_168 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_169;
  assign dataGroup_lo_hi_169 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_170;
  assign dataGroup_lo_hi_170 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_171;
  assign dataGroup_lo_hi_171 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_172;
  assign dataGroup_lo_hi_172 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_173;
  assign dataGroup_lo_hi_173 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_174;
  assign dataGroup_lo_hi_174 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_175;
  assign dataGroup_lo_hi_175 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_176;
  assign dataGroup_lo_hi_176 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_177;
  assign dataGroup_lo_hi_177 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_178;
  assign dataGroup_lo_hi_178 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_179;
  assign dataGroup_lo_hi_179 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_180;
  assign dataGroup_lo_hi_180 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_181;
  assign dataGroup_lo_hi_181 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_182;
  assign dataGroup_lo_hi_182 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_183;
  assign dataGroup_lo_hi_183 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_184;
  assign dataGroup_lo_hi_184 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_185;
  assign dataGroup_lo_hi_185 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_186;
  assign dataGroup_lo_hi_186 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_187;
  assign dataGroup_lo_hi_187 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_188;
  assign dataGroup_lo_hi_188 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_189;
  assign dataGroup_lo_hi_189 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_190;
  assign dataGroup_lo_hi_190 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_191;
  assign dataGroup_lo_hi_191 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_192;
  assign dataGroup_lo_hi_192 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_193;
  assign dataGroup_lo_hi_193 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_194;
  assign dataGroup_lo_hi_194 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_195;
  assign dataGroup_lo_hi_195 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_196;
  assign dataGroup_lo_hi_196 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_197;
  assign dataGroup_lo_hi_197 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_198;
  assign dataGroup_lo_hi_198 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_199;
  assign dataGroup_lo_hi_199 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_200;
  assign dataGroup_lo_hi_200 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_201;
  assign dataGroup_lo_hi_201 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_202;
  assign dataGroup_lo_hi_202 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_203;
  assign dataGroup_lo_hi_203 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_204;
  assign dataGroup_lo_hi_204 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_205;
  assign dataGroup_lo_hi_205 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_206;
  assign dataGroup_lo_hi_206 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_207;
  assign dataGroup_lo_hi_207 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_208;
  assign dataGroup_lo_hi_208 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_209;
  assign dataGroup_lo_hi_209 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_210;
  assign dataGroup_lo_hi_210 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_211;
  assign dataGroup_lo_hi_211 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_212;
  assign dataGroup_lo_hi_212 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_213;
  assign dataGroup_lo_hi_213 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_214;
  assign dataGroup_lo_hi_214 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_215;
  assign dataGroup_lo_hi_215 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_216;
  assign dataGroup_lo_hi_216 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_217;
  assign dataGroup_lo_hi_217 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_218;
  assign dataGroup_lo_hi_218 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_219;
  assign dataGroup_lo_hi_219 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_220;
  assign dataGroup_lo_hi_220 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_221;
  assign dataGroup_lo_hi_221 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_222;
  assign dataGroup_lo_hi_222 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_223;
  assign dataGroup_lo_hi_223 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_224;
  assign dataGroup_lo_hi_224 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_225;
  assign dataGroup_lo_hi_225 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_226;
  assign dataGroup_lo_hi_226 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_227;
  assign dataGroup_lo_hi_227 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_228;
  assign dataGroup_lo_hi_228 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_229;
  assign dataGroup_lo_hi_229 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_230;
  assign dataGroup_lo_hi_230 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_231;
  assign dataGroup_lo_hi_231 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_232;
  assign dataGroup_lo_hi_232 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_233;
  assign dataGroup_lo_hi_233 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_234;
  assign dataGroup_lo_hi_234 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_235;
  assign dataGroup_lo_hi_235 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_236;
  assign dataGroup_lo_hi_236 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_237;
  assign dataGroup_lo_hi_237 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_238;
  assign dataGroup_lo_hi_238 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_239;
  assign dataGroup_lo_hi_239 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_240;
  assign dataGroup_lo_hi_240 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_241;
  assign dataGroup_lo_hi_241 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_242;
  assign dataGroup_lo_hi_242 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_243;
  assign dataGroup_lo_hi_243 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_244;
  assign dataGroup_lo_hi_244 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_245;
  assign dataGroup_lo_hi_245 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_246;
  assign dataGroup_lo_hi_246 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_247;
  assign dataGroup_lo_hi_247 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_248;
  assign dataGroup_lo_hi_248 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_249;
  assign dataGroup_lo_hi_249 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_250;
  assign dataGroup_lo_hi_250 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_251;
  assign dataGroup_lo_hi_251 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_252;
  assign dataGroup_lo_hi_252 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_253;
  assign dataGroup_lo_hi_253 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_254;
  assign dataGroup_lo_hi_254 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_255;
  assign dataGroup_lo_hi_255 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_256;
  assign dataGroup_lo_hi_256 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_257;
  assign dataGroup_lo_hi_257 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_258;
  assign dataGroup_lo_hi_258 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_259;
  assign dataGroup_lo_hi_259 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_260;
  assign dataGroup_lo_hi_260 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_261;
  assign dataGroup_lo_hi_261 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_262;
  assign dataGroup_lo_hi_262 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_263;
  assign dataGroup_lo_hi_263 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_264;
  assign dataGroup_lo_hi_264 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_265;
  assign dataGroup_lo_hi_265 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_266;
  assign dataGroup_lo_hi_266 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_267;
  assign dataGroup_lo_hi_267 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_268;
  assign dataGroup_lo_hi_268 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_269;
  assign dataGroup_lo_hi_269 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_270;
  assign dataGroup_lo_hi_270 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_271;
  assign dataGroup_lo_hi_271 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_272;
  assign dataGroup_lo_hi_272 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_273;
  assign dataGroup_lo_hi_273 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_274;
  assign dataGroup_lo_hi_274 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_275;
  assign dataGroup_lo_hi_275 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_276;
  assign dataGroup_lo_hi_276 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_277;
  assign dataGroup_lo_hi_277 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_278;
  assign dataGroup_lo_hi_278 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_279;
  assign dataGroup_lo_hi_279 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_280;
  assign dataGroup_lo_hi_280 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_281;
  assign dataGroup_lo_hi_281 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_282;
  assign dataGroup_lo_hi_282 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_283;
  assign dataGroup_lo_hi_283 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_284;
  assign dataGroup_lo_hi_284 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_285;
  assign dataGroup_lo_hi_285 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_286;
  assign dataGroup_lo_hi_286 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_287;
  assign dataGroup_lo_hi_287 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_288;
  assign dataGroup_lo_hi_288 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_289;
  assign dataGroup_lo_hi_289 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_290;
  assign dataGroup_lo_hi_290 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_291;
  assign dataGroup_lo_hi_291 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_292;
  assign dataGroup_lo_hi_292 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_293;
  assign dataGroup_lo_hi_293 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_294;
  assign dataGroup_lo_hi_294 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_295;
  assign dataGroup_lo_hi_295 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_296;
  assign dataGroup_lo_hi_296 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_297;
  assign dataGroup_lo_hi_297 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_298;
  assign dataGroup_lo_hi_298 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_299;
  assign dataGroup_lo_hi_299 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_300;
  assign dataGroup_lo_hi_300 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_301;
  assign dataGroup_lo_hi_301 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_302;
  assign dataGroup_lo_hi_302 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_303;
  assign dataGroup_lo_hi_303 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_304;
  assign dataGroup_lo_hi_304 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_305;
  assign dataGroup_lo_hi_305 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_306;
  assign dataGroup_lo_hi_306 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_307;
  assign dataGroup_lo_hi_307 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_308;
  assign dataGroup_lo_hi_308 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_309;
  assign dataGroup_lo_hi_309 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_310;
  assign dataGroup_lo_hi_310 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_311;
  assign dataGroup_lo_hi_311 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_312;
  assign dataGroup_lo_hi_312 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_313;
  assign dataGroup_lo_hi_313 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_314;
  assign dataGroup_lo_hi_314 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_315;
  assign dataGroup_lo_hi_315 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_316;
  assign dataGroup_lo_hi_316 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_317;
  assign dataGroup_lo_hi_317 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_318;
  assign dataGroup_lo_hi_318 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_319;
  assign dataGroup_lo_hi_319 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_320;
  assign dataGroup_lo_hi_320 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_321;
  assign dataGroup_lo_hi_321 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_322;
  assign dataGroup_lo_hi_322 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_323;
  assign dataGroup_lo_hi_323 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_324;
  assign dataGroup_lo_hi_324 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_325;
  assign dataGroup_lo_hi_325 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_326;
  assign dataGroup_lo_hi_326 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_327;
  assign dataGroup_lo_hi_327 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_328;
  assign dataGroup_lo_hi_328 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_329;
  assign dataGroup_lo_hi_329 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_330;
  assign dataGroup_lo_hi_330 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_331;
  assign dataGroup_lo_hi_331 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_332;
  assign dataGroup_lo_hi_332 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_333;
  assign dataGroup_lo_hi_333 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_334;
  assign dataGroup_lo_hi_334 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_335;
  assign dataGroup_lo_hi_335 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_336;
  assign dataGroup_lo_hi_336 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_337;
  assign dataGroup_lo_hi_337 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_338;
  assign dataGroup_lo_hi_338 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_339;
  assign dataGroup_lo_hi_339 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_340;
  assign dataGroup_lo_hi_340 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_341;
  assign dataGroup_lo_hi_341 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_342;
  assign dataGroup_lo_hi_342 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_343;
  assign dataGroup_lo_hi_343 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_344;
  assign dataGroup_lo_hi_344 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_345;
  assign dataGroup_lo_hi_345 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_346;
  assign dataGroup_lo_hi_346 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_347;
  assign dataGroup_lo_hi_347 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_348;
  assign dataGroup_lo_hi_348 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_349;
  assign dataGroup_lo_hi_349 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_350;
  assign dataGroup_lo_hi_350 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_351;
  assign dataGroup_lo_hi_351 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_352;
  assign dataGroup_lo_hi_352 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_353;
  assign dataGroup_lo_hi_353 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_354;
  assign dataGroup_lo_hi_354 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_355;
  assign dataGroup_lo_hi_355 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_356;
  assign dataGroup_lo_hi_356 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_357;
  assign dataGroup_lo_hi_357 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_358;
  assign dataGroup_lo_hi_358 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_359;
  assign dataGroup_lo_hi_359 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_360;
  assign dataGroup_lo_hi_360 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_361;
  assign dataGroup_lo_hi_361 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_362;
  assign dataGroup_lo_hi_362 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_363;
  assign dataGroup_lo_hi_363 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_364;
  assign dataGroup_lo_hi_364 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_365;
  assign dataGroup_lo_hi_365 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_366;
  assign dataGroup_lo_hi_366 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_367;
  assign dataGroup_lo_hi_367 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_368;
  assign dataGroup_lo_hi_368 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_369;
  assign dataGroup_lo_hi_369 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_370;
  assign dataGroup_lo_hi_370 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_371;
  assign dataGroup_lo_hi_371 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_372;
  assign dataGroup_lo_hi_372 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_373;
  assign dataGroup_lo_hi_373 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_374;
  assign dataGroup_lo_hi_374 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_375;
  assign dataGroup_lo_hi_375 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_376;
  assign dataGroup_lo_hi_376 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_377;
  assign dataGroup_lo_hi_377 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_378;
  assign dataGroup_lo_hi_378 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_379;
  assign dataGroup_lo_hi_379 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_380;
  assign dataGroup_lo_hi_380 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_381;
  assign dataGroup_lo_hi_381 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_382;
  assign dataGroup_lo_hi_382 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_383;
  assign dataGroup_lo_hi_383 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_384;
  assign dataGroup_lo_hi_384 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_385;
  assign dataGroup_lo_hi_385 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_386;
  assign dataGroup_lo_hi_386 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_387;
  assign dataGroup_lo_hi_387 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_388;
  assign dataGroup_lo_hi_388 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_389;
  assign dataGroup_lo_hi_389 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_390;
  assign dataGroup_lo_hi_390 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_391;
  assign dataGroup_lo_hi_391 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_392;
  assign dataGroup_lo_hi_392 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_393;
  assign dataGroup_lo_hi_393 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_394;
  assign dataGroup_lo_hi_394 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_395;
  assign dataGroup_lo_hi_395 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_396;
  assign dataGroup_lo_hi_396 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_397;
  assign dataGroup_lo_hi_397 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_398;
  assign dataGroup_lo_hi_398 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_399;
  assign dataGroup_lo_hi_399 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_400;
  assign dataGroup_lo_hi_400 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_401;
  assign dataGroup_lo_hi_401 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_402;
  assign dataGroup_lo_hi_402 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_403;
  assign dataGroup_lo_hi_403 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_404;
  assign dataGroup_lo_hi_404 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_405;
  assign dataGroup_lo_hi_405 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_406;
  assign dataGroup_lo_hi_406 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_407;
  assign dataGroup_lo_hi_407 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_408;
  assign dataGroup_lo_hi_408 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_409;
  assign dataGroup_lo_hi_409 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_410;
  assign dataGroup_lo_hi_410 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_411;
  assign dataGroup_lo_hi_411 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_412;
  assign dataGroup_lo_hi_412 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_413;
  assign dataGroup_lo_hi_413 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_414;
  assign dataGroup_lo_hi_414 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_415;
  assign dataGroup_lo_hi_415 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_416;
  assign dataGroup_lo_hi_416 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_417;
  assign dataGroup_lo_hi_417 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_418;
  assign dataGroup_lo_hi_418 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_419;
  assign dataGroup_lo_hi_419 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_420;
  assign dataGroup_lo_hi_420 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_421;
  assign dataGroup_lo_hi_421 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_422;
  assign dataGroup_lo_hi_422 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_423;
  assign dataGroup_lo_hi_423 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_424;
  assign dataGroup_lo_hi_424 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_425;
  assign dataGroup_lo_hi_425 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_426;
  assign dataGroup_lo_hi_426 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_427;
  assign dataGroup_lo_hi_427 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_428;
  assign dataGroup_lo_hi_428 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_429;
  assign dataGroup_lo_hi_429 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_430;
  assign dataGroup_lo_hi_430 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_431;
  assign dataGroup_lo_hi_431 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_432;
  assign dataGroup_lo_hi_432 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_433;
  assign dataGroup_lo_hi_433 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_434;
  assign dataGroup_lo_hi_434 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_435;
  assign dataGroup_lo_hi_435 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_436;
  assign dataGroup_lo_hi_436 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_437;
  assign dataGroup_lo_hi_437 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_438;
  assign dataGroup_lo_hi_438 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_439;
  assign dataGroup_lo_hi_439 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_440;
  assign dataGroup_lo_hi_440 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_441;
  assign dataGroup_lo_hi_441 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_442;
  assign dataGroup_lo_hi_442 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_443;
  assign dataGroup_lo_hi_443 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_444;
  assign dataGroup_lo_hi_444 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_445;
  assign dataGroup_lo_hi_445 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_446;
  assign dataGroup_lo_hi_446 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_447;
  assign dataGroup_lo_hi_447 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_448;
  assign dataGroup_lo_hi_448 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_449;
  assign dataGroup_lo_hi_449 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_450;
  assign dataGroup_lo_hi_450 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_451;
  assign dataGroup_lo_hi_451 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_452;
  assign dataGroup_lo_hi_452 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_453;
  assign dataGroup_lo_hi_453 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_454;
  assign dataGroup_lo_hi_454 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_455;
  assign dataGroup_lo_hi_455 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_456;
  assign dataGroup_lo_hi_456 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_457;
  assign dataGroup_lo_hi_457 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_458;
  assign dataGroup_lo_hi_458 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_459;
  assign dataGroup_lo_hi_459 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_460;
  assign dataGroup_lo_hi_460 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_461;
  assign dataGroup_lo_hi_461 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_462;
  assign dataGroup_lo_hi_462 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_463;
  assign dataGroup_lo_hi_463 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_464;
  assign dataGroup_lo_hi_464 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_465;
  assign dataGroup_lo_hi_465 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_466;
  assign dataGroup_lo_hi_466 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_467;
  assign dataGroup_lo_hi_467 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_468;
  assign dataGroup_lo_hi_468 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_469;
  assign dataGroup_lo_hi_469 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_470;
  assign dataGroup_lo_hi_470 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_471;
  assign dataGroup_lo_hi_471 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_472;
  assign dataGroup_lo_hi_472 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_473;
  assign dataGroup_lo_hi_473 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_474;
  assign dataGroup_lo_hi_474 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_475;
  assign dataGroup_lo_hi_475 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_476;
  assign dataGroup_lo_hi_476 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_477;
  assign dataGroup_lo_hi_477 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_478;
  assign dataGroup_lo_hi_478 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_479;
  assign dataGroup_lo_hi_479 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_480;
  assign dataGroup_lo_hi_480 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_481;
  assign dataGroup_lo_hi_481 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_482;
  assign dataGroup_lo_hi_482 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_483;
  assign dataGroup_lo_hi_483 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_484;
  assign dataGroup_lo_hi_484 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_485;
  assign dataGroup_lo_hi_485 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_486;
  assign dataGroup_lo_hi_486 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_487;
  assign dataGroup_lo_hi_487 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_488;
  assign dataGroup_lo_hi_488 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_489;
  assign dataGroup_lo_hi_489 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_490;
  assign dataGroup_lo_hi_490 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_491;
  assign dataGroup_lo_hi_491 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_492;
  assign dataGroup_lo_hi_492 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_493;
  assign dataGroup_lo_hi_493 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_494;
  assign dataGroup_lo_hi_494 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_495;
  assign dataGroup_lo_hi_495 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_496;
  assign dataGroup_lo_hi_496 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_497;
  assign dataGroup_lo_hi_497 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_498;
  assign dataGroup_lo_hi_498 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_499;
  assign dataGroup_lo_hi_499 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_500;
  assign dataGroup_lo_hi_500 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_501;
  assign dataGroup_lo_hi_501 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_502;
  assign dataGroup_lo_hi_502 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_503;
  assign dataGroup_lo_hi_503 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_504;
  assign dataGroup_lo_hi_504 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_505;
  assign dataGroup_lo_hi_505 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_506;
  assign dataGroup_lo_hi_506 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_507;
  assign dataGroup_lo_hi_507 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_508;
  assign dataGroup_lo_hi_508 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_509;
  assign dataGroup_lo_hi_509 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_510;
  assign dataGroup_lo_hi_510 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_511;
  assign dataGroup_lo_hi_511 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_512;
  assign dataGroup_lo_hi_512 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_513;
  assign dataGroup_lo_hi_513 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_514;
  assign dataGroup_lo_hi_514 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_515;
  assign dataGroup_lo_hi_515 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_516;
  assign dataGroup_lo_hi_516 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_517;
  assign dataGroup_lo_hi_517 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_518;
  assign dataGroup_lo_hi_518 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_519;
  assign dataGroup_lo_hi_519 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_520;
  assign dataGroup_lo_hi_520 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_521;
  assign dataGroup_lo_hi_521 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_522;
  assign dataGroup_lo_hi_522 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_523;
  assign dataGroup_lo_hi_523 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_524;
  assign dataGroup_lo_hi_524 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_525;
  assign dataGroup_lo_hi_525 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_526;
  assign dataGroup_lo_hi_526 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_527;
  assign dataGroup_lo_hi_527 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_528;
  assign dataGroup_lo_hi_528 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_529;
  assign dataGroup_lo_hi_529 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_530;
  assign dataGroup_lo_hi_530 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_531;
  assign dataGroup_lo_hi_531 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_532;
  assign dataGroup_lo_hi_532 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_533;
  assign dataGroup_lo_hi_533 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_534;
  assign dataGroup_lo_hi_534 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_535;
  assign dataGroup_lo_hi_535 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_536;
  assign dataGroup_lo_hi_536 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_537;
  assign dataGroup_lo_hi_537 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_538;
  assign dataGroup_lo_hi_538 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_539;
  assign dataGroup_lo_hi_539 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_540;
  assign dataGroup_lo_hi_540 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_541;
  assign dataGroup_lo_hi_541 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_542;
  assign dataGroup_lo_hi_542 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_543;
  assign dataGroup_lo_hi_543 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_544;
  assign dataGroup_lo_hi_544 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_545;
  assign dataGroup_lo_hi_545 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_546;
  assign dataGroup_lo_hi_546 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_547;
  assign dataGroup_lo_hi_547 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_548;
  assign dataGroup_lo_hi_548 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_549;
  assign dataGroup_lo_hi_549 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_550;
  assign dataGroup_lo_hi_550 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_551;
  assign dataGroup_lo_hi_551 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_552;
  assign dataGroup_lo_hi_552 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_553;
  assign dataGroup_lo_hi_553 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_554;
  assign dataGroup_lo_hi_554 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_555;
  assign dataGroup_lo_hi_555 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_556;
  assign dataGroup_lo_hi_556 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_557;
  assign dataGroup_lo_hi_557 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_558;
  assign dataGroup_lo_hi_558 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_559;
  assign dataGroup_lo_hi_559 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_560;
  assign dataGroup_lo_hi_560 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_561;
  assign dataGroup_lo_hi_561 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_562;
  assign dataGroup_lo_hi_562 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_563;
  assign dataGroup_lo_hi_563 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_564;
  assign dataGroup_lo_hi_564 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_565;
  assign dataGroup_lo_hi_565 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_566;
  assign dataGroup_lo_hi_566 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_567;
  assign dataGroup_lo_hi_567 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_568;
  assign dataGroup_lo_hi_568 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_569;
  assign dataGroup_lo_hi_569 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_570;
  assign dataGroup_lo_hi_570 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_571;
  assign dataGroup_lo_hi_571 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_572;
  assign dataGroup_lo_hi_572 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_573;
  assign dataGroup_lo_hi_573 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_574;
  assign dataGroup_lo_hi_574 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_575;
  assign dataGroup_lo_hi_575 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_576;
  assign dataGroup_lo_hi_576 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_577;
  assign dataGroup_lo_hi_577 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_578;
  assign dataGroup_lo_hi_578 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_579;
  assign dataGroup_lo_hi_579 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_580;
  assign dataGroup_lo_hi_580 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_581;
  assign dataGroup_lo_hi_581 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_582;
  assign dataGroup_lo_hi_582 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_583;
  assign dataGroup_lo_hi_583 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_584;
  assign dataGroup_lo_hi_584 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_585;
  assign dataGroup_lo_hi_585 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_586;
  assign dataGroup_lo_hi_586 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_587;
  assign dataGroup_lo_hi_587 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_588;
  assign dataGroup_lo_hi_588 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_589;
  assign dataGroup_lo_hi_589 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_590;
  assign dataGroup_lo_hi_590 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_591;
  assign dataGroup_lo_hi_591 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_592;
  assign dataGroup_lo_hi_592 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_593;
  assign dataGroup_lo_hi_593 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_594;
  assign dataGroup_lo_hi_594 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_595;
  assign dataGroup_lo_hi_595 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_596;
  assign dataGroup_lo_hi_596 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_597;
  assign dataGroup_lo_hi_597 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_598;
  assign dataGroup_lo_hi_598 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_599;
  assign dataGroup_lo_hi_599 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_600;
  assign dataGroup_lo_hi_600 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_601;
  assign dataGroup_lo_hi_601 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_602;
  assign dataGroup_lo_hi_602 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_603;
  assign dataGroup_lo_hi_603 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_604;
  assign dataGroup_lo_hi_604 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_605;
  assign dataGroup_lo_hi_605 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_606;
  assign dataGroup_lo_hi_606 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_607;
  assign dataGroup_lo_hi_607 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_608;
  assign dataGroup_lo_hi_608 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_609;
  assign dataGroup_lo_hi_609 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_610;
  assign dataGroup_lo_hi_610 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_611;
  assign dataGroup_lo_hi_611 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_612;
  assign dataGroup_lo_hi_612 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_613;
  assign dataGroup_lo_hi_613 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_614;
  assign dataGroup_lo_hi_614 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_615;
  assign dataGroup_lo_hi_615 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_616;
  assign dataGroup_lo_hi_616 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_617;
  assign dataGroup_lo_hi_617 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_618;
  assign dataGroup_lo_hi_618 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_619;
  assign dataGroup_lo_hi_619 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_620;
  assign dataGroup_lo_hi_620 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_621;
  assign dataGroup_lo_hi_621 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_622;
  assign dataGroup_lo_hi_622 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_623;
  assign dataGroup_lo_hi_623 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_624;
  assign dataGroup_lo_hi_624 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_625;
  assign dataGroup_lo_hi_625 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_626;
  assign dataGroup_lo_hi_626 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_627;
  assign dataGroup_lo_hi_627 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_628;
  assign dataGroup_lo_hi_628 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_629;
  assign dataGroup_lo_hi_629 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_630;
  assign dataGroup_lo_hi_630 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_631;
  assign dataGroup_lo_hi_631 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_632;
  assign dataGroup_lo_hi_632 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_633;
  assign dataGroup_lo_hi_633 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_634;
  assign dataGroup_lo_hi_634 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_635;
  assign dataGroup_lo_hi_635 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_636;
  assign dataGroup_lo_hi_636 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_637;
  assign dataGroup_lo_hi_637 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_638;
  assign dataGroup_lo_hi_638 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_639;
  assign dataGroup_lo_hi_639 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_640;
  assign dataGroup_lo_hi_640 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_641;
  assign dataGroup_lo_hi_641 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_642;
  assign dataGroup_lo_hi_642 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_643;
  assign dataGroup_lo_hi_643 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_644;
  assign dataGroup_lo_hi_644 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_645;
  assign dataGroup_lo_hi_645 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_646;
  assign dataGroup_lo_hi_646 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_647;
  assign dataGroup_lo_hi_647 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_648;
  assign dataGroup_lo_hi_648 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_649;
  assign dataGroup_lo_hi_649 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_650;
  assign dataGroup_lo_hi_650 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_651;
  assign dataGroup_lo_hi_651 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_652;
  assign dataGroup_lo_hi_652 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_653;
  assign dataGroup_lo_hi_653 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_654;
  assign dataGroup_lo_hi_654 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_655;
  assign dataGroup_lo_hi_655 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_656;
  assign dataGroup_lo_hi_656 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_657;
  assign dataGroup_lo_hi_657 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_658;
  assign dataGroup_lo_hi_658 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_659;
  assign dataGroup_lo_hi_659 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_660;
  assign dataGroup_lo_hi_660 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_661;
  assign dataGroup_lo_hi_661 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_662;
  assign dataGroup_lo_hi_662 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_663;
  assign dataGroup_lo_hi_663 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_664;
  assign dataGroup_lo_hi_664 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_665;
  assign dataGroup_lo_hi_665 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_666;
  assign dataGroup_lo_hi_666 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_667;
  assign dataGroup_lo_hi_667 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_668;
  assign dataGroup_lo_hi_668 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_669;
  assign dataGroup_lo_hi_669 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_670;
  assign dataGroup_lo_hi_670 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_671;
  assign dataGroup_lo_hi_671 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_672;
  assign dataGroup_lo_hi_672 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_673;
  assign dataGroup_lo_hi_673 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_674;
  assign dataGroup_lo_hi_674 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_675;
  assign dataGroup_lo_hi_675 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_676;
  assign dataGroup_lo_hi_676 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_677;
  assign dataGroup_lo_hi_677 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_678;
  assign dataGroup_lo_hi_678 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_679;
  assign dataGroup_lo_hi_679 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_680;
  assign dataGroup_lo_hi_680 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_681;
  assign dataGroup_lo_hi_681 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_682;
  assign dataGroup_lo_hi_682 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_683;
  assign dataGroup_lo_hi_683 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_684;
  assign dataGroup_lo_hi_684 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_685;
  assign dataGroup_lo_hi_685 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_686;
  assign dataGroup_lo_hi_686 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_687;
  assign dataGroup_lo_hi_687 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_688;
  assign dataGroup_lo_hi_688 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_689;
  assign dataGroup_lo_hi_689 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_690;
  assign dataGroup_lo_hi_690 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_691;
  assign dataGroup_lo_hi_691 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_692;
  assign dataGroup_lo_hi_692 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_693;
  assign dataGroup_lo_hi_693 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_694;
  assign dataGroup_lo_hi_694 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_695;
  assign dataGroup_lo_hi_695 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_696;
  assign dataGroup_lo_hi_696 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_697;
  assign dataGroup_lo_hi_697 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_698;
  assign dataGroup_lo_hi_698 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_699;
  assign dataGroup_lo_hi_699 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_700;
  assign dataGroup_lo_hi_700 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_701;
  assign dataGroup_lo_hi_701 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_702;
  assign dataGroup_lo_hi_702 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_703;
  assign dataGroup_lo_hi_703 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_704;
  assign dataGroup_lo_hi_704 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_705;
  assign dataGroup_lo_hi_705 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_706;
  assign dataGroup_lo_hi_706 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_707;
  assign dataGroup_lo_hi_707 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_708;
  assign dataGroup_lo_hi_708 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_709;
  assign dataGroup_lo_hi_709 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_710;
  assign dataGroup_lo_hi_710 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_711;
  assign dataGroup_lo_hi_711 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_712;
  assign dataGroup_lo_hi_712 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_713;
  assign dataGroup_lo_hi_713 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_714;
  assign dataGroup_lo_hi_714 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_715;
  assign dataGroup_lo_hi_715 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_716;
  assign dataGroup_lo_hi_716 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_717;
  assign dataGroup_lo_hi_717 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_718;
  assign dataGroup_lo_hi_718 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_719;
  assign dataGroup_lo_hi_719 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_720;
  assign dataGroup_lo_hi_720 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_721;
  assign dataGroup_lo_hi_721 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_722;
  assign dataGroup_lo_hi_722 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_723;
  assign dataGroup_lo_hi_723 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_724;
  assign dataGroup_lo_hi_724 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_725;
  assign dataGroup_lo_hi_725 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_726;
  assign dataGroup_lo_hi_726 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_727;
  assign dataGroup_lo_hi_727 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_728;
  assign dataGroup_lo_hi_728 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_729;
  assign dataGroup_lo_hi_729 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_730;
  assign dataGroup_lo_hi_730 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_731;
  assign dataGroup_lo_hi_731 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_732;
  assign dataGroup_lo_hi_732 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_733;
  assign dataGroup_lo_hi_733 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_734;
  assign dataGroup_lo_hi_734 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_735;
  assign dataGroup_lo_hi_735 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_736;
  assign dataGroup_lo_hi_736 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_737;
  assign dataGroup_lo_hi_737 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_738;
  assign dataGroup_lo_hi_738 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_739;
  assign dataGroup_lo_hi_739 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_740;
  assign dataGroup_lo_hi_740 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_741;
  assign dataGroup_lo_hi_741 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_742;
  assign dataGroup_lo_hi_742 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_743;
  assign dataGroup_lo_hi_743 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_744;
  assign dataGroup_lo_hi_744 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_745;
  assign dataGroup_lo_hi_745 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_746;
  assign dataGroup_lo_hi_746 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_747;
  assign dataGroup_lo_hi_747 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_748;
  assign dataGroup_lo_hi_748 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_749;
  assign dataGroup_lo_hi_749 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_750;
  assign dataGroup_lo_hi_750 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_751;
  assign dataGroup_lo_hi_751 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_752;
  assign dataGroup_lo_hi_752 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_753;
  assign dataGroup_lo_hi_753 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_754;
  assign dataGroup_lo_hi_754 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_755;
  assign dataGroup_lo_hi_755 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_756;
  assign dataGroup_lo_hi_756 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_757;
  assign dataGroup_lo_hi_757 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_758;
  assign dataGroup_lo_hi_758 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_759;
  assign dataGroup_lo_hi_759 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_760;
  assign dataGroup_lo_hi_760 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_761;
  assign dataGroup_lo_hi_761 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_762;
  assign dataGroup_lo_hi_762 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_763;
  assign dataGroup_lo_hi_763 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_764;
  assign dataGroup_lo_hi_764 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_765;
  assign dataGroup_lo_hi_765 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_766;
  assign dataGroup_lo_hi_766 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_767;
  assign dataGroup_lo_hi_767 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_768;
  assign dataGroup_lo_hi_768 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_769;
  assign dataGroup_lo_hi_769 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_770;
  assign dataGroup_lo_hi_770 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_771;
  assign dataGroup_lo_hi_771 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_772;
  assign dataGroup_lo_hi_772 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_773;
  assign dataGroup_lo_hi_773 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_774;
  assign dataGroup_lo_hi_774 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_775;
  assign dataGroup_lo_hi_775 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_776;
  assign dataGroup_lo_hi_776 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_777;
  assign dataGroup_lo_hi_777 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_778;
  assign dataGroup_lo_hi_778 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_779;
  assign dataGroup_lo_hi_779 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_780;
  assign dataGroup_lo_hi_780 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_781;
  assign dataGroup_lo_hi_781 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_782;
  assign dataGroup_lo_hi_782 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_783;
  assign dataGroup_lo_hi_783 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_784;
  assign dataGroup_lo_hi_784 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_785;
  assign dataGroup_lo_hi_785 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_786;
  assign dataGroup_lo_hi_786 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_787;
  assign dataGroup_lo_hi_787 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_788;
  assign dataGroup_lo_hi_788 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_789;
  assign dataGroup_lo_hi_789 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_790;
  assign dataGroup_lo_hi_790 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_791;
  assign dataGroup_lo_hi_791 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_792;
  assign dataGroup_lo_hi_792 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_793;
  assign dataGroup_lo_hi_793 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_794;
  assign dataGroup_lo_hi_794 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_795;
  assign dataGroup_lo_hi_795 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_796;
  assign dataGroup_lo_hi_796 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_797;
  assign dataGroup_lo_hi_797 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_798;
  assign dataGroup_lo_hi_798 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_799;
  assign dataGroup_lo_hi_799 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_800;
  assign dataGroup_lo_hi_800 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_801;
  assign dataGroup_lo_hi_801 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_802;
  assign dataGroup_lo_hi_802 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_803;
  assign dataGroup_lo_hi_803 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_804;
  assign dataGroup_lo_hi_804 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_805;
  assign dataGroup_lo_hi_805 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_806;
  assign dataGroup_lo_hi_806 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_807;
  assign dataGroup_lo_hi_807 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_808;
  assign dataGroup_lo_hi_808 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_809;
  assign dataGroup_lo_hi_809 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_810;
  assign dataGroup_lo_hi_810 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_811;
  assign dataGroup_lo_hi_811 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_812;
  assign dataGroup_lo_hi_812 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_813;
  assign dataGroup_lo_hi_813 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_814;
  assign dataGroup_lo_hi_814 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_815;
  assign dataGroup_lo_hi_815 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_816;
  assign dataGroup_lo_hi_816 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_817;
  assign dataGroup_lo_hi_817 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_818;
  assign dataGroup_lo_hi_818 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_819;
  assign dataGroup_lo_hi_819 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_820;
  assign dataGroup_lo_hi_820 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_821;
  assign dataGroup_lo_hi_821 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_822;
  assign dataGroup_lo_hi_822 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_823;
  assign dataGroup_lo_hi_823 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_824;
  assign dataGroup_lo_hi_824 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_825;
  assign dataGroup_lo_hi_825 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_826;
  assign dataGroup_lo_hi_826 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_827;
  assign dataGroup_lo_hi_827 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_828;
  assign dataGroup_lo_hi_828 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_829;
  assign dataGroup_lo_hi_829 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_830;
  assign dataGroup_lo_hi_830 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_831;
  assign dataGroup_lo_hi_831 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_832;
  assign dataGroup_lo_hi_832 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_833;
  assign dataGroup_lo_hi_833 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_834;
  assign dataGroup_lo_hi_834 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_835;
  assign dataGroup_lo_hi_835 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_836;
  assign dataGroup_lo_hi_836 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_837;
  assign dataGroup_lo_hi_837 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_838;
  assign dataGroup_lo_hi_838 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_839;
  assign dataGroup_lo_hi_839 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_840;
  assign dataGroup_lo_hi_840 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_841;
  assign dataGroup_lo_hi_841 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_842;
  assign dataGroup_lo_hi_842 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_843;
  assign dataGroup_lo_hi_843 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_844;
  assign dataGroup_lo_hi_844 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_845;
  assign dataGroup_lo_hi_845 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_846;
  assign dataGroup_lo_hi_846 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_847;
  assign dataGroup_lo_hi_847 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_848;
  assign dataGroup_lo_hi_848 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_849;
  assign dataGroup_lo_hi_849 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_850;
  assign dataGroup_lo_hi_850 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_851;
  assign dataGroup_lo_hi_851 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_852;
  assign dataGroup_lo_hi_852 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_853;
  assign dataGroup_lo_hi_853 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_854;
  assign dataGroup_lo_hi_854 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_855;
  assign dataGroup_lo_hi_855 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_856;
  assign dataGroup_lo_hi_856 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_857;
  assign dataGroup_lo_hi_857 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_858;
  assign dataGroup_lo_hi_858 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_859;
  assign dataGroup_lo_hi_859 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_860;
  assign dataGroup_lo_hi_860 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_861;
  assign dataGroup_lo_hi_861 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_862;
  assign dataGroup_lo_hi_862 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_863;
  assign dataGroup_lo_hi_863 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_864;
  assign dataGroup_lo_hi_864 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_865;
  assign dataGroup_lo_hi_865 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_866;
  assign dataGroup_lo_hi_866 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_867;
  assign dataGroup_lo_hi_867 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_868;
  assign dataGroup_lo_hi_868 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_869;
  assign dataGroup_lo_hi_869 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_870;
  assign dataGroup_lo_hi_870 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_871;
  assign dataGroup_lo_hi_871 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_872;
  assign dataGroup_lo_hi_872 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_873;
  assign dataGroup_lo_hi_873 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_874;
  assign dataGroup_lo_hi_874 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_875;
  assign dataGroup_lo_hi_875 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_876;
  assign dataGroup_lo_hi_876 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_877;
  assign dataGroup_lo_hi_877 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_878;
  assign dataGroup_lo_hi_878 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_879;
  assign dataGroup_lo_hi_879 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_880;
  assign dataGroup_lo_hi_880 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_881;
  assign dataGroup_lo_hi_881 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_882;
  assign dataGroup_lo_hi_882 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_883;
  assign dataGroup_lo_hi_883 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_884;
  assign dataGroup_lo_hi_884 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_885;
  assign dataGroup_lo_hi_885 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_886;
  assign dataGroup_lo_hi_886 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_887;
  assign dataGroup_lo_hi_887 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_888;
  assign dataGroup_lo_hi_888 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_889;
  assign dataGroup_lo_hi_889 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_890;
  assign dataGroup_lo_hi_890 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_891;
  assign dataGroup_lo_hi_891 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_892;
  assign dataGroup_lo_hi_892 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_893;
  assign dataGroup_lo_hi_893 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_894;
  assign dataGroup_lo_hi_894 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_895;
  assign dataGroup_lo_hi_895 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_896;
  assign dataGroup_lo_hi_896 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_897;
  assign dataGroup_lo_hi_897 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_898;
  assign dataGroup_lo_hi_898 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_899;
  assign dataGroup_lo_hi_899 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_900;
  assign dataGroup_lo_hi_900 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_901;
  assign dataGroup_lo_hi_901 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_902;
  assign dataGroup_lo_hi_902 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_903;
  assign dataGroup_lo_hi_903 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_904;
  assign dataGroup_lo_hi_904 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_905;
  assign dataGroup_lo_hi_905 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_906;
  assign dataGroup_lo_hi_906 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_907;
  assign dataGroup_lo_hi_907 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_908;
  assign dataGroup_lo_hi_908 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_909;
  assign dataGroup_lo_hi_909 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_910;
  assign dataGroup_lo_hi_910 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_911;
  assign dataGroup_lo_hi_911 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_912;
  assign dataGroup_lo_hi_912 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_913;
  assign dataGroup_lo_hi_913 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_914;
  assign dataGroup_lo_hi_914 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_915;
  assign dataGroup_lo_hi_915 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_916;
  assign dataGroup_lo_hi_916 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_917;
  assign dataGroup_lo_hi_917 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_918;
  assign dataGroup_lo_hi_918 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_919;
  assign dataGroup_lo_hi_919 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_920;
  assign dataGroup_lo_hi_920 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_921;
  assign dataGroup_lo_hi_921 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_922;
  assign dataGroup_lo_hi_922 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_923;
  assign dataGroup_lo_hi_923 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_924;
  assign dataGroup_lo_hi_924 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_925;
  assign dataGroup_lo_hi_925 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_926;
  assign dataGroup_lo_hi_926 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_927;
  assign dataGroup_lo_hi_927 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_928;
  assign dataGroup_lo_hi_928 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_929;
  assign dataGroup_lo_hi_929 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_930;
  assign dataGroup_lo_hi_930 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_931;
  assign dataGroup_lo_hi_931 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_932;
  assign dataGroup_lo_hi_932 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_933;
  assign dataGroup_lo_hi_933 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_934;
  assign dataGroup_lo_hi_934 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_935;
  assign dataGroup_lo_hi_935 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_936;
  assign dataGroup_lo_hi_936 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_937;
  assign dataGroup_lo_hi_937 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_938;
  assign dataGroup_lo_hi_938 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_939;
  assign dataGroup_lo_hi_939 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_940;
  assign dataGroup_lo_hi_940 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_941;
  assign dataGroup_lo_hi_941 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_942;
  assign dataGroup_lo_hi_942 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_943;
  assign dataGroup_lo_hi_943 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_944;
  assign dataGroup_lo_hi_944 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_945;
  assign dataGroup_lo_hi_945 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_946;
  assign dataGroup_lo_hi_946 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_947;
  assign dataGroup_lo_hi_947 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_948;
  assign dataGroup_lo_hi_948 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_949;
  assign dataGroup_lo_hi_949 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_950;
  assign dataGroup_lo_hi_950 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_951;
  assign dataGroup_lo_hi_951 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_952;
  assign dataGroup_lo_hi_952 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_953;
  assign dataGroup_lo_hi_953 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_954;
  assign dataGroup_lo_hi_954 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_955;
  assign dataGroup_lo_hi_955 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_956;
  assign dataGroup_lo_hi_956 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_957;
  assign dataGroup_lo_hi_957 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_958;
  assign dataGroup_lo_hi_958 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_959;
  assign dataGroup_lo_hi_959 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_960;
  assign dataGroup_lo_hi_960 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_961;
  assign dataGroup_lo_hi_961 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_962;
  assign dataGroup_lo_hi_962 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_963;
  assign dataGroup_lo_hi_963 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_964;
  assign dataGroup_lo_hi_964 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_965;
  assign dataGroup_lo_hi_965 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_966;
  assign dataGroup_lo_hi_966 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_967;
  assign dataGroup_lo_hi_967 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_968;
  assign dataGroup_lo_hi_968 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_969;
  assign dataGroup_lo_hi_969 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_970;
  assign dataGroup_lo_hi_970 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_971;
  assign dataGroup_lo_hi_971 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_972;
  assign dataGroup_lo_hi_972 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_973;
  assign dataGroup_lo_hi_973 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_974;
  assign dataGroup_lo_hi_974 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_975;
  assign dataGroup_lo_hi_975 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_976;
  assign dataGroup_lo_hi_976 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_977;
  assign dataGroup_lo_hi_977 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_978;
  assign dataGroup_lo_hi_978 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_979;
  assign dataGroup_lo_hi_979 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_980;
  assign dataGroup_lo_hi_980 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_981;
  assign dataGroup_lo_hi_981 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_982;
  assign dataGroup_lo_hi_982 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_983;
  assign dataGroup_lo_hi_983 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_984;
  assign dataGroup_lo_hi_984 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_985;
  assign dataGroup_lo_hi_985 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_986;
  assign dataGroup_lo_hi_986 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_987;
  assign dataGroup_lo_hi_987 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_988;
  assign dataGroup_lo_hi_988 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_989;
  assign dataGroup_lo_hi_989 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_990;
  assign dataGroup_lo_hi_990 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_991;
  assign dataGroup_lo_hi_991 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_992;
  assign dataGroup_lo_hi_992 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_993;
  assign dataGroup_lo_hi_993 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_994;
  assign dataGroup_lo_hi_994 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_995;
  assign dataGroup_lo_hi_995 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_996;
  assign dataGroup_lo_hi_996 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_997;
  assign dataGroup_lo_hi_997 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_998;
  assign dataGroup_lo_hi_998 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_999;
  assign dataGroup_lo_hi_999 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1000;
  assign dataGroup_lo_hi_1000 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1001;
  assign dataGroup_lo_hi_1001 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1002;
  assign dataGroup_lo_hi_1002 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1003;
  assign dataGroup_lo_hi_1003 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1004;
  assign dataGroup_lo_hi_1004 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1005;
  assign dataGroup_lo_hi_1005 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1006;
  assign dataGroup_lo_hi_1006 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1007;
  assign dataGroup_lo_hi_1007 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1008;
  assign dataGroup_lo_hi_1008 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1009;
  assign dataGroup_lo_hi_1009 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1010;
  assign dataGroup_lo_hi_1010 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1011;
  assign dataGroup_lo_hi_1011 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1012;
  assign dataGroup_lo_hi_1012 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1013;
  assign dataGroup_lo_hi_1013 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1014;
  assign dataGroup_lo_hi_1014 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1015;
  assign dataGroup_lo_hi_1015 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1016;
  assign dataGroup_lo_hi_1016 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1017;
  assign dataGroup_lo_hi_1017 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1018;
  assign dataGroup_lo_hi_1018 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1019;
  assign dataGroup_lo_hi_1019 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1020;
  assign dataGroup_lo_hi_1020 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1021;
  assign dataGroup_lo_hi_1021 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1022;
  assign dataGroup_lo_hi_1022 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1023;
  assign dataGroup_lo_hi_1023 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1024;
  assign dataGroup_lo_hi_1024 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1025;
  assign dataGroup_lo_hi_1025 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1026;
  assign dataGroup_lo_hi_1026 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1027;
  assign dataGroup_lo_hi_1027 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1028;
  assign dataGroup_lo_hi_1028 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1029;
  assign dataGroup_lo_hi_1029 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1030;
  assign dataGroup_lo_hi_1030 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1031;
  assign dataGroup_lo_hi_1031 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1032;
  assign dataGroup_lo_hi_1032 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1033;
  assign dataGroup_lo_hi_1033 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1034;
  assign dataGroup_lo_hi_1034 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1035;
  assign dataGroup_lo_hi_1035 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1036;
  assign dataGroup_lo_hi_1036 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1037;
  assign dataGroup_lo_hi_1037 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1038;
  assign dataGroup_lo_hi_1038 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1039;
  assign dataGroup_lo_hi_1039 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1040;
  assign dataGroup_lo_hi_1040 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1041;
  assign dataGroup_lo_hi_1041 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1042;
  assign dataGroup_lo_hi_1042 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1043;
  assign dataGroup_lo_hi_1043 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1044;
  assign dataGroup_lo_hi_1044 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1045;
  assign dataGroup_lo_hi_1045 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1046;
  assign dataGroup_lo_hi_1046 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1047;
  assign dataGroup_lo_hi_1047 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1048;
  assign dataGroup_lo_hi_1048 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1049;
  assign dataGroup_lo_hi_1049 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1050;
  assign dataGroup_lo_hi_1050 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1051;
  assign dataGroup_lo_hi_1051 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1052;
  assign dataGroup_lo_hi_1052 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1053;
  assign dataGroup_lo_hi_1053 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1054;
  assign dataGroup_lo_hi_1054 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1055;
  assign dataGroup_lo_hi_1055 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1056;
  assign dataGroup_lo_hi_1056 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1057;
  assign dataGroup_lo_hi_1057 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1058;
  assign dataGroup_lo_hi_1058 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1059;
  assign dataGroup_lo_hi_1059 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1060;
  assign dataGroup_lo_hi_1060 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1061;
  assign dataGroup_lo_hi_1061 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1062;
  assign dataGroup_lo_hi_1062 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1063;
  assign dataGroup_lo_hi_1063 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1064;
  assign dataGroup_lo_hi_1064 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1065;
  assign dataGroup_lo_hi_1065 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1066;
  assign dataGroup_lo_hi_1066 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1067;
  assign dataGroup_lo_hi_1067 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1068;
  assign dataGroup_lo_hi_1068 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1069;
  assign dataGroup_lo_hi_1069 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1070;
  assign dataGroup_lo_hi_1070 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1071;
  assign dataGroup_lo_hi_1071 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1072;
  assign dataGroup_lo_hi_1072 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1073;
  assign dataGroup_lo_hi_1073 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1074;
  assign dataGroup_lo_hi_1074 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1075;
  assign dataGroup_lo_hi_1075 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1076;
  assign dataGroup_lo_hi_1076 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1077;
  assign dataGroup_lo_hi_1077 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1078;
  assign dataGroup_lo_hi_1078 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1079;
  assign dataGroup_lo_hi_1079 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1080;
  assign dataGroup_lo_hi_1080 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1081;
  assign dataGroup_lo_hi_1081 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1082;
  assign dataGroup_lo_hi_1082 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1083;
  assign dataGroup_lo_hi_1083 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1084;
  assign dataGroup_lo_hi_1084 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1085;
  assign dataGroup_lo_hi_1085 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1086;
  assign dataGroup_lo_hi_1086 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1087;
  assign dataGroup_lo_hi_1087 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1088;
  assign dataGroup_lo_hi_1088 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1089;
  assign dataGroup_lo_hi_1089 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1090;
  assign dataGroup_lo_hi_1090 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1091;
  assign dataGroup_lo_hi_1091 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1092;
  assign dataGroup_lo_hi_1092 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1093;
  assign dataGroup_lo_hi_1093 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1094;
  assign dataGroup_lo_hi_1094 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1095;
  assign dataGroup_lo_hi_1095 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1096;
  assign dataGroup_lo_hi_1096 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1097;
  assign dataGroup_lo_hi_1097 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1098;
  assign dataGroup_lo_hi_1098 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1099;
  assign dataGroup_lo_hi_1099 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1100;
  assign dataGroup_lo_hi_1100 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1101;
  assign dataGroup_lo_hi_1101 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1102;
  assign dataGroup_lo_hi_1102 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1103;
  assign dataGroup_lo_hi_1103 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1104;
  assign dataGroup_lo_hi_1104 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1105;
  assign dataGroup_lo_hi_1105 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1106;
  assign dataGroup_lo_hi_1106 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1107;
  assign dataGroup_lo_hi_1107 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1108;
  assign dataGroup_lo_hi_1108 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1109;
  assign dataGroup_lo_hi_1109 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1110;
  assign dataGroup_lo_hi_1110 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1111;
  assign dataGroup_lo_hi_1111 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1112;
  assign dataGroup_lo_hi_1112 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1113;
  assign dataGroup_lo_hi_1113 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1114;
  assign dataGroup_lo_hi_1114 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1115;
  assign dataGroup_lo_hi_1115 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1116;
  assign dataGroup_lo_hi_1116 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1117;
  assign dataGroup_lo_hi_1117 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1118;
  assign dataGroup_lo_hi_1118 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1119;
  assign dataGroup_lo_hi_1119 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1120;
  assign dataGroup_lo_hi_1120 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1121;
  assign dataGroup_lo_hi_1121 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1122;
  assign dataGroup_lo_hi_1122 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1123;
  assign dataGroup_lo_hi_1123 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1124;
  assign dataGroup_lo_hi_1124 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1125;
  assign dataGroup_lo_hi_1125 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1126;
  assign dataGroup_lo_hi_1126 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1127;
  assign dataGroup_lo_hi_1127 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1128;
  assign dataGroup_lo_hi_1128 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1129;
  assign dataGroup_lo_hi_1129 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1130;
  assign dataGroup_lo_hi_1130 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1131;
  assign dataGroup_lo_hi_1131 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1132;
  assign dataGroup_lo_hi_1132 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1133;
  assign dataGroup_lo_hi_1133 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1134;
  assign dataGroup_lo_hi_1134 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1135;
  assign dataGroup_lo_hi_1135 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1136;
  assign dataGroup_lo_hi_1136 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1137;
  assign dataGroup_lo_hi_1137 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1138;
  assign dataGroup_lo_hi_1138 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1139;
  assign dataGroup_lo_hi_1139 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1140;
  assign dataGroup_lo_hi_1140 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1141;
  assign dataGroup_lo_hi_1141 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1142;
  assign dataGroup_lo_hi_1142 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1143;
  assign dataGroup_lo_hi_1143 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1144;
  assign dataGroup_lo_hi_1144 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1145;
  assign dataGroup_lo_hi_1145 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1146;
  assign dataGroup_lo_hi_1146 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1147;
  assign dataGroup_lo_hi_1147 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1148;
  assign dataGroup_lo_hi_1148 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1149;
  assign dataGroup_lo_hi_1149 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1150;
  assign dataGroup_lo_hi_1150 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1151;
  assign dataGroup_lo_hi_1151 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1152;
  assign dataGroup_lo_hi_1152 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1153;
  assign dataGroup_lo_hi_1153 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1154;
  assign dataGroup_lo_hi_1154 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1155;
  assign dataGroup_lo_hi_1155 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1156;
  assign dataGroup_lo_hi_1156 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1157;
  assign dataGroup_lo_hi_1157 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1158;
  assign dataGroup_lo_hi_1158 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1159;
  assign dataGroup_lo_hi_1159 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1160;
  assign dataGroup_lo_hi_1160 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1161;
  assign dataGroup_lo_hi_1161 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1162;
  assign dataGroup_lo_hi_1162 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1163;
  assign dataGroup_lo_hi_1163 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1164;
  assign dataGroup_lo_hi_1164 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1165;
  assign dataGroup_lo_hi_1165 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1166;
  assign dataGroup_lo_hi_1166 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1167;
  assign dataGroup_lo_hi_1167 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1168;
  assign dataGroup_lo_hi_1168 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1169;
  assign dataGroup_lo_hi_1169 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1170;
  assign dataGroup_lo_hi_1170 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1171;
  assign dataGroup_lo_hi_1171 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1172;
  assign dataGroup_lo_hi_1172 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1173;
  assign dataGroup_lo_hi_1173 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1174;
  assign dataGroup_lo_hi_1174 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1175;
  assign dataGroup_lo_hi_1175 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1176;
  assign dataGroup_lo_hi_1176 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1177;
  assign dataGroup_lo_hi_1177 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1178;
  assign dataGroup_lo_hi_1178 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1179;
  assign dataGroup_lo_hi_1179 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1180;
  assign dataGroup_lo_hi_1180 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1181;
  assign dataGroup_lo_hi_1181 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1182;
  assign dataGroup_lo_hi_1182 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1183;
  assign dataGroup_lo_hi_1183 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1184;
  assign dataGroup_lo_hi_1184 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1185;
  assign dataGroup_lo_hi_1185 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1186;
  assign dataGroup_lo_hi_1186 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1187;
  assign dataGroup_lo_hi_1187 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1188;
  assign dataGroup_lo_hi_1188 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1189;
  assign dataGroup_lo_hi_1189 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1190;
  assign dataGroup_lo_hi_1190 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1191;
  assign dataGroup_lo_hi_1191 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1192;
  assign dataGroup_lo_hi_1192 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1193;
  assign dataGroup_lo_hi_1193 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1194;
  assign dataGroup_lo_hi_1194 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1195;
  assign dataGroup_lo_hi_1195 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1196;
  assign dataGroup_lo_hi_1196 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1197;
  assign dataGroup_lo_hi_1197 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1198;
  assign dataGroup_lo_hi_1198 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1199;
  assign dataGroup_lo_hi_1199 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1200;
  assign dataGroup_lo_hi_1200 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1201;
  assign dataGroup_lo_hi_1201 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1202;
  assign dataGroup_lo_hi_1202 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1203;
  assign dataGroup_lo_hi_1203 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1204;
  assign dataGroup_lo_hi_1204 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1205;
  assign dataGroup_lo_hi_1205 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1206;
  assign dataGroup_lo_hi_1206 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1207;
  assign dataGroup_lo_hi_1207 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1208;
  assign dataGroup_lo_hi_1208 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1209;
  assign dataGroup_lo_hi_1209 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1210;
  assign dataGroup_lo_hi_1210 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1211;
  assign dataGroup_lo_hi_1211 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1212;
  assign dataGroup_lo_hi_1212 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1213;
  assign dataGroup_lo_hi_1213 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1214;
  assign dataGroup_lo_hi_1214 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1215;
  assign dataGroup_lo_hi_1215 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1216;
  assign dataGroup_lo_hi_1216 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1217;
  assign dataGroup_lo_hi_1217 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1218;
  assign dataGroup_lo_hi_1218 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1219;
  assign dataGroup_lo_hi_1219 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1220;
  assign dataGroup_lo_hi_1220 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1221;
  assign dataGroup_lo_hi_1221 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1222;
  assign dataGroup_lo_hi_1222 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1223;
  assign dataGroup_lo_hi_1223 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1224;
  assign dataGroup_lo_hi_1224 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1225;
  assign dataGroup_lo_hi_1225 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1226;
  assign dataGroup_lo_hi_1226 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1227;
  assign dataGroup_lo_hi_1227 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1228;
  assign dataGroup_lo_hi_1228 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1229;
  assign dataGroup_lo_hi_1229 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1230;
  assign dataGroup_lo_hi_1230 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1231;
  assign dataGroup_lo_hi_1231 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1232;
  assign dataGroup_lo_hi_1232 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1233;
  assign dataGroup_lo_hi_1233 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1234;
  assign dataGroup_lo_hi_1234 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1235;
  assign dataGroup_lo_hi_1235 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1236;
  assign dataGroup_lo_hi_1236 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1237;
  assign dataGroup_lo_hi_1237 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1238;
  assign dataGroup_lo_hi_1238 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1239;
  assign dataGroup_lo_hi_1239 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1240;
  assign dataGroup_lo_hi_1240 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1241;
  assign dataGroup_lo_hi_1241 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1242;
  assign dataGroup_lo_hi_1242 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1243;
  assign dataGroup_lo_hi_1243 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1244;
  assign dataGroup_lo_hi_1244 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1245;
  assign dataGroup_lo_hi_1245 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1246;
  assign dataGroup_lo_hi_1246 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1247;
  assign dataGroup_lo_hi_1247 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1248;
  assign dataGroup_lo_hi_1248 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1249;
  assign dataGroup_lo_hi_1249 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1250;
  assign dataGroup_lo_hi_1250 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1251;
  assign dataGroup_lo_hi_1251 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1252;
  assign dataGroup_lo_hi_1252 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1253;
  assign dataGroup_lo_hi_1253 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1254;
  assign dataGroup_lo_hi_1254 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1255;
  assign dataGroup_lo_hi_1255 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1256;
  assign dataGroup_lo_hi_1256 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1257;
  assign dataGroup_lo_hi_1257 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1258;
  assign dataGroup_lo_hi_1258 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1259;
  assign dataGroup_lo_hi_1259 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1260;
  assign dataGroup_lo_hi_1260 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1261;
  assign dataGroup_lo_hi_1261 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1262;
  assign dataGroup_lo_hi_1262 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1263;
  assign dataGroup_lo_hi_1263 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1264;
  assign dataGroup_lo_hi_1264 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1265;
  assign dataGroup_lo_hi_1265 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1266;
  assign dataGroup_lo_hi_1266 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1267;
  assign dataGroup_lo_hi_1267 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1268;
  assign dataGroup_lo_hi_1268 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1269;
  assign dataGroup_lo_hi_1269 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1270;
  assign dataGroup_lo_hi_1270 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1271;
  assign dataGroup_lo_hi_1271 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1272;
  assign dataGroup_lo_hi_1272 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1273;
  assign dataGroup_lo_hi_1273 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1274;
  assign dataGroup_lo_hi_1274 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1275;
  assign dataGroup_lo_hi_1275 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1276;
  assign dataGroup_lo_hi_1276 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1277;
  assign dataGroup_lo_hi_1277 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1278;
  assign dataGroup_lo_hi_1278 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1279;
  assign dataGroup_lo_hi_1279 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1280;
  assign dataGroup_lo_hi_1280 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1281;
  assign dataGroup_lo_hi_1281 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1282;
  assign dataGroup_lo_hi_1282 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1283;
  assign dataGroup_lo_hi_1283 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1284;
  assign dataGroup_lo_hi_1284 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1285;
  assign dataGroup_lo_hi_1285 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1286;
  assign dataGroup_lo_hi_1286 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1287;
  assign dataGroup_lo_hi_1287 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1288;
  assign dataGroup_lo_hi_1288 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1289;
  assign dataGroup_lo_hi_1289 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1290;
  assign dataGroup_lo_hi_1290 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1291;
  assign dataGroup_lo_hi_1291 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1292;
  assign dataGroup_lo_hi_1292 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1293;
  assign dataGroup_lo_hi_1293 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1294;
  assign dataGroup_lo_hi_1294 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1295;
  assign dataGroup_lo_hi_1295 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1296;
  assign dataGroup_lo_hi_1296 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1297;
  assign dataGroup_lo_hi_1297 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1298;
  assign dataGroup_lo_hi_1298 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1299;
  assign dataGroup_lo_hi_1299 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1300;
  assign dataGroup_lo_hi_1300 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1301;
  assign dataGroup_lo_hi_1301 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1302;
  assign dataGroup_lo_hi_1302 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1303;
  assign dataGroup_lo_hi_1303 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1304;
  assign dataGroup_lo_hi_1304 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1305;
  assign dataGroup_lo_hi_1305 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1306;
  assign dataGroup_lo_hi_1306 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1307;
  assign dataGroup_lo_hi_1307 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1308;
  assign dataGroup_lo_hi_1308 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1309;
  assign dataGroup_lo_hi_1309 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1310;
  assign dataGroup_lo_hi_1310 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1311;
  assign dataGroup_lo_hi_1311 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1312;
  assign dataGroup_lo_hi_1312 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1313;
  assign dataGroup_lo_hi_1313 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1314;
  assign dataGroup_lo_hi_1314 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1315;
  assign dataGroup_lo_hi_1315 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1316;
  assign dataGroup_lo_hi_1316 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1317;
  assign dataGroup_lo_hi_1317 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1318;
  assign dataGroup_lo_hi_1318 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1319;
  assign dataGroup_lo_hi_1319 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1320;
  assign dataGroup_lo_hi_1320 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1321;
  assign dataGroup_lo_hi_1321 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1322;
  assign dataGroup_lo_hi_1322 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1323;
  assign dataGroup_lo_hi_1323 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1324;
  assign dataGroup_lo_hi_1324 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1325;
  assign dataGroup_lo_hi_1325 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1326;
  assign dataGroup_lo_hi_1326 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1327;
  assign dataGroup_lo_hi_1327 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1328;
  assign dataGroup_lo_hi_1328 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1329;
  assign dataGroup_lo_hi_1329 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1330;
  assign dataGroup_lo_hi_1330 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1331;
  assign dataGroup_lo_hi_1331 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1332;
  assign dataGroup_lo_hi_1332 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1333;
  assign dataGroup_lo_hi_1333 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1334;
  assign dataGroup_lo_hi_1334 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1335;
  assign dataGroup_lo_hi_1335 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1336;
  assign dataGroup_lo_hi_1336 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1337;
  assign dataGroup_lo_hi_1337 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1338;
  assign dataGroup_lo_hi_1338 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1339;
  assign dataGroup_lo_hi_1339 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1340;
  assign dataGroup_lo_hi_1340 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1341;
  assign dataGroup_lo_hi_1341 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1342;
  assign dataGroup_lo_hi_1342 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1343;
  assign dataGroup_lo_hi_1343 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1344;
  assign dataGroup_lo_hi_1344 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1345;
  assign dataGroup_lo_hi_1345 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1346;
  assign dataGroup_lo_hi_1346 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1347;
  assign dataGroup_lo_hi_1347 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1348;
  assign dataGroup_lo_hi_1348 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1349;
  assign dataGroup_lo_hi_1349 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1350;
  assign dataGroup_lo_hi_1350 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1351;
  assign dataGroup_lo_hi_1351 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1352;
  assign dataGroup_lo_hi_1352 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1353;
  assign dataGroup_lo_hi_1353 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1354;
  assign dataGroup_lo_hi_1354 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1355;
  assign dataGroup_lo_hi_1355 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1356;
  assign dataGroup_lo_hi_1356 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1357;
  assign dataGroup_lo_hi_1357 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1358;
  assign dataGroup_lo_hi_1358 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1359;
  assign dataGroup_lo_hi_1359 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1360;
  assign dataGroup_lo_hi_1360 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1361;
  assign dataGroup_lo_hi_1361 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1362;
  assign dataGroup_lo_hi_1362 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1363;
  assign dataGroup_lo_hi_1363 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1364;
  assign dataGroup_lo_hi_1364 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1365;
  assign dataGroup_lo_hi_1365 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1366;
  assign dataGroup_lo_hi_1366 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1367;
  assign dataGroup_lo_hi_1367 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1368;
  assign dataGroup_lo_hi_1368 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1369;
  assign dataGroup_lo_hi_1369 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1370;
  assign dataGroup_lo_hi_1370 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1371;
  assign dataGroup_lo_hi_1371 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1372;
  assign dataGroup_lo_hi_1372 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1373;
  assign dataGroup_lo_hi_1373 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1374;
  assign dataGroup_lo_hi_1374 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1375;
  assign dataGroup_lo_hi_1375 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1376;
  assign dataGroup_lo_hi_1376 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1377;
  assign dataGroup_lo_hi_1377 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1378;
  assign dataGroup_lo_hi_1378 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1379;
  assign dataGroup_lo_hi_1379 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1380;
  assign dataGroup_lo_hi_1380 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1381;
  assign dataGroup_lo_hi_1381 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1382;
  assign dataGroup_lo_hi_1382 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1383;
  assign dataGroup_lo_hi_1383 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1384;
  assign dataGroup_lo_hi_1384 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1385;
  assign dataGroup_lo_hi_1385 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1386;
  assign dataGroup_lo_hi_1386 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1387;
  assign dataGroup_lo_hi_1387 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1388;
  assign dataGroup_lo_hi_1388 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1389;
  assign dataGroup_lo_hi_1389 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1390;
  assign dataGroup_lo_hi_1390 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1391;
  assign dataGroup_lo_hi_1391 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1392;
  assign dataGroup_lo_hi_1392 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1393;
  assign dataGroup_lo_hi_1393 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1394;
  assign dataGroup_lo_hi_1394 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1395;
  assign dataGroup_lo_hi_1395 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1396;
  assign dataGroup_lo_hi_1396 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1397;
  assign dataGroup_lo_hi_1397 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1398;
  assign dataGroup_lo_hi_1398 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1399;
  assign dataGroup_lo_hi_1399 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1400;
  assign dataGroup_lo_hi_1400 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1401;
  assign dataGroup_lo_hi_1401 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1402;
  assign dataGroup_lo_hi_1402 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1403;
  assign dataGroup_lo_hi_1403 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1404;
  assign dataGroup_lo_hi_1404 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1405;
  assign dataGroup_lo_hi_1405 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1406;
  assign dataGroup_lo_hi_1406 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1407;
  assign dataGroup_lo_hi_1407 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1408;
  assign dataGroup_lo_hi_1408 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1409;
  assign dataGroup_lo_hi_1409 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1410;
  assign dataGroup_lo_hi_1410 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1411;
  assign dataGroup_lo_hi_1411 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1412;
  assign dataGroup_lo_hi_1412 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1413;
  assign dataGroup_lo_hi_1413 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1414;
  assign dataGroup_lo_hi_1414 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1415;
  assign dataGroup_lo_hi_1415 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1416;
  assign dataGroup_lo_hi_1416 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1417;
  assign dataGroup_lo_hi_1417 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1418;
  assign dataGroup_lo_hi_1418 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1419;
  assign dataGroup_lo_hi_1419 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1420;
  assign dataGroup_lo_hi_1420 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1421;
  assign dataGroup_lo_hi_1421 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1422;
  assign dataGroup_lo_hi_1422 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1423;
  assign dataGroup_lo_hi_1423 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1424;
  assign dataGroup_lo_hi_1424 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1425;
  assign dataGroup_lo_hi_1425 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1426;
  assign dataGroup_lo_hi_1426 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1427;
  assign dataGroup_lo_hi_1427 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1428;
  assign dataGroup_lo_hi_1428 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1429;
  assign dataGroup_lo_hi_1429 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1430;
  assign dataGroup_lo_hi_1430 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1431;
  assign dataGroup_lo_hi_1431 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1432;
  assign dataGroup_lo_hi_1432 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1433;
  assign dataGroup_lo_hi_1433 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1434;
  assign dataGroup_lo_hi_1434 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1435;
  assign dataGroup_lo_hi_1435 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1436;
  assign dataGroup_lo_hi_1436 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1437;
  assign dataGroup_lo_hi_1437 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1438;
  assign dataGroup_lo_hi_1438 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1439;
  assign dataGroup_lo_hi_1439 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1440;
  assign dataGroup_lo_hi_1440 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1441;
  assign dataGroup_lo_hi_1441 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1442;
  assign dataGroup_lo_hi_1442 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1443;
  assign dataGroup_lo_hi_1443 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1444;
  assign dataGroup_lo_hi_1444 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1445;
  assign dataGroup_lo_hi_1445 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1446;
  assign dataGroup_lo_hi_1446 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1447;
  assign dataGroup_lo_hi_1447 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1448;
  assign dataGroup_lo_hi_1448 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1449;
  assign dataGroup_lo_hi_1449 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1450;
  assign dataGroup_lo_hi_1450 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1451;
  assign dataGroup_lo_hi_1451 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1452;
  assign dataGroup_lo_hi_1452 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1453;
  assign dataGroup_lo_hi_1453 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1454;
  assign dataGroup_lo_hi_1454 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1455;
  assign dataGroup_lo_hi_1455 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1456;
  assign dataGroup_lo_hi_1456 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1457;
  assign dataGroup_lo_hi_1457 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1458;
  assign dataGroup_lo_hi_1458 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1459;
  assign dataGroup_lo_hi_1459 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1460;
  assign dataGroup_lo_hi_1460 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1461;
  assign dataGroup_lo_hi_1461 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1462;
  assign dataGroup_lo_hi_1462 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1463;
  assign dataGroup_lo_hi_1463 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1464;
  assign dataGroup_lo_hi_1464 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1465;
  assign dataGroup_lo_hi_1465 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1466;
  assign dataGroup_lo_hi_1466 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1467;
  assign dataGroup_lo_hi_1467 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1468;
  assign dataGroup_lo_hi_1468 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1469;
  assign dataGroup_lo_hi_1469 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1470;
  assign dataGroup_lo_hi_1470 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1471;
  assign dataGroup_lo_hi_1471 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1472;
  assign dataGroup_lo_hi_1472 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1473;
  assign dataGroup_lo_hi_1473 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1474;
  assign dataGroup_lo_hi_1474 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1475;
  assign dataGroup_lo_hi_1475 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1476;
  assign dataGroup_lo_hi_1476 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1477;
  assign dataGroup_lo_hi_1477 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1478;
  assign dataGroup_lo_hi_1478 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1479;
  assign dataGroup_lo_hi_1479 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1480;
  assign dataGroup_lo_hi_1480 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1481;
  assign dataGroup_lo_hi_1481 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1482;
  assign dataGroup_lo_hi_1482 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1483;
  assign dataGroup_lo_hi_1483 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1484;
  assign dataGroup_lo_hi_1484 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1485;
  assign dataGroup_lo_hi_1485 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1486;
  assign dataGroup_lo_hi_1486 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1487;
  assign dataGroup_lo_hi_1487 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1488;
  assign dataGroup_lo_hi_1488 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1489;
  assign dataGroup_lo_hi_1489 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1490;
  assign dataGroup_lo_hi_1490 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1491;
  assign dataGroup_lo_hi_1491 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1492;
  assign dataGroup_lo_hi_1492 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1493;
  assign dataGroup_lo_hi_1493 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1494;
  assign dataGroup_lo_hi_1494 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1495;
  assign dataGroup_lo_hi_1495 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1496;
  assign dataGroup_lo_hi_1496 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1497;
  assign dataGroup_lo_hi_1497 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1498;
  assign dataGroup_lo_hi_1498 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1499;
  assign dataGroup_lo_hi_1499 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1500;
  assign dataGroup_lo_hi_1500 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1501;
  assign dataGroup_lo_hi_1501 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1502;
  assign dataGroup_lo_hi_1502 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1503;
  assign dataGroup_lo_hi_1503 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1504;
  assign dataGroup_lo_hi_1504 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1505;
  assign dataGroup_lo_hi_1505 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1506;
  assign dataGroup_lo_hi_1506 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1507;
  assign dataGroup_lo_hi_1507 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1508;
  assign dataGroup_lo_hi_1508 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1509;
  assign dataGroup_lo_hi_1509 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1510;
  assign dataGroup_lo_hi_1510 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1511;
  assign dataGroup_lo_hi_1511 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1512;
  assign dataGroup_lo_hi_1512 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1513;
  assign dataGroup_lo_hi_1513 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1514;
  assign dataGroup_lo_hi_1514 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1515;
  assign dataGroup_lo_hi_1515 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1516;
  assign dataGroup_lo_hi_1516 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1517;
  assign dataGroup_lo_hi_1517 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1518;
  assign dataGroup_lo_hi_1518 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1519;
  assign dataGroup_lo_hi_1519 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1520;
  assign dataGroup_lo_hi_1520 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1521;
  assign dataGroup_lo_hi_1521 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1522;
  assign dataGroup_lo_hi_1522 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1523;
  assign dataGroup_lo_hi_1523 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1524;
  assign dataGroup_lo_hi_1524 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1525;
  assign dataGroup_lo_hi_1525 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1526;
  assign dataGroup_lo_hi_1526 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1527;
  assign dataGroup_lo_hi_1527 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1528;
  assign dataGroup_lo_hi_1528 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1529;
  assign dataGroup_lo_hi_1529 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1530;
  assign dataGroup_lo_hi_1530 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1531;
  assign dataGroup_lo_hi_1531 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1532;
  assign dataGroup_lo_hi_1532 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1533;
  assign dataGroup_lo_hi_1533 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1534;
  assign dataGroup_lo_hi_1534 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1535;
  assign dataGroup_lo_hi_1535 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1536;
  assign dataGroup_lo_hi_1536 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1537;
  assign dataGroup_lo_hi_1537 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1538;
  assign dataGroup_lo_hi_1538 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1539;
  assign dataGroup_lo_hi_1539 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1540;
  assign dataGroup_lo_hi_1540 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1541;
  assign dataGroup_lo_hi_1541 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1542;
  assign dataGroup_lo_hi_1542 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1543;
  assign dataGroup_lo_hi_1543 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1544;
  assign dataGroup_lo_hi_1544 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1545;
  assign dataGroup_lo_hi_1545 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1546;
  assign dataGroup_lo_hi_1546 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1547;
  assign dataGroup_lo_hi_1547 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1548;
  assign dataGroup_lo_hi_1548 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1549;
  assign dataGroup_lo_hi_1549 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1550;
  assign dataGroup_lo_hi_1550 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1551;
  assign dataGroup_lo_hi_1551 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1552;
  assign dataGroup_lo_hi_1552 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1553;
  assign dataGroup_lo_hi_1553 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1554;
  assign dataGroup_lo_hi_1554 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1555;
  assign dataGroup_lo_hi_1555 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1556;
  assign dataGroup_lo_hi_1556 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1557;
  assign dataGroup_lo_hi_1557 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1558;
  assign dataGroup_lo_hi_1558 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1559;
  assign dataGroup_lo_hi_1559 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1560;
  assign dataGroup_lo_hi_1560 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1561;
  assign dataGroup_lo_hi_1561 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1562;
  assign dataGroup_lo_hi_1562 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1563;
  assign dataGroup_lo_hi_1563 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1564;
  assign dataGroup_lo_hi_1564 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1565;
  assign dataGroup_lo_hi_1565 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1566;
  assign dataGroup_lo_hi_1566 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1567;
  assign dataGroup_lo_hi_1567 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1568;
  assign dataGroup_lo_hi_1568 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1569;
  assign dataGroup_lo_hi_1569 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1570;
  assign dataGroup_lo_hi_1570 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1571;
  assign dataGroup_lo_hi_1571 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1572;
  assign dataGroup_lo_hi_1572 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1573;
  assign dataGroup_lo_hi_1573 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1574;
  assign dataGroup_lo_hi_1574 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1575;
  assign dataGroup_lo_hi_1575 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1576;
  assign dataGroup_lo_hi_1576 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1577;
  assign dataGroup_lo_hi_1577 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1578;
  assign dataGroup_lo_hi_1578 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1579;
  assign dataGroup_lo_hi_1579 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1580;
  assign dataGroup_lo_hi_1580 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1581;
  assign dataGroup_lo_hi_1581 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1582;
  assign dataGroup_lo_hi_1582 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1583;
  assign dataGroup_lo_hi_1583 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1584;
  assign dataGroup_lo_hi_1584 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1585;
  assign dataGroup_lo_hi_1585 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1586;
  assign dataGroup_lo_hi_1586 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1587;
  assign dataGroup_lo_hi_1587 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1588;
  assign dataGroup_lo_hi_1588 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1589;
  assign dataGroup_lo_hi_1589 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1590;
  assign dataGroup_lo_hi_1590 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1591;
  assign dataGroup_lo_hi_1591 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1592;
  assign dataGroup_lo_hi_1592 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1593;
  assign dataGroup_lo_hi_1593 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1594;
  assign dataGroup_lo_hi_1594 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1595;
  assign dataGroup_lo_hi_1595 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1596;
  assign dataGroup_lo_hi_1596 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1597;
  assign dataGroup_lo_hi_1597 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1598;
  assign dataGroup_lo_hi_1598 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1599;
  assign dataGroup_lo_hi_1599 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1600;
  assign dataGroup_lo_hi_1600 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1601;
  assign dataGroup_lo_hi_1601 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1602;
  assign dataGroup_lo_hi_1602 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1603;
  assign dataGroup_lo_hi_1603 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1604;
  assign dataGroup_lo_hi_1604 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1605;
  assign dataGroup_lo_hi_1605 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1606;
  assign dataGroup_lo_hi_1606 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1607;
  assign dataGroup_lo_hi_1607 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1608;
  assign dataGroup_lo_hi_1608 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1609;
  assign dataGroup_lo_hi_1609 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1610;
  assign dataGroup_lo_hi_1610 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1611;
  assign dataGroup_lo_hi_1611 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1612;
  assign dataGroup_lo_hi_1612 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1613;
  assign dataGroup_lo_hi_1613 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1614;
  assign dataGroup_lo_hi_1614 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1615;
  assign dataGroup_lo_hi_1615 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1616;
  assign dataGroup_lo_hi_1616 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1617;
  assign dataGroup_lo_hi_1617 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1618;
  assign dataGroup_lo_hi_1618 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1619;
  assign dataGroup_lo_hi_1619 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1620;
  assign dataGroup_lo_hi_1620 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1621;
  assign dataGroup_lo_hi_1621 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1622;
  assign dataGroup_lo_hi_1622 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1623;
  assign dataGroup_lo_hi_1623 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1624;
  assign dataGroup_lo_hi_1624 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1625;
  assign dataGroup_lo_hi_1625 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1626;
  assign dataGroup_lo_hi_1626 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1627;
  assign dataGroup_lo_hi_1627 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1628;
  assign dataGroup_lo_hi_1628 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1629;
  assign dataGroup_lo_hi_1629 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1630;
  assign dataGroup_lo_hi_1630 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1631;
  assign dataGroup_lo_hi_1631 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1632;
  assign dataGroup_lo_hi_1632 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1633;
  assign dataGroup_lo_hi_1633 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1634;
  assign dataGroup_lo_hi_1634 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1635;
  assign dataGroup_lo_hi_1635 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1636;
  assign dataGroup_lo_hi_1636 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1637;
  assign dataGroup_lo_hi_1637 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1638;
  assign dataGroup_lo_hi_1638 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1639;
  assign dataGroup_lo_hi_1639 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1640;
  assign dataGroup_lo_hi_1640 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1641;
  assign dataGroup_lo_hi_1641 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1642;
  assign dataGroup_lo_hi_1642 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1643;
  assign dataGroup_lo_hi_1643 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1644;
  assign dataGroup_lo_hi_1644 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1645;
  assign dataGroup_lo_hi_1645 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1646;
  assign dataGroup_lo_hi_1646 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1647;
  assign dataGroup_lo_hi_1647 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1648;
  assign dataGroup_lo_hi_1648 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1649;
  assign dataGroup_lo_hi_1649 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1650;
  assign dataGroup_lo_hi_1650 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1651;
  assign dataGroup_lo_hi_1651 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1652;
  assign dataGroup_lo_hi_1652 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1653;
  assign dataGroup_lo_hi_1653 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1654;
  assign dataGroup_lo_hi_1654 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1655;
  assign dataGroup_lo_hi_1655 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1656;
  assign dataGroup_lo_hi_1656 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1657;
  assign dataGroup_lo_hi_1657 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1658;
  assign dataGroup_lo_hi_1658 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1659;
  assign dataGroup_lo_hi_1659 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1660;
  assign dataGroup_lo_hi_1660 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1661;
  assign dataGroup_lo_hi_1661 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1662;
  assign dataGroup_lo_hi_1662 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1663;
  assign dataGroup_lo_hi_1663 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1664;
  assign dataGroup_lo_hi_1664 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1665;
  assign dataGroup_lo_hi_1665 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1666;
  assign dataGroup_lo_hi_1666 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1667;
  assign dataGroup_lo_hi_1667 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1668;
  assign dataGroup_lo_hi_1668 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1669;
  assign dataGroup_lo_hi_1669 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1670;
  assign dataGroup_lo_hi_1670 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1671;
  assign dataGroup_lo_hi_1671 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1672;
  assign dataGroup_lo_hi_1672 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1673;
  assign dataGroup_lo_hi_1673 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1674;
  assign dataGroup_lo_hi_1674 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1675;
  assign dataGroup_lo_hi_1675 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1676;
  assign dataGroup_lo_hi_1676 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1677;
  assign dataGroup_lo_hi_1677 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1678;
  assign dataGroup_lo_hi_1678 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1679;
  assign dataGroup_lo_hi_1679 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1680;
  assign dataGroup_lo_hi_1680 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1681;
  assign dataGroup_lo_hi_1681 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1682;
  assign dataGroup_lo_hi_1682 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1683;
  assign dataGroup_lo_hi_1683 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1684;
  assign dataGroup_lo_hi_1684 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1685;
  assign dataGroup_lo_hi_1685 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1686;
  assign dataGroup_lo_hi_1686 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1687;
  assign dataGroup_lo_hi_1687 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1688;
  assign dataGroup_lo_hi_1688 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1689;
  assign dataGroup_lo_hi_1689 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1690;
  assign dataGroup_lo_hi_1690 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1691;
  assign dataGroup_lo_hi_1691 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1692;
  assign dataGroup_lo_hi_1692 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1693;
  assign dataGroup_lo_hi_1693 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1694;
  assign dataGroup_lo_hi_1694 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1695;
  assign dataGroup_lo_hi_1695 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1696;
  assign dataGroup_lo_hi_1696 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1697;
  assign dataGroup_lo_hi_1697 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1698;
  assign dataGroup_lo_hi_1698 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1699;
  assign dataGroup_lo_hi_1699 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1700;
  assign dataGroup_lo_hi_1700 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1701;
  assign dataGroup_lo_hi_1701 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1702;
  assign dataGroup_lo_hi_1702 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1703;
  assign dataGroup_lo_hi_1703 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1704;
  assign dataGroup_lo_hi_1704 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1705;
  assign dataGroup_lo_hi_1705 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1706;
  assign dataGroup_lo_hi_1706 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1707;
  assign dataGroup_lo_hi_1707 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1708;
  assign dataGroup_lo_hi_1708 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1709;
  assign dataGroup_lo_hi_1709 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1710;
  assign dataGroup_lo_hi_1710 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1711;
  assign dataGroup_lo_hi_1711 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1712;
  assign dataGroup_lo_hi_1712 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1713;
  assign dataGroup_lo_hi_1713 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1714;
  assign dataGroup_lo_hi_1714 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1715;
  assign dataGroup_lo_hi_1715 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1716;
  assign dataGroup_lo_hi_1716 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1717;
  assign dataGroup_lo_hi_1717 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1718;
  assign dataGroup_lo_hi_1718 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1719;
  assign dataGroup_lo_hi_1719 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1720;
  assign dataGroup_lo_hi_1720 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1721;
  assign dataGroup_lo_hi_1721 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1722;
  assign dataGroup_lo_hi_1722 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1723;
  assign dataGroup_lo_hi_1723 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1724;
  assign dataGroup_lo_hi_1724 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1725;
  assign dataGroup_lo_hi_1725 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1726;
  assign dataGroup_lo_hi_1726 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1727;
  assign dataGroup_lo_hi_1727 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1728;
  assign dataGroup_lo_hi_1728 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1729;
  assign dataGroup_lo_hi_1729 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1730;
  assign dataGroup_lo_hi_1730 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1731;
  assign dataGroup_lo_hi_1731 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1732;
  assign dataGroup_lo_hi_1732 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1733;
  assign dataGroup_lo_hi_1733 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1734;
  assign dataGroup_lo_hi_1734 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1735;
  assign dataGroup_lo_hi_1735 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1736;
  assign dataGroup_lo_hi_1736 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1737;
  assign dataGroup_lo_hi_1737 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1738;
  assign dataGroup_lo_hi_1738 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1739;
  assign dataGroup_lo_hi_1739 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1740;
  assign dataGroup_lo_hi_1740 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1741;
  assign dataGroup_lo_hi_1741 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1742;
  assign dataGroup_lo_hi_1742 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1743;
  assign dataGroup_lo_hi_1743 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1744;
  assign dataGroup_lo_hi_1744 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1745;
  assign dataGroup_lo_hi_1745 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1746;
  assign dataGroup_lo_hi_1746 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1747;
  assign dataGroup_lo_hi_1747 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1748;
  assign dataGroup_lo_hi_1748 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1749;
  assign dataGroup_lo_hi_1749 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1750;
  assign dataGroup_lo_hi_1750 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1751;
  assign dataGroup_lo_hi_1751 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1752;
  assign dataGroup_lo_hi_1752 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1753;
  assign dataGroup_lo_hi_1753 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1754;
  assign dataGroup_lo_hi_1754 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1755;
  assign dataGroup_lo_hi_1755 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1756;
  assign dataGroup_lo_hi_1756 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1757;
  assign dataGroup_lo_hi_1757 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1758;
  assign dataGroup_lo_hi_1758 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1759;
  assign dataGroup_lo_hi_1759 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1760;
  assign dataGroup_lo_hi_1760 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1761;
  assign dataGroup_lo_hi_1761 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1762;
  assign dataGroup_lo_hi_1762 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1763;
  assign dataGroup_lo_hi_1763 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1764;
  assign dataGroup_lo_hi_1764 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1765;
  assign dataGroup_lo_hi_1765 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1766;
  assign dataGroup_lo_hi_1766 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1767;
  assign dataGroup_lo_hi_1767 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1768;
  assign dataGroup_lo_hi_1768 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1769;
  assign dataGroup_lo_hi_1769 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1770;
  assign dataGroup_lo_hi_1770 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1771;
  assign dataGroup_lo_hi_1771 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1772;
  assign dataGroup_lo_hi_1772 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1773;
  assign dataGroup_lo_hi_1773 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1774;
  assign dataGroup_lo_hi_1774 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1775;
  assign dataGroup_lo_hi_1775 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1776;
  assign dataGroup_lo_hi_1776 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1777;
  assign dataGroup_lo_hi_1777 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1778;
  assign dataGroup_lo_hi_1778 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1779;
  assign dataGroup_lo_hi_1779 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1780;
  assign dataGroup_lo_hi_1780 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1781;
  assign dataGroup_lo_hi_1781 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1782;
  assign dataGroup_lo_hi_1782 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1783;
  assign dataGroup_lo_hi_1783 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1784;
  assign dataGroup_lo_hi_1784 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1785;
  assign dataGroup_lo_hi_1785 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1786;
  assign dataGroup_lo_hi_1786 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1787;
  assign dataGroup_lo_hi_1787 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1788;
  assign dataGroup_lo_hi_1788 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1789;
  assign dataGroup_lo_hi_1789 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1790;
  assign dataGroup_lo_hi_1790 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1791;
  assign dataGroup_lo_hi_1791 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1792;
  assign dataGroup_lo_hi_1792 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1793;
  assign dataGroup_lo_hi_1793 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1794;
  assign dataGroup_lo_hi_1794 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1795;
  assign dataGroup_lo_hi_1795 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1796;
  assign dataGroup_lo_hi_1796 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1797;
  assign dataGroup_lo_hi_1797 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1798;
  assign dataGroup_lo_hi_1798 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1799;
  assign dataGroup_lo_hi_1799 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1800;
  assign dataGroup_lo_hi_1800 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1801;
  assign dataGroup_lo_hi_1801 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1802;
  assign dataGroup_lo_hi_1802 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1803;
  assign dataGroup_lo_hi_1803 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1804;
  assign dataGroup_lo_hi_1804 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1805;
  assign dataGroup_lo_hi_1805 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1806;
  assign dataGroup_lo_hi_1806 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1807;
  assign dataGroup_lo_hi_1807 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1808;
  assign dataGroup_lo_hi_1808 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1809;
  assign dataGroup_lo_hi_1809 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1810;
  assign dataGroup_lo_hi_1810 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1811;
  assign dataGroup_lo_hi_1811 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1812;
  assign dataGroup_lo_hi_1812 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1813;
  assign dataGroup_lo_hi_1813 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1814;
  assign dataGroup_lo_hi_1814 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1815;
  assign dataGroup_lo_hi_1815 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1816;
  assign dataGroup_lo_hi_1816 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1817;
  assign dataGroup_lo_hi_1817 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1818;
  assign dataGroup_lo_hi_1818 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1819;
  assign dataGroup_lo_hi_1819 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1820;
  assign dataGroup_lo_hi_1820 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1821;
  assign dataGroup_lo_hi_1821 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1822;
  assign dataGroup_lo_hi_1822 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1823;
  assign dataGroup_lo_hi_1823 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1824;
  assign dataGroup_lo_hi_1824 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1825;
  assign dataGroup_lo_hi_1825 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1826;
  assign dataGroup_lo_hi_1826 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1827;
  assign dataGroup_lo_hi_1827 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1828;
  assign dataGroup_lo_hi_1828 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1829;
  assign dataGroup_lo_hi_1829 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1830;
  assign dataGroup_lo_hi_1830 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1831;
  assign dataGroup_lo_hi_1831 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1832;
  assign dataGroup_lo_hi_1832 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1833;
  assign dataGroup_lo_hi_1833 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1834;
  assign dataGroup_lo_hi_1834 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1835;
  assign dataGroup_lo_hi_1835 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1836;
  assign dataGroup_lo_hi_1836 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1837;
  assign dataGroup_lo_hi_1837 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1838;
  assign dataGroup_lo_hi_1838 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1839;
  assign dataGroup_lo_hi_1839 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1840;
  assign dataGroup_lo_hi_1840 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1841;
  assign dataGroup_lo_hi_1841 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1842;
  assign dataGroup_lo_hi_1842 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1843;
  assign dataGroup_lo_hi_1843 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1844;
  assign dataGroup_lo_hi_1844 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1845;
  assign dataGroup_lo_hi_1845 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1846;
  assign dataGroup_lo_hi_1846 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1847;
  assign dataGroup_lo_hi_1847 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1848;
  assign dataGroup_lo_hi_1848 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1849;
  assign dataGroup_lo_hi_1849 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1850;
  assign dataGroup_lo_hi_1850 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1851;
  assign dataGroup_lo_hi_1851 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1852;
  assign dataGroup_lo_hi_1852 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1853;
  assign dataGroup_lo_hi_1853 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1854;
  assign dataGroup_lo_hi_1854 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1855;
  assign dataGroup_lo_hi_1855 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1856;
  assign dataGroup_lo_hi_1856 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1857;
  assign dataGroup_lo_hi_1857 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1858;
  assign dataGroup_lo_hi_1858 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1859;
  assign dataGroup_lo_hi_1859 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1860;
  assign dataGroup_lo_hi_1860 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1861;
  assign dataGroup_lo_hi_1861 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1862;
  assign dataGroup_lo_hi_1862 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1863;
  assign dataGroup_lo_hi_1863 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1864;
  assign dataGroup_lo_hi_1864 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1865;
  assign dataGroup_lo_hi_1865 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1866;
  assign dataGroup_lo_hi_1866 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1867;
  assign dataGroup_lo_hi_1867 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1868;
  assign dataGroup_lo_hi_1868 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1869;
  assign dataGroup_lo_hi_1869 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1870;
  assign dataGroup_lo_hi_1870 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1871;
  assign dataGroup_lo_hi_1871 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1872;
  assign dataGroup_lo_hi_1872 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1873;
  assign dataGroup_lo_hi_1873 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1874;
  assign dataGroup_lo_hi_1874 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1875;
  assign dataGroup_lo_hi_1875 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1876;
  assign dataGroup_lo_hi_1876 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1877;
  assign dataGroup_lo_hi_1877 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1878;
  assign dataGroup_lo_hi_1878 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1879;
  assign dataGroup_lo_hi_1879 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1880;
  assign dataGroup_lo_hi_1880 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1881;
  assign dataGroup_lo_hi_1881 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1882;
  assign dataGroup_lo_hi_1882 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1883;
  assign dataGroup_lo_hi_1883 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1884;
  assign dataGroup_lo_hi_1884 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1885;
  assign dataGroup_lo_hi_1885 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1886;
  assign dataGroup_lo_hi_1886 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1887;
  assign dataGroup_lo_hi_1887 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1888;
  assign dataGroup_lo_hi_1888 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1889;
  assign dataGroup_lo_hi_1889 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1890;
  assign dataGroup_lo_hi_1890 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1891;
  assign dataGroup_lo_hi_1891 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1892;
  assign dataGroup_lo_hi_1892 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1893;
  assign dataGroup_lo_hi_1893 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1894;
  assign dataGroup_lo_hi_1894 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1895;
  assign dataGroup_lo_hi_1895 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1896;
  assign dataGroup_lo_hi_1896 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1897;
  assign dataGroup_lo_hi_1897 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1898;
  assign dataGroup_lo_hi_1898 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1899;
  assign dataGroup_lo_hi_1899 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1900;
  assign dataGroup_lo_hi_1900 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1901;
  assign dataGroup_lo_hi_1901 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1902;
  assign dataGroup_lo_hi_1902 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1903;
  assign dataGroup_lo_hi_1903 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1904;
  assign dataGroup_lo_hi_1904 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1905;
  assign dataGroup_lo_hi_1905 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1906;
  assign dataGroup_lo_hi_1906 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1907;
  assign dataGroup_lo_hi_1907 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1908;
  assign dataGroup_lo_hi_1908 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1909;
  assign dataGroup_lo_hi_1909 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1910;
  assign dataGroup_lo_hi_1910 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1911;
  assign dataGroup_lo_hi_1911 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1912;
  assign dataGroup_lo_hi_1912 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1913;
  assign dataGroup_lo_hi_1913 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1914;
  assign dataGroup_lo_hi_1914 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1915;
  assign dataGroup_lo_hi_1915 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1916;
  assign dataGroup_lo_hi_1916 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1917;
  assign dataGroup_lo_hi_1917 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1918;
  assign dataGroup_lo_hi_1918 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1919;
  assign dataGroup_lo_hi_1919 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1920;
  assign dataGroup_lo_hi_1920 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1921;
  assign dataGroup_lo_hi_1921 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1922;
  assign dataGroup_lo_hi_1922 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1923;
  assign dataGroup_lo_hi_1923 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1924;
  assign dataGroup_lo_hi_1924 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1925;
  assign dataGroup_lo_hi_1925 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1926;
  assign dataGroup_lo_hi_1926 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1927;
  assign dataGroup_lo_hi_1927 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1928;
  assign dataGroup_lo_hi_1928 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1929;
  assign dataGroup_lo_hi_1929 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1930;
  assign dataGroup_lo_hi_1930 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1931;
  assign dataGroup_lo_hi_1931 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1932;
  assign dataGroup_lo_hi_1932 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1933;
  assign dataGroup_lo_hi_1933 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1934;
  assign dataGroup_lo_hi_1934 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1935;
  assign dataGroup_lo_hi_1935 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1936;
  assign dataGroup_lo_hi_1936 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1937;
  assign dataGroup_lo_hi_1937 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1938;
  assign dataGroup_lo_hi_1938 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1939;
  assign dataGroup_lo_hi_1939 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1940;
  assign dataGroup_lo_hi_1940 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1941;
  assign dataGroup_lo_hi_1941 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1942;
  assign dataGroup_lo_hi_1942 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1943;
  assign dataGroup_lo_hi_1943 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1944;
  assign dataGroup_lo_hi_1944 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1945;
  assign dataGroup_lo_hi_1945 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1946;
  assign dataGroup_lo_hi_1946 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1947;
  assign dataGroup_lo_hi_1947 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1948;
  assign dataGroup_lo_hi_1948 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1949;
  assign dataGroup_lo_hi_1949 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1950;
  assign dataGroup_lo_hi_1950 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1951;
  assign dataGroup_lo_hi_1951 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1952;
  assign dataGroup_lo_hi_1952 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1953;
  assign dataGroup_lo_hi_1953 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1954;
  assign dataGroup_lo_hi_1954 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1955;
  assign dataGroup_lo_hi_1955 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1956;
  assign dataGroup_lo_hi_1956 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1957;
  assign dataGroup_lo_hi_1957 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1958;
  assign dataGroup_lo_hi_1958 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1959;
  assign dataGroup_lo_hi_1959 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1960;
  assign dataGroup_lo_hi_1960 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1961;
  assign dataGroup_lo_hi_1961 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1962;
  assign dataGroup_lo_hi_1962 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1963;
  assign dataGroup_lo_hi_1963 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1964;
  assign dataGroup_lo_hi_1964 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1965;
  assign dataGroup_lo_hi_1965 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1966;
  assign dataGroup_lo_hi_1966 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1967;
  assign dataGroup_lo_hi_1967 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1968;
  assign dataGroup_lo_hi_1968 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1969;
  assign dataGroup_lo_hi_1969 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1970;
  assign dataGroup_lo_hi_1970 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1971;
  assign dataGroup_lo_hi_1971 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1972;
  assign dataGroup_lo_hi_1972 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1973;
  assign dataGroup_lo_hi_1973 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1974;
  assign dataGroup_lo_hi_1974 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1975;
  assign dataGroup_lo_hi_1975 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1976;
  assign dataGroup_lo_hi_1976 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1977;
  assign dataGroup_lo_hi_1977 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1978;
  assign dataGroup_lo_hi_1978 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1979;
  assign dataGroup_lo_hi_1979 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1980;
  assign dataGroup_lo_hi_1980 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1981;
  assign dataGroup_lo_hi_1981 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1982;
  assign dataGroup_lo_hi_1982 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1983;
  assign dataGroup_lo_hi_1983 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1984;
  assign dataGroup_lo_hi_1984 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1985;
  assign dataGroup_lo_hi_1985 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1986;
  assign dataGroup_lo_hi_1986 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1987;
  assign dataGroup_lo_hi_1987 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1988;
  assign dataGroup_lo_hi_1988 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1989;
  assign dataGroup_lo_hi_1989 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1990;
  assign dataGroup_lo_hi_1990 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1991;
  assign dataGroup_lo_hi_1991 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1992;
  assign dataGroup_lo_hi_1992 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1993;
  assign dataGroup_lo_hi_1993 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1994;
  assign dataGroup_lo_hi_1994 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1995;
  assign dataGroup_lo_hi_1995 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1996;
  assign dataGroup_lo_hi_1996 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1997;
  assign dataGroup_lo_hi_1997 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1998;
  assign dataGroup_lo_hi_1998 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_1999;
  assign dataGroup_lo_hi_1999 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2000;
  assign dataGroup_lo_hi_2000 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2001;
  assign dataGroup_lo_hi_2001 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2002;
  assign dataGroup_lo_hi_2002 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2003;
  assign dataGroup_lo_hi_2003 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2004;
  assign dataGroup_lo_hi_2004 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2005;
  assign dataGroup_lo_hi_2005 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2006;
  assign dataGroup_lo_hi_2006 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2007;
  assign dataGroup_lo_hi_2007 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2008;
  assign dataGroup_lo_hi_2008 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2009;
  assign dataGroup_lo_hi_2009 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2010;
  assign dataGroup_lo_hi_2010 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2011;
  assign dataGroup_lo_hi_2011 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2012;
  assign dataGroup_lo_hi_2012 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2013;
  assign dataGroup_lo_hi_2013 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2014;
  assign dataGroup_lo_hi_2014 = _GEN_5;
  wire [511:0]  dataGroup_lo_hi_2015;
  assign dataGroup_lo_hi_2015 = _GEN_5;
  wire [1023:0] dataGroup_lo = {dataGroup_lo_hi, dataGroup_lo_lo};
  wire [511:0]  _GEN_6 = {dataSelect_5, dataSelect_4};
  wire [511:0]  dataGroup_hi_lo;
  assign dataGroup_hi_lo = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1;
  assign dataGroup_hi_lo_1 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2;
  assign dataGroup_hi_lo_2 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_3;
  assign dataGroup_hi_lo_3 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_4;
  assign dataGroup_hi_lo_4 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_5;
  assign dataGroup_hi_lo_5 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_6;
  assign dataGroup_hi_lo_6 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_7;
  assign dataGroup_hi_lo_7 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_8;
  assign dataGroup_hi_lo_8 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_9;
  assign dataGroup_hi_lo_9 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_10;
  assign dataGroup_hi_lo_10 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_11;
  assign dataGroup_hi_lo_11 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_12;
  assign dataGroup_hi_lo_12 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_13;
  assign dataGroup_hi_lo_13 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_14;
  assign dataGroup_hi_lo_14 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_15;
  assign dataGroup_hi_lo_15 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_16;
  assign dataGroup_hi_lo_16 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_17;
  assign dataGroup_hi_lo_17 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_18;
  assign dataGroup_hi_lo_18 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_19;
  assign dataGroup_hi_lo_19 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_20;
  assign dataGroup_hi_lo_20 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_21;
  assign dataGroup_hi_lo_21 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_22;
  assign dataGroup_hi_lo_22 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_23;
  assign dataGroup_hi_lo_23 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_24;
  assign dataGroup_hi_lo_24 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_25;
  assign dataGroup_hi_lo_25 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_26;
  assign dataGroup_hi_lo_26 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_27;
  assign dataGroup_hi_lo_27 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_28;
  assign dataGroup_hi_lo_28 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_29;
  assign dataGroup_hi_lo_29 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_30;
  assign dataGroup_hi_lo_30 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_31;
  assign dataGroup_hi_lo_31 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_32;
  assign dataGroup_hi_lo_32 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_33;
  assign dataGroup_hi_lo_33 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_34;
  assign dataGroup_hi_lo_34 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_35;
  assign dataGroup_hi_lo_35 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_36;
  assign dataGroup_hi_lo_36 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_37;
  assign dataGroup_hi_lo_37 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_38;
  assign dataGroup_hi_lo_38 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_39;
  assign dataGroup_hi_lo_39 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_40;
  assign dataGroup_hi_lo_40 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_41;
  assign dataGroup_hi_lo_41 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_42;
  assign dataGroup_hi_lo_42 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_43;
  assign dataGroup_hi_lo_43 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_44;
  assign dataGroup_hi_lo_44 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_45;
  assign dataGroup_hi_lo_45 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_46;
  assign dataGroup_hi_lo_46 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_47;
  assign dataGroup_hi_lo_47 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_48;
  assign dataGroup_hi_lo_48 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_49;
  assign dataGroup_hi_lo_49 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_50;
  assign dataGroup_hi_lo_50 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_51;
  assign dataGroup_hi_lo_51 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_52;
  assign dataGroup_hi_lo_52 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_53;
  assign dataGroup_hi_lo_53 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_54;
  assign dataGroup_hi_lo_54 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_55;
  assign dataGroup_hi_lo_55 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_56;
  assign dataGroup_hi_lo_56 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_57;
  assign dataGroup_hi_lo_57 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_58;
  assign dataGroup_hi_lo_58 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_59;
  assign dataGroup_hi_lo_59 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_60;
  assign dataGroup_hi_lo_60 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_61;
  assign dataGroup_hi_lo_61 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_62;
  assign dataGroup_hi_lo_62 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_63;
  assign dataGroup_hi_lo_63 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_64;
  assign dataGroup_hi_lo_64 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_65;
  assign dataGroup_hi_lo_65 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_66;
  assign dataGroup_hi_lo_66 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_67;
  assign dataGroup_hi_lo_67 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_68;
  assign dataGroup_hi_lo_68 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_69;
  assign dataGroup_hi_lo_69 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_70;
  assign dataGroup_hi_lo_70 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_71;
  assign dataGroup_hi_lo_71 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_72;
  assign dataGroup_hi_lo_72 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_73;
  assign dataGroup_hi_lo_73 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_74;
  assign dataGroup_hi_lo_74 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_75;
  assign dataGroup_hi_lo_75 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_76;
  assign dataGroup_hi_lo_76 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_77;
  assign dataGroup_hi_lo_77 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_78;
  assign dataGroup_hi_lo_78 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_79;
  assign dataGroup_hi_lo_79 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_80;
  assign dataGroup_hi_lo_80 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_81;
  assign dataGroup_hi_lo_81 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_82;
  assign dataGroup_hi_lo_82 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_83;
  assign dataGroup_hi_lo_83 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_84;
  assign dataGroup_hi_lo_84 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_85;
  assign dataGroup_hi_lo_85 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_86;
  assign dataGroup_hi_lo_86 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_87;
  assign dataGroup_hi_lo_87 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_88;
  assign dataGroup_hi_lo_88 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_89;
  assign dataGroup_hi_lo_89 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_90;
  assign dataGroup_hi_lo_90 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_91;
  assign dataGroup_hi_lo_91 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_92;
  assign dataGroup_hi_lo_92 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_93;
  assign dataGroup_hi_lo_93 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_94;
  assign dataGroup_hi_lo_94 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_95;
  assign dataGroup_hi_lo_95 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_96;
  assign dataGroup_hi_lo_96 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_97;
  assign dataGroup_hi_lo_97 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_98;
  assign dataGroup_hi_lo_98 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_99;
  assign dataGroup_hi_lo_99 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_100;
  assign dataGroup_hi_lo_100 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_101;
  assign dataGroup_hi_lo_101 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_102;
  assign dataGroup_hi_lo_102 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_103;
  assign dataGroup_hi_lo_103 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_104;
  assign dataGroup_hi_lo_104 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_105;
  assign dataGroup_hi_lo_105 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_106;
  assign dataGroup_hi_lo_106 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_107;
  assign dataGroup_hi_lo_107 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_108;
  assign dataGroup_hi_lo_108 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_109;
  assign dataGroup_hi_lo_109 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_110;
  assign dataGroup_hi_lo_110 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_111;
  assign dataGroup_hi_lo_111 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_112;
  assign dataGroup_hi_lo_112 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_113;
  assign dataGroup_hi_lo_113 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_114;
  assign dataGroup_hi_lo_114 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_115;
  assign dataGroup_hi_lo_115 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_116;
  assign dataGroup_hi_lo_116 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_117;
  assign dataGroup_hi_lo_117 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_118;
  assign dataGroup_hi_lo_118 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_119;
  assign dataGroup_hi_lo_119 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_120;
  assign dataGroup_hi_lo_120 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_121;
  assign dataGroup_hi_lo_121 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_122;
  assign dataGroup_hi_lo_122 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_123;
  assign dataGroup_hi_lo_123 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_124;
  assign dataGroup_hi_lo_124 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_125;
  assign dataGroup_hi_lo_125 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_126;
  assign dataGroup_hi_lo_126 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_127;
  assign dataGroup_hi_lo_127 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_128;
  assign dataGroup_hi_lo_128 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_129;
  assign dataGroup_hi_lo_129 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_130;
  assign dataGroup_hi_lo_130 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_131;
  assign dataGroup_hi_lo_131 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_132;
  assign dataGroup_hi_lo_132 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_133;
  assign dataGroup_hi_lo_133 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_134;
  assign dataGroup_hi_lo_134 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_135;
  assign dataGroup_hi_lo_135 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_136;
  assign dataGroup_hi_lo_136 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_137;
  assign dataGroup_hi_lo_137 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_138;
  assign dataGroup_hi_lo_138 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_139;
  assign dataGroup_hi_lo_139 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_140;
  assign dataGroup_hi_lo_140 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_141;
  assign dataGroup_hi_lo_141 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_142;
  assign dataGroup_hi_lo_142 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_143;
  assign dataGroup_hi_lo_143 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_144;
  assign dataGroup_hi_lo_144 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_145;
  assign dataGroup_hi_lo_145 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_146;
  assign dataGroup_hi_lo_146 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_147;
  assign dataGroup_hi_lo_147 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_148;
  assign dataGroup_hi_lo_148 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_149;
  assign dataGroup_hi_lo_149 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_150;
  assign dataGroup_hi_lo_150 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_151;
  assign dataGroup_hi_lo_151 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_152;
  assign dataGroup_hi_lo_152 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_153;
  assign dataGroup_hi_lo_153 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_154;
  assign dataGroup_hi_lo_154 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_155;
  assign dataGroup_hi_lo_155 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_156;
  assign dataGroup_hi_lo_156 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_157;
  assign dataGroup_hi_lo_157 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_158;
  assign dataGroup_hi_lo_158 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_159;
  assign dataGroup_hi_lo_159 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_160;
  assign dataGroup_hi_lo_160 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_161;
  assign dataGroup_hi_lo_161 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_162;
  assign dataGroup_hi_lo_162 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_163;
  assign dataGroup_hi_lo_163 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_164;
  assign dataGroup_hi_lo_164 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_165;
  assign dataGroup_hi_lo_165 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_166;
  assign dataGroup_hi_lo_166 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_167;
  assign dataGroup_hi_lo_167 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_168;
  assign dataGroup_hi_lo_168 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_169;
  assign dataGroup_hi_lo_169 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_170;
  assign dataGroup_hi_lo_170 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_171;
  assign dataGroup_hi_lo_171 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_172;
  assign dataGroup_hi_lo_172 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_173;
  assign dataGroup_hi_lo_173 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_174;
  assign dataGroup_hi_lo_174 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_175;
  assign dataGroup_hi_lo_175 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_176;
  assign dataGroup_hi_lo_176 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_177;
  assign dataGroup_hi_lo_177 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_178;
  assign dataGroup_hi_lo_178 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_179;
  assign dataGroup_hi_lo_179 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_180;
  assign dataGroup_hi_lo_180 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_181;
  assign dataGroup_hi_lo_181 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_182;
  assign dataGroup_hi_lo_182 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_183;
  assign dataGroup_hi_lo_183 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_184;
  assign dataGroup_hi_lo_184 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_185;
  assign dataGroup_hi_lo_185 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_186;
  assign dataGroup_hi_lo_186 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_187;
  assign dataGroup_hi_lo_187 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_188;
  assign dataGroup_hi_lo_188 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_189;
  assign dataGroup_hi_lo_189 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_190;
  assign dataGroup_hi_lo_190 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_191;
  assign dataGroup_hi_lo_191 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_192;
  assign dataGroup_hi_lo_192 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_193;
  assign dataGroup_hi_lo_193 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_194;
  assign dataGroup_hi_lo_194 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_195;
  assign dataGroup_hi_lo_195 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_196;
  assign dataGroup_hi_lo_196 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_197;
  assign dataGroup_hi_lo_197 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_198;
  assign dataGroup_hi_lo_198 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_199;
  assign dataGroup_hi_lo_199 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_200;
  assign dataGroup_hi_lo_200 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_201;
  assign dataGroup_hi_lo_201 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_202;
  assign dataGroup_hi_lo_202 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_203;
  assign dataGroup_hi_lo_203 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_204;
  assign dataGroup_hi_lo_204 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_205;
  assign dataGroup_hi_lo_205 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_206;
  assign dataGroup_hi_lo_206 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_207;
  assign dataGroup_hi_lo_207 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_208;
  assign dataGroup_hi_lo_208 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_209;
  assign dataGroup_hi_lo_209 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_210;
  assign dataGroup_hi_lo_210 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_211;
  assign dataGroup_hi_lo_211 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_212;
  assign dataGroup_hi_lo_212 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_213;
  assign dataGroup_hi_lo_213 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_214;
  assign dataGroup_hi_lo_214 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_215;
  assign dataGroup_hi_lo_215 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_216;
  assign dataGroup_hi_lo_216 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_217;
  assign dataGroup_hi_lo_217 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_218;
  assign dataGroup_hi_lo_218 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_219;
  assign dataGroup_hi_lo_219 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_220;
  assign dataGroup_hi_lo_220 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_221;
  assign dataGroup_hi_lo_221 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_222;
  assign dataGroup_hi_lo_222 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_223;
  assign dataGroup_hi_lo_223 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_224;
  assign dataGroup_hi_lo_224 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_225;
  assign dataGroup_hi_lo_225 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_226;
  assign dataGroup_hi_lo_226 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_227;
  assign dataGroup_hi_lo_227 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_228;
  assign dataGroup_hi_lo_228 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_229;
  assign dataGroup_hi_lo_229 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_230;
  assign dataGroup_hi_lo_230 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_231;
  assign dataGroup_hi_lo_231 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_232;
  assign dataGroup_hi_lo_232 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_233;
  assign dataGroup_hi_lo_233 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_234;
  assign dataGroup_hi_lo_234 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_235;
  assign dataGroup_hi_lo_235 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_236;
  assign dataGroup_hi_lo_236 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_237;
  assign dataGroup_hi_lo_237 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_238;
  assign dataGroup_hi_lo_238 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_239;
  assign dataGroup_hi_lo_239 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_240;
  assign dataGroup_hi_lo_240 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_241;
  assign dataGroup_hi_lo_241 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_242;
  assign dataGroup_hi_lo_242 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_243;
  assign dataGroup_hi_lo_243 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_244;
  assign dataGroup_hi_lo_244 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_245;
  assign dataGroup_hi_lo_245 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_246;
  assign dataGroup_hi_lo_246 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_247;
  assign dataGroup_hi_lo_247 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_248;
  assign dataGroup_hi_lo_248 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_249;
  assign dataGroup_hi_lo_249 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_250;
  assign dataGroup_hi_lo_250 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_251;
  assign dataGroup_hi_lo_251 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_252;
  assign dataGroup_hi_lo_252 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_253;
  assign dataGroup_hi_lo_253 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_254;
  assign dataGroup_hi_lo_254 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_255;
  assign dataGroup_hi_lo_255 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_256;
  assign dataGroup_hi_lo_256 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_257;
  assign dataGroup_hi_lo_257 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_258;
  assign dataGroup_hi_lo_258 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_259;
  assign dataGroup_hi_lo_259 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_260;
  assign dataGroup_hi_lo_260 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_261;
  assign dataGroup_hi_lo_261 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_262;
  assign dataGroup_hi_lo_262 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_263;
  assign dataGroup_hi_lo_263 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_264;
  assign dataGroup_hi_lo_264 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_265;
  assign dataGroup_hi_lo_265 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_266;
  assign dataGroup_hi_lo_266 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_267;
  assign dataGroup_hi_lo_267 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_268;
  assign dataGroup_hi_lo_268 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_269;
  assign dataGroup_hi_lo_269 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_270;
  assign dataGroup_hi_lo_270 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_271;
  assign dataGroup_hi_lo_271 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_272;
  assign dataGroup_hi_lo_272 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_273;
  assign dataGroup_hi_lo_273 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_274;
  assign dataGroup_hi_lo_274 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_275;
  assign dataGroup_hi_lo_275 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_276;
  assign dataGroup_hi_lo_276 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_277;
  assign dataGroup_hi_lo_277 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_278;
  assign dataGroup_hi_lo_278 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_279;
  assign dataGroup_hi_lo_279 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_280;
  assign dataGroup_hi_lo_280 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_281;
  assign dataGroup_hi_lo_281 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_282;
  assign dataGroup_hi_lo_282 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_283;
  assign dataGroup_hi_lo_283 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_284;
  assign dataGroup_hi_lo_284 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_285;
  assign dataGroup_hi_lo_285 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_286;
  assign dataGroup_hi_lo_286 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_287;
  assign dataGroup_hi_lo_287 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_288;
  assign dataGroup_hi_lo_288 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_289;
  assign dataGroup_hi_lo_289 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_290;
  assign dataGroup_hi_lo_290 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_291;
  assign dataGroup_hi_lo_291 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_292;
  assign dataGroup_hi_lo_292 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_293;
  assign dataGroup_hi_lo_293 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_294;
  assign dataGroup_hi_lo_294 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_295;
  assign dataGroup_hi_lo_295 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_296;
  assign dataGroup_hi_lo_296 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_297;
  assign dataGroup_hi_lo_297 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_298;
  assign dataGroup_hi_lo_298 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_299;
  assign dataGroup_hi_lo_299 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_300;
  assign dataGroup_hi_lo_300 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_301;
  assign dataGroup_hi_lo_301 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_302;
  assign dataGroup_hi_lo_302 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_303;
  assign dataGroup_hi_lo_303 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_304;
  assign dataGroup_hi_lo_304 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_305;
  assign dataGroup_hi_lo_305 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_306;
  assign dataGroup_hi_lo_306 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_307;
  assign dataGroup_hi_lo_307 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_308;
  assign dataGroup_hi_lo_308 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_309;
  assign dataGroup_hi_lo_309 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_310;
  assign dataGroup_hi_lo_310 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_311;
  assign dataGroup_hi_lo_311 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_312;
  assign dataGroup_hi_lo_312 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_313;
  assign dataGroup_hi_lo_313 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_314;
  assign dataGroup_hi_lo_314 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_315;
  assign dataGroup_hi_lo_315 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_316;
  assign dataGroup_hi_lo_316 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_317;
  assign dataGroup_hi_lo_317 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_318;
  assign dataGroup_hi_lo_318 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_319;
  assign dataGroup_hi_lo_319 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_320;
  assign dataGroup_hi_lo_320 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_321;
  assign dataGroup_hi_lo_321 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_322;
  assign dataGroup_hi_lo_322 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_323;
  assign dataGroup_hi_lo_323 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_324;
  assign dataGroup_hi_lo_324 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_325;
  assign dataGroup_hi_lo_325 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_326;
  assign dataGroup_hi_lo_326 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_327;
  assign dataGroup_hi_lo_327 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_328;
  assign dataGroup_hi_lo_328 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_329;
  assign dataGroup_hi_lo_329 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_330;
  assign dataGroup_hi_lo_330 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_331;
  assign dataGroup_hi_lo_331 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_332;
  assign dataGroup_hi_lo_332 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_333;
  assign dataGroup_hi_lo_333 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_334;
  assign dataGroup_hi_lo_334 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_335;
  assign dataGroup_hi_lo_335 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_336;
  assign dataGroup_hi_lo_336 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_337;
  assign dataGroup_hi_lo_337 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_338;
  assign dataGroup_hi_lo_338 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_339;
  assign dataGroup_hi_lo_339 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_340;
  assign dataGroup_hi_lo_340 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_341;
  assign dataGroup_hi_lo_341 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_342;
  assign dataGroup_hi_lo_342 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_343;
  assign dataGroup_hi_lo_343 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_344;
  assign dataGroup_hi_lo_344 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_345;
  assign dataGroup_hi_lo_345 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_346;
  assign dataGroup_hi_lo_346 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_347;
  assign dataGroup_hi_lo_347 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_348;
  assign dataGroup_hi_lo_348 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_349;
  assign dataGroup_hi_lo_349 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_350;
  assign dataGroup_hi_lo_350 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_351;
  assign dataGroup_hi_lo_351 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_352;
  assign dataGroup_hi_lo_352 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_353;
  assign dataGroup_hi_lo_353 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_354;
  assign dataGroup_hi_lo_354 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_355;
  assign dataGroup_hi_lo_355 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_356;
  assign dataGroup_hi_lo_356 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_357;
  assign dataGroup_hi_lo_357 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_358;
  assign dataGroup_hi_lo_358 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_359;
  assign dataGroup_hi_lo_359 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_360;
  assign dataGroup_hi_lo_360 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_361;
  assign dataGroup_hi_lo_361 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_362;
  assign dataGroup_hi_lo_362 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_363;
  assign dataGroup_hi_lo_363 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_364;
  assign dataGroup_hi_lo_364 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_365;
  assign dataGroup_hi_lo_365 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_366;
  assign dataGroup_hi_lo_366 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_367;
  assign dataGroup_hi_lo_367 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_368;
  assign dataGroup_hi_lo_368 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_369;
  assign dataGroup_hi_lo_369 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_370;
  assign dataGroup_hi_lo_370 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_371;
  assign dataGroup_hi_lo_371 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_372;
  assign dataGroup_hi_lo_372 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_373;
  assign dataGroup_hi_lo_373 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_374;
  assign dataGroup_hi_lo_374 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_375;
  assign dataGroup_hi_lo_375 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_376;
  assign dataGroup_hi_lo_376 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_377;
  assign dataGroup_hi_lo_377 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_378;
  assign dataGroup_hi_lo_378 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_379;
  assign dataGroup_hi_lo_379 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_380;
  assign dataGroup_hi_lo_380 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_381;
  assign dataGroup_hi_lo_381 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_382;
  assign dataGroup_hi_lo_382 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_383;
  assign dataGroup_hi_lo_383 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_384;
  assign dataGroup_hi_lo_384 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_385;
  assign dataGroup_hi_lo_385 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_386;
  assign dataGroup_hi_lo_386 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_387;
  assign dataGroup_hi_lo_387 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_388;
  assign dataGroup_hi_lo_388 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_389;
  assign dataGroup_hi_lo_389 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_390;
  assign dataGroup_hi_lo_390 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_391;
  assign dataGroup_hi_lo_391 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_392;
  assign dataGroup_hi_lo_392 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_393;
  assign dataGroup_hi_lo_393 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_394;
  assign dataGroup_hi_lo_394 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_395;
  assign dataGroup_hi_lo_395 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_396;
  assign dataGroup_hi_lo_396 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_397;
  assign dataGroup_hi_lo_397 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_398;
  assign dataGroup_hi_lo_398 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_399;
  assign dataGroup_hi_lo_399 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_400;
  assign dataGroup_hi_lo_400 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_401;
  assign dataGroup_hi_lo_401 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_402;
  assign dataGroup_hi_lo_402 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_403;
  assign dataGroup_hi_lo_403 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_404;
  assign dataGroup_hi_lo_404 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_405;
  assign dataGroup_hi_lo_405 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_406;
  assign dataGroup_hi_lo_406 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_407;
  assign dataGroup_hi_lo_407 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_408;
  assign dataGroup_hi_lo_408 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_409;
  assign dataGroup_hi_lo_409 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_410;
  assign dataGroup_hi_lo_410 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_411;
  assign dataGroup_hi_lo_411 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_412;
  assign dataGroup_hi_lo_412 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_413;
  assign dataGroup_hi_lo_413 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_414;
  assign dataGroup_hi_lo_414 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_415;
  assign dataGroup_hi_lo_415 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_416;
  assign dataGroup_hi_lo_416 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_417;
  assign dataGroup_hi_lo_417 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_418;
  assign dataGroup_hi_lo_418 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_419;
  assign dataGroup_hi_lo_419 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_420;
  assign dataGroup_hi_lo_420 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_421;
  assign dataGroup_hi_lo_421 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_422;
  assign dataGroup_hi_lo_422 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_423;
  assign dataGroup_hi_lo_423 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_424;
  assign dataGroup_hi_lo_424 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_425;
  assign dataGroup_hi_lo_425 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_426;
  assign dataGroup_hi_lo_426 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_427;
  assign dataGroup_hi_lo_427 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_428;
  assign dataGroup_hi_lo_428 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_429;
  assign dataGroup_hi_lo_429 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_430;
  assign dataGroup_hi_lo_430 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_431;
  assign dataGroup_hi_lo_431 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_432;
  assign dataGroup_hi_lo_432 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_433;
  assign dataGroup_hi_lo_433 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_434;
  assign dataGroup_hi_lo_434 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_435;
  assign dataGroup_hi_lo_435 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_436;
  assign dataGroup_hi_lo_436 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_437;
  assign dataGroup_hi_lo_437 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_438;
  assign dataGroup_hi_lo_438 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_439;
  assign dataGroup_hi_lo_439 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_440;
  assign dataGroup_hi_lo_440 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_441;
  assign dataGroup_hi_lo_441 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_442;
  assign dataGroup_hi_lo_442 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_443;
  assign dataGroup_hi_lo_443 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_444;
  assign dataGroup_hi_lo_444 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_445;
  assign dataGroup_hi_lo_445 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_446;
  assign dataGroup_hi_lo_446 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_447;
  assign dataGroup_hi_lo_447 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_448;
  assign dataGroup_hi_lo_448 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_449;
  assign dataGroup_hi_lo_449 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_450;
  assign dataGroup_hi_lo_450 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_451;
  assign dataGroup_hi_lo_451 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_452;
  assign dataGroup_hi_lo_452 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_453;
  assign dataGroup_hi_lo_453 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_454;
  assign dataGroup_hi_lo_454 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_455;
  assign dataGroup_hi_lo_455 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_456;
  assign dataGroup_hi_lo_456 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_457;
  assign dataGroup_hi_lo_457 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_458;
  assign dataGroup_hi_lo_458 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_459;
  assign dataGroup_hi_lo_459 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_460;
  assign dataGroup_hi_lo_460 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_461;
  assign dataGroup_hi_lo_461 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_462;
  assign dataGroup_hi_lo_462 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_463;
  assign dataGroup_hi_lo_463 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_464;
  assign dataGroup_hi_lo_464 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_465;
  assign dataGroup_hi_lo_465 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_466;
  assign dataGroup_hi_lo_466 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_467;
  assign dataGroup_hi_lo_467 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_468;
  assign dataGroup_hi_lo_468 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_469;
  assign dataGroup_hi_lo_469 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_470;
  assign dataGroup_hi_lo_470 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_471;
  assign dataGroup_hi_lo_471 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_472;
  assign dataGroup_hi_lo_472 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_473;
  assign dataGroup_hi_lo_473 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_474;
  assign dataGroup_hi_lo_474 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_475;
  assign dataGroup_hi_lo_475 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_476;
  assign dataGroup_hi_lo_476 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_477;
  assign dataGroup_hi_lo_477 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_478;
  assign dataGroup_hi_lo_478 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_479;
  assign dataGroup_hi_lo_479 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_480;
  assign dataGroup_hi_lo_480 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_481;
  assign dataGroup_hi_lo_481 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_482;
  assign dataGroup_hi_lo_482 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_483;
  assign dataGroup_hi_lo_483 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_484;
  assign dataGroup_hi_lo_484 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_485;
  assign dataGroup_hi_lo_485 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_486;
  assign dataGroup_hi_lo_486 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_487;
  assign dataGroup_hi_lo_487 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_488;
  assign dataGroup_hi_lo_488 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_489;
  assign dataGroup_hi_lo_489 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_490;
  assign dataGroup_hi_lo_490 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_491;
  assign dataGroup_hi_lo_491 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_492;
  assign dataGroup_hi_lo_492 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_493;
  assign dataGroup_hi_lo_493 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_494;
  assign dataGroup_hi_lo_494 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_495;
  assign dataGroup_hi_lo_495 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_496;
  assign dataGroup_hi_lo_496 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_497;
  assign dataGroup_hi_lo_497 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_498;
  assign dataGroup_hi_lo_498 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_499;
  assign dataGroup_hi_lo_499 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_500;
  assign dataGroup_hi_lo_500 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_501;
  assign dataGroup_hi_lo_501 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_502;
  assign dataGroup_hi_lo_502 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_503;
  assign dataGroup_hi_lo_503 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_504;
  assign dataGroup_hi_lo_504 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_505;
  assign dataGroup_hi_lo_505 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_506;
  assign dataGroup_hi_lo_506 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_507;
  assign dataGroup_hi_lo_507 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_508;
  assign dataGroup_hi_lo_508 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_509;
  assign dataGroup_hi_lo_509 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_510;
  assign dataGroup_hi_lo_510 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_511;
  assign dataGroup_hi_lo_511 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_512;
  assign dataGroup_hi_lo_512 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_513;
  assign dataGroup_hi_lo_513 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_514;
  assign dataGroup_hi_lo_514 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_515;
  assign dataGroup_hi_lo_515 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_516;
  assign dataGroup_hi_lo_516 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_517;
  assign dataGroup_hi_lo_517 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_518;
  assign dataGroup_hi_lo_518 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_519;
  assign dataGroup_hi_lo_519 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_520;
  assign dataGroup_hi_lo_520 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_521;
  assign dataGroup_hi_lo_521 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_522;
  assign dataGroup_hi_lo_522 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_523;
  assign dataGroup_hi_lo_523 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_524;
  assign dataGroup_hi_lo_524 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_525;
  assign dataGroup_hi_lo_525 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_526;
  assign dataGroup_hi_lo_526 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_527;
  assign dataGroup_hi_lo_527 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_528;
  assign dataGroup_hi_lo_528 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_529;
  assign dataGroup_hi_lo_529 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_530;
  assign dataGroup_hi_lo_530 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_531;
  assign dataGroup_hi_lo_531 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_532;
  assign dataGroup_hi_lo_532 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_533;
  assign dataGroup_hi_lo_533 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_534;
  assign dataGroup_hi_lo_534 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_535;
  assign dataGroup_hi_lo_535 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_536;
  assign dataGroup_hi_lo_536 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_537;
  assign dataGroup_hi_lo_537 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_538;
  assign dataGroup_hi_lo_538 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_539;
  assign dataGroup_hi_lo_539 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_540;
  assign dataGroup_hi_lo_540 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_541;
  assign dataGroup_hi_lo_541 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_542;
  assign dataGroup_hi_lo_542 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_543;
  assign dataGroup_hi_lo_543 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_544;
  assign dataGroup_hi_lo_544 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_545;
  assign dataGroup_hi_lo_545 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_546;
  assign dataGroup_hi_lo_546 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_547;
  assign dataGroup_hi_lo_547 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_548;
  assign dataGroup_hi_lo_548 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_549;
  assign dataGroup_hi_lo_549 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_550;
  assign dataGroup_hi_lo_550 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_551;
  assign dataGroup_hi_lo_551 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_552;
  assign dataGroup_hi_lo_552 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_553;
  assign dataGroup_hi_lo_553 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_554;
  assign dataGroup_hi_lo_554 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_555;
  assign dataGroup_hi_lo_555 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_556;
  assign dataGroup_hi_lo_556 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_557;
  assign dataGroup_hi_lo_557 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_558;
  assign dataGroup_hi_lo_558 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_559;
  assign dataGroup_hi_lo_559 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_560;
  assign dataGroup_hi_lo_560 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_561;
  assign dataGroup_hi_lo_561 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_562;
  assign dataGroup_hi_lo_562 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_563;
  assign dataGroup_hi_lo_563 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_564;
  assign dataGroup_hi_lo_564 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_565;
  assign dataGroup_hi_lo_565 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_566;
  assign dataGroup_hi_lo_566 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_567;
  assign dataGroup_hi_lo_567 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_568;
  assign dataGroup_hi_lo_568 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_569;
  assign dataGroup_hi_lo_569 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_570;
  assign dataGroup_hi_lo_570 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_571;
  assign dataGroup_hi_lo_571 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_572;
  assign dataGroup_hi_lo_572 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_573;
  assign dataGroup_hi_lo_573 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_574;
  assign dataGroup_hi_lo_574 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_575;
  assign dataGroup_hi_lo_575 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_576;
  assign dataGroup_hi_lo_576 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_577;
  assign dataGroup_hi_lo_577 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_578;
  assign dataGroup_hi_lo_578 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_579;
  assign dataGroup_hi_lo_579 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_580;
  assign dataGroup_hi_lo_580 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_581;
  assign dataGroup_hi_lo_581 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_582;
  assign dataGroup_hi_lo_582 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_583;
  assign dataGroup_hi_lo_583 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_584;
  assign dataGroup_hi_lo_584 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_585;
  assign dataGroup_hi_lo_585 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_586;
  assign dataGroup_hi_lo_586 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_587;
  assign dataGroup_hi_lo_587 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_588;
  assign dataGroup_hi_lo_588 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_589;
  assign dataGroup_hi_lo_589 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_590;
  assign dataGroup_hi_lo_590 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_591;
  assign dataGroup_hi_lo_591 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_592;
  assign dataGroup_hi_lo_592 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_593;
  assign dataGroup_hi_lo_593 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_594;
  assign dataGroup_hi_lo_594 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_595;
  assign dataGroup_hi_lo_595 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_596;
  assign dataGroup_hi_lo_596 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_597;
  assign dataGroup_hi_lo_597 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_598;
  assign dataGroup_hi_lo_598 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_599;
  assign dataGroup_hi_lo_599 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_600;
  assign dataGroup_hi_lo_600 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_601;
  assign dataGroup_hi_lo_601 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_602;
  assign dataGroup_hi_lo_602 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_603;
  assign dataGroup_hi_lo_603 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_604;
  assign dataGroup_hi_lo_604 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_605;
  assign dataGroup_hi_lo_605 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_606;
  assign dataGroup_hi_lo_606 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_607;
  assign dataGroup_hi_lo_607 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_608;
  assign dataGroup_hi_lo_608 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_609;
  assign dataGroup_hi_lo_609 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_610;
  assign dataGroup_hi_lo_610 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_611;
  assign dataGroup_hi_lo_611 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_612;
  assign dataGroup_hi_lo_612 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_613;
  assign dataGroup_hi_lo_613 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_614;
  assign dataGroup_hi_lo_614 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_615;
  assign dataGroup_hi_lo_615 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_616;
  assign dataGroup_hi_lo_616 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_617;
  assign dataGroup_hi_lo_617 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_618;
  assign dataGroup_hi_lo_618 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_619;
  assign dataGroup_hi_lo_619 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_620;
  assign dataGroup_hi_lo_620 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_621;
  assign dataGroup_hi_lo_621 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_622;
  assign dataGroup_hi_lo_622 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_623;
  assign dataGroup_hi_lo_623 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_624;
  assign dataGroup_hi_lo_624 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_625;
  assign dataGroup_hi_lo_625 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_626;
  assign dataGroup_hi_lo_626 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_627;
  assign dataGroup_hi_lo_627 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_628;
  assign dataGroup_hi_lo_628 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_629;
  assign dataGroup_hi_lo_629 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_630;
  assign dataGroup_hi_lo_630 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_631;
  assign dataGroup_hi_lo_631 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_632;
  assign dataGroup_hi_lo_632 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_633;
  assign dataGroup_hi_lo_633 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_634;
  assign dataGroup_hi_lo_634 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_635;
  assign dataGroup_hi_lo_635 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_636;
  assign dataGroup_hi_lo_636 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_637;
  assign dataGroup_hi_lo_637 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_638;
  assign dataGroup_hi_lo_638 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_639;
  assign dataGroup_hi_lo_639 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_640;
  assign dataGroup_hi_lo_640 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_641;
  assign dataGroup_hi_lo_641 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_642;
  assign dataGroup_hi_lo_642 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_643;
  assign dataGroup_hi_lo_643 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_644;
  assign dataGroup_hi_lo_644 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_645;
  assign dataGroup_hi_lo_645 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_646;
  assign dataGroup_hi_lo_646 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_647;
  assign dataGroup_hi_lo_647 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_648;
  assign dataGroup_hi_lo_648 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_649;
  assign dataGroup_hi_lo_649 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_650;
  assign dataGroup_hi_lo_650 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_651;
  assign dataGroup_hi_lo_651 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_652;
  assign dataGroup_hi_lo_652 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_653;
  assign dataGroup_hi_lo_653 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_654;
  assign dataGroup_hi_lo_654 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_655;
  assign dataGroup_hi_lo_655 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_656;
  assign dataGroup_hi_lo_656 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_657;
  assign dataGroup_hi_lo_657 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_658;
  assign dataGroup_hi_lo_658 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_659;
  assign dataGroup_hi_lo_659 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_660;
  assign dataGroup_hi_lo_660 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_661;
  assign dataGroup_hi_lo_661 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_662;
  assign dataGroup_hi_lo_662 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_663;
  assign dataGroup_hi_lo_663 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_664;
  assign dataGroup_hi_lo_664 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_665;
  assign dataGroup_hi_lo_665 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_666;
  assign dataGroup_hi_lo_666 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_667;
  assign dataGroup_hi_lo_667 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_668;
  assign dataGroup_hi_lo_668 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_669;
  assign dataGroup_hi_lo_669 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_670;
  assign dataGroup_hi_lo_670 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_671;
  assign dataGroup_hi_lo_671 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_672;
  assign dataGroup_hi_lo_672 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_673;
  assign dataGroup_hi_lo_673 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_674;
  assign dataGroup_hi_lo_674 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_675;
  assign dataGroup_hi_lo_675 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_676;
  assign dataGroup_hi_lo_676 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_677;
  assign dataGroup_hi_lo_677 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_678;
  assign dataGroup_hi_lo_678 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_679;
  assign dataGroup_hi_lo_679 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_680;
  assign dataGroup_hi_lo_680 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_681;
  assign dataGroup_hi_lo_681 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_682;
  assign dataGroup_hi_lo_682 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_683;
  assign dataGroup_hi_lo_683 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_684;
  assign dataGroup_hi_lo_684 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_685;
  assign dataGroup_hi_lo_685 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_686;
  assign dataGroup_hi_lo_686 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_687;
  assign dataGroup_hi_lo_687 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_688;
  assign dataGroup_hi_lo_688 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_689;
  assign dataGroup_hi_lo_689 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_690;
  assign dataGroup_hi_lo_690 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_691;
  assign dataGroup_hi_lo_691 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_692;
  assign dataGroup_hi_lo_692 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_693;
  assign dataGroup_hi_lo_693 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_694;
  assign dataGroup_hi_lo_694 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_695;
  assign dataGroup_hi_lo_695 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_696;
  assign dataGroup_hi_lo_696 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_697;
  assign dataGroup_hi_lo_697 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_698;
  assign dataGroup_hi_lo_698 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_699;
  assign dataGroup_hi_lo_699 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_700;
  assign dataGroup_hi_lo_700 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_701;
  assign dataGroup_hi_lo_701 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_702;
  assign dataGroup_hi_lo_702 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_703;
  assign dataGroup_hi_lo_703 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_704;
  assign dataGroup_hi_lo_704 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_705;
  assign dataGroup_hi_lo_705 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_706;
  assign dataGroup_hi_lo_706 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_707;
  assign dataGroup_hi_lo_707 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_708;
  assign dataGroup_hi_lo_708 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_709;
  assign dataGroup_hi_lo_709 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_710;
  assign dataGroup_hi_lo_710 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_711;
  assign dataGroup_hi_lo_711 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_712;
  assign dataGroup_hi_lo_712 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_713;
  assign dataGroup_hi_lo_713 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_714;
  assign dataGroup_hi_lo_714 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_715;
  assign dataGroup_hi_lo_715 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_716;
  assign dataGroup_hi_lo_716 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_717;
  assign dataGroup_hi_lo_717 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_718;
  assign dataGroup_hi_lo_718 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_719;
  assign dataGroup_hi_lo_719 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_720;
  assign dataGroup_hi_lo_720 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_721;
  assign dataGroup_hi_lo_721 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_722;
  assign dataGroup_hi_lo_722 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_723;
  assign dataGroup_hi_lo_723 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_724;
  assign dataGroup_hi_lo_724 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_725;
  assign dataGroup_hi_lo_725 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_726;
  assign dataGroup_hi_lo_726 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_727;
  assign dataGroup_hi_lo_727 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_728;
  assign dataGroup_hi_lo_728 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_729;
  assign dataGroup_hi_lo_729 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_730;
  assign dataGroup_hi_lo_730 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_731;
  assign dataGroup_hi_lo_731 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_732;
  assign dataGroup_hi_lo_732 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_733;
  assign dataGroup_hi_lo_733 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_734;
  assign dataGroup_hi_lo_734 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_735;
  assign dataGroup_hi_lo_735 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_736;
  assign dataGroup_hi_lo_736 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_737;
  assign dataGroup_hi_lo_737 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_738;
  assign dataGroup_hi_lo_738 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_739;
  assign dataGroup_hi_lo_739 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_740;
  assign dataGroup_hi_lo_740 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_741;
  assign dataGroup_hi_lo_741 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_742;
  assign dataGroup_hi_lo_742 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_743;
  assign dataGroup_hi_lo_743 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_744;
  assign dataGroup_hi_lo_744 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_745;
  assign dataGroup_hi_lo_745 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_746;
  assign dataGroup_hi_lo_746 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_747;
  assign dataGroup_hi_lo_747 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_748;
  assign dataGroup_hi_lo_748 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_749;
  assign dataGroup_hi_lo_749 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_750;
  assign dataGroup_hi_lo_750 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_751;
  assign dataGroup_hi_lo_751 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_752;
  assign dataGroup_hi_lo_752 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_753;
  assign dataGroup_hi_lo_753 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_754;
  assign dataGroup_hi_lo_754 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_755;
  assign dataGroup_hi_lo_755 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_756;
  assign dataGroup_hi_lo_756 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_757;
  assign dataGroup_hi_lo_757 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_758;
  assign dataGroup_hi_lo_758 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_759;
  assign dataGroup_hi_lo_759 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_760;
  assign dataGroup_hi_lo_760 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_761;
  assign dataGroup_hi_lo_761 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_762;
  assign dataGroup_hi_lo_762 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_763;
  assign dataGroup_hi_lo_763 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_764;
  assign dataGroup_hi_lo_764 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_765;
  assign dataGroup_hi_lo_765 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_766;
  assign dataGroup_hi_lo_766 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_767;
  assign dataGroup_hi_lo_767 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_768;
  assign dataGroup_hi_lo_768 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_769;
  assign dataGroup_hi_lo_769 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_770;
  assign dataGroup_hi_lo_770 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_771;
  assign dataGroup_hi_lo_771 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_772;
  assign dataGroup_hi_lo_772 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_773;
  assign dataGroup_hi_lo_773 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_774;
  assign dataGroup_hi_lo_774 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_775;
  assign dataGroup_hi_lo_775 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_776;
  assign dataGroup_hi_lo_776 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_777;
  assign dataGroup_hi_lo_777 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_778;
  assign dataGroup_hi_lo_778 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_779;
  assign dataGroup_hi_lo_779 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_780;
  assign dataGroup_hi_lo_780 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_781;
  assign dataGroup_hi_lo_781 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_782;
  assign dataGroup_hi_lo_782 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_783;
  assign dataGroup_hi_lo_783 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_784;
  assign dataGroup_hi_lo_784 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_785;
  assign dataGroup_hi_lo_785 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_786;
  assign dataGroup_hi_lo_786 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_787;
  assign dataGroup_hi_lo_787 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_788;
  assign dataGroup_hi_lo_788 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_789;
  assign dataGroup_hi_lo_789 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_790;
  assign dataGroup_hi_lo_790 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_791;
  assign dataGroup_hi_lo_791 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_792;
  assign dataGroup_hi_lo_792 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_793;
  assign dataGroup_hi_lo_793 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_794;
  assign dataGroup_hi_lo_794 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_795;
  assign dataGroup_hi_lo_795 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_796;
  assign dataGroup_hi_lo_796 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_797;
  assign dataGroup_hi_lo_797 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_798;
  assign dataGroup_hi_lo_798 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_799;
  assign dataGroup_hi_lo_799 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_800;
  assign dataGroup_hi_lo_800 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_801;
  assign dataGroup_hi_lo_801 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_802;
  assign dataGroup_hi_lo_802 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_803;
  assign dataGroup_hi_lo_803 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_804;
  assign dataGroup_hi_lo_804 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_805;
  assign dataGroup_hi_lo_805 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_806;
  assign dataGroup_hi_lo_806 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_807;
  assign dataGroup_hi_lo_807 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_808;
  assign dataGroup_hi_lo_808 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_809;
  assign dataGroup_hi_lo_809 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_810;
  assign dataGroup_hi_lo_810 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_811;
  assign dataGroup_hi_lo_811 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_812;
  assign dataGroup_hi_lo_812 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_813;
  assign dataGroup_hi_lo_813 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_814;
  assign dataGroup_hi_lo_814 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_815;
  assign dataGroup_hi_lo_815 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_816;
  assign dataGroup_hi_lo_816 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_817;
  assign dataGroup_hi_lo_817 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_818;
  assign dataGroup_hi_lo_818 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_819;
  assign dataGroup_hi_lo_819 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_820;
  assign dataGroup_hi_lo_820 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_821;
  assign dataGroup_hi_lo_821 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_822;
  assign dataGroup_hi_lo_822 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_823;
  assign dataGroup_hi_lo_823 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_824;
  assign dataGroup_hi_lo_824 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_825;
  assign dataGroup_hi_lo_825 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_826;
  assign dataGroup_hi_lo_826 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_827;
  assign dataGroup_hi_lo_827 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_828;
  assign dataGroup_hi_lo_828 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_829;
  assign dataGroup_hi_lo_829 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_830;
  assign dataGroup_hi_lo_830 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_831;
  assign dataGroup_hi_lo_831 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_832;
  assign dataGroup_hi_lo_832 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_833;
  assign dataGroup_hi_lo_833 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_834;
  assign dataGroup_hi_lo_834 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_835;
  assign dataGroup_hi_lo_835 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_836;
  assign dataGroup_hi_lo_836 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_837;
  assign dataGroup_hi_lo_837 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_838;
  assign dataGroup_hi_lo_838 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_839;
  assign dataGroup_hi_lo_839 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_840;
  assign dataGroup_hi_lo_840 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_841;
  assign dataGroup_hi_lo_841 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_842;
  assign dataGroup_hi_lo_842 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_843;
  assign dataGroup_hi_lo_843 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_844;
  assign dataGroup_hi_lo_844 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_845;
  assign dataGroup_hi_lo_845 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_846;
  assign dataGroup_hi_lo_846 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_847;
  assign dataGroup_hi_lo_847 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_848;
  assign dataGroup_hi_lo_848 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_849;
  assign dataGroup_hi_lo_849 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_850;
  assign dataGroup_hi_lo_850 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_851;
  assign dataGroup_hi_lo_851 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_852;
  assign dataGroup_hi_lo_852 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_853;
  assign dataGroup_hi_lo_853 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_854;
  assign dataGroup_hi_lo_854 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_855;
  assign dataGroup_hi_lo_855 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_856;
  assign dataGroup_hi_lo_856 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_857;
  assign dataGroup_hi_lo_857 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_858;
  assign dataGroup_hi_lo_858 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_859;
  assign dataGroup_hi_lo_859 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_860;
  assign dataGroup_hi_lo_860 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_861;
  assign dataGroup_hi_lo_861 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_862;
  assign dataGroup_hi_lo_862 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_863;
  assign dataGroup_hi_lo_863 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_864;
  assign dataGroup_hi_lo_864 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_865;
  assign dataGroup_hi_lo_865 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_866;
  assign dataGroup_hi_lo_866 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_867;
  assign dataGroup_hi_lo_867 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_868;
  assign dataGroup_hi_lo_868 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_869;
  assign dataGroup_hi_lo_869 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_870;
  assign dataGroup_hi_lo_870 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_871;
  assign dataGroup_hi_lo_871 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_872;
  assign dataGroup_hi_lo_872 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_873;
  assign dataGroup_hi_lo_873 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_874;
  assign dataGroup_hi_lo_874 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_875;
  assign dataGroup_hi_lo_875 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_876;
  assign dataGroup_hi_lo_876 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_877;
  assign dataGroup_hi_lo_877 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_878;
  assign dataGroup_hi_lo_878 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_879;
  assign dataGroup_hi_lo_879 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_880;
  assign dataGroup_hi_lo_880 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_881;
  assign dataGroup_hi_lo_881 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_882;
  assign dataGroup_hi_lo_882 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_883;
  assign dataGroup_hi_lo_883 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_884;
  assign dataGroup_hi_lo_884 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_885;
  assign dataGroup_hi_lo_885 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_886;
  assign dataGroup_hi_lo_886 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_887;
  assign dataGroup_hi_lo_887 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_888;
  assign dataGroup_hi_lo_888 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_889;
  assign dataGroup_hi_lo_889 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_890;
  assign dataGroup_hi_lo_890 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_891;
  assign dataGroup_hi_lo_891 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_892;
  assign dataGroup_hi_lo_892 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_893;
  assign dataGroup_hi_lo_893 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_894;
  assign dataGroup_hi_lo_894 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_895;
  assign dataGroup_hi_lo_895 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_896;
  assign dataGroup_hi_lo_896 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_897;
  assign dataGroup_hi_lo_897 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_898;
  assign dataGroup_hi_lo_898 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_899;
  assign dataGroup_hi_lo_899 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_900;
  assign dataGroup_hi_lo_900 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_901;
  assign dataGroup_hi_lo_901 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_902;
  assign dataGroup_hi_lo_902 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_903;
  assign dataGroup_hi_lo_903 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_904;
  assign dataGroup_hi_lo_904 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_905;
  assign dataGroup_hi_lo_905 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_906;
  assign dataGroup_hi_lo_906 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_907;
  assign dataGroup_hi_lo_907 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_908;
  assign dataGroup_hi_lo_908 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_909;
  assign dataGroup_hi_lo_909 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_910;
  assign dataGroup_hi_lo_910 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_911;
  assign dataGroup_hi_lo_911 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_912;
  assign dataGroup_hi_lo_912 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_913;
  assign dataGroup_hi_lo_913 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_914;
  assign dataGroup_hi_lo_914 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_915;
  assign dataGroup_hi_lo_915 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_916;
  assign dataGroup_hi_lo_916 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_917;
  assign dataGroup_hi_lo_917 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_918;
  assign dataGroup_hi_lo_918 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_919;
  assign dataGroup_hi_lo_919 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_920;
  assign dataGroup_hi_lo_920 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_921;
  assign dataGroup_hi_lo_921 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_922;
  assign dataGroup_hi_lo_922 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_923;
  assign dataGroup_hi_lo_923 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_924;
  assign dataGroup_hi_lo_924 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_925;
  assign dataGroup_hi_lo_925 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_926;
  assign dataGroup_hi_lo_926 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_927;
  assign dataGroup_hi_lo_927 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_928;
  assign dataGroup_hi_lo_928 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_929;
  assign dataGroup_hi_lo_929 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_930;
  assign dataGroup_hi_lo_930 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_931;
  assign dataGroup_hi_lo_931 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_932;
  assign dataGroup_hi_lo_932 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_933;
  assign dataGroup_hi_lo_933 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_934;
  assign dataGroup_hi_lo_934 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_935;
  assign dataGroup_hi_lo_935 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_936;
  assign dataGroup_hi_lo_936 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_937;
  assign dataGroup_hi_lo_937 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_938;
  assign dataGroup_hi_lo_938 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_939;
  assign dataGroup_hi_lo_939 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_940;
  assign dataGroup_hi_lo_940 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_941;
  assign dataGroup_hi_lo_941 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_942;
  assign dataGroup_hi_lo_942 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_943;
  assign dataGroup_hi_lo_943 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_944;
  assign dataGroup_hi_lo_944 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_945;
  assign dataGroup_hi_lo_945 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_946;
  assign dataGroup_hi_lo_946 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_947;
  assign dataGroup_hi_lo_947 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_948;
  assign dataGroup_hi_lo_948 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_949;
  assign dataGroup_hi_lo_949 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_950;
  assign dataGroup_hi_lo_950 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_951;
  assign dataGroup_hi_lo_951 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_952;
  assign dataGroup_hi_lo_952 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_953;
  assign dataGroup_hi_lo_953 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_954;
  assign dataGroup_hi_lo_954 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_955;
  assign dataGroup_hi_lo_955 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_956;
  assign dataGroup_hi_lo_956 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_957;
  assign dataGroup_hi_lo_957 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_958;
  assign dataGroup_hi_lo_958 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_959;
  assign dataGroup_hi_lo_959 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_960;
  assign dataGroup_hi_lo_960 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_961;
  assign dataGroup_hi_lo_961 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_962;
  assign dataGroup_hi_lo_962 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_963;
  assign dataGroup_hi_lo_963 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_964;
  assign dataGroup_hi_lo_964 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_965;
  assign dataGroup_hi_lo_965 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_966;
  assign dataGroup_hi_lo_966 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_967;
  assign dataGroup_hi_lo_967 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_968;
  assign dataGroup_hi_lo_968 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_969;
  assign dataGroup_hi_lo_969 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_970;
  assign dataGroup_hi_lo_970 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_971;
  assign dataGroup_hi_lo_971 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_972;
  assign dataGroup_hi_lo_972 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_973;
  assign dataGroup_hi_lo_973 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_974;
  assign dataGroup_hi_lo_974 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_975;
  assign dataGroup_hi_lo_975 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_976;
  assign dataGroup_hi_lo_976 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_977;
  assign dataGroup_hi_lo_977 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_978;
  assign dataGroup_hi_lo_978 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_979;
  assign dataGroup_hi_lo_979 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_980;
  assign dataGroup_hi_lo_980 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_981;
  assign dataGroup_hi_lo_981 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_982;
  assign dataGroup_hi_lo_982 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_983;
  assign dataGroup_hi_lo_983 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_984;
  assign dataGroup_hi_lo_984 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_985;
  assign dataGroup_hi_lo_985 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_986;
  assign dataGroup_hi_lo_986 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_987;
  assign dataGroup_hi_lo_987 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_988;
  assign dataGroup_hi_lo_988 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_989;
  assign dataGroup_hi_lo_989 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_990;
  assign dataGroup_hi_lo_990 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_991;
  assign dataGroup_hi_lo_991 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_992;
  assign dataGroup_hi_lo_992 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_993;
  assign dataGroup_hi_lo_993 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_994;
  assign dataGroup_hi_lo_994 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_995;
  assign dataGroup_hi_lo_995 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_996;
  assign dataGroup_hi_lo_996 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_997;
  assign dataGroup_hi_lo_997 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_998;
  assign dataGroup_hi_lo_998 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_999;
  assign dataGroup_hi_lo_999 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1000;
  assign dataGroup_hi_lo_1000 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1001;
  assign dataGroup_hi_lo_1001 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1002;
  assign dataGroup_hi_lo_1002 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1003;
  assign dataGroup_hi_lo_1003 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1004;
  assign dataGroup_hi_lo_1004 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1005;
  assign dataGroup_hi_lo_1005 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1006;
  assign dataGroup_hi_lo_1006 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1007;
  assign dataGroup_hi_lo_1007 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1008;
  assign dataGroup_hi_lo_1008 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1009;
  assign dataGroup_hi_lo_1009 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1010;
  assign dataGroup_hi_lo_1010 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1011;
  assign dataGroup_hi_lo_1011 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1012;
  assign dataGroup_hi_lo_1012 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1013;
  assign dataGroup_hi_lo_1013 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1014;
  assign dataGroup_hi_lo_1014 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1015;
  assign dataGroup_hi_lo_1015 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1016;
  assign dataGroup_hi_lo_1016 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1017;
  assign dataGroup_hi_lo_1017 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1018;
  assign dataGroup_hi_lo_1018 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1019;
  assign dataGroup_hi_lo_1019 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1020;
  assign dataGroup_hi_lo_1020 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1021;
  assign dataGroup_hi_lo_1021 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1022;
  assign dataGroup_hi_lo_1022 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1023;
  assign dataGroup_hi_lo_1023 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1024;
  assign dataGroup_hi_lo_1024 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1025;
  assign dataGroup_hi_lo_1025 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1026;
  assign dataGroup_hi_lo_1026 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1027;
  assign dataGroup_hi_lo_1027 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1028;
  assign dataGroup_hi_lo_1028 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1029;
  assign dataGroup_hi_lo_1029 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1030;
  assign dataGroup_hi_lo_1030 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1031;
  assign dataGroup_hi_lo_1031 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1032;
  assign dataGroup_hi_lo_1032 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1033;
  assign dataGroup_hi_lo_1033 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1034;
  assign dataGroup_hi_lo_1034 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1035;
  assign dataGroup_hi_lo_1035 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1036;
  assign dataGroup_hi_lo_1036 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1037;
  assign dataGroup_hi_lo_1037 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1038;
  assign dataGroup_hi_lo_1038 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1039;
  assign dataGroup_hi_lo_1039 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1040;
  assign dataGroup_hi_lo_1040 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1041;
  assign dataGroup_hi_lo_1041 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1042;
  assign dataGroup_hi_lo_1042 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1043;
  assign dataGroup_hi_lo_1043 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1044;
  assign dataGroup_hi_lo_1044 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1045;
  assign dataGroup_hi_lo_1045 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1046;
  assign dataGroup_hi_lo_1046 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1047;
  assign dataGroup_hi_lo_1047 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1048;
  assign dataGroup_hi_lo_1048 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1049;
  assign dataGroup_hi_lo_1049 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1050;
  assign dataGroup_hi_lo_1050 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1051;
  assign dataGroup_hi_lo_1051 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1052;
  assign dataGroup_hi_lo_1052 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1053;
  assign dataGroup_hi_lo_1053 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1054;
  assign dataGroup_hi_lo_1054 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1055;
  assign dataGroup_hi_lo_1055 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1056;
  assign dataGroup_hi_lo_1056 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1057;
  assign dataGroup_hi_lo_1057 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1058;
  assign dataGroup_hi_lo_1058 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1059;
  assign dataGroup_hi_lo_1059 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1060;
  assign dataGroup_hi_lo_1060 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1061;
  assign dataGroup_hi_lo_1061 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1062;
  assign dataGroup_hi_lo_1062 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1063;
  assign dataGroup_hi_lo_1063 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1064;
  assign dataGroup_hi_lo_1064 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1065;
  assign dataGroup_hi_lo_1065 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1066;
  assign dataGroup_hi_lo_1066 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1067;
  assign dataGroup_hi_lo_1067 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1068;
  assign dataGroup_hi_lo_1068 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1069;
  assign dataGroup_hi_lo_1069 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1070;
  assign dataGroup_hi_lo_1070 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1071;
  assign dataGroup_hi_lo_1071 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1072;
  assign dataGroup_hi_lo_1072 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1073;
  assign dataGroup_hi_lo_1073 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1074;
  assign dataGroup_hi_lo_1074 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1075;
  assign dataGroup_hi_lo_1075 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1076;
  assign dataGroup_hi_lo_1076 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1077;
  assign dataGroup_hi_lo_1077 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1078;
  assign dataGroup_hi_lo_1078 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1079;
  assign dataGroup_hi_lo_1079 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1080;
  assign dataGroup_hi_lo_1080 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1081;
  assign dataGroup_hi_lo_1081 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1082;
  assign dataGroup_hi_lo_1082 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1083;
  assign dataGroup_hi_lo_1083 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1084;
  assign dataGroup_hi_lo_1084 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1085;
  assign dataGroup_hi_lo_1085 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1086;
  assign dataGroup_hi_lo_1086 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1087;
  assign dataGroup_hi_lo_1087 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1088;
  assign dataGroup_hi_lo_1088 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1089;
  assign dataGroup_hi_lo_1089 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1090;
  assign dataGroup_hi_lo_1090 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1091;
  assign dataGroup_hi_lo_1091 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1092;
  assign dataGroup_hi_lo_1092 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1093;
  assign dataGroup_hi_lo_1093 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1094;
  assign dataGroup_hi_lo_1094 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1095;
  assign dataGroup_hi_lo_1095 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1096;
  assign dataGroup_hi_lo_1096 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1097;
  assign dataGroup_hi_lo_1097 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1098;
  assign dataGroup_hi_lo_1098 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1099;
  assign dataGroup_hi_lo_1099 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1100;
  assign dataGroup_hi_lo_1100 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1101;
  assign dataGroup_hi_lo_1101 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1102;
  assign dataGroup_hi_lo_1102 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1103;
  assign dataGroup_hi_lo_1103 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1104;
  assign dataGroup_hi_lo_1104 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1105;
  assign dataGroup_hi_lo_1105 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1106;
  assign dataGroup_hi_lo_1106 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1107;
  assign dataGroup_hi_lo_1107 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1108;
  assign dataGroup_hi_lo_1108 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1109;
  assign dataGroup_hi_lo_1109 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1110;
  assign dataGroup_hi_lo_1110 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1111;
  assign dataGroup_hi_lo_1111 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1112;
  assign dataGroup_hi_lo_1112 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1113;
  assign dataGroup_hi_lo_1113 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1114;
  assign dataGroup_hi_lo_1114 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1115;
  assign dataGroup_hi_lo_1115 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1116;
  assign dataGroup_hi_lo_1116 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1117;
  assign dataGroup_hi_lo_1117 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1118;
  assign dataGroup_hi_lo_1118 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1119;
  assign dataGroup_hi_lo_1119 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1120;
  assign dataGroup_hi_lo_1120 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1121;
  assign dataGroup_hi_lo_1121 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1122;
  assign dataGroup_hi_lo_1122 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1123;
  assign dataGroup_hi_lo_1123 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1124;
  assign dataGroup_hi_lo_1124 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1125;
  assign dataGroup_hi_lo_1125 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1126;
  assign dataGroup_hi_lo_1126 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1127;
  assign dataGroup_hi_lo_1127 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1128;
  assign dataGroup_hi_lo_1128 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1129;
  assign dataGroup_hi_lo_1129 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1130;
  assign dataGroup_hi_lo_1130 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1131;
  assign dataGroup_hi_lo_1131 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1132;
  assign dataGroup_hi_lo_1132 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1133;
  assign dataGroup_hi_lo_1133 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1134;
  assign dataGroup_hi_lo_1134 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1135;
  assign dataGroup_hi_lo_1135 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1136;
  assign dataGroup_hi_lo_1136 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1137;
  assign dataGroup_hi_lo_1137 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1138;
  assign dataGroup_hi_lo_1138 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1139;
  assign dataGroup_hi_lo_1139 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1140;
  assign dataGroup_hi_lo_1140 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1141;
  assign dataGroup_hi_lo_1141 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1142;
  assign dataGroup_hi_lo_1142 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1143;
  assign dataGroup_hi_lo_1143 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1144;
  assign dataGroup_hi_lo_1144 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1145;
  assign dataGroup_hi_lo_1145 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1146;
  assign dataGroup_hi_lo_1146 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1147;
  assign dataGroup_hi_lo_1147 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1148;
  assign dataGroup_hi_lo_1148 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1149;
  assign dataGroup_hi_lo_1149 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1150;
  assign dataGroup_hi_lo_1150 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1151;
  assign dataGroup_hi_lo_1151 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1152;
  assign dataGroup_hi_lo_1152 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1153;
  assign dataGroup_hi_lo_1153 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1154;
  assign dataGroup_hi_lo_1154 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1155;
  assign dataGroup_hi_lo_1155 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1156;
  assign dataGroup_hi_lo_1156 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1157;
  assign dataGroup_hi_lo_1157 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1158;
  assign dataGroup_hi_lo_1158 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1159;
  assign dataGroup_hi_lo_1159 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1160;
  assign dataGroup_hi_lo_1160 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1161;
  assign dataGroup_hi_lo_1161 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1162;
  assign dataGroup_hi_lo_1162 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1163;
  assign dataGroup_hi_lo_1163 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1164;
  assign dataGroup_hi_lo_1164 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1165;
  assign dataGroup_hi_lo_1165 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1166;
  assign dataGroup_hi_lo_1166 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1167;
  assign dataGroup_hi_lo_1167 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1168;
  assign dataGroup_hi_lo_1168 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1169;
  assign dataGroup_hi_lo_1169 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1170;
  assign dataGroup_hi_lo_1170 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1171;
  assign dataGroup_hi_lo_1171 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1172;
  assign dataGroup_hi_lo_1172 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1173;
  assign dataGroup_hi_lo_1173 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1174;
  assign dataGroup_hi_lo_1174 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1175;
  assign dataGroup_hi_lo_1175 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1176;
  assign dataGroup_hi_lo_1176 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1177;
  assign dataGroup_hi_lo_1177 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1178;
  assign dataGroup_hi_lo_1178 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1179;
  assign dataGroup_hi_lo_1179 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1180;
  assign dataGroup_hi_lo_1180 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1181;
  assign dataGroup_hi_lo_1181 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1182;
  assign dataGroup_hi_lo_1182 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1183;
  assign dataGroup_hi_lo_1183 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1184;
  assign dataGroup_hi_lo_1184 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1185;
  assign dataGroup_hi_lo_1185 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1186;
  assign dataGroup_hi_lo_1186 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1187;
  assign dataGroup_hi_lo_1187 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1188;
  assign dataGroup_hi_lo_1188 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1189;
  assign dataGroup_hi_lo_1189 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1190;
  assign dataGroup_hi_lo_1190 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1191;
  assign dataGroup_hi_lo_1191 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1192;
  assign dataGroup_hi_lo_1192 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1193;
  assign dataGroup_hi_lo_1193 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1194;
  assign dataGroup_hi_lo_1194 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1195;
  assign dataGroup_hi_lo_1195 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1196;
  assign dataGroup_hi_lo_1196 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1197;
  assign dataGroup_hi_lo_1197 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1198;
  assign dataGroup_hi_lo_1198 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1199;
  assign dataGroup_hi_lo_1199 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1200;
  assign dataGroup_hi_lo_1200 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1201;
  assign dataGroup_hi_lo_1201 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1202;
  assign dataGroup_hi_lo_1202 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1203;
  assign dataGroup_hi_lo_1203 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1204;
  assign dataGroup_hi_lo_1204 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1205;
  assign dataGroup_hi_lo_1205 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1206;
  assign dataGroup_hi_lo_1206 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1207;
  assign dataGroup_hi_lo_1207 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1208;
  assign dataGroup_hi_lo_1208 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1209;
  assign dataGroup_hi_lo_1209 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1210;
  assign dataGroup_hi_lo_1210 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1211;
  assign dataGroup_hi_lo_1211 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1212;
  assign dataGroup_hi_lo_1212 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1213;
  assign dataGroup_hi_lo_1213 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1214;
  assign dataGroup_hi_lo_1214 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1215;
  assign dataGroup_hi_lo_1215 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1216;
  assign dataGroup_hi_lo_1216 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1217;
  assign dataGroup_hi_lo_1217 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1218;
  assign dataGroup_hi_lo_1218 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1219;
  assign dataGroup_hi_lo_1219 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1220;
  assign dataGroup_hi_lo_1220 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1221;
  assign dataGroup_hi_lo_1221 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1222;
  assign dataGroup_hi_lo_1222 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1223;
  assign dataGroup_hi_lo_1223 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1224;
  assign dataGroup_hi_lo_1224 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1225;
  assign dataGroup_hi_lo_1225 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1226;
  assign dataGroup_hi_lo_1226 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1227;
  assign dataGroup_hi_lo_1227 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1228;
  assign dataGroup_hi_lo_1228 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1229;
  assign dataGroup_hi_lo_1229 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1230;
  assign dataGroup_hi_lo_1230 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1231;
  assign dataGroup_hi_lo_1231 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1232;
  assign dataGroup_hi_lo_1232 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1233;
  assign dataGroup_hi_lo_1233 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1234;
  assign dataGroup_hi_lo_1234 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1235;
  assign dataGroup_hi_lo_1235 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1236;
  assign dataGroup_hi_lo_1236 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1237;
  assign dataGroup_hi_lo_1237 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1238;
  assign dataGroup_hi_lo_1238 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1239;
  assign dataGroup_hi_lo_1239 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1240;
  assign dataGroup_hi_lo_1240 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1241;
  assign dataGroup_hi_lo_1241 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1242;
  assign dataGroup_hi_lo_1242 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1243;
  assign dataGroup_hi_lo_1243 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1244;
  assign dataGroup_hi_lo_1244 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1245;
  assign dataGroup_hi_lo_1245 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1246;
  assign dataGroup_hi_lo_1246 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1247;
  assign dataGroup_hi_lo_1247 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1248;
  assign dataGroup_hi_lo_1248 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1249;
  assign dataGroup_hi_lo_1249 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1250;
  assign dataGroup_hi_lo_1250 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1251;
  assign dataGroup_hi_lo_1251 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1252;
  assign dataGroup_hi_lo_1252 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1253;
  assign dataGroup_hi_lo_1253 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1254;
  assign dataGroup_hi_lo_1254 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1255;
  assign dataGroup_hi_lo_1255 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1256;
  assign dataGroup_hi_lo_1256 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1257;
  assign dataGroup_hi_lo_1257 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1258;
  assign dataGroup_hi_lo_1258 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1259;
  assign dataGroup_hi_lo_1259 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1260;
  assign dataGroup_hi_lo_1260 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1261;
  assign dataGroup_hi_lo_1261 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1262;
  assign dataGroup_hi_lo_1262 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1263;
  assign dataGroup_hi_lo_1263 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1264;
  assign dataGroup_hi_lo_1264 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1265;
  assign dataGroup_hi_lo_1265 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1266;
  assign dataGroup_hi_lo_1266 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1267;
  assign dataGroup_hi_lo_1267 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1268;
  assign dataGroup_hi_lo_1268 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1269;
  assign dataGroup_hi_lo_1269 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1270;
  assign dataGroup_hi_lo_1270 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1271;
  assign dataGroup_hi_lo_1271 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1272;
  assign dataGroup_hi_lo_1272 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1273;
  assign dataGroup_hi_lo_1273 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1274;
  assign dataGroup_hi_lo_1274 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1275;
  assign dataGroup_hi_lo_1275 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1276;
  assign dataGroup_hi_lo_1276 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1277;
  assign dataGroup_hi_lo_1277 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1278;
  assign dataGroup_hi_lo_1278 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1279;
  assign dataGroup_hi_lo_1279 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1280;
  assign dataGroup_hi_lo_1280 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1281;
  assign dataGroup_hi_lo_1281 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1282;
  assign dataGroup_hi_lo_1282 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1283;
  assign dataGroup_hi_lo_1283 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1284;
  assign dataGroup_hi_lo_1284 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1285;
  assign dataGroup_hi_lo_1285 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1286;
  assign dataGroup_hi_lo_1286 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1287;
  assign dataGroup_hi_lo_1287 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1288;
  assign dataGroup_hi_lo_1288 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1289;
  assign dataGroup_hi_lo_1289 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1290;
  assign dataGroup_hi_lo_1290 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1291;
  assign dataGroup_hi_lo_1291 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1292;
  assign dataGroup_hi_lo_1292 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1293;
  assign dataGroup_hi_lo_1293 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1294;
  assign dataGroup_hi_lo_1294 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1295;
  assign dataGroup_hi_lo_1295 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1296;
  assign dataGroup_hi_lo_1296 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1297;
  assign dataGroup_hi_lo_1297 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1298;
  assign dataGroup_hi_lo_1298 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1299;
  assign dataGroup_hi_lo_1299 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1300;
  assign dataGroup_hi_lo_1300 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1301;
  assign dataGroup_hi_lo_1301 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1302;
  assign dataGroup_hi_lo_1302 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1303;
  assign dataGroup_hi_lo_1303 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1304;
  assign dataGroup_hi_lo_1304 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1305;
  assign dataGroup_hi_lo_1305 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1306;
  assign dataGroup_hi_lo_1306 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1307;
  assign dataGroup_hi_lo_1307 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1308;
  assign dataGroup_hi_lo_1308 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1309;
  assign dataGroup_hi_lo_1309 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1310;
  assign dataGroup_hi_lo_1310 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1311;
  assign dataGroup_hi_lo_1311 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1312;
  assign dataGroup_hi_lo_1312 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1313;
  assign dataGroup_hi_lo_1313 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1314;
  assign dataGroup_hi_lo_1314 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1315;
  assign dataGroup_hi_lo_1315 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1316;
  assign dataGroup_hi_lo_1316 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1317;
  assign dataGroup_hi_lo_1317 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1318;
  assign dataGroup_hi_lo_1318 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1319;
  assign dataGroup_hi_lo_1319 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1320;
  assign dataGroup_hi_lo_1320 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1321;
  assign dataGroup_hi_lo_1321 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1322;
  assign dataGroup_hi_lo_1322 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1323;
  assign dataGroup_hi_lo_1323 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1324;
  assign dataGroup_hi_lo_1324 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1325;
  assign dataGroup_hi_lo_1325 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1326;
  assign dataGroup_hi_lo_1326 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1327;
  assign dataGroup_hi_lo_1327 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1328;
  assign dataGroup_hi_lo_1328 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1329;
  assign dataGroup_hi_lo_1329 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1330;
  assign dataGroup_hi_lo_1330 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1331;
  assign dataGroup_hi_lo_1331 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1332;
  assign dataGroup_hi_lo_1332 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1333;
  assign dataGroup_hi_lo_1333 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1334;
  assign dataGroup_hi_lo_1334 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1335;
  assign dataGroup_hi_lo_1335 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1336;
  assign dataGroup_hi_lo_1336 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1337;
  assign dataGroup_hi_lo_1337 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1338;
  assign dataGroup_hi_lo_1338 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1339;
  assign dataGroup_hi_lo_1339 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1340;
  assign dataGroup_hi_lo_1340 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1341;
  assign dataGroup_hi_lo_1341 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1342;
  assign dataGroup_hi_lo_1342 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1343;
  assign dataGroup_hi_lo_1343 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1344;
  assign dataGroup_hi_lo_1344 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1345;
  assign dataGroup_hi_lo_1345 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1346;
  assign dataGroup_hi_lo_1346 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1347;
  assign dataGroup_hi_lo_1347 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1348;
  assign dataGroup_hi_lo_1348 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1349;
  assign dataGroup_hi_lo_1349 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1350;
  assign dataGroup_hi_lo_1350 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1351;
  assign dataGroup_hi_lo_1351 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1352;
  assign dataGroup_hi_lo_1352 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1353;
  assign dataGroup_hi_lo_1353 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1354;
  assign dataGroup_hi_lo_1354 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1355;
  assign dataGroup_hi_lo_1355 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1356;
  assign dataGroup_hi_lo_1356 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1357;
  assign dataGroup_hi_lo_1357 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1358;
  assign dataGroup_hi_lo_1358 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1359;
  assign dataGroup_hi_lo_1359 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1360;
  assign dataGroup_hi_lo_1360 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1361;
  assign dataGroup_hi_lo_1361 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1362;
  assign dataGroup_hi_lo_1362 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1363;
  assign dataGroup_hi_lo_1363 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1364;
  assign dataGroup_hi_lo_1364 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1365;
  assign dataGroup_hi_lo_1365 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1366;
  assign dataGroup_hi_lo_1366 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1367;
  assign dataGroup_hi_lo_1367 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1368;
  assign dataGroup_hi_lo_1368 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1369;
  assign dataGroup_hi_lo_1369 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1370;
  assign dataGroup_hi_lo_1370 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1371;
  assign dataGroup_hi_lo_1371 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1372;
  assign dataGroup_hi_lo_1372 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1373;
  assign dataGroup_hi_lo_1373 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1374;
  assign dataGroup_hi_lo_1374 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1375;
  assign dataGroup_hi_lo_1375 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1376;
  assign dataGroup_hi_lo_1376 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1377;
  assign dataGroup_hi_lo_1377 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1378;
  assign dataGroup_hi_lo_1378 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1379;
  assign dataGroup_hi_lo_1379 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1380;
  assign dataGroup_hi_lo_1380 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1381;
  assign dataGroup_hi_lo_1381 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1382;
  assign dataGroup_hi_lo_1382 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1383;
  assign dataGroup_hi_lo_1383 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1384;
  assign dataGroup_hi_lo_1384 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1385;
  assign dataGroup_hi_lo_1385 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1386;
  assign dataGroup_hi_lo_1386 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1387;
  assign dataGroup_hi_lo_1387 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1388;
  assign dataGroup_hi_lo_1388 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1389;
  assign dataGroup_hi_lo_1389 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1390;
  assign dataGroup_hi_lo_1390 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1391;
  assign dataGroup_hi_lo_1391 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1392;
  assign dataGroup_hi_lo_1392 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1393;
  assign dataGroup_hi_lo_1393 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1394;
  assign dataGroup_hi_lo_1394 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1395;
  assign dataGroup_hi_lo_1395 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1396;
  assign dataGroup_hi_lo_1396 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1397;
  assign dataGroup_hi_lo_1397 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1398;
  assign dataGroup_hi_lo_1398 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1399;
  assign dataGroup_hi_lo_1399 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1400;
  assign dataGroup_hi_lo_1400 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1401;
  assign dataGroup_hi_lo_1401 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1402;
  assign dataGroup_hi_lo_1402 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1403;
  assign dataGroup_hi_lo_1403 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1404;
  assign dataGroup_hi_lo_1404 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1405;
  assign dataGroup_hi_lo_1405 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1406;
  assign dataGroup_hi_lo_1406 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1407;
  assign dataGroup_hi_lo_1407 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1408;
  assign dataGroup_hi_lo_1408 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1409;
  assign dataGroup_hi_lo_1409 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1410;
  assign dataGroup_hi_lo_1410 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1411;
  assign dataGroup_hi_lo_1411 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1412;
  assign dataGroup_hi_lo_1412 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1413;
  assign dataGroup_hi_lo_1413 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1414;
  assign dataGroup_hi_lo_1414 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1415;
  assign dataGroup_hi_lo_1415 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1416;
  assign dataGroup_hi_lo_1416 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1417;
  assign dataGroup_hi_lo_1417 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1418;
  assign dataGroup_hi_lo_1418 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1419;
  assign dataGroup_hi_lo_1419 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1420;
  assign dataGroup_hi_lo_1420 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1421;
  assign dataGroup_hi_lo_1421 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1422;
  assign dataGroup_hi_lo_1422 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1423;
  assign dataGroup_hi_lo_1423 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1424;
  assign dataGroup_hi_lo_1424 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1425;
  assign dataGroup_hi_lo_1425 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1426;
  assign dataGroup_hi_lo_1426 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1427;
  assign dataGroup_hi_lo_1427 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1428;
  assign dataGroup_hi_lo_1428 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1429;
  assign dataGroup_hi_lo_1429 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1430;
  assign dataGroup_hi_lo_1430 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1431;
  assign dataGroup_hi_lo_1431 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1432;
  assign dataGroup_hi_lo_1432 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1433;
  assign dataGroup_hi_lo_1433 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1434;
  assign dataGroup_hi_lo_1434 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1435;
  assign dataGroup_hi_lo_1435 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1436;
  assign dataGroup_hi_lo_1436 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1437;
  assign dataGroup_hi_lo_1437 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1438;
  assign dataGroup_hi_lo_1438 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1439;
  assign dataGroup_hi_lo_1439 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1440;
  assign dataGroup_hi_lo_1440 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1441;
  assign dataGroup_hi_lo_1441 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1442;
  assign dataGroup_hi_lo_1442 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1443;
  assign dataGroup_hi_lo_1443 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1444;
  assign dataGroup_hi_lo_1444 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1445;
  assign dataGroup_hi_lo_1445 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1446;
  assign dataGroup_hi_lo_1446 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1447;
  assign dataGroup_hi_lo_1447 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1448;
  assign dataGroup_hi_lo_1448 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1449;
  assign dataGroup_hi_lo_1449 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1450;
  assign dataGroup_hi_lo_1450 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1451;
  assign dataGroup_hi_lo_1451 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1452;
  assign dataGroup_hi_lo_1452 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1453;
  assign dataGroup_hi_lo_1453 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1454;
  assign dataGroup_hi_lo_1454 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1455;
  assign dataGroup_hi_lo_1455 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1456;
  assign dataGroup_hi_lo_1456 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1457;
  assign dataGroup_hi_lo_1457 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1458;
  assign dataGroup_hi_lo_1458 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1459;
  assign dataGroup_hi_lo_1459 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1460;
  assign dataGroup_hi_lo_1460 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1461;
  assign dataGroup_hi_lo_1461 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1462;
  assign dataGroup_hi_lo_1462 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1463;
  assign dataGroup_hi_lo_1463 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1464;
  assign dataGroup_hi_lo_1464 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1465;
  assign dataGroup_hi_lo_1465 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1466;
  assign dataGroup_hi_lo_1466 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1467;
  assign dataGroup_hi_lo_1467 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1468;
  assign dataGroup_hi_lo_1468 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1469;
  assign dataGroup_hi_lo_1469 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1470;
  assign dataGroup_hi_lo_1470 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1471;
  assign dataGroup_hi_lo_1471 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1472;
  assign dataGroup_hi_lo_1472 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1473;
  assign dataGroup_hi_lo_1473 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1474;
  assign dataGroup_hi_lo_1474 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1475;
  assign dataGroup_hi_lo_1475 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1476;
  assign dataGroup_hi_lo_1476 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1477;
  assign dataGroup_hi_lo_1477 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1478;
  assign dataGroup_hi_lo_1478 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1479;
  assign dataGroup_hi_lo_1479 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1480;
  assign dataGroup_hi_lo_1480 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1481;
  assign dataGroup_hi_lo_1481 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1482;
  assign dataGroup_hi_lo_1482 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1483;
  assign dataGroup_hi_lo_1483 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1484;
  assign dataGroup_hi_lo_1484 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1485;
  assign dataGroup_hi_lo_1485 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1486;
  assign dataGroup_hi_lo_1486 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1487;
  assign dataGroup_hi_lo_1487 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1488;
  assign dataGroup_hi_lo_1488 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1489;
  assign dataGroup_hi_lo_1489 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1490;
  assign dataGroup_hi_lo_1490 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1491;
  assign dataGroup_hi_lo_1491 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1492;
  assign dataGroup_hi_lo_1492 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1493;
  assign dataGroup_hi_lo_1493 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1494;
  assign dataGroup_hi_lo_1494 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1495;
  assign dataGroup_hi_lo_1495 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1496;
  assign dataGroup_hi_lo_1496 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1497;
  assign dataGroup_hi_lo_1497 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1498;
  assign dataGroup_hi_lo_1498 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1499;
  assign dataGroup_hi_lo_1499 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1500;
  assign dataGroup_hi_lo_1500 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1501;
  assign dataGroup_hi_lo_1501 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1502;
  assign dataGroup_hi_lo_1502 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1503;
  assign dataGroup_hi_lo_1503 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1504;
  assign dataGroup_hi_lo_1504 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1505;
  assign dataGroup_hi_lo_1505 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1506;
  assign dataGroup_hi_lo_1506 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1507;
  assign dataGroup_hi_lo_1507 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1508;
  assign dataGroup_hi_lo_1508 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1509;
  assign dataGroup_hi_lo_1509 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1510;
  assign dataGroup_hi_lo_1510 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1511;
  assign dataGroup_hi_lo_1511 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1512;
  assign dataGroup_hi_lo_1512 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1513;
  assign dataGroup_hi_lo_1513 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1514;
  assign dataGroup_hi_lo_1514 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1515;
  assign dataGroup_hi_lo_1515 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1516;
  assign dataGroup_hi_lo_1516 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1517;
  assign dataGroup_hi_lo_1517 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1518;
  assign dataGroup_hi_lo_1518 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1519;
  assign dataGroup_hi_lo_1519 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1520;
  assign dataGroup_hi_lo_1520 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1521;
  assign dataGroup_hi_lo_1521 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1522;
  assign dataGroup_hi_lo_1522 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1523;
  assign dataGroup_hi_lo_1523 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1524;
  assign dataGroup_hi_lo_1524 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1525;
  assign dataGroup_hi_lo_1525 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1526;
  assign dataGroup_hi_lo_1526 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1527;
  assign dataGroup_hi_lo_1527 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1528;
  assign dataGroup_hi_lo_1528 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1529;
  assign dataGroup_hi_lo_1529 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1530;
  assign dataGroup_hi_lo_1530 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1531;
  assign dataGroup_hi_lo_1531 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1532;
  assign dataGroup_hi_lo_1532 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1533;
  assign dataGroup_hi_lo_1533 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1534;
  assign dataGroup_hi_lo_1534 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1535;
  assign dataGroup_hi_lo_1535 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1536;
  assign dataGroup_hi_lo_1536 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1537;
  assign dataGroup_hi_lo_1537 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1538;
  assign dataGroup_hi_lo_1538 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1539;
  assign dataGroup_hi_lo_1539 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1540;
  assign dataGroup_hi_lo_1540 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1541;
  assign dataGroup_hi_lo_1541 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1542;
  assign dataGroup_hi_lo_1542 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1543;
  assign dataGroup_hi_lo_1543 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1544;
  assign dataGroup_hi_lo_1544 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1545;
  assign dataGroup_hi_lo_1545 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1546;
  assign dataGroup_hi_lo_1546 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1547;
  assign dataGroup_hi_lo_1547 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1548;
  assign dataGroup_hi_lo_1548 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1549;
  assign dataGroup_hi_lo_1549 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1550;
  assign dataGroup_hi_lo_1550 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1551;
  assign dataGroup_hi_lo_1551 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1552;
  assign dataGroup_hi_lo_1552 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1553;
  assign dataGroup_hi_lo_1553 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1554;
  assign dataGroup_hi_lo_1554 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1555;
  assign dataGroup_hi_lo_1555 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1556;
  assign dataGroup_hi_lo_1556 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1557;
  assign dataGroup_hi_lo_1557 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1558;
  assign dataGroup_hi_lo_1558 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1559;
  assign dataGroup_hi_lo_1559 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1560;
  assign dataGroup_hi_lo_1560 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1561;
  assign dataGroup_hi_lo_1561 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1562;
  assign dataGroup_hi_lo_1562 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1563;
  assign dataGroup_hi_lo_1563 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1564;
  assign dataGroup_hi_lo_1564 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1565;
  assign dataGroup_hi_lo_1565 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1566;
  assign dataGroup_hi_lo_1566 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1567;
  assign dataGroup_hi_lo_1567 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1568;
  assign dataGroup_hi_lo_1568 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1569;
  assign dataGroup_hi_lo_1569 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1570;
  assign dataGroup_hi_lo_1570 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1571;
  assign dataGroup_hi_lo_1571 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1572;
  assign dataGroup_hi_lo_1572 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1573;
  assign dataGroup_hi_lo_1573 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1574;
  assign dataGroup_hi_lo_1574 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1575;
  assign dataGroup_hi_lo_1575 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1576;
  assign dataGroup_hi_lo_1576 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1577;
  assign dataGroup_hi_lo_1577 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1578;
  assign dataGroup_hi_lo_1578 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1579;
  assign dataGroup_hi_lo_1579 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1580;
  assign dataGroup_hi_lo_1580 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1581;
  assign dataGroup_hi_lo_1581 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1582;
  assign dataGroup_hi_lo_1582 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1583;
  assign dataGroup_hi_lo_1583 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1584;
  assign dataGroup_hi_lo_1584 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1585;
  assign dataGroup_hi_lo_1585 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1586;
  assign dataGroup_hi_lo_1586 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1587;
  assign dataGroup_hi_lo_1587 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1588;
  assign dataGroup_hi_lo_1588 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1589;
  assign dataGroup_hi_lo_1589 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1590;
  assign dataGroup_hi_lo_1590 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1591;
  assign dataGroup_hi_lo_1591 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1592;
  assign dataGroup_hi_lo_1592 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1593;
  assign dataGroup_hi_lo_1593 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1594;
  assign dataGroup_hi_lo_1594 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1595;
  assign dataGroup_hi_lo_1595 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1596;
  assign dataGroup_hi_lo_1596 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1597;
  assign dataGroup_hi_lo_1597 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1598;
  assign dataGroup_hi_lo_1598 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1599;
  assign dataGroup_hi_lo_1599 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1600;
  assign dataGroup_hi_lo_1600 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1601;
  assign dataGroup_hi_lo_1601 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1602;
  assign dataGroup_hi_lo_1602 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1603;
  assign dataGroup_hi_lo_1603 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1604;
  assign dataGroup_hi_lo_1604 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1605;
  assign dataGroup_hi_lo_1605 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1606;
  assign dataGroup_hi_lo_1606 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1607;
  assign dataGroup_hi_lo_1607 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1608;
  assign dataGroup_hi_lo_1608 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1609;
  assign dataGroup_hi_lo_1609 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1610;
  assign dataGroup_hi_lo_1610 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1611;
  assign dataGroup_hi_lo_1611 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1612;
  assign dataGroup_hi_lo_1612 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1613;
  assign dataGroup_hi_lo_1613 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1614;
  assign dataGroup_hi_lo_1614 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1615;
  assign dataGroup_hi_lo_1615 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1616;
  assign dataGroup_hi_lo_1616 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1617;
  assign dataGroup_hi_lo_1617 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1618;
  assign dataGroup_hi_lo_1618 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1619;
  assign dataGroup_hi_lo_1619 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1620;
  assign dataGroup_hi_lo_1620 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1621;
  assign dataGroup_hi_lo_1621 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1622;
  assign dataGroup_hi_lo_1622 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1623;
  assign dataGroup_hi_lo_1623 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1624;
  assign dataGroup_hi_lo_1624 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1625;
  assign dataGroup_hi_lo_1625 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1626;
  assign dataGroup_hi_lo_1626 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1627;
  assign dataGroup_hi_lo_1627 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1628;
  assign dataGroup_hi_lo_1628 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1629;
  assign dataGroup_hi_lo_1629 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1630;
  assign dataGroup_hi_lo_1630 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1631;
  assign dataGroup_hi_lo_1631 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1632;
  assign dataGroup_hi_lo_1632 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1633;
  assign dataGroup_hi_lo_1633 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1634;
  assign dataGroup_hi_lo_1634 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1635;
  assign dataGroup_hi_lo_1635 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1636;
  assign dataGroup_hi_lo_1636 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1637;
  assign dataGroup_hi_lo_1637 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1638;
  assign dataGroup_hi_lo_1638 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1639;
  assign dataGroup_hi_lo_1639 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1640;
  assign dataGroup_hi_lo_1640 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1641;
  assign dataGroup_hi_lo_1641 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1642;
  assign dataGroup_hi_lo_1642 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1643;
  assign dataGroup_hi_lo_1643 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1644;
  assign dataGroup_hi_lo_1644 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1645;
  assign dataGroup_hi_lo_1645 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1646;
  assign dataGroup_hi_lo_1646 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1647;
  assign dataGroup_hi_lo_1647 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1648;
  assign dataGroup_hi_lo_1648 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1649;
  assign dataGroup_hi_lo_1649 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1650;
  assign dataGroup_hi_lo_1650 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1651;
  assign dataGroup_hi_lo_1651 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1652;
  assign dataGroup_hi_lo_1652 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1653;
  assign dataGroup_hi_lo_1653 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1654;
  assign dataGroup_hi_lo_1654 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1655;
  assign dataGroup_hi_lo_1655 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1656;
  assign dataGroup_hi_lo_1656 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1657;
  assign dataGroup_hi_lo_1657 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1658;
  assign dataGroup_hi_lo_1658 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1659;
  assign dataGroup_hi_lo_1659 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1660;
  assign dataGroup_hi_lo_1660 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1661;
  assign dataGroup_hi_lo_1661 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1662;
  assign dataGroup_hi_lo_1662 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1663;
  assign dataGroup_hi_lo_1663 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1664;
  assign dataGroup_hi_lo_1664 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1665;
  assign dataGroup_hi_lo_1665 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1666;
  assign dataGroup_hi_lo_1666 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1667;
  assign dataGroup_hi_lo_1667 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1668;
  assign dataGroup_hi_lo_1668 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1669;
  assign dataGroup_hi_lo_1669 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1670;
  assign dataGroup_hi_lo_1670 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1671;
  assign dataGroup_hi_lo_1671 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1672;
  assign dataGroup_hi_lo_1672 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1673;
  assign dataGroup_hi_lo_1673 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1674;
  assign dataGroup_hi_lo_1674 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1675;
  assign dataGroup_hi_lo_1675 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1676;
  assign dataGroup_hi_lo_1676 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1677;
  assign dataGroup_hi_lo_1677 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1678;
  assign dataGroup_hi_lo_1678 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1679;
  assign dataGroup_hi_lo_1679 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1680;
  assign dataGroup_hi_lo_1680 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1681;
  assign dataGroup_hi_lo_1681 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1682;
  assign dataGroup_hi_lo_1682 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1683;
  assign dataGroup_hi_lo_1683 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1684;
  assign dataGroup_hi_lo_1684 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1685;
  assign dataGroup_hi_lo_1685 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1686;
  assign dataGroup_hi_lo_1686 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1687;
  assign dataGroup_hi_lo_1687 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1688;
  assign dataGroup_hi_lo_1688 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1689;
  assign dataGroup_hi_lo_1689 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1690;
  assign dataGroup_hi_lo_1690 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1691;
  assign dataGroup_hi_lo_1691 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1692;
  assign dataGroup_hi_lo_1692 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1693;
  assign dataGroup_hi_lo_1693 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1694;
  assign dataGroup_hi_lo_1694 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1695;
  assign dataGroup_hi_lo_1695 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1696;
  assign dataGroup_hi_lo_1696 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1697;
  assign dataGroup_hi_lo_1697 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1698;
  assign dataGroup_hi_lo_1698 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1699;
  assign dataGroup_hi_lo_1699 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1700;
  assign dataGroup_hi_lo_1700 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1701;
  assign dataGroup_hi_lo_1701 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1702;
  assign dataGroup_hi_lo_1702 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1703;
  assign dataGroup_hi_lo_1703 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1704;
  assign dataGroup_hi_lo_1704 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1705;
  assign dataGroup_hi_lo_1705 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1706;
  assign dataGroup_hi_lo_1706 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1707;
  assign dataGroup_hi_lo_1707 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1708;
  assign dataGroup_hi_lo_1708 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1709;
  assign dataGroup_hi_lo_1709 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1710;
  assign dataGroup_hi_lo_1710 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1711;
  assign dataGroup_hi_lo_1711 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1712;
  assign dataGroup_hi_lo_1712 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1713;
  assign dataGroup_hi_lo_1713 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1714;
  assign dataGroup_hi_lo_1714 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1715;
  assign dataGroup_hi_lo_1715 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1716;
  assign dataGroup_hi_lo_1716 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1717;
  assign dataGroup_hi_lo_1717 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1718;
  assign dataGroup_hi_lo_1718 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1719;
  assign dataGroup_hi_lo_1719 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1720;
  assign dataGroup_hi_lo_1720 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1721;
  assign dataGroup_hi_lo_1721 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1722;
  assign dataGroup_hi_lo_1722 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1723;
  assign dataGroup_hi_lo_1723 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1724;
  assign dataGroup_hi_lo_1724 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1725;
  assign dataGroup_hi_lo_1725 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1726;
  assign dataGroup_hi_lo_1726 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1727;
  assign dataGroup_hi_lo_1727 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1728;
  assign dataGroup_hi_lo_1728 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1729;
  assign dataGroup_hi_lo_1729 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1730;
  assign dataGroup_hi_lo_1730 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1731;
  assign dataGroup_hi_lo_1731 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1732;
  assign dataGroup_hi_lo_1732 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1733;
  assign dataGroup_hi_lo_1733 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1734;
  assign dataGroup_hi_lo_1734 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1735;
  assign dataGroup_hi_lo_1735 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1736;
  assign dataGroup_hi_lo_1736 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1737;
  assign dataGroup_hi_lo_1737 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1738;
  assign dataGroup_hi_lo_1738 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1739;
  assign dataGroup_hi_lo_1739 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1740;
  assign dataGroup_hi_lo_1740 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1741;
  assign dataGroup_hi_lo_1741 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1742;
  assign dataGroup_hi_lo_1742 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1743;
  assign dataGroup_hi_lo_1743 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1744;
  assign dataGroup_hi_lo_1744 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1745;
  assign dataGroup_hi_lo_1745 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1746;
  assign dataGroup_hi_lo_1746 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1747;
  assign dataGroup_hi_lo_1747 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1748;
  assign dataGroup_hi_lo_1748 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1749;
  assign dataGroup_hi_lo_1749 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1750;
  assign dataGroup_hi_lo_1750 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1751;
  assign dataGroup_hi_lo_1751 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1752;
  assign dataGroup_hi_lo_1752 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1753;
  assign dataGroup_hi_lo_1753 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1754;
  assign dataGroup_hi_lo_1754 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1755;
  assign dataGroup_hi_lo_1755 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1756;
  assign dataGroup_hi_lo_1756 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1757;
  assign dataGroup_hi_lo_1757 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1758;
  assign dataGroup_hi_lo_1758 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1759;
  assign dataGroup_hi_lo_1759 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1760;
  assign dataGroup_hi_lo_1760 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1761;
  assign dataGroup_hi_lo_1761 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1762;
  assign dataGroup_hi_lo_1762 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1763;
  assign dataGroup_hi_lo_1763 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1764;
  assign dataGroup_hi_lo_1764 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1765;
  assign dataGroup_hi_lo_1765 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1766;
  assign dataGroup_hi_lo_1766 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1767;
  assign dataGroup_hi_lo_1767 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1768;
  assign dataGroup_hi_lo_1768 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1769;
  assign dataGroup_hi_lo_1769 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1770;
  assign dataGroup_hi_lo_1770 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1771;
  assign dataGroup_hi_lo_1771 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1772;
  assign dataGroup_hi_lo_1772 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1773;
  assign dataGroup_hi_lo_1773 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1774;
  assign dataGroup_hi_lo_1774 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1775;
  assign dataGroup_hi_lo_1775 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1776;
  assign dataGroup_hi_lo_1776 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1777;
  assign dataGroup_hi_lo_1777 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1778;
  assign dataGroup_hi_lo_1778 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1779;
  assign dataGroup_hi_lo_1779 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1780;
  assign dataGroup_hi_lo_1780 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1781;
  assign dataGroup_hi_lo_1781 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1782;
  assign dataGroup_hi_lo_1782 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1783;
  assign dataGroup_hi_lo_1783 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1784;
  assign dataGroup_hi_lo_1784 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1785;
  assign dataGroup_hi_lo_1785 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1786;
  assign dataGroup_hi_lo_1786 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1787;
  assign dataGroup_hi_lo_1787 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1788;
  assign dataGroup_hi_lo_1788 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1789;
  assign dataGroup_hi_lo_1789 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1790;
  assign dataGroup_hi_lo_1790 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1791;
  assign dataGroup_hi_lo_1791 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1792;
  assign dataGroup_hi_lo_1792 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1793;
  assign dataGroup_hi_lo_1793 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1794;
  assign dataGroup_hi_lo_1794 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1795;
  assign dataGroup_hi_lo_1795 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1796;
  assign dataGroup_hi_lo_1796 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1797;
  assign dataGroup_hi_lo_1797 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1798;
  assign dataGroup_hi_lo_1798 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1799;
  assign dataGroup_hi_lo_1799 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1800;
  assign dataGroup_hi_lo_1800 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1801;
  assign dataGroup_hi_lo_1801 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1802;
  assign dataGroup_hi_lo_1802 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1803;
  assign dataGroup_hi_lo_1803 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1804;
  assign dataGroup_hi_lo_1804 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1805;
  assign dataGroup_hi_lo_1805 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1806;
  assign dataGroup_hi_lo_1806 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1807;
  assign dataGroup_hi_lo_1807 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1808;
  assign dataGroup_hi_lo_1808 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1809;
  assign dataGroup_hi_lo_1809 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1810;
  assign dataGroup_hi_lo_1810 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1811;
  assign dataGroup_hi_lo_1811 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1812;
  assign dataGroup_hi_lo_1812 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1813;
  assign dataGroup_hi_lo_1813 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1814;
  assign dataGroup_hi_lo_1814 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1815;
  assign dataGroup_hi_lo_1815 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1816;
  assign dataGroup_hi_lo_1816 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1817;
  assign dataGroup_hi_lo_1817 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1818;
  assign dataGroup_hi_lo_1818 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1819;
  assign dataGroup_hi_lo_1819 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1820;
  assign dataGroup_hi_lo_1820 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1821;
  assign dataGroup_hi_lo_1821 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1822;
  assign dataGroup_hi_lo_1822 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1823;
  assign dataGroup_hi_lo_1823 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1824;
  assign dataGroup_hi_lo_1824 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1825;
  assign dataGroup_hi_lo_1825 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1826;
  assign dataGroup_hi_lo_1826 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1827;
  assign dataGroup_hi_lo_1827 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1828;
  assign dataGroup_hi_lo_1828 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1829;
  assign dataGroup_hi_lo_1829 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1830;
  assign dataGroup_hi_lo_1830 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1831;
  assign dataGroup_hi_lo_1831 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1832;
  assign dataGroup_hi_lo_1832 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1833;
  assign dataGroup_hi_lo_1833 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1834;
  assign dataGroup_hi_lo_1834 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1835;
  assign dataGroup_hi_lo_1835 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1836;
  assign dataGroup_hi_lo_1836 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1837;
  assign dataGroup_hi_lo_1837 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1838;
  assign dataGroup_hi_lo_1838 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1839;
  assign dataGroup_hi_lo_1839 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1840;
  assign dataGroup_hi_lo_1840 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1841;
  assign dataGroup_hi_lo_1841 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1842;
  assign dataGroup_hi_lo_1842 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1843;
  assign dataGroup_hi_lo_1843 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1844;
  assign dataGroup_hi_lo_1844 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1845;
  assign dataGroup_hi_lo_1845 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1846;
  assign dataGroup_hi_lo_1846 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1847;
  assign dataGroup_hi_lo_1847 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1848;
  assign dataGroup_hi_lo_1848 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1849;
  assign dataGroup_hi_lo_1849 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1850;
  assign dataGroup_hi_lo_1850 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1851;
  assign dataGroup_hi_lo_1851 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1852;
  assign dataGroup_hi_lo_1852 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1853;
  assign dataGroup_hi_lo_1853 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1854;
  assign dataGroup_hi_lo_1854 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1855;
  assign dataGroup_hi_lo_1855 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1856;
  assign dataGroup_hi_lo_1856 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1857;
  assign dataGroup_hi_lo_1857 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1858;
  assign dataGroup_hi_lo_1858 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1859;
  assign dataGroup_hi_lo_1859 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1860;
  assign dataGroup_hi_lo_1860 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1861;
  assign dataGroup_hi_lo_1861 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1862;
  assign dataGroup_hi_lo_1862 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1863;
  assign dataGroup_hi_lo_1863 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1864;
  assign dataGroup_hi_lo_1864 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1865;
  assign dataGroup_hi_lo_1865 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1866;
  assign dataGroup_hi_lo_1866 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1867;
  assign dataGroup_hi_lo_1867 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1868;
  assign dataGroup_hi_lo_1868 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1869;
  assign dataGroup_hi_lo_1869 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1870;
  assign dataGroup_hi_lo_1870 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1871;
  assign dataGroup_hi_lo_1871 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1872;
  assign dataGroup_hi_lo_1872 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1873;
  assign dataGroup_hi_lo_1873 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1874;
  assign dataGroup_hi_lo_1874 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1875;
  assign dataGroup_hi_lo_1875 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1876;
  assign dataGroup_hi_lo_1876 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1877;
  assign dataGroup_hi_lo_1877 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1878;
  assign dataGroup_hi_lo_1878 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1879;
  assign dataGroup_hi_lo_1879 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1880;
  assign dataGroup_hi_lo_1880 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1881;
  assign dataGroup_hi_lo_1881 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1882;
  assign dataGroup_hi_lo_1882 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1883;
  assign dataGroup_hi_lo_1883 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1884;
  assign dataGroup_hi_lo_1884 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1885;
  assign dataGroup_hi_lo_1885 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1886;
  assign dataGroup_hi_lo_1886 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1887;
  assign dataGroup_hi_lo_1887 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1888;
  assign dataGroup_hi_lo_1888 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1889;
  assign dataGroup_hi_lo_1889 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1890;
  assign dataGroup_hi_lo_1890 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1891;
  assign dataGroup_hi_lo_1891 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1892;
  assign dataGroup_hi_lo_1892 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1893;
  assign dataGroup_hi_lo_1893 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1894;
  assign dataGroup_hi_lo_1894 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1895;
  assign dataGroup_hi_lo_1895 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1896;
  assign dataGroup_hi_lo_1896 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1897;
  assign dataGroup_hi_lo_1897 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1898;
  assign dataGroup_hi_lo_1898 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1899;
  assign dataGroup_hi_lo_1899 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1900;
  assign dataGroup_hi_lo_1900 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1901;
  assign dataGroup_hi_lo_1901 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1902;
  assign dataGroup_hi_lo_1902 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1903;
  assign dataGroup_hi_lo_1903 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1904;
  assign dataGroup_hi_lo_1904 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1905;
  assign dataGroup_hi_lo_1905 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1906;
  assign dataGroup_hi_lo_1906 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1907;
  assign dataGroup_hi_lo_1907 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1908;
  assign dataGroup_hi_lo_1908 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1909;
  assign dataGroup_hi_lo_1909 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1910;
  assign dataGroup_hi_lo_1910 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1911;
  assign dataGroup_hi_lo_1911 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1912;
  assign dataGroup_hi_lo_1912 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1913;
  assign dataGroup_hi_lo_1913 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1914;
  assign dataGroup_hi_lo_1914 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1915;
  assign dataGroup_hi_lo_1915 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1916;
  assign dataGroup_hi_lo_1916 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1917;
  assign dataGroup_hi_lo_1917 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1918;
  assign dataGroup_hi_lo_1918 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1919;
  assign dataGroup_hi_lo_1919 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1920;
  assign dataGroup_hi_lo_1920 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1921;
  assign dataGroup_hi_lo_1921 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1922;
  assign dataGroup_hi_lo_1922 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1923;
  assign dataGroup_hi_lo_1923 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1924;
  assign dataGroup_hi_lo_1924 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1925;
  assign dataGroup_hi_lo_1925 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1926;
  assign dataGroup_hi_lo_1926 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1927;
  assign dataGroup_hi_lo_1927 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1928;
  assign dataGroup_hi_lo_1928 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1929;
  assign dataGroup_hi_lo_1929 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1930;
  assign dataGroup_hi_lo_1930 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1931;
  assign dataGroup_hi_lo_1931 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1932;
  assign dataGroup_hi_lo_1932 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1933;
  assign dataGroup_hi_lo_1933 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1934;
  assign dataGroup_hi_lo_1934 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1935;
  assign dataGroup_hi_lo_1935 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1936;
  assign dataGroup_hi_lo_1936 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1937;
  assign dataGroup_hi_lo_1937 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1938;
  assign dataGroup_hi_lo_1938 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1939;
  assign dataGroup_hi_lo_1939 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1940;
  assign dataGroup_hi_lo_1940 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1941;
  assign dataGroup_hi_lo_1941 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1942;
  assign dataGroup_hi_lo_1942 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1943;
  assign dataGroup_hi_lo_1943 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1944;
  assign dataGroup_hi_lo_1944 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1945;
  assign dataGroup_hi_lo_1945 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1946;
  assign dataGroup_hi_lo_1946 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1947;
  assign dataGroup_hi_lo_1947 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1948;
  assign dataGroup_hi_lo_1948 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1949;
  assign dataGroup_hi_lo_1949 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1950;
  assign dataGroup_hi_lo_1950 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1951;
  assign dataGroup_hi_lo_1951 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1952;
  assign dataGroup_hi_lo_1952 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1953;
  assign dataGroup_hi_lo_1953 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1954;
  assign dataGroup_hi_lo_1954 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1955;
  assign dataGroup_hi_lo_1955 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1956;
  assign dataGroup_hi_lo_1956 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1957;
  assign dataGroup_hi_lo_1957 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1958;
  assign dataGroup_hi_lo_1958 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1959;
  assign dataGroup_hi_lo_1959 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1960;
  assign dataGroup_hi_lo_1960 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1961;
  assign dataGroup_hi_lo_1961 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1962;
  assign dataGroup_hi_lo_1962 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1963;
  assign dataGroup_hi_lo_1963 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1964;
  assign dataGroup_hi_lo_1964 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1965;
  assign dataGroup_hi_lo_1965 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1966;
  assign dataGroup_hi_lo_1966 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1967;
  assign dataGroup_hi_lo_1967 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1968;
  assign dataGroup_hi_lo_1968 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1969;
  assign dataGroup_hi_lo_1969 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1970;
  assign dataGroup_hi_lo_1970 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1971;
  assign dataGroup_hi_lo_1971 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1972;
  assign dataGroup_hi_lo_1972 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1973;
  assign dataGroup_hi_lo_1973 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1974;
  assign dataGroup_hi_lo_1974 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1975;
  assign dataGroup_hi_lo_1975 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1976;
  assign dataGroup_hi_lo_1976 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1977;
  assign dataGroup_hi_lo_1977 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1978;
  assign dataGroup_hi_lo_1978 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1979;
  assign dataGroup_hi_lo_1979 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1980;
  assign dataGroup_hi_lo_1980 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1981;
  assign dataGroup_hi_lo_1981 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1982;
  assign dataGroup_hi_lo_1982 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1983;
  assign dataGroup_hi_lo_1983 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1984;
  assign dataGroup_hi_lo_1984 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1985;
  assign dataGroup_hi_lo_1985 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1986;
  assign dataGroup_hi_lo_1986 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1987;
  assign dataGroup_hi_lo_1987 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1988;
  assign dataGroup_hi_lo_1988 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1989;
  assign dataGroup_hi_lo_1989 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1990;
  assign dataGroup_hi_lo_1990 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1991;
  assign dataGroup_hi_lo_1991 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1992;
  assign dataGroup_hi_lo_1992 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1993;
  assign dataGroup_hi_lo_1993 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1994;
  assign dataGroup_hi_lo_1994 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1995;
  assign dataGroup_hi_lo_1995 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1996;
  assign dataGroup_hi_lo_1996 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1997;
  assign dataGroup_hi_lo_1997 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1998;
  assign dataGroup_hi_lo_1998 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_1999;
  assign dataGroup_hi_lo_1999 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2000;
  assign dataGroup_hi_lo_2000 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2001;
  assign dataGroup_hi_lo_2001 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2002;
  assign dataGroup_hi_lo_2002 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2003;
  assign dataGroup_hi_lo_2003 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2004;
  assign dataGroup_hi_lo_2004 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2005;
  assign dataGroup_hi_lo_2005 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2006;
  assign dataGroup_hi_lo_2006 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2007;
  assign dataGroup_hi_lo_2007 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2008;
  assign dataGroup_hi_lo_2008 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2009;
  assign dataGroup_hi_lo_2009 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2010;
  assign dataGroup_hi_lo_2010 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2011;
  assign dataGroup_hi_lo_2011 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2012;
  assign dataGroup_hi_lo_2012 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2013;
  assign dataGroup_hi_lo_2013 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2014;
  assign dataGroup_hi_lo_2014 = _GEN_6;
  wire [511:0]  dataGroup_hi_lo_2015;
  assign dataGroup_hi_lo_2015 = _GEN_6;
  wire [511:0]  _GEN_7 = {dataSelect_7, dataSelect_6};
  wire [511:0]  dataGroup_hi_hi;
  assign dataGroup_hi_hi = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1;
  assign dataGroup_hi_hi_1 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2;
  assign dataGroup_hi_hi_2 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_3;
  assign dataGroup_hi_hi_3 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_4;
  assign dataGroup_hi_hi_4 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_5;
  assign dataGroup_hi_hi_5 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_6;
  assign dataGroup_hi_hi_6 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_7;
  assign dataGroup_hi_hi_7 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_8;
  assign dataGroup_hi_hi_8 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_9;
  assign dataGroup_hi_hi_9 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_10;
  assign dataGroup_hi_hi_10 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_11;
  assign dataGroup_hi_hi_11 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_12;
  assign dataGroup_hi_hi_12 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_13;
  assign dataGroup_hi_hi_13 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_14;
  assign dataGroup_hi_hi_14 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_15;
  assign dataGroup_hi_hi_15 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_16;
  assign dataGroup_hi_hi_16 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_17;
  assign dataGroup_hi_hi_17 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_18;
  assign dataGroup_hi_hi_18 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_19;
  assign dataGroup_hi_hi_19 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_20;
  assign dataGroup_hi_hi_20 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_21;
  assign dataGroup_hi_hi_21 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_22;
  assign dataGroup_hi_hi_22 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_23;
  assign dataGroup_hi_hi_23 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_24;
  assign dataGroup_hi_hi_24 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_25;
  assign dataGroup_hi_hi_25 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_26;
  assign dataGroup_hi_hi_26 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_27;
  assign dataGroup_hi_hi_27 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_28;
  assign dataGroup_hi_hi_28 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_29;
  assign dataGroup_hi_hi_29 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_30;
  assign dataGroup_hi_hi_30 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_31;
  assign dataGroup_hi_hi_31 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_32;
  assign dataGroup_hi_hi_32 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_33;
  assign dataGroup_hi_hi_33 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_34;
  assign dataGroup_hi_hi_34 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_35;
  assign dataGroup_hi_hi_35 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_36;
  assign dataGroup_hi_hi_36 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_37;
  assign dataGroup_hi_hi_37 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_38;
  assign dataGroup_hi_hi_38 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_39;
  assign dataGroup_hi_hi_39 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_40;
  assign dataGroup_hi_hi_40 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_41;
  assign dataGroup_hi_hi_41 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_42;
  assign dataGroup_hi_hi_42 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_43;
  assign dataGroup_hi_hi_43 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_44;
  assign dataGroup_hi_hi_44 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_45;
  assign dataGroup_hi_hi_45 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_46;
  assign dataGroup_hi_hi_46 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_47;
  assign dataGroup_hi_hi_47 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_48;
  assign dataGroup_hi_hi_48 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_49;
  assign dataGroup_hi_hi_49 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_50;
  assign dataGroup_hi_hi_50 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_51;
  assign dataGroup_hi_hi_51 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_52;
  assign dataGroup_hi_hi_52 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_53;
  assign dataGroup_hi_hi_53 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_54;
  assign dataGroup_hi_hi_54 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_55;
  assign dataGroup_hi_hi_55 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_56;
  assign dataGroup_hi_hi_56 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_57;
  assign dataGroup_hi_hi_57 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_58;
  assign dataGroup_hi_hi_58 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_59;
  assign dataGroup_hi_hi_59 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_60;
  assign dataGroup_hi_hi_60 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_61;
  assign dataGroup_hi_hi_61 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_62;
  assign dataGroup_hi_hi_62 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_63;
  assign dataGroup_hi_hi_63 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_64;
  assign dataGroup_hi_hi_64 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_65;
  assign dataGroup_hi_hi_65 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_66;
  assign dataGroup_hi_hi_66 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_67;
  assign dataGroup_hi_hi_67 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_68;
  assign dataGroup_hi_hi_68 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_69;
  assign dataGroup_hi_hi_69 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_70;
  assign dataGroup_hi_hi_70 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_71;
  assign dataGroup_hi_hi_71 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_72;
  assign dataGroup_hi_hi_72 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_73;
  assign dataGroup_hi_hi_73 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_74;
  assign dataGroup_hi_hi_74 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_75;
  assign dataGroup_hi_hi_75 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_76;
  assign dataGroup_hi_hi_76 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_77;
  assign dataGroup_hi_hi_77 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_78;
  assign dataGroup_hi_hi_78 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_79;
  assign dataGroup_hi_hi_79 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_80;
  assign dataGroup_hi_hi_80 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_81;
  assign dataGroup_hi_hi_81 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_82;
  assign dataGroup_hi_hi_82 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_83;
  assign dataGroup_hi_hi_83 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_84;
  assign dataGroup_hi_hi_84 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_85;
  assign dataGroup_hi_hi_85 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_86;
  assign dataGroup_hi_hi_86 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_87;
  assign dataGroup_hi_hi_87 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_88;
  assign dataGroup_hi_hi_88 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_89;
  assign dataGroup_hi_hi_89 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_90;
  assign dataGroup_hi_hi_90 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_91;
  assign dataGroup_hi_hi_91 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_92;
  assign dataGroup_hi_hi_92 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_93;
  assign dataGroup_hi_hi_93 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_94;
  assign dataGroup_hi_hi_94 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_95;
  assign dataGroup_hi_hi_95 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_96;
  assign dataGroup_hi_hi_96 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_97;
  assign dataGroup_hi_hi_97 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_98;
  assign dataGroup_hi_hi_98 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_99;
  assign dataGroup_hi_hi_99 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_100;
  assign dataGroup_hi_hi_100 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_101;
  assign dataGroup_hi_hi_101 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_102;
  assign dataGroup_hi_hi_102 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_103;
  assign dataGroup_hi_hi_103 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_104;
  assign dataGroup_hi_hi_104 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_105;
  assign dataGroup_hi_hi_105 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_106;
  assign dataGroup_hi_hi_106 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_107;
  assign dataGroup_hi_hi_107 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_108;
  assign dataGroup_hi_hi_108 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_109;
  assign dataGroup_hi_hi_109 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_110;
  assign dataGroup_hi_hi_110 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_111;
  assign dataGroup_hi_hi_111 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_112;
  assign dataGroup_hi_hi_112 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_113;
  assign dataGroup_hi_hi_113 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_114;
  assign dataGroup_hi_hi_114 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_115;
  assign dataGroup_hi_hi_115 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_116;
  assign dataGroup_hi_hi_116 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_117;
  assign dataGroup_hi_hi_117 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_118;
  assign dataGroup_hi_hi_118 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_119;
  assign dataGroup_hi_hi_119 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_120;
  assign dataGroup_hi_hi_120 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_121;
  assign dataGroup_hi_hi_121 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_122;
  assign dataGroup_hi_hi_122 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_123;
  assign dataGroup_hi_hi_123 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_124;
  assign dataGroup_hi_hi_124 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_125;
  assign dataGroup_hi_hi_125 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_126;
  assign dataGroup_hi_hi_126 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_127;
  assign dataGroup_hi_hi_127 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_128;
  assign dataGroup_hi_hi_128 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_129;
  assign dataGroup_hi_hi_129 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_130;
  assign dataGroup_hi_hi_130 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_131;
  assign dataGroup_hi_hi_131 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_132;
  assign dataGroup_hi_hi_132 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_133;
  assign dataGroup_hi_hi_133 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_134;
  assign dataGroup_hi_hi_134 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_135;
  assign dataGroup_hi_hi_135 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_136;
  assign dataGroup_hi_hi_136 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_137;
  assign dataGroup_hi_hi_137 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_138;
  assign dataGroup_hi_hi_138 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_139;
  assign dataGroup_hi_hi_139 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_140;
  assign dataGroup_hi_hi_140 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_141;
  assign dataGroup_hi_hi_141 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_142;
  assign dataGroup_hi_hi_142 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_143;
  assign dataGroup_hi_hi_143 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_144;
  assign dataGroup_hi_hi_144 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_145;
  assign dataGroup_hi_hi_145 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_146;
  assign dataGroup_hi_hi_146 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_147;
  assign dataGroup_hi_hi_147 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_148;
  assign dataGroup_hi_hi_148 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_149;
  assign dataGroup_hi_hi_149 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_150;
  assign dataGroup_hi_hi_150 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_151;
  assign dataGroup_hi_hi_151 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_152;
  assign dataGroup_hi_hi_152 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_153;
  assign dataGroup_hi_hi_153 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_154;
  assign dataGroup_hi_hi_154 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_155;
  assign dataGroup_hi_hi_155 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_156;
  assign dataGroup_hi_hi_156 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_157;
  assign dataGroup_hi_hi_157 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_158;
  assign dataGroup_hi_hi_158 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_159;
  assign dataGroup_hi_hi_159 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_160;
  assign dataGroup_hi_hi_160 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_161;
  assign dataGroup_hi_hi_161 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_162;
  assign dataGroup_hi_hi_162 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_163;
  assign dataGroup_hi_hi_163 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_164;
  assign dataGroup_hi_hi_164 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_165;
  assign dataGroup_hi_hi_165 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_166;
  assign dataGroup_hi_hi_166 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_167;
  assign dataGroup_hi_hi_167 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_168;
  assign dataGroup_hi_hi_168 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_169;
  assign dataGroup_hi_hi_169 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_170;
  assign dataGroup_hi_hi_170 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_171;
  assign dataGroup_hi_hi_171 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_172;
  assign dataGroup_hi_hi_172 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_173;
  assign dataGroup_hi_hi_173 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_174;
  assign dataGroup_hi_hi_174 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_175;
  assign dataGroup_hi_hi_175 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_176;
  assign dataGroup_hi_hi_176 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_177;
  assign dataGroup_hi_hi_177 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_178;
  assign dataGroup_hi_hi_178 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_179;
  assign dataGroup_hi_hi_179 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_180;
  assign dataGroup_hi_hi_180 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_181;
  assign dataGroup_hi_hi_181 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_182;
  assign dataGroup_hi_hi_182 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_183;
  assign dataGroup_hi_hi_183 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_184;
  assign dataGroup_hi_hi_184 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_185;
  assign dataGroup_hi_hi_185 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_186;
  assign dataGroup_hi_hi_186 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_187;
  assign dataGroup_hi_hi_187 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_188;
  assign dataGroup_hi_hi_188 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_189;
  assign dataGroup_hi_hi_189 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_190;
  assign dataGroup_hi_hi_190 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_191;
  assign dataGroup_hi_hi_191 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_192;
  assign dataGroup_hi_hi_192 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_193;
  assign dataGroup_hi_hi_193 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_194;
  assign dataGroup_hi_hi_194 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_195;
  assign dataGroup_hi_hi_195 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_196;
  assign dataGroup_hi_hi_196 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_197;
  assign dataGroup_hi_hi_197 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_198;
  assign dataGroup_hi_hi_198 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_199;
  assign dataGroup_hi_hi_199 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_200;
  assign dataGroup_hi_hi_200 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_201;
  assign dataGroup_hi_hi_201 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_202;
  assign dataGroup_hi_hi_202 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_203;
  assign dataGroup_hi_hi_203 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_204;
  assign dataGroup_hi_hi_204 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_205;
  assign dataGroup_hi_hi_205 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_206;
  assign dataGroup_hi_hi_206 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_207;
  assign dataGroup_hi_hi_207 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_208;
  assign dataGroup_hi_hi_208 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_209;
  assign dataGroup_hi_hi_209 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_210;
  assign dataGroup_hi_hi_210 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_211;
  assign dataGroup_hi_hi_211 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_212;
  assign dataGroup_hi_hi_212 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_213;
  assign dataGroup_hi_hi_213 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_214;
  assign dataGroup_hi_hi_214 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_215;
  assign dataGroup_hi_hi_215 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_216;
  assign dataGroup_hi_hi_216 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_217;
  assign dataGroup_hi_hi_217 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_218;
  assign dataGroup_hi_hi_218 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_219;
  assign dataGroup_hi_hi_219 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_220;
  assign dataGroup_hi_hi_220 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_221;
  assign dataGroup_hi_hi_221 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_222;
  assign dataGroup_hi_hi_222 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_223;
  assign dataGroup_hi_hi_223 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_224;
  assign dataGroup_hi_hi_224 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_225;
  assign dataGroup_hi_hi_225 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_226;
  assign dataGroup_hi_hi_226 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_227;
  assign dataGroup_hi_hi_227 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_228;
  assign dataGroup_hi_hi_228 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_229;
  assign dataGroup_hi_hi_229 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_230;
  assign dataGroup_hi_hi_230 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_231;
  assign dataGroup_hi_hi_231 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_232;
  assign dataGroup_hi_hi_232 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_233;
  assign dataGroup_hi_hi_233 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_234;
  assign dataGroup_hi_hi_234 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_235;
  assign dataGroup_hi_hi_235 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_236;
  assign dataGroup_hi_hi_236 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_237;
  assign dataGroup_hi_hi_237 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_238;
  assign dataGroup_hi_hi_238 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_239;
  assign dataGroup_hi_hi_239 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_240;
  assign dataGroup_hi_hi_240 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_241;
  assign dataGroup_hi_hi_241 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_242;
  assign dataGroup_hi_hi_242 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_243;
  assign dataGroup_hi_hi_243 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_244;
  assign dataGroup_hi_hi_244 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_245;
  assign dataGroup_hi_hi_245 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_246;
  assign dataGroup_hi_hi_246 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_247;
  assign dataGroup_hi_hi_247 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_248;
  assign dataGroup_hi_hi_248 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_249;
  assign dataGroup_hi_hi_249 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_250;
  assign dataGroup_hi_hi_250 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_251;
  assign dataGroup_hi_hi_251 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_252;
  assign dataGroup_hi_hi_252 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_253;
  assign dataGroup_hi_hi_253 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_254;
  assign dataGroup_hi_hi_254 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_255;
  assign dataGroup_hi_hi_255 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_256;
  assign dataGroup_hi_hi_256 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_257;
  assign dataGroup_hi_hi_257 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_258;
  assign dataGroup_hi_hi_258 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_259;
  assign dataGroup_hi_hi_259 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_260;
  assign dataGroup_hi_hi_260 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_261;
  assign dataGroup_hi_hi_261 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_262;
  assign dataGroup_hi_hi_262 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_263;
  assign dataGroup_hi_hi_263 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_264;
  assign dataGroup_hi_hi_264 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_265;
  assign dataGroup_hi_hi_265 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_266;
  assign dataGroup_hi_hi_266 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_267;
  assign dataGroup_hi_hi_267 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_268;
  assign dataGroup_hi_hi_268 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_269;
  assign dataGroup_hi_hi_269 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_270;
  assign dataGroup_hi_hi_270 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_271;
  assign dataGroup_hi_hi_271 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_272;
  assign dataGroup_hi_hi_272 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_273;
  assign dataGroup_hi_hi_273 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_274;
  assign dataGroup_hi_hi_274 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_275;
  assign dataGroup_hi_hi_275 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_276;
  assign dataGroup_hi_hi_276 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_277;
  assign dataGroup_hi_hi_277 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_278;
  assign dataGroup_hi_hi_278 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_279;
  assign dataGroup_hi_hi_279 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_280;
  assign dataGroup_hi_hi_280 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_281;
  assign dataGroup_hi_hi_281 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_282;
  assign dataGroup_hi_hi_282 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_283;
  assign dataGroup_hi_hi_283 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_284;
  assign dataGroup_hi_hi_284 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_285;
  assign dataGroup_hi_hi_285 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_286;
  assign dataGroup_hi_hi_286 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_287;
  assign dataGroup_hi_hi_287 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_288;
  assign dataGroup_hi_hi_288 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_289;
  assign dataGroup_hi_hi_289 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_290;
  assign dataGroup_hi_hi_290 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_291;
  assign dataGroup_hi_hi_291 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_292;
  assign dataGroup_hi_hi_292 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_293;
  assign dataGroup_hi_hi_293 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_294;
  assign dataGroup_hi_hi_294 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_295;
  assign dataGroup_hi_hi_295 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_296;
  assign dataGroup_hi_hi_296 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_297;
  assign dataGroup_hi_hi_297 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_298;
  assign dataGroup_hi_hi_298 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_299;
  assign dataGroup_hi_hi_299 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_300;
  assign dataGroup_hi_hi_300 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_301;
  assign dataGroup_hi_hi_301 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_302;
  assign dataGroup_hi_hi_302 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_303;
  assign dataGroup_hi_hi_303 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_304;
  assign dataGroup_hi_hi_304 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_305;
  assign dataGroup_hi_hi_305 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_306;
  assign dataGroup_hi_hi_306 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_307;
  assign dataGroup_hi_hi_307 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_308;
  assign dataGroup_hi_hi_308 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_309;
  assign dataGroup_hi_hi_309 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_310;
  assign dataGroup_hi_hi_310 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_311;
  assign dataGroup_hi_hi_311 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_312;
  assign dataGroup_hi_hi_312 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_313;
  assign dataGroup_hi_hi_313 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_314;
  assign dataGroup_hi_hi_314 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_315;
  assign dataGroup_hi_hi_315 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_316;
  assign dataGroup_hi_hi_316 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_317;
  assign dataGroup_hi_hi_317 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_318;
  assign dataGroup_hi_hi_318 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_319;
  assign dataGroup_hi_hi_319 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_320;
  assign dataGroup_hi_hi_320 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_321;
  assign dataGroup_hi_hi_321 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_322;
  assign dataGroup_hi_hi_322 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_323;
  assign dataGroup_hi_hi_323 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_324;
  assign dataGroup_hi_hi_324 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_325;
  assign dataGroup_hi_hi_325 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_326;
  assign dataGroup_hi_hi_326 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_327;
  assign dataGroup_hi_hi_327 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_328;
  assign dataGroup_hi_hi_328 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_329;
  assign dataGroup_hi_hi_329 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_330;
  assign dataGroup_hi_hi_330 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_331;
  assign dataGroup_hi_hi_331 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_332;
  assign dataGroup_hi_hi_332 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_333;
  assign dataGroup_hi_hi_333 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_334;
  assign dataGroup_hi_hi_334 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_335;
  assign dataGroup_hi_hi_335 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_336;
  assign dataGroup_hi_hi_336 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_337;
  assign dataGroup_hi_hi_337 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_338;
  assign dataGroup_hi_hi_338 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_339;
  assign dataGroup_hi_hi_339 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_340;
  assign dataGroup_hi_hi_340 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_341;
  assign dataGroup_hi_hi_341 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_342;
  assign dataGroup_hi_hi_342 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_343;
  assign dataGroup_hi_hi_343 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_344;
  assign dataGroup_hi_hi_344 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_345;
  assign dataGroup_hi_hi_345 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_346;
  assign dataGroup_hi_hi_346 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_347;
  assign dataGroup_hi_hi_347 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_348;
  assign dataGroup_hi_hi_348 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_349;
  assign dataGroup_hi_hi_349 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_350;
  assign dataGroup_hi_hi_350 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_351;
  assign dataGroup_hi_hi_351 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_352;
  assign dataGroup_hi_hi_352 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_353;
  assign dataGroup_hi_hi_353 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_354;
  assign dataGroup_hi_hi_354 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_355;
  assign dataGroup_hi_hi_355 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_356;
  assign dataGroup_hi_hi_356 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_357;
  assign dataGroup_hi_hi_357 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_358;
  assign dataGroup_hi_hi_358 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_359;
  assign dataGroup_hi_hi_359 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_360;
  assign dataGroup_hi_hi_360 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_361;
  assign dataGroup_hi_hi_361 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_362;
  assign dataGroup_hi_hi_362 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_363;
  assign dataGroup_hi_hi_363 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_364;
  assign dataGroup_hi_hi_364 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_365;
  assign dataGroup_hi_hi_365 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_366;
  assign dataGroup_hi_hi_366 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_367;
  assign dataGroup_hi_hi_367 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_368;
  assign dataGroup_hi_hi_368 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_369;
  assign dataGroup_hi_hi_369 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_370;
  assign dataGroup_hi_hi_370 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_371;
  assign dataGroup_hi_hi_371 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_372;
  assign dataGroup_hi_hi_372 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_373;
  assign dataGroup_hi_hi_373 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_374;
  assign dataGroup_hi_hi_374 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_375;
  assign dataGroup_hi_hi_375 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_376;
  assign dataGroup_hi_hi_376 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_377;
  assign dataGroup_hi_hi_377 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_378;
  assign dataGroup_hi_hi_378 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_379;
  assign dataGroup_hi_hi_379 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_380;
  assign dataGroup_hi_hi_380 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_381;
  assign dataGroup_hi_hi_381 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_382;
  assign dataGroup_hi_hi_382 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_383;
  assign dataGroup_hi_hi_383 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_384;
  assign dataGroup_hi_hi_384 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_385;
  assign dataGroup_hi_hi_385 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_386;
  assign dataGroup_hi_hi_386 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_387;
  assign dataGroup_hi_hi_387 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_388;
  assign dataGroup_hi_hi_388 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_389;
  assign dataGroup_hi_hi_389 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_390;
  assign dataGroup_hi_hi_390 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_391;
  assign dataGroup_hi_hi_391 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_392;
  assign dataGroup_hi_hi_392 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_393;
  assign dataGroup_hi_hi_393 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_394;
  assign dataGroup_hi_hi_394 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_395;
  assign dataGroup_hi_hi_395 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_396;
  assign dataGroup_hi_hi_396 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_397;
  assign dataGroup_hi_hi_397 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_398;
  assign dataGroup_hi_hi_398 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_399;
  assign dataGroup_hi_hi_399 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_400;
  assign dataGroup_hi_hi_400 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_401;
  assign dataGroup_hi_hi_401 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_402;
  assign dataGroup_hi_hi_402 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_403;
  assign dataGroup_hi_hi_403 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_404;
  assign dataGroup_hi_hi_404 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_405;
  assign dataGroup_hi_hi_405 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_406;
  assign dataGroup_hi_hi_406 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_407;
  assign dataGroup_hi_hi_407 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_408;
  assign dataGroup_hi_hi_408 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_409;
  assign dataGroup_hi_hi_409 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_410;
  assign dataGroup_hi_hi_410 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_411;
  assign dataGroup_hi_hi_411 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_412;
  assign dataGroup_hi_hi_412 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_413;
  assign dataGroup_hi_hi_413 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_414;
  assign dataGroup_hi_hi_414 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_415;
  assign dataGroup_hi_hi_415 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_416;
  assign dataGroup_hi_hi_416 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_417;
  assign dataGroup_hi_hi_417 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_418;
  assign dataGroup_hi_hi_418 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_419;
  assign dataGroup_hi_hi_419 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_420;
  assign dataGroup_hi_hi_420 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_421;
  assign dataGroup_hi_hi_421 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_422;
  assign dataGroup_hi_hi_422 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_423;
  assign dataGroup_hi_hi_423 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_424;
  assign dataGroup_hi_hi_424 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_425;
  assign dataGroup_hi_hi_425 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_426;
  assign dataGroup_hi_hi_426 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_427;
  assign dataGroup_hi_hi_427 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_428;
  assign dataGroup_hi_hi_428 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_429;
  assign dataGroup_hi_hi_429 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_430;
  assign dataGroup_hi_hi_430 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_431;
  assign dataGroup_hi_hi_431 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_432;
  assign dataGroup_hi_hi_432 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_433;
  assign dataGroup_hi_hi_433 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_434;
  assign dataGroup_hi_hi_434 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_435;
  assign dataGroup_hi_hi_435 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_436;
  assign dataGroup_hi_hi_436 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_437;
  assign dataGroup_hi_hi_437 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_438;
  assign dataGroup_hi_hi_438 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_439;
  assign dataGroup_hi_hi_439 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_440;
  assign dataGroup_hi_hi_440 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_441;
  assign dataGroup_hi_hi_441 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_442;
  assign dataGroup_hi_hi_442 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_443;
  assign dataGroup_hi_hi_443 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_444;
  assign dataGroup_hi_hi_444 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_445;
  assign dataGroup_hi_hi_445 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_446;
  assign dataGroup_hi_hi_446 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_447;
  assign dataGroup_hi_hi_447 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_448;
  assign dataGroup_hi_hi_448 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_449;
  assign dataGroup_hi_hi_449 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_450;
  assign dataGroup_hi_hi_450 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_451;
  assign dataGroup_hi_hi_451 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_452;
  assign dataGroup_hi_hi_452 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_453;
  assign dataGroup_hi_hi_453 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_454;
  assign dataGroup_hi_hi_454 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_455;
  assign dataGroup_hi_hi_455 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_456;
  assign dataGroup_hi_hi_456 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_457;
  assign dataGroup_hi_hi_457 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_458;
  assign dataGroup_hi_hi_458 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_459;
  assign dataGroup_hi_hi_459 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_460;
  assign dataGroup_hi_hi_460 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_461;
  assign dataGroup_hi_hi_461 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_462;
  assign dataGroup_hi_hi_462 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_463;
  assign dataGroup_hi_hi_463 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_464;
  assign dataGroup_hi_hi_464 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_465;
  assign dataGroup_hi_hi_465 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_466;
  assign dataGroup_hi_hi_466 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_467;
  assign dataGroup_hi_hi_467 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_468;
  assign dataGroup_hi_hi_468 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_469;
  assign dataGroup_hi_hi_469 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_470;
  assign dataGroup_hi_hi_470 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_471;
  assign dataGroup_hi_hi_471 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_472;
  assign dataGroup_hi_hi_472 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_473;
  assign dataGroup_hi_hi_473 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_474;
  assign dataGroup_hi_hi_474 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_475;
  assign dataGroup_hi_hi_475 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_476;
  assign dataGroup_hi_hi_476 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_477;
  assign dataGroup_hi_hi_477 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_478;
  assign dataGroup_hi_hi_478 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_479;
  assign dataGroup_hi_hi_479 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_480;
  assign dataGroup_hi_hi_480 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_481;
  assign dataGroup_hi_hi_481 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_482;
  assign dataGroup_hi_hi_482 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_483;
  assign dataGroup_hi_hi_483 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_484;
  assign dataGroup_hi_hi_484 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_485;
  assign dataGroup_hi_hi_485 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_486;
  assign dataGroup_hi_hi_486 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_487;
  assign dataGroup_hi_hi_487 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_488;
  assign dataGroup_hi_hi_488 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_489;
  assign dataGroup_hi_hi_489 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_490;
  assign dataGroup_hi_hi_490 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_491;
  assign dataGroup_hi_hi_491 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_492;
  assign dataGroup_hi_hi_492 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_493;
  assign dataGroup_hi_hi_493 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_494;
  assign dataGroup_hi_hi_494 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_495;
  assign dataGroup_hi_hi_495 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_496;
  assign dataGroup_hi_hi_496 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_497;
  assign dataGroup_hi_hi_497 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_498;
  assign dataGroup_hi_hi_498 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_499;
  assign dataGroup_hi_hi_499 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_500;
  assign dataGroup_hi_hi_500 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_501;
  assign dataGroup_hi_hi_501 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_502;
  assign dataGroup_hi_hi_502 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_503;
  assign dataGroup_hi_hi_503 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_504;
  assign dataGroup_hi_hi_504 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_505;
  assign dataGroup_hi_hi_505 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_506;
  assign dataGroup_hi_hi_506 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_507;
  assign dataGroup_hi_hi_507 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_508;
  assign dataGroup_hi_hi_508 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_509;
  assign dataGroup_hi_hi_509 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_510;
  assign dataGroup_hi_hi_510 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_511;
  assign dataGroup_hi_hi_511 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_512;
  assign dataGroup_hi_hi_512 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_513;
  assign dataGroup_hi_hi_513 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_514;
  assign dataGroup_hi_hi_514 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_515;
  assign dataGroup_hi_hi_515 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_516;
  assign dataGroup_hi_hi_516 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_517;
  assign dataGroup_hi_hi_517 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_518;
  assign dataGroup_hi_hi_518 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_519;
  assign dataGroup_hi_hi_519 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_520;
  assign dataGroup_hi_hi_520 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_521;
  assign dataGroup_hi_hi_521 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_522;
  assign dataGroup_hi_hi_522 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_523;
  assign dataGroup_hi_hi_523 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_524;
  assign dataGroup_hi_hi_524 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_525;
  assign dataGroup_hi_hi_525 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_526;
  assign dataGroup_hi_hi_526 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_527;
  assign dataGroup_hi_hi_527 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_528;
  assign dataGroup_hi_hi_528 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_529;
  assign dataGroup_hi_hi_529 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_530;
  assign dataGroup_hi_hi_530 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_531;
  assign dataGroup_hi_hi_531 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_532;
  assign dataGroup_hi_hi_532 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_533;
  assign dataGroup_hi_hi_533 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_534;
  assign dataGroup_hi_hi_534 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_535;
  assign dataGroup_hi_hi_535 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_536;
  assign dataGroup_hi_hi_536 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_537;
  assign dataGroup_hi_hi_537 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_538;
  assign dataGroup_hi_hi_538 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_539;
  assign dataGroup_hi_hi_539 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_540;
  assign dataGroup_hi_hi_540 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_541;
  assign dataGroup_hi_hi_541 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_542;
  assign dataGroup_hi_hi_542 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_543;
  assign dataGroup_hi_hi_543 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_544;
  assign dataGroup_hi_hi_544 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_545;
  assign dataGroup_hi_hi_545 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_546;
  assign dataGroup_hi_hi_546 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_547;
  assign dataGroup_hi_hi_547 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_548;
  assign dataGroup_hi_hi_548 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_549;
  assign dataGroup_hi_hi_549 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_550;
  assign dataGroup_hi_hi_550 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_551;
  assign dataGroup_hi_hi_551 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_552;
  assign dataGroup_hi_hi_552 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_553;
  assign dataGroup_hi_hi_553 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_554;
  assign dataGroup_hi_hi_554 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_555;
  assign dataGroup_hi_hi_555 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_556;
  assign dataGroup_hi_hi_556 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_557;
  assign dataGroup_hi_hi_557 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_558;
  assign dataGroup_hi_hi_558 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_559;
  assign dataGroup_hi_hi_559 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_560;
  assign dataGroup_hi_hi_560 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_561;
  assign dataGroup_hi_hi_561 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_562;
  assign dataGroup_hi_hi_562 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_563;
  assign dataGroup_hi_hi_563 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_564;
  assign dataGroup_hi_hi_564 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_565;
  assign dataGroup_hi_hi_565 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_566;
  assign dataGroup_hi_hi_566 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_567;
  assign dataGroup_hi_hi_567 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_568;
  assign dataGroup_hi_hi_568 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_569;
  assign dataGroup_hi_hi_569 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_570;
  assign dataGroup_hi_hi_570 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_571;
  assign dataGroup_hi_hi_571 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_572;
  assign dataGroup_hi_hi_572 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_573;
  assign dataGroup_hi_hi_573 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_574;
  assign dataGroup_hi_hi_574 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_575;
  assign dataGroup_hi_hi_575 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_576;
  assign dataGroup_hi_hi_576 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_577;
  assign dataGroup_hi_hi_577 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_578;
  assign dataGroup_hi_hi_578 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_579;
  assign dataGroup_hi_hi_579 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_580;
  assign dataGroup_hi_hi_580 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_581;
  assign dataGroup_hi_hi_581 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_582;
  assign dataGroup_hi_hi_582 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_583;
  assign dataGroup_hi_hi_583 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_584;
  assign dataGroup_hi_hi_584 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_585;
  assign dataGroup_hi_hi_585 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_586;
  assign dataGroup_hi_hi_586 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_587;
  assign dataGroup_hi_hi_587 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_588;
  assign dataGroup_hi_hi_588 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_589;
  assign dataGroup_hi_hi_589 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_590;
  assign dataGroup_hi_hi_590 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_591;
  assign dataGroup_hi_hi_591 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_592;
  assign dataGroup_hi_hi_592 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_593;
  assign dataGroup_hi_hi_593 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_594;
  assign dataGroup_hi_hi_594 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_595;
  assign dataGroup_hi_hi_595 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_596;
  assign dataGroup_hi_hi_596 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_597;
  assign dataGroup_hi_hi_597 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_598;
  assign dataGroup_hi_hi_598 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_599;
  assign dataGroup_hi_hi_599 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_600;
  assign dataGroup_hi_hi_600 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_601;
  assign dataGroup_hi_hi_601 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_602;
  assign dataGroup_hi_hi_602 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_603;
  assign dataGroup_hi_hi_603 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_604;
  assign dataGroup_hi_hi_604 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_605;
  assign dataGroup_hi_hi_605 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_606;
  assign dataGroup_hi_hi_606 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_607;
  assign dataGroup_hi_hi_607 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_608;
  assign dataGroup_hi_hi_608 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_609;
  assign dataGroup_hi_hi_609 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_610;
  assign dataGroup_hi_hi_610 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_611;
  assign dataGroup_hi_hi_611 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_612;
  assign dataGroup_hi_hi_612 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_613;
  assign dataGroup_hi_hi_613 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_614;
  assign dataGroup_hi_hi_614 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_615;
  assign dataGroup_hi_hi_615 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_616;
  assign dataGroup_hi_hi_616 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_617;
  assign dataGroup_hi_hi_617 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_618;
  assign dataGroup_hi_hi_618 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_619;
  assign dataGroup_hi_hi_619 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_620;
  assign dataGroup_hi_hi_620 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_621;
  assign dataGroup_hi_hi_621 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_622;
  assign dataGroup_hi_hi_622 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_623;
  assign dataGroup_hi_hi_623 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_624;
  assign dataGroup_hi_hi_624 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_625;
  assign dataGroup_hi_hi_625 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_626;
  assign dataGroup_hi_hi_626 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_627;
  assign dataGroup_hi_hi_627 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_628;
  assign dataGroup_hi_hi_628 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_629;
  assign dataGroup_hi_hi_629 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_630;
  assign dataGroup_hi_hi_630 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_631;
  assign dataGroup_hi_hi_631 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_632;
  assign dataGroup_hi_hi_632 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_633;
  assign dataGroup_hi_hi_633 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_634;
  assign dataGroup_hi_hi_634 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_635;
  assign dataGroup_hi_hi_635 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_636;
  assign dataGroup_hi_hi_636 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_637;
  assign dataGroup_hi_hi_637 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_638;
  assign dataGroup_hi_hi_638 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_639;
  assign dataGroup_hi_hi_639 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_640;
  assign dataGroup_hi_hi_640 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_641;
  assign dataGroup_hi_hi_641 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_642;
  assign dataGroup_hi_hi_642 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_643;
  assign dataGroup_hi_hi_643 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_644;
  assign dataGroup_hi_hi_644 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_645;
  assign dataGroup_hi_hi_645 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_646;
  assign dataGroup_hi_hi_646 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_647;
  assign dataGroup_hi_hi_647 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_648;
  assign dataGroup_hi_hi_648 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_649;
  assign dataGroup_hi_hi_649 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_650;
  assign dataGroup_hi_hi_650 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_651;
  assign dataGroup_hi_hi_651 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_652;
  assign dataGroup_hi_hi_652 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_653;
  assign dataGroup_hi_hi_653 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_654;
  assign dataGroup_hi_hi_654 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_655;
  assign dataGroup_hi_hi_655 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_656;
  assign dataGroup_hi_hi_656 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_657;
  assign dataGroup_hi_hi_657 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_658;
  assign dataGroup_hi_hi_658 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_659;
  assign dataGroup_hi_hi_659 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_660;
  assign dataGroup_hi_hi_660 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_661;
  assign dataGroup_hi_hi_661 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_662;
  assign dataGroup_hi_hi_662 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_663;
  assign dataGroup_hi_hi_663 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_664;
  assign dataGroup_hi_hi_664 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_665;
  assign dataGroup_hi_hi_665 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_666;
  assign dataGroup_hi_hi_666 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_667;
  assign dataGroup_hi_hi_667 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_668;
  assign dataGroup_hi_hi_668 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_669;
  assign dataGroup_hi_hi_669 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_670;
  assign dataGroup_hi_hi_670 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_671;
  assign dataGroup_hi_hi_671 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_672;
  assign dataGroup_hi_hi_672 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_673;
  assign dataGroup_hi_hi_673 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_674;
  assign dataGroup_hi_hi_674 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_675;
  assign dataGroup_hi_hi_675 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_676;
  assign dataGroup_hi_hi_676 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_677;
  assign dataGroup_hi_hi_677 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_678;
  assign dataGroup_hi_hi_678 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_679;
  assign dataGroup_hi_hi_679 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_680;
  assign dataGroup_hi_hi_680 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_681;
  assign dataGroup_hi_hi_681 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_682;
  assign dataGroup_hi_hi_682 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_683;
  assign dataGroup_hi_hi_683 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_684;
  assign dataGroup_hi_hi_684 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_685;
  assign dataGroup_hi_hi_685 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_686;
  assign dataGroup_hi_hi_686 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_687;
  assign dataGroup_hi_hi_687 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_688;
  assign dataGroup_hi_hi_688 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_689;
  assign dataGroup_hi_hi_689 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_690;
  assign dataGroup_hi_hi_690 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_691;
  assign dataGroup_hi_hi_691 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_692;
  assign dataGroup_hi_hi_692 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_693;
  assign dataGroup_hi_hi_693 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_694;
  assign dataGroup_hi_hi_694 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_695;
  assign dataGroup_hi_hi_695 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_696;
  assign dataGroup_hi_hi_696 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_697;
  assign dataGroup_hi_hi_697 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_698;
  assign dataGroup_hi_hi_698 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_699;
  assign dataGroup_hi_hi_699 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_700;
  assign dataGroup_hi_hi_700 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_701;
  assign dataGroup_hi_hi_701 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_702;
  assign dataGroup_hi_hi_702 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_703;
  assign dataGroup_hi_hi_703 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_704;
  assign dataGroup_hi_hi_704 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_705;
  assign dataGroup_hi_hi_705 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_706;
  assign dataGroup_hi_hi_706 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_707;
  assign dataGroup_hi_hi_707 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_708;
  assign dataGroup_hi_hi_708 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_709;
  assign dataGroup_hi_hi_709 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_710;
  assign dataGroup_hi_hi_710 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_711;
  assign dataGroup_hi_hi_711 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_712;
  assign dataGroup_hi_hi_712 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_713;
  assign dataGroup_hi_hi_713 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_714;
  assign dataGroup_hi_hi_714 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_715;
  assign dataGroup_hi_hi_715 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_716;
  assign dataGroup_hi_hi_716 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_717;
  assign dataGroup_hi_hi_717 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_718;
  assign dataGroup_hi_hi_718 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_719;
  assign dataGroup_hi_hi_719 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_720;
  assign dataGroup_hi_hi_720 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_721;
  assign dataGroup_hi_hi_721 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_722;
  assign dataGroup_hi_hi_722 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_723;
  assign dataGroup_hi_hi_723 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_724;
  assign dataGroup_hi_hi_724 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_725;
  assign dataGroup_hi_hi_725 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_726;
  assign dataGroup_hi_hi_726 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_727;
  assign dataGroup_hi_hi_727 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_728;
  assign dataGroup_hi_hi_728 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_729;
  assign dataGroup_hi_hi_729 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_730;
  assign dataGroup_hi_hi_730 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_731;
  assign dataGroup_hi_hi_731 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_732;
  assign dataGroup_hi_hi_732 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_733;
  assign dataGroup_hi_hi_733 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_734;
  assign dataGroup_hi_hi_734 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_735;
  assign dataGroup_hi_hi_735 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_736;
  assign dataGroup_hi_hi_736 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_737;
  assign dataGroup_hi_hi_737 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_738;
  assign dataGroup_hi_hi_738 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_739;
  assign dataGroup_hi_hi_739 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_740;
  assign dataGroup_hi_hi_740 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_741;
  assign dataGroup_hi_hi_741 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_742;
  assign dataGroup_hi_hi_742 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_743;
  assign dataGroup_hi_hi_743 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_744;
  assign dataGroup_hi_hi_744 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_745;
  assign dataGroup_hi_hi_745 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_746;
  assign dataGroup_hi_hi_746 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_747;
  assign dataGroup_hi_hi_747 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_748;
  assign dataGroup_hi_hi_748 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_749;
  assign dataGroup_hi_hi_749 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_750;
  assign dataGroup_hi_hi_750 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_751;
  assign dataGroup_hi_hi_751 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_752;
  assign dataGroup_hi_hi_752 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_753;
  assign dataGroup_hi_hi_753 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_754;
  assign dataGroup_hi_hi_754 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_755;
  assign dataGroup_hi_hi_755 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_756;
  assign dataGroup_hi_hi_756 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_757;
  assign dataGroup_hi_hi_757 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_758;
  assign dataGroup_hi_hi_758 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_759;
  assign dataGroup_hi_hi_759 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_760;
  assign dataGroup_hi_hi_760 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_761;
  assign dataGroup_hi_hi_761 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_762;
  assign dataGroup_hi_hi_762 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_763;
  assign dataGroup_hi_hi_763 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_764;
  assign dataGroup_hi_hi_764 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_765;
  assign dataGroup_hi_hi_765 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_766;
  assign dataGroup_hi_hi_766 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_767;
  assign dataGroup_hi_hi_767 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_768;
  assign dataGroup_hi_hi_768 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_769;
  assign dataGroup_hi_hi_769 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_770;
  assign dataGroup_hi_hi_770 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_771;
  assign dataGroup_hi_hi_771 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_772;
  assign dataGroup_hi_hi_772 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_773;
  assign dataGroup_hi_hi_773 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_774;
  assign dataGroup_hi_hi_774 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_775;
  assign dataGroup_hi_hi_775 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_776;
  assign dataGroup_hi_hi_776 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_777;
  assign dataGroup_hi_hi_777 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_778;
  assign dataGroup_hi_hi_778 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_779;
  assign dataGroup_hi_hi_779 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_780;
  assign dataGroup_hi_hi_780 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_781;
  assign dataGroup_hi_hi_781 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_782;
  assign dataGroup_hi_hi_782 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_783;
  assign dataGroup_hi_hi_783 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_784;
  assign dataGroup_hi_hi_784 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_785;
  assign dataGroup_hi_hi_785 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_786;
  assign dataGroup_hi_hi_786 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_787;
  assign dataGroup_hi_hi_787 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_788;
  assign dataGroup_hi_hi_788 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_789;
  assign dataGroup_hi_hi_789 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_790;
  assign dataGroup_hi_hi_790 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_791;
  assign dataGroup_hi_hi_791 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_792;
  assign dataGroup_hi_hi_792 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_793;
  assign dataGroup_hi_hi_793 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_794;
  assign dataGroup_hi_hi_794 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_795;
  assign dataGroup_hi_hi_795 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_796;
  assign dataGroup_hi_hi_796 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_797;
  assign dataGroup_hi_hi_797 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_798;
  assign dataGroup_hi_hi_798 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_799;
  assign dataGroup_hi_hi_799 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_800;
  assign dataGroup_hi_hi_800 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_801;
  assign dataGroup_hi_hi_801 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_802;
  assign dataGroup_hi_hi_802 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_803;
  assign dataGroup_hi_hi_803 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_804;
  assign dataGroup_hi_hi_804 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_805;
  assign dataGroup_hi_hi_805 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_806;
  assign dataGroup_hi_hi_806 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_807;
  assign dataGroup_hi_hi_807 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_808;
  assign dataGroup_hi_hi_808 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_809;
  assign dataGroup_hi_hi_809 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_810;
  assign dataGroup_hi_hi_810 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_811;
  assign dataGroup_hi_hi_811 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_812;
  assign dataGroup_hi_hi_812 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_813;
  assign dataGroup_hi_hi_813 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_814;
  assign dataGroup_hi_hi_814 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_815;
  assign dataGroup_hi_hi_815 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_816;
  assign dataGroup_hi_hi_816 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_817;
  assign dataGroup_hi_hi_817 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_818;
  assign dataGroup_hi_hi_818 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_819;
  assign dataGroup_hi_hi_819 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_820;
  assign dataGroup_hi_hi_820 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_821;
  assign dataGroup_hi_hi_821 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_822;
  assign dataGroup_hi_hi_822 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_823;
  assign dataGroup_hi_hi_823 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_824;
  assign dataGroup_hi_hi_824 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_825;
  assign dataGroup_hi_hi_825 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_826;
  assign dataGroup_hi_hi_826 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_827;
  assign dataGroup_hi_hi_827 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_828;
  assign dataGroup_hi_hi_828 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_829;
  assign dataGroup_hi_hi_829 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_830;
  assign dataGroup_hi_hi_830 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_831;
  assign dataGroup_hi_hi_831 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_832;
  assign dataGroup_hi_hi_832 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_833;
  assign dataGroup_hi_hi_833 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_834;
  assign dataGroup_hi_hi_834 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_835;
  assign dataGroup_hi_hi_835 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_836;
  assign dataGroup_hi_hi_836 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_837;
  assign dataGroup_hi_hi_837 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_838;
  assign dataGroup_hi_hi_838 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_839;
  assign dataGroup_hi_hi_839 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_840;
  assign dataGroup_hi_hi_840 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_841;
  assign dataGroup_hi_hi_841 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_842;
  assign dataGroup_hi_hi_842 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_843;
  assign dataGroup_hi_hi_843 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_844;
  assign dataGroup_hi_hi_844 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_845;
  assign dataGroup_hi_hi_845 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_846;
  assign dataGroup_hi_hi_846 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_847;
  assign dataGroup_hi_hi_847 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_848;
  assign dataGroup_hi_hi_848 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_849;
  assign dataGroup_hi_hi_849 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_850;
  assign dataGroup_hi_hi_850 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_851;
  assign dataGroup_hi_hi_851 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_852;
  assign dataGroup_hi_hi_852 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_853;
  assign dataGroup_hi_hi_853 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_854;
  assign dataGroup_hi_hi_854 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_855;
  assign dataGroup_hi_hi_855 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_856;
  assign dataGroup_hi_hi_856 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_857;
  assign dataGroup_hi_hi_857 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_858;
  assign dataGroup_hi_hi_858 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_859;
  assign dataGroup_hi_hi_859 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_860;
  assign dataGroup_hi_hi_860 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_861;
  assign dataGroup_hi_hi_861 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_862;
  assign dataGroup_hi_hi_862 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_863;
  assign dataGroup_hi_hi_863 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_864;
  assign dataGroup_hi_hi_864 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_865;
  assign dataGroup_hi_hi_865 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_866;
  assign dataGroup_hi_hi_866 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_867;
  assign dataGroup_hi_hi_867 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_868;
  assign dataGroup_hi_hi_868 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_869;
  assign dataGroup_hi_hi_869 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_870;
  assign dataGroup_hi_hi_870 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_871;
  assign dataGroup_hi_hi_871 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_872;
  assign dataGroup_hi_hi_872 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_873;
  assign dataGroup_hi_hi_873 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_874;
  assign dataGroup_hi_hi_874 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_875;
  assign dataGroup_hi_hi_875 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_876;
  assign dataGroup_hi_hi_876 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_877;
  assign dataGroup_hi_hi_877 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_878;
  assign dataGroup_hi_hi_878 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_879;
  assign dataGroup_hi_hi_879 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_880;
  assign dataGroup_hi_hi_880 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_881;
  assign dataGroup_hi_hi_881 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_882;
  assign dataGroup_hi_hi_882 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_883;
  assign dataGroup_hi_hi_883 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_884;
  assign dataGroup_hi_hi_884 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_885;
  assign dataGroup_hi_hi_885 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_886;
  assign dataGroup_hi_hi_886 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_887;
  assign dataGroup_hi_hi_887 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_888;
  assign dataGroup_hi_hi_888 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_889;
  assign dataGroup_hi_hi_889 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_890;
  assign dataGroup_hi_hi_890 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_891;
  assign dataGroup_hi_hi_891 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_892;
  assign dataGroup_hi_hi_892 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_893;
  assign dataGroup_hi_hi_893 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_894;
  assign dataGroup_hi_hi_894 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_895;
  assign dataGroup_hi_hi_895 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_896;
  assign dataGroup_hi_hi_896 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_897;
  assign dataGroup_hi_hi_897 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_898;
  assign dataGroup_hi_hi_898 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_899;
  assign dataGroup_hi_hi_899 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_900;
  assign dataGroup_hi_hi_900 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_901;
  assign dataGroup_hi_hi_901 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_902;
  assign dataGroup_hi_hi_902 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_903;
  assign dataGroup_hi_hi_903 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_904;
  assign dataGroup_hi_hi_904 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_905;
  assign dataGroup_hi_hi_905 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_906;
  assign dataGroup_hi_hi_906 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_907;
  assign dataGroup_hi_hi_907 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_908;
  assign dataGroup_hi_hi_908 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_909;
  assign dataGroup_hi_hi_909 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_910;
  assign dataGroup_hi_hi_910 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_911;
  assign dataGroup_hi_hi_911 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_912;
  assign dataGroup_hi_hi_912 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_913;
  assign dataGroup_hi_hi_913 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_914;
  assign dataGroup_hi_hi_914 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_915;
  assign dataGroup_hi_hi_915 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_916;
  assign dataGroup_hi_hi_916 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_917;
  assign dataGroup_hi_hi_917 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_918;
  assign dataGroup_hi_hi_918 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_919;
  assign dataGroup_hi_hi_919 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_920;
  assign dataGroup_hi_hi_920 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_921;
  assign dataGroup_hi_hi_921 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_922;
  assign dataGroup_hi_hi_922 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_923;
  assign dataGroup_hi_hi_923 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_924;
  assign dataGroup_hi_hi_924 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_925;
  assign dataGroup_hi_hi_925 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_926;
  assign dataGroup_hi_hi_926 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_927;
  assign dataGroup_hi_hi_927 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_928;
  assign dataGroup_hi_hi_928 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_929;
  assign dataGroup_hi_hi_929 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_930;
  assign dataGroup_hi_hi_930 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_931;
  assign dataGroup_hi_hi_931 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_932;
  assign dataGroup_hi_hi_932 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_933;
  assign dataGroup_hi_hi_933 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_934;
  assign dataGroup_hi_hi_934 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_935;
  assign dataGroup_hi_hi_935 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_936;
  assign dataGroup_hi_hi_936 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_937;
  assign dataGroup_hi_hi_937 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_938;
  assign dataGroup_hi_hi_938 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_939;
  assign dataGroup_hi_hi_939 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_940;
  assign dataGroup_hi_hi_940 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_941;
  assign dataGroup_hi_hi_941 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_942;
  assign dataGroup_hi_hi_942 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_943;
  assign dataGroup_hi_hi_943 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_944;
  assign dataGroup_hi_hi_944 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_945;
  assign dataGroup_hi_hi_945 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_946;
  assign dataGroup_hi_hi_946 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_947;
  assign dataGroup_hi_hi_947 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_948;
  assign dataGroup_hi_hi_948 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_949;
  assign dataGroup_hi_hi_949 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_950;
  assign dataGroup_hi_hi_950 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_951;
  assign dataGroup_hi_hi_951 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_952;
  assign dataGroup_hi_hi_952 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_953;
  assign dataGroup_hi_hi_953 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_954;
  assign dataGroup_hi_hi_954 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_955;
  assign dataGroup_hi_hi_955 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_956;
  assign dataGroup_hi_hi_956 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_957;
  assign dataGroup_hi_hi_957 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_958;
  assign dataGroup_hi_hi_958 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_959;
  assign dataGroup_hi_hi_959 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_960;
  assign dataGroup_hi_hi_960 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_961;
  assign dataGroup_hi_hi_961 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_962;
  assign dataGroup_hi_hi_962 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_963;
  assign dataGroup_hi_hi_963 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_964;
  assign dataGroup_hi_hi_964 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_965;
  assign dataGroup_hi_hi_965 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_966;
  assign dataGroup_hi_hi_966 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_967;
  assign dataGroup_hi_hi_967 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_968;
  assign dataGroup_hi_hi_968 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_969;
  assign dataGroup_hi_hi_969 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_970;
  assign dataGroup_hi_hi_970 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_971;
  assign dataGroup_hi_hi_971 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_972;
  assign dataGroup_hi_hi_972 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_973;
  assign dataGroup_hi_hi_973 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_974;
  assign dataGroup_hi_hi_974 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_975;
  assign dataGroup_hi_hi_975 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_976;
  assign dataGroup_hi_hi_976 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_977;
  assign dataGroup_hi_hi_977 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_978;
  assign dataGroup_hi_hi_978 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_979;
  assign dataGroup_hi_hi_979 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_980;
  assign dataGroup_hi_hi_980 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_981;
  assign dataGroup_hi_hi_981 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_982;
  assign dataGroup_hi_hi_982 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_983;
  assign dataGroup_hi_hi_983 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_984;
  assign dataGroup_hi_hi_984 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_985;
  assign dataGroup_hi_hi_985 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_986;
  assign dataGroup_hi_hi_986 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_987;
  assign dataGroup_hi_hi_987 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_988;
  assign dataGroup_hi_hi_988 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_989;
  assign dataGroup_hi_hi_989 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_990;
  assign dataGroup_hi_hi_990 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_991;
  assign dataGroup_hi_hi_991 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_992;
  assign dataGroup_hi_hi_992 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_993;
  assign dataGroup_hi_hi_993 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_994;
  assign dataGroup_hi_hi_994 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_995;
  assign dataGroup_hi_hi_995 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_996;
  assign dataGroup_hi_hi_996 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_997;
  assign dataGroup_hi_hi_997 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_998;
  assign dataGroup_hi_hi_998 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_999;
  assign dataGroup_hi_hi_999 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1000;
  assign dataGroup_hi_hi_1000 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1001;
  assign dataGroup_hi_hi_1001 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1002;
  assign dataGroup_hi_hi_1002 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1003;
  assign dataGroup_hi_hi_1003 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1004;
  assign dataGroup_hi_hi_1004 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1005;
  assign dataGroup_hi_hi_1005 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1006;
  assign dataGroup_hi_hi_1006 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1007;
  assign dataGroup_hi_hi_1007 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1008;
  assign dataGroup_hi_hi_1008 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1009;
  assign dataGroup_hi_hi_1009 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1010;
  assign dataGroup_hi_hi_1010 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1011;
  assign dataGroup_hi_hi_1011 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1012;
  assign dataGroup_hi_hi_1012 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1013;
  assign dataGroup_hi_hi_1013 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1014;
  assign dataGroup_hi_hi_1014 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1015;
  assign dataGroup_hi_hi_1015 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1016;
  assign dataGroup_hi_hi_1016 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1017;
  assign dataGroup_hi_hi_1017 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1018;
  assign dataGroup_hi_hi_1018 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1019;
  assign dataGroup_hi_hi_1019 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1020;
  assign dataGroup_hi_hi_1020 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1021;
  assign dataGroup_hi_hi_1021 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1022;
  assign dataGroup_hi_hi_1022 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1023;
  assign dataGroup_hi_hi_1023 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1024;
  assign dataGroup_hi_hi_1024 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1025;
  assign dataGroup_hi_hi_1025 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1026;
  assign dataGroup_hi_hi_1026 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1027;
  assign dataGroup_hi_hi_1027 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1028;
  assign dataGroup_hi_hi_1028 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1029;
  assign dataGroup_hi_hi_1029 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1030;
  assign dataGroup_hi_hi_1030 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1031;
  assign dataGroup_hi_hi_1031 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1032;
  assign dataGroup_hi_hi_1032 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1033;
  assign dataGroup_hi_hi_1033 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1034;
  assign dataGroup_hi_hi_1034 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1035;
  assign dataGroup_hi_hi_1035 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1036;
  assign dataGroup_hi_hi_1036 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1037;
  assign dataGroup_hi_hi_1037 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1038;
  assign dataGroup_hi_hi_1038 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1039;
  assign dataGroup_hi_hi_1039 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1040;
  assign dataGroup_hi_hi_1040 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1041;
  assign dataGroup_hi_hi_1041 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1042;
  assign dataGroup_hi_hi_1042 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1043;
  assign dataGroup_hi_hi_1043 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1044;
  assign dataGroup_hi_hi_1044 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1045;
  assign dataGroup_hi_hi_1045 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1046;
  assign dataGroup_hi_hi_1046 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1047;
  assign dataGroup_hi_hi_1047 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1048;
  assign dataGroup_hi_hi_1048 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1049;
  assign dataGroup_hi_hi_1049 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1050;
  assign dataGroup_hi_hi_1050 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1051;
  assign dataGroup_hi_hi_1051 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1052;
  assign dataGroup_hi_hi_1052 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1053;
  assign dataGroup_hi_hi_1053 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1054;
  assign dataGroup_hi_hi_1054 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1055;
  assign dataGroup_hi_hi_1055 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1056;
  assign dataGroup_hi_hi_1056 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1057;
  assign dataGroup_hi_hi_1057 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1058;
  assign dataGroup_hi_hi_1058 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1059;
  assign dataGroup_hi_hi_1059 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1060;
  assign dataGroup_hi_hi_1060 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1061;
  assign dataGroup_hi_hi_1061 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1062;
  assign dataGroup_hi_hi_1062 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1063;
  assign dataGroup_hi_hi_1063 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1064;
  assign dataGroup_hi_hi_1064 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1065;
  assign dataGroup_hi_hi_1065 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1066;
  assign dataGroup_hi_hi_1066 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1067;
  assign dataGroup_hi_hi_1067 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1068;
  assign dataGroup_hi_hi_1068 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1069;
  assign dataGroup_hi_hi_1069 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1070;
  assign dataGroup_hi_hi_1070 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1071;
  assign dataGroup_hi_hi_1071 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1072;
  assign dataGroup_hi_hi_1072 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1073;
  assign dataGroup_hi_hi_1073 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1074;
  assign dataGroup_hi_hi_1074 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1075;
  assign dataGroup_hi_hi_1075 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1076;
  assign dataGroup_hi_hi_1076 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1077;
  assign dataGroup_hi_hi_1077 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1078;
  assign dataGroup_hi_hi_1078 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1079;
  assign dataGroup_hi_hi_1079 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1080;
  assign dataGroup_hi_hi_1080 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1081;
  assign dataGroup_hi_hi_1081 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1082;
  assign dataGroup_hi_hi_1082 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1083;
  assign dataGroup_hi_hi_1083 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1084;
  assign dataGroup_hi_hi_1084 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1085;
  assign dataGroup_hi_hi_1085 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1086;
  assign dataGroup_hi_hi_1086 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1087;
  assign dataGroup_hi_hi_1087 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1088;
  assign dataGroup_hi_hi_1088 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1089;
  assign dataGroup_hi_hi_1089 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1090;
  assign dataGroup_hi_hi_1090 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1091;
  assign dataGroup_hi_hi_1091 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1092;
  assign dataGroup_hi_hi_1092 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1093;
  assign dataGroup_hi_hi_1093 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1094;
  assign dataGroup_hi_hi_1094 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1095;
  assign dataGroup_hi_hi_1095 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1096;
  assign dataGroup_hi_hi_1096 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1097;
  assign dataGroup_hi_hi_1097 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1098;
  assign dataGroup_hi_hi_1098 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1099;
  assign dataGroup_hi_hi_1099 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1100;
  assign dataGroup_hi_hi_1100 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1101;
  assign dataGroup_hi_hi_1101 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1102;
  assign dataGroup_hi_hi_1102 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1103;
  assign dataGroup_hi_hi_1103 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1104;
  assign dataGroup_hi_hi_1104 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1105;
  assign dataGroup_hi_hi_1105 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1106;
  assign dataGroup_hi_hi_1106 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1107;
  assign dataGroup_hi_hi_1107 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1108;
  assign dataGroup_hi_hi_1108 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1109;
  assign dataGroup_hi_hi_1109 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1110;
  assign dataGroup_hi_hi_1110 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1111;
  assign dataGroup_hi_hi_1111 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1112;
  assign dataGroup_hi_hi_1112 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1113;
  assign dataGroup_hi_hi_1113 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1114;
  assign dataGroup_hi_hi_1114 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1115;
  assign dataGroup_hi_hi_1115 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1116;
  assign dataGroup_hi_hi_1116 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1117;
  assign dataGroup_hi_hi_1117 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1118;
  assign dataGroup_hi_hi_1118 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1119;
  assign dataGroup_hi_hi_1119 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1120;
  assign dataGroup_hi_hi_1120 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1121;
  assign dataGroup_hi_hi_1121 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1122;
  assign dataGroup_hi_hi_1122 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1123;
  assign dataGroup_hi_hi_1123 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1124;
  assign dataGroup_hi_hi_1124 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1125;
  assign dataGroup_hi_hi_1125 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1126;
  assign dataGroup_hi_hi_1126 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1127;
  assign dataGroup_hi_hi_1127 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1128;
  assign dataGroup_hi_hi_1128 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1129;
  assign dataGroup_hi_hi_1129 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1130;
  assign dataGroup_hi_hi_1130 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1131;
  assign dataGroup_hi_hi_1131 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1132;
  assign dataGroup_hi_hi_1132 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1133;
  assign dataGroup_hi_hi_1133 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1134;
  assign dataGroup_hi_hi_1134 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1135;
  assign dataGroup_hi_hi_1135 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1136;
  assign dataGroup_hi_hi_1136 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1137;
  assign dataGroup_hi_hi_1137 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1138;
  assign dataGroup_hi_hi_1138 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1139;
  assign dataGroup_hi_hi_1139 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1140;
  assign dataGroup_hi_hi_1140 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1141;
  assign dataGroup_hi_hi_1141 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1142;
  assign dataGroup_hi_hi_1142 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1143;
  assign dataGroup_hi_hi_1143 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1144;
  assign dataGroup_hi_hi_1144 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1145;
  assign dataGroup_hi_hi_1145 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1146;
  assign dataGroup_hi_hi_1146 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1147;
  assign dataGroup_hi_hi_1147 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1148;
  assign dataGroup_hi_hi_1148 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1149;
  assign dataGroup_hi_hi_1149 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1150;
  assign dataGroup_hi_hi_1150 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1151;
  assign dataGroup_hi_hi_1151 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1152;
  assign dataGroup_hi_hi_1152 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1153;
  assign dataGroup_hi_hi_1153 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1154;
  assign dataGroup_hi_hi_1154 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1155;
  assign dataGroup_hi_hi_1155 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1156;
  assign dataGroup_hi_hi_1156 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1157;
  assign dataGroup_hi_hi_1157 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1158;
  assign dataGroup_hi_hi_1158 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1159;
  assign dataGroup_hi_hi_1159 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1160;
  assign dataGroup_hi_hi_1160 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1161;
  assign dataGroup_hi_hi_1161 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1162;
  assign dataGroup_hi_hi_1162 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1163;
  assign dataGroup_hi_hi_1163 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1164;
  assign dataGroup_hi_hi_1164 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1165;
  assign dataGroup_hi_hi_1165 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1166;
  assign dataGroup_hi_hi_1166 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1167;
  assign dataGroup_hi_hi_1167 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1168;
  assign dataGroup_hi_hi_1168 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1169;
  assign dataGroup_hi_hi_1169 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1170;
  assign dataGroup_hi_hi_1170 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1171;
  assign dataGroup_hi_hi_1171 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1172;
  assign dataGroup_hi_hi_1172 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1173;
  assign dataGroup_hi_hi_1173 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1174;
  assign dataGroup_hi_hi_1174 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1175;
  assign dataGroup_hi_hi_1175 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1176;
  assign dataGroup_hi_hi_1176 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1177;
  assign dataGroup_hi_hi_1177 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1178;
  assign dataGroup_hi_hi_1178 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1179;
  assign dataGroup_hi_hi_1179 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1180;
  assign dataGroup_hi_hi_1180 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1181;
  assign dataGroup_hi_hi_1181 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1182;
  assign dataGroup_hi_hi_1182 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1183;
  assign dataGroup_hi_hi_1183 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1184;
  assign dataGroup_hi_hi_1184 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1185;
  assign dataGroup_hi_hi_1185 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1186;
  assign dataGroup_hi_hi_1186 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1187;
  assign dataGroup_hi_hi_1187 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1188;
  assign dataGroup_hi_hi_1188 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1189;
  assign dataGroup_hi_hi_1189 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1190;
  assign dataGroup_hi_hi_1190 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1191;
  assign dataGroup_hi_hi_1191 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1192;
  assign dataGroup_hi_hi_1192 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1193;
  assign dataGroup_hi_hi_1193 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1194;
  assign dataGroup_hi_hi_1194 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1195;
  assign dataGroup_hi_hi_1195 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1196;
  assign dataGroup_hi_hi_1196 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1197;
  assign dataGroup_hi_hi_1197 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1198;
  assign dataGroup_hi_hi_1198 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1199;
  assign dataGroup_hi_hi_1199 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1200;
  assign dataGroup_hi_hi_1200 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1201;
  assign dataGroup_hi_hi_1201 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1202;
  assign dataGroup_hi_hi_1202 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1203;
  assign dataGroup_hi_hi_1203 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1204;
  assign dataGroup_hi_hi_1204 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1205;
  assign dataGroup_hi_hi_1205 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1206;
  assign dataGroup_hi_hi_1206 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1207;
  assign dataGroup_hi_hi_1207 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1208;
  assign dataGroup_hi_hi_1208 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1209;
  assign dataGroup_hi_hi_1209 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1210;
  assign dataGroup_hi_hi_1210 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1211;
  assign dataGroup_hi_hi_1211 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1212;
  assign dataGroup_hi_hi_1212 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1213;
  assign dataGroup_hi_hi_1213 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1214;
  assign dataGroup_hi_hi_1214 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1215;
  assign dataGroup_hi_hi_1215 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1216;
  assign dataGroup_hi_hi_1216 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1217;
  assign dataGroup_hi_hi_1217 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1218;
  assign dataGroup_hi_hi_1218 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1219;
  assign dataGroup_hi_hi_1219 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1220;
  assign dataGroup_hi_hi_1220 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1221;
  assign dataGroup_hi_hi_1221 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1222;
  assign dataGroup_hi_hi_1222 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1223;
  assign dataGroup_hi_hi_1223 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1224;
  assign dataGroup_hi_hi_1224 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1225;
  assign dataGroup_hi_hi_1225 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1226;
  assign dataGroup_hi_hi_1226 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1227;
  assign dataGroup_hi_hi_1227 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1228;
  assign dataGroup_hi_hi_1228 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1229;
  assign dataGroup_hi_hi_1229 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1230;
  assign dataGroup_hi_hi_1230 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1231;
  assign dataGroup_hi_hi_1231 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1232;
  assign dataGroup_hi_hi_1232 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1233;
  assign dataGroup_hi_hi_1233 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1234;
  assign dataGroup_hi_hi_1234 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1235;
  assign dataGroup_hi_hi_1235 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1236;
  assign dataGroup_hi_hi_1236 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1237;
  assign dataGroup_hi_hi_1237 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1238;
  assign dataGroup_hi_hi_1238 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1239;
  assign dataGroup_hi_hi_1239 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1240;
  assign dataGroup_hi_hi_1240 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1241;
  assign dataGroup_hi_hi_1241 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1242;
  assign dataGroup_hi_hi_1242 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1243;
  assign dataGroup_hi_hi_1243 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1244;
  assign dataGroup_hi_hi_1244 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1245;
  assign dataGroup_hi_hi_1245 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1246;
  assign dataGroup_hi_hi_1246 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1247;
  assign dataGroup_hi_hi_1247 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1248;
  assign dataGroup_hi_hi_1248 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1249;
  assign dataGroup_hi_hi_1249 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1250;
  assign dataGroup_hi_hi_1250 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1251;
  assign dataGroup_hi_hi_1251 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1252;
  assign dataGroup_hi_hi_1252 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1253;
  assign dataGroup_hi_hi_1253 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1254;
  assign dataGroup_hi_hi_1254 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1255;
  assign dataGroup_hi_hi_1255 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1256;
  assign dataGroup_hi_hi_1256 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1257;
  assign dataGroup_hi_hi_1257 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1258;
  assign dataGroup_hi_hi_1258 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1259;
  assign dataGroup_hi_hi_1259 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1260;
  assign dataGroup_hi_hi_1260 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1261;
  assign dataGroup_hi_hi_1261 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1262;
  assign dataGroup_hi_hi_1262 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1263;
  assign dataGroup_hi_hi_1263 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1264;
  assign dataGroup_hi_hi_1264 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1265;
  assign dataGroup_hi_hi_1265 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1266;
  assign dataGroup_hi_hi_1266 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1267;
  assign dataGroup_hi_hi_1267 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1268;
  assign dataGroup_hi_hi_1268 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1269;
  assign dataGroup_hi_hi_1269 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1270;
  assign dataGroup_hi_hi_1270 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1271;
  assign dataGroup_hi_hi_1271 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1272;
  assign dataGroup_hi_hi_1272 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1273;
  assign dataGroup_hi_hi_1273 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1274;
  assign dataGroup_hi_hi_1274 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1275;
  assign dataGroup_hi_hi_1275 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1276;
  assign dataGroup_hi_hi_1276 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1277;
  assign dataGroup_hi_hi_1277 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1278;
  assign dataGroup_hi_hi_1278 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1279;
  assign dataGroup_hi_hi_1279 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1280;
  assign dataGroup_hi_hi_1280 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1281;
  assign dataGroup_hi_hi_1281 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1282;
  assign dataGroup_hi_hi_1282 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1283;
  assign dataGroup_hi_hi_1283 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1284;
  assign dataGroup_hi_hi_1284 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1285;
  assign dataGroup_hi_hi_1285 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1286;
  assign dataGroup_hi_hi_1286 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1287;
  assign dataGroup_hi_hi_1287 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1288;
  assign dataGroup_hi_hi_1288 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1289;
  assign dataGroup_hi_hi_1289 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1290;
  assign dataGroup_hi_hi_1290 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1291;
  assign dataGroup_hi_hi_1291 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1292;
  assign dataGroup_hi_hi_1292 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1293;
  assign dataGroup_hi_hi_1293 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1294;
  assign dataGroup_hi_hi_1294 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1295;
  assign dataGroup_hi_hi_1295 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1296;
  assign dataGroup_hi_hi_1296 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1297;
  assign dataGroup_hi_hi_1297 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1298;
  assign dataGroup_hi_hi_1298 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1299;
  assign dataGroup_hi_hi_1299 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1300;
  assign dataGroup_hi_hi_1300 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1301;
  assign dataGroup_hi_hi_1301 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1302;
  assign dataGroup_hi_hi_1302 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1303;
  assign dataGroup_hi_hi_1303 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1304;
  assign dataGroup_hi_hi_1304 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1305;
  assign dataGroup_hi_hi_1305 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1306;
  assign dataGroup_hi_hi_1306 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1307;
  assign dataGroup_hi_hi_1307 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1308;
  assign dataGroup_hi_hi_1308 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1309;
  assign dataGroup_hi_hi_1309 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1310;
  assign dataGroup_hi_hi_1310 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1311;
  assign dataGroup_hi_hi_1311 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1312;
  assign dataGroup_hi_hi_1312 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1313;
  assign dataGroup_hi_hi_1313 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1314;
  assign dataGroup_hi_hi_1314 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1315;
  assign dataGroup_hi_hi_1315 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1316;
  assign dataGroup_hi_hi_1316 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1317;
  assign dataGroup_hi_hi_1317 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1318;
  assign dataGroup_hi_hi_1318 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1319;
  assign dataGroup_hi_hi_1319 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1320;
  assign dataGroup_hi_hi_1320 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1321;
  assign dataGroup_hi_hi_1321 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1322;
  assign dataGroup_hi_hi_1322 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1323;
  assign dataGroup_hi_hi_1323 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1324;
  assign dataGroup_hi_hi_1324 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1325;
  assign dataGroup_hi_hi_1325 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1326;
  assign dataGroup_hi_hi_1326 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1327;
  assign dataGroup_hi_hi_1327 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1328;
  assign dataGroup_hi_hi_1328 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1329;
  assign dataGroup_hi_hi_1329 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1330;
  assign dataGroup_hi_hi_1330 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1331;
  assign dataGroup_hi_hi_1331 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1332;
  assign dataGroup_hi_hi_1332 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1333;
  assign dataGroup_hi_hi_1333 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1334;
  assign dataGroup_hi_hi_1334 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1335;
  assign dataGroup_hi_hi_1335 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1336;
  assign dataGroup_hi_hi_1336 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1337;
  assign dataGroup_hi_hi_1337 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1338;
  assign dataGroup_hi_hi_1338 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1339;
  assign dataGroup_hi_hi_1339 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1340;
  assign dataGroup_hi_hi_1340 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1341;
  assign dataGroup_hi_hi_1341 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1342;
  assign dataGroup_hi_hi_1342 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1343;
  assign dataGroup_hi_hi_1343 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1344;
  assign dataGroup_hi_hi_1344 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1345;
  assign dataGroup_hi_hi_1345 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1346;
  assign dataGroup_hi_hi_1346 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1347;
  assign dataGroup_hi_hi_1347 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1348;
  assign dataGroup_hi_hi_1348 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1349;
  assign dataGroup_hi_hi_1349 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1350;
  assign dataGroup_hi_hi_1350 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1351;
  assign dataGroup_hi_hi_1351 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1352;
  assign dataGroup_hi_hi_1352 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1353;
  assign dataGroup_hi_hi_1353 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1354;
  assign dataGroup_hi_hi_1354 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1355;
  assign dataGroup_hi_hi_1355 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1356;
  assign dataGroup_hi_hi_1356 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1357;
  assign dataGroup_hi_hi_1357 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1358;
  assign dataGroup_hi_hi_1358 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1359;
  assign dataGroup_hi_hi_1359 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1360;
  assign dataGroup_hi_hi_1360 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1361;
  assign dataGroup_hi_hi_1361 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1362;
  assign dataGroup_hi_hi_1362 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1363;
  assign dataGroup_hi_hi_1363 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1364;
  assign dataGroup_hi_hi_1364 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1365;
  assign dataGroup_hi_hi_1365 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1366;
  assign dataGroup_hi_hi_1366 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1367;
  assign dataGroup_hi_hi_1367 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1368;
  assign dataGroup_hi_hi_1368 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1369;
  assign dataGroup_hi_hi_1369 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1370;
  assign dataGroup_hi_hi_1370 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1371;
  assign dataGroup_hi_hi_1371 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1372;
  assign dataGroup_hi_hi_1372 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1373;
  assign dataGroup_hi_hi_1373 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1374;
  assign dataGroup_hi_hi_1374 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1375;
  assign dataGroup_hi_hi_1375 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1376;
  assign dataGroup_hi_hi_1376 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1377;
  assign dataGroup_hi_hi_1377 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1378;
  assign dataGroup_hi_hi_1378 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1379;
  assign dataGroup_hi_hi_1379 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1380;
  assign dataGroup_hi_hi_1380 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1381;
  assign dataGroup_hi_hi_1381 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1382;
  assign dataGroup_hi_hi_1382 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1383;
  assign dataGroup_hi_hi_1383 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1384;
  assign dataGroup_hi_hi_1384 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1385;
  assign dataGroup_hi_hi_1385 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1386;
  assign dataGroup_hi_hi_1386 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1387;
  assign dataGroup_hi_hi_1387 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1388;
  assign dataGroup_hi_hi_1388 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1389;
  assign dataGroup_hi_hi_1389 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1390;
  assign dataGroup_hi_hi_1390 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1391;
  assign dataGroup_hi_hi_1391 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1392;
  assign dataGroup_hi_hi_1392 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1393;
  assign dataGroup_hi_hi_1393 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1394;
  assign dataGroup_hi_hi_1394 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1395;
  assign dataGroup_hi_hi_1395 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1396;
  assign dataGroup_hi_hi_1396 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1397;
  assign dataGroup_hi_hi_1397 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1398;
  assign dataGroup_hi_hi_1398 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1399;
  assign dataGroup_hi_hi_1399 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1400;
  assign dataGroup_hi_hi_1400 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1401;
  assign dataGroup_hi_hi_1401 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1402;
  assign dataGroup_hi_hi_1402 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1403;
  assign dataGroup_hi_hi_1403 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1404;
  assign dataGroup_hi_hi_1404 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1405;
  assign dataGroup_hi_hi_1405 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1406;
  assign dataGroup_hi_hi_1406 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1407;
  assign dataGroup_hi_hi_1407 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1408;
  assign dataGroup_hi_hi_1408 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1409;
  assign dataGroup_hi_hi_1409 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1410;
  assign dataGroup_hi_hi_1410 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1411;
  assign dataGroup_hi_hi_1411 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1412;
  assign dataGroup_hi_hi_1412 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1413;
  assign dataGroup_hi_hi_1413 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1414;
  assign dataGroup_hi_hi_1414 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1415;
  assign dataGroup_hi_hi_1415 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1416;
  assign dataGroup_hi_hi_1416 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1417;
  assign dataGroup_hi_hi_1417 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1418;
  assign dataGroup_hi_hi_1418 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1419;
  assign dataGroup_hi_hi_1419 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1420;
  assign dataGroup_hi_hi_1420 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1421;
  assign dataGroup_hi_hi_1421 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1422;
  assign dataGroup_hi_hi_1422 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1423;
  assign dataGroup_hi_hi_1423 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1424;
  assign dataGroup_hi_hi_1424 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1425;
  assign dataGroup_hi_hi_1425 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1426;
  assign dataGroup_hi_hi_1426 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1427;
  assign dataGroup_hi_hi_1427 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1428;
  assign dataGroup_hi_hi_1428 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1429;
  assign dataGroup_hi_hi_1429 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1430;
  assign dataGroup_hi_hi_1430 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1431;
  assign dataGroup_hi_hi_1431 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1432;
  assign dataGroup_hi_hi_1432 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1433;
  assign dataGroup_hi_hi_1433 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1434;
  assign dataGroup_hi_hi_1434 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1435;
  assign dataGroup_hi_hi_1435 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1436;
  assign dataGroup_hi_hi_1436 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1437;
  assign dataGroup_hi_hi_1437 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1438;
  assign dataGroup_hi_hi_1438 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1439;
  assign dataGroup_hi_hi_1439 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1440;
  assign dataGroup_hi_hi_1440 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1441;
  assign dataGroup_hi_hi_1441 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1442;
  assign dataGroup_hi_hi_1442 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1443;
  assign dataGroup_hi_hi_1443 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1444;
  assign dataGroup_hi_hi_1444 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1445;
  assign dataGroup_hi_hi_1445 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1446;
  assign dataGroup_hi_hi_1446 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1447;
  assign dataGroup_hi_hi_1447 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1448;
  assign dataGroup_hi_hi_1448 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1449;
  assign dataGroup_hi_hi_1449 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1450;
  assign dataGroup_hi_hi_1450 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1451;
  assign dataGroup_hi_hi_1451 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1452;
  assign dataGroup_hi_hi_1452 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1453;
  assign dataGroup_hi_hi_1453 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1454;
  assign dataGroup_hi_hi_1454 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1455;
  assign dataGroup_hi_hi_1455 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1456;
  assign dataGroup_hi_hi_1456 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1457;
  assign dataGroup_hi_hi_1457 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1458;
  assign dataGroup_hi_hi_1458 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1459;
  assign dataGroup_hi_hi_1459 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1460;
  assign dataGroup_hi_hi_1460 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1461;
  assign dataGroup_hi_hi_1461 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1462;
  assign dataGroup_hi_hi_1462 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1463;
  assign dataGroup_hi_hi_1463 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1464;
  assign dataGroup_hi_hi_1464 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1465;
  assign dataGroup_hi_hi_1465 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1466;
  assign dataGroup_hi_hi_1466 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1467;
  assign dataGroup_hi_hi_1467 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1468;
  assign dataGroup_hi_hi_1468 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1469;
  assign dataGroup_hi_hi_1469 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1470;
  assign dataGroup_hi_hi_1470 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1471;
  assign dataGroup_hi_hi_1471 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1472;
  assign dataGroup_hi_hi_1472 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1473;
  assign dataGroup_hi_hi_1473 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1474;
  assign dataGroup_hi_hi_1474 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1475;
  assign dataGroup_hi_hi_1475 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1476;
  assign dataGroup_hi_hi_1476 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1477;
  assign dataGroup_hi_hi_1477 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1478;
  assign dataGroup_hi_hi_1478 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1479;
  assign dataGroup_hi_hi_1479 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1480;
  assign dataGroup_hi_hi_1480 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1481;
  assign dataGroup_hi_hi_1481 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1482;
  assign dataGroup_hi_hi_1482 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1483;
  assign dataGroup_hi_hi_1483 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1484;
  assign dataGroup_hi_hi_1484 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1485;
  assign dataGroup_hi_hi_1485 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1486;
  assign dataGroup_hi_hi_1486 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1487;
  assign dataGroup_hi_hi_1487 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1488;
  assign dataGroup_hi_hi_1488 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1489;
  assign dataGroup_hi_hi_1489 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1490;
  assign dataGroup_hi_hi_1490 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1491;
  assign dataGroup_hi_hi_1491 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1492;
  assign dataGroup_hi_hi_1492 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1493;
  assign dataGroup_hi_hi_1493 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1494;
  assign dataGroup_hi_hi_1494 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1495;
  assign dataGroup_hi_hi_1495 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1496;
  assign dataGroup_hi_hi_1496 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1497;
  assign dataGroup_hi_hi_1497 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1498;
  assign dataGroup_hi_hi_1498 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1499;
  assign dataGroup_hi_hi_1499 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1500;
  assign dataGroup_hi_hi_1500 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1501;
  assign dataGroup_hi_hi_1501 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1502;
  assign dataGroup_hi_hi_1502 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1503;
  assign dataGroup_hi_hi_1503 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1504;
  assign dataGroup_hi_hi_1504 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1505;
  assign dataGroup_hi_hi_1505 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1506;
  assign dataGroup_hi_hi_1506 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1507;
  assign dataGroup_hi_hi_1507 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1508;
  assign dataGroup_hi_hi_1508 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1509;
  assign dataGroup_hi_hi_1509 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1510;
  assign dataGroup_hi_hi_1510 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1511;
  assign dataGroup_hi_hi_1511 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1512;
  assign dataGroup_hi_hi_1512 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1513;
  assign dataGroup_hi_hi_1513 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1514;
  assign dataGroup_hi_hi_1514 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1515;
  assign dataGroup_hi_hi_1515 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1516;
  assign dataGroup_hi_hi_1516 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1517;
  assign dataGroup_hi_hi_1517 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1518;
  assign dataGroup_hi_hi_1518 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1519;
  assign dataGroup_hi_hi_1519 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1520;
  assign dataGroup_hi_hi_1520 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1521;
  assign dataGroup_hi_hi_1521 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1522;
  assign dataGroup_hi_hi_1522 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1523;
  assign dataGroup_hi_hi_1523 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1524;
  assign dataGroup_hi_hi_1524 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1525;
  assign dataGroup_hi_hi_1525 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1526;
  assign dataGroup_hi_hi_1526 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1527;
  assign dataGroup_hi_hi_1527 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1528;
  assign dataGroup_hi_hi_1528 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1529;
  assign dataGroup_hi_hi_1529 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1530;
  assign dataGroup_hi_hi_1530 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1531;
  assign dataGroup_hi_hi_1531 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1532;
  assign dataGroup_hi_hi_1532 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1533;
  assign dataGroup_hi_hi_1533 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1534;
  assign dataGroup_hi_hi_1534 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1535;
  assign dataGroup_hi_hi_1535 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1536;
  assign dataGroup_hi_hi_1536 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1537;
  assign dataGroup_hi_hi_1537 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1538;
  assign dataGroup_hi_hi_1538 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1539;
  assign dataGroup_hi_hi_1539 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1540;
  assign dataGroup_hi_hi_1540 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1541;
  assign dataGroup_hi_hi_1541 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1542;
  assign dataGroup_hi_hi_1542 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1543;
  assign dataGroup_hi_hi_1543 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1544;
  assign dataGroup_hi_hi_1544 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1545;
  assign dataGroup_hi_hi_1545 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1546;
  assign dataGroup_hi_hi_1546 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1547;
  assign dataGroup_hi_hi_1547 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1548;
  assign dataGroup_hi_hi_1548 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1549;
  assign dataGroup_hi_hi_1549 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1550;
  assign dataGroup_hi_hi_1550 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1551;
  assign dataGroup_hi_hi_1551 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1552;
  assign dataGroup_hi_hi_1552 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1553;
  assign dataGroup_hi_hi_1553 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1554;
  assign dataGroup_hi_hi_1554 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1555;
  assign dataGroup_hi_hi_1555 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1556;
  assign dataGroup_hi_hi_1556 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1557;
  assign dataGroup_hi_hi_1557 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1558;
  assign dataGroup_hi_hi_1558 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1559;
  assign dataGroup_hi_hi_1559 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1560;
  assign dataGroup_hi_hi_1560 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1561;
  assign dataGroup_hi_hi_1561 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1562;
  assign dataGroup_hi_hi_1562 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1563;
  assign dataGroup_hi_hi_1563 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1564;
  assign dataGroup_hi_hi_1564 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1565;
  assign dataGroup_hi_hi_1565 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1566;
  assign dataGroup_hi_hi_1566 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1567;
  assign dataGroup_hi_hi_1567 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1568;
  assign dataGroup_hi_hi_1568 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1569;
  assign dataGroup_hi_hi_1569 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1570;
  assign dataGroup_hi_hi_1570 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1571;
  assign dataGroup_hi_hi_1571 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1572;
  assign dataGroup_hi_hi_1572 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1573;
  assign dataGroup_hi_hi_1573 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1574;
  assign dataGroup_hi_hi_1574 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1575;
  assign dataGroup_hi_hi_1575 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1576;
  assign dataGroup_hi_hi_1576 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1577;
  assign dataGroup_hi_hi_1577 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1578;
  assign dataGroup_hi_hi_1578 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1579;
  assign dataGroup_hi_hi_1579 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1580;
  assign dataGroup_hi_hi_1580 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1581;
  assign dataGroup_hi_hi_1581 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1582;
  assign dataGroup_hi_hi_1582 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1583;
  assign dataGroup_hi_hi_1583 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1584;
  assign dataGroup_hi_hi_1584 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1585;
  assign dataGroup_hi_hi_1585 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1586;
  assign dataGroup_hi_hi_1586 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1587;
  assign dataGroup_hi_hi_1587 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1588;
  assign dataGroup_hi_hi_1588 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1589;
  assign dataGroup_hi_hi_1589 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1590;
  assign dataGroup_hi_hi_1590 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1591;
  assign dataGroup_hi_hi_1591 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1592;
  assign dataGroup_hi_hi_1592 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1593;
  assign dataGroup_hi_hi_1593 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1594;
  assign dataGroup_hi_hi_1594 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1595;
  assign dataGroup_hi_hi_1595 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1596;
  assign dataGroup_hi_hi_1596 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1597;
  assign dataGroup_hi_hi_1597 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1598;
  assign dataGroup_hi_hi_1598 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1599;
  assign dataGroup_hi_hi_1599 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1600;
  assign dataGroup_hi_hi_1600 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1601;
  assign dataGroup_hi_hi_1601 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1602;
  assign dataGroup_hi_hi_1602 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1603;
  assign dataGroup_hi_hi_1603 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1604;
  assign dataGroup_hi_hi_1604 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1605;
  assign dataGroup_hi_hi_1605 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1606;
  assign dataGroup_hi_hi_1606 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1607;
  assign dataGroup_hi_hi_1607 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1608;
  assign dataGroup_hi_hi_1608 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1609;
  assign dataGroup_hi_hi_1609 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1610;
  assign dataGroup_hi_hi_1610 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1611;
  assign dataGroup_hi_hi_1611 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1612;
  assign dataGroup_hi_hi_1612 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1613;
  assign dataGroup_hi_hi_1613 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1614;
  assign dataGroup_hi_hi_1614 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1615;
  assign dataGroup_hi_hi_1615 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1616;
  assign dataGroup_hi_hi_1616 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1617;
  assign dataGroup_hi_hi_1617 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1618;
  assign dataGroup_hi_hi_1618 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1619;
  assign dataGroup_hi_hi_1619 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1620;
  assign dataGroup_hi_hi_1620 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1621;
  assign dataGroup_hi_hi_1621 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1622;
  assign dataGroup_hi_hi_1622 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1623;
  assign dataGroup_hi_hi_1623 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1624;
  assign dataGroup_hi_hi_1624 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1625;
  assign dataGroup_hi_hi_1625 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1626;
  assign dataGroup_hi_hi_1626 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1627;
  assign dataGroup_hi_hi_1627 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1628;
  assign dataGroup_hi_hi_1628 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1629;
  assign dataGroup_hi_hi_1629 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1630;
  assign dataGroup_hi_hi_1630 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1631;
  assign dataGroup_hi_hi_1631 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1632;
  assign dataGroup_hi_hi_1632 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1633;
  assign dataGroup_hi_hi_1633 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1634;
  assign dataGroup_hi_hi_1634 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1635;
  assign dataGroup_hi_hi_1635 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1636;
  assign dataGroup_hi_hi_1636 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1637;
  assign dataGroup_hi_hi_1637 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1638;
  assign dataGroup_hi_hi_1638 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1639;
  assign dataGroup_hi_hi_1639 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1640;
  assign dataGroup_hi_hi_1640 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1641;
  assign dataGroup_hi_hi_1641 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1642;
  assign dataGroup_hi_hi_1642 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1643;
  assign dataGroup_hi_hi_1643 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1644;
  assign dataGroup_hi_hi_1644 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1645;
  assign dataGroup_hi_hi_1645 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1646;
  assign dataGroup_hi_hi_1646 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1647;
  assign dataGroup_hi_hi_1647 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1648;
  assign dataGroup_hi_hi_1648 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1649;
  assign dataGroup_hi_hi_1649 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1650;
  assign dataGroup_hi_hi_1650 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1651;
  assign dataGroup_hi_hi_1651 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1652;
  assign dataGroup_hi_hi_1652 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1653;
  assign dataGroup_hi_hi_1653 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1654;
  assign dataGroup_hi_hi_1654 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1655;
  assign dataGroup_hi_hi_1655 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1656;
  assign dataGroup_hi_hi_1656 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1657;
  assign dataGroup_hi_hi_1657 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1658;
  assign dataGroup_hi_hi_1658 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1659;
  assign dataGroup_hi_hi_1659 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1660;
  assign dataGroup_hi_hi_1660 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1661;
  assign dataGroup_hi_hi_1661 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1662;
  assign dataGroup_hi_hi_1662 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1663;
  assign dataGroup_hi_hi_1663 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1664;
  assign dataGroup_hi_hi_1664 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1665;
  assign dataGroup_hi_hi_1665 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1666;
  assign dataGroup_hi_hi_1666 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1667;
  assign dataGroup_hi_hi_1667 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1668;
  assign dataGroup_hi_hi_1668 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1669;
  assign dataGroup_hi_hi_1669 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1670;
  assign dataGroup_hi_hi_1670 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1671;
  assign dataGroup_hi_hi_1671 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1672;
  assign dataGroup_hi_hi_1672 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1673;
  assign dataGroup_hi_hi_1673 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1674;
  assign dataGroup_hi_hi_1674 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1675;
  assign dataGroup_hi_hi_1675 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1676;
  assign dataGroup_hi_hi_1676 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1677;
  assign dataGroup_hi_hi_1677 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1678;
  assign dataGroup_hi_hi_1678 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1679;
  assign dataGroup_hi_hi_1679 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1680;
  assign dataGroup_hi_hi_1680 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1681;
  assign dataGroup_hi_hi_1681 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1682;
  assign dataGroup_hi_hi_1682 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1683;
  assign dataGroup_hi_hi_1683 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1684;
  assign dataGroup_hi_hi_1684 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1685;
  assign dataGroup_hi_hi_1685 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1686;
  assign dataGroup_hi_hi_1686 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1687;
  assign dataGroup_hi_hi_1687 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1688;
  assign dataGroup_hi_hi_1688 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1689;
  assign dataGroup_hi_hi_1689 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1690;
  assign dataGroup_hi_hi_1690 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1691;
  assign dataGroup_hi_hi_1691 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1692;
  assign dataGroup_hi_hi_1692 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1693;
  assign dataGroup_hi_hi_1693 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1694;
  assign dataGroup_hi_hi_1694 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1695;
  assign dataGroup_hi_hi_1695 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1696;
  assign dataGroup_hi_hi_1696 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1697;
  assign dataGroup_hi_hi_1697 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1698;
  assign dataGroup_hi_hi_1698 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1699;
  assign dataGroup_hi_hi_1699 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1700;
  assign dataGroup_hi_hi_1700 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1701;
  assign dataGroup_hi_hi_1701 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1702;
  assign dataGroup_hi_hi_1702 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1703;
  assign dataGroup_hi_hi_1703 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1704;
  assign dataGroup_hi_hi_1704 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1705;
  assign dataGroup_hi_hi_1705 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1706;
  assign dataGroup_hi_hi_1706 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1707;
  assign dataGroup_hi_hi_1707 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1708;
  assign dataGroup_hi_hi_1708 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1709;
  assign dataGroup_hi_hi_1709 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1710;
  assign dataGroup_hi_hi_1710 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1711;
  assign dataGroup_hi_hi_1711 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1712;
  assign dataGroup_hi_hi_1712 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1713;
  assign dataGroup_hi_hi_1713 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1714;
  assign dataGroup_hi_hi_1714 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1715;
  assign dataGroup_hi_hi_1715 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1716;
  assign dataGroup_hi_hi_1716 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1717;
  assign dataGroup_hi_hi_1717 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1718;
  assign dataGroup_hi_hi_1718 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1719;
  assign dataGroup_hi_hi_1719 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1720;
  assign dataGroup_hi_hi_1720 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1721;
  assign dataGroup_hi_hi_1721 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1722;
  assign dataGroup_hi_hi_1722 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1723;
  assign dataGroup_hi_hi_1723 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1724;
  assign dataGroup_hi_hi_1724 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1725;
  assign dataGroup_hi_hi_1725 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1726;
  assign dataGroup_hi_hi_1726 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1727;
  assign dataGroup_hi_hi_1727 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1728;
  assign dataGroup_hi_hi_1728 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1729;
  assign dataGroup_hi_hi_1729 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1730;
  assign dataGroup_hi_hi_1730 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1731;
  assign dataGroup_hi_hi_1731 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1732;
  assign dataGroup_hi_hi_1732 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1733;
  assign dataGroup_hi_hi_1733 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1734;
  assign dataGroup_hi_hi_1734 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1735;
  assign dataGroup_hi_hi_1735 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1736;
  assign dataGroup_hi_hi_1736 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1737;
  assign dataGroup_hi_hi_1737 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1738;
  assign dataGroup_hi_hi_1738 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1739;
  assign dataGroup_hi_hi_1739 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1740;
  assign dataGroup_hi_hi_1740 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1741;
  assign dataGroup_hi_hi_1741 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1742;
  assign dataGroup_hi_hi_1742 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1743;
  assign dataGroup_hi_hi_1743 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1744;
  assign dataGroup_hi_hi_1744 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1745;
  assign dataGroup_hi_hi_1745 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1746;
  assign dataGroup_hi_hi_1746 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1747;
  assign dataGroup_hi_hi_1747 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1748;
  assign dataGroup_hi_hi_1748 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1749;
  assign dataGroup_hi_hi_1749 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1750;
  assign dataGroup_hi_hi_1750 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1751;
  assign dataGroup_hi_hi_1751 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1752;
  assign dataGroup_hi_hi_1752 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1753;
  assign dataGroup_hi_hi_1753 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1754;
  assign dataGroup_hi_hi_1754 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1755;
  assign dataGroup_hi_hi_1755 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1756;
  assign dataGroup_hi_hi_1756 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1757;
  assign dataGroup_hi_hi_1757 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1758;
  assign dataGroup_hi_hi_1758 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1759;
  assign dataGroup_hi_hi_1759 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1760;
  assign dataGroup_hi_hi_1760 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1761;
  assign dataGroup_hi_hi_1761 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1762;
  assign dataGroup_hi_hi_1762 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1763;
  assign dataGroup_hi_hi_1763 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1764;
  assign dataGroup_hi_hi_1764 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1765;
  assign dataGroup_hi_hi_1765 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1766;
  assign dataGroup_hi_hi_1766 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1767;
  assign dataGroup_hi_hi_1767 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1768;
  assign dataGroup_hi_hi_1768 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1769;
  assign dataGroup_hi_hi_1769 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1770;
  assign dataGroup_hi_hi_1770 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1771;
  assign dataGroup_hi_hi_1771 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1772;
  assign dataGroup_hi_hi_1772 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1773;
  assign dataGroup_hi_hi_1773 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1774;
  assign dataGroup_hi_hi_1774 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1775;
  assign dataGroup_hi_hi_1775 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1776;
  assign dataGroup_hi_hi_1776 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1777;
  assign dataGroup_hi_hi_1777 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1778;
  assign dataGroup_hi_hi_1778 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1779;
  assign dataGroup_hi_hi_1779 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1780;
  assign dataGroup_hi_hi_1780 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1781;
  assign dataGroup_hi_hi_1781 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1782;
  assign dataGroup_hi_hi_1782 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1783;
  assign dataGroup_hi_hi_1783 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1784;
  assign dataGroup_hi_hi_1784 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1785;
  assign dataGroup_hi_hi_1785 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1786;
  assign dataGroup_hi_hi_1786 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1787;
  assign dataGroup_hi_hi_1787 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1788;
  assign dataGroup_hi_hi_1788 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1789;
  assign dataGroup_hi_hi_1789 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1790;
  assign dataGroup_hi_hi_1790 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1791;
  assign dataGroup_hi_hi_1791 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1792;
  assign dataGroup_hi_hi_1792 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1793;
  assign dataGroup_hi_hi_1793 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1794;
  assign dataGroup_hi_hi_1794 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1795;
  assign dataGroup_hi_hi_1795 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1796;
  assign dataGroup_hi_hi_1796 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1797;
  assign dataGroup_hi_hi_1797 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1798;
  assign dataGroup_hi_hi_1798 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1799;
  assign dataGroup_hi_hi_1799 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1800;
  assign dataGroup_hi_hi_1800 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1801;
  assign dataGroup_hi_hi_1801 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1802;
  assign dataGroup_hi_hi_1802 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1803;
  assign dataGroup_hi_hi_1803 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1804;
  assign dataGroup_hi_hi_1804 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1805;
  assign dataGroup_hi_hi_1805 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1806;
  assign dataGroup_hi_hi_1806 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1807;
  assign dataGroup_hi_hi_1807 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1808;
  assign dataGroup_hi_hi_1808 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1809;
  assign dataGroup_hi_hi_1809 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1810;
  assign dataGroup_hi_hi_1810 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1811;
  assign dataGroup_hi_hi_1811 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1812;
  assign dataGroup_hi_hi_1812 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1813;
  assign dataGroup_hi_hi_1813 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1814;
  assign dataGroup_hi_hi_1814 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1815;
  assign dataGroup_hi_hi_1815 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1816;
  assign dataGroup_hi_hi_1816 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1817;
  assign dataGroup_hi_hi_1817 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1818;
  assign dataGroup_hi_hi_1818 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1819;
  assign dataGroup_hi_hi_1819 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1820;
  assign dataGroup_hi_hi_1820 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1821;
  assign dataGroup_hi_hi_1821 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1822;
  assign dataGroup_hi_hi_1822 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1823;
  assign dataGroup_hi_hi_1823 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1824;
  assign dataGroup_hi_hi_1824 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1825;
  assign dataGroup_hi_hi_1825 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1826;
  assign dataGroup_hi_hi_1826 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1827;
  assign dataGroup_hi_hi_1827 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1828;
  assign dataGroup_hi_hi_1828 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1829;
  assign dataGroup_hi_hi_1829 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1830;
  assign dataGroup_hi_hi_1830 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1831;
  assign dataGroup_hi_hi_1831 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1832;
  assign dataGroup_hi_hi_1832 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1833;
  assign dataGroup_hi_hi_1833 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1834;
  assign dataGroup_hi_hi_1834 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1835;
  assign dataGroup_hi_hi_1835 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1836;
  assign dataGroup_hi_hi_1836 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1837;
  assign dataGroup_hi_hi_1837 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1838;
  assign dataGroup_hi_hi_1838 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1839;
  assign dataGroup_hi_hi_1839 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1840;
  assign dataGroup_hi_hi_1840 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1841;
  assign dataGroup_hi_hi_1841 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1842;
  assign dataGroup_hi_hi_1842 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1843;
  assign dataGroup_hi_hi_1843 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1844;
  assign dataGroup_hi_hi_1844 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1845;
  assign dataGroup_hi_hi_1845 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1846;
  assign dataGroup_hi_hi_1846 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1847;
  assign dataGroup_hi_hi_1847 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1848;
  assign dataGroup_hi_hi_1848 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1849;
  assign dataGroup_hi_hi_1849 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1850;
  assign dataGroup_hi_hi_1850 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1851;
  assign dataGroup_hi_hi_1851 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1852;
  assign dataGroup_hi_hi_1852 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1853;
  assign dataGroup_hi_hi_1853 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1854;
  assign dataGroup_hi_hi_1854 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1855;
  assign dataGroup_hi_hi_1855 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1856;
  assign dataGroup_hi_hi_1856 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1857;
  assign dataGroup_hi_hi_1857 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1858;
  assign dataGroup_hi_hi_1858 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1859;
  assign dataGroup_hi_hi_1859 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1860;
  assign dataGroup_hi_hi_1860 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1861;
  assign dataGroup_hi_hi_1861 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1862;
  assign dataGroup_hi_hi_1862 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1863;
  assign dataGroup_hi_hi_1863 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1864;
  assign dataGroup_hi_hi_1864 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1865;
  assign dataGroup_hi_hi_1865 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1866;
  assign dataGroup_hi_hi_1866 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1867;
  assign dataGroup_hi_hi_1867 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1868;
  assign dataGroup_hi_hi_1868 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1869;
  assign dataGroup_hi_hi_1869 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1870;
  assign dataGroup_hi_hi_1870 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1871;
  assign dataGroup_hi_hi_1871 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1872;
  assign dataGroup_hi_hi_1872 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1873;
  assign dataGroup_hi_hi_1873 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1874;
  assign dataGroup_hi_hi_1874 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1875;
  assign dataGroup_hi_hi_1875 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1876;
  assign dataGroup_hi_hi_1876 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1877;
  assign dataGroup_hi_hi_1877 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1878;
  assign dataGroup_hi_hi_1878 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1879;
  assign dataGroup_hi_hi_1879 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1880;
  assign dataGroup_hi_hi_1880 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1881;
  assign dataGroup_hi_hi_1881 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1882;
  assign dataGroup_hi_hi_1882 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1883;
  assign dataGroup_hi_hi_1883 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1884;
  assign dataGroup_hi_hi_1884 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1885;
  assign dataGroup_hi_hi_1885 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1886;
  assign dataGroup_hi_hi_1886 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1887;
  assign dataGroup_hi_hi_1887 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1888;
  assign dataGroup_hi_hi_1888 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1889;
  assign dataGroup_hi_hi_1889 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1890;
  assign dataGroup_hi_hi_1890 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1891;
  assign dataGroup_hi_hi_1891 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1892;
  assign dataGroup_hi_hi_1892 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1893;
  assign dataGroup_hi_hi_1893 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1894;
  assign dataGroup_hi_hi_1894 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1895;
  assign dataGroup_hi_hi_1895 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1896;
  assign dataGroup_hi_hi_1896 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1897;
  assign dataGroup_hi_hi_1897 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1898;
  assign dataGroup_hi_hi_1898 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1899;
  assign dataGroup_hi_hi_1899 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1900;
  assign dataGroup_hi_hi_1900 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1901;
  assign dataGroup_hi_hi_1901 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1902;
  assign dataGroup_hi_hi_1902 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1903;
  assign dataGroup_hi_hi_1903 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1904;
  assign dataGroup_hi_hi_1904 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1905;
  assign dataGroup_hi_hi_1905 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1906;
  assign dataGroup_hi_hi_1906 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1907;
  assign dataGroup_hi_hi_1907 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1908;
  assign dataGroup_hi_hi_1908 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1909;
  assign dataGroup_hi_hi_1909 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1910;
  assign dataGroup_hi_hi_1910 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1911;
  assign dataGroup_hi_hi_1911 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1912;
  assign dataGroup_hi_hi_1912 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1913;
  assign dataGroup_hi_hi_1913 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1914;
  assign dataGroup_hi_hi_1914 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1915;
  assign dataGroup_hi_hi_1915 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1916;
  assign dataGroup_hi_hi_1916 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1917;
  assign dataGroup_hi_hi_1917 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1918;
  assign dataGroup_hi_hi_1918 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1919;
  assign dataGroup_hi_hi_1919 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1920;
  assign dataGroup_hi_hi_1920 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1921;
  assign dataGroup_hi_hi_1921 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1922;
  assign dataGroup_hi_hi_1922 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1923;
  assign dataGroup_hi_hi_1923 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1924;
  assign dataGroup_hi_hi_1924 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1925;
  assign dataGroup_hi_hi_1925 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1926;
  assign dataGroup_hi_hi_1926 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1927;
  assign dataGroup_hi_hi_1927 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1928;
  assign dataGroup_hi_hi_1928 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1929;
  assign dataGroup_hi_hi_1929 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1930;
  assign dataGroup_hi_hi_1930 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1931;
  assign dataGroup_hi_hi_1931 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1932;
  assign dataGroup_hi_hi_1932 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1933;
  assign dataGroup_hi_hi_1933 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1934;
  assign dataGroup_hi_hi_1934 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1935;
  assign dataGroup_hi_hi_1935 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1936;
  assign dataGroup_hi_hi_1936 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1937;
  assign dataGroup_hi_hi_1937 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1938;
  assign dataGroup_hi_hi_1938 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1939;
  assign dataGroup_hi_hi_1939 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1940;
  assign dataGroup_hi_hi_1940 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1941;
  assign dataGroup_hi_hi_1941 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1942;
  assign dataGroup_hi_hi_1942 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1943;
  assign dataGroup_hi_hi_1943 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1944;
  assign dataGroup_hi_hi_1944 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1945;
  assign dataGroup_hi_hi_1945 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1946;
  assign dataGroup_hi_hi_1946 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1947;
  assign dataGroup_hi_hi_1947 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1948;
  assign dataGroup_hi_hi_1948 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1949;
  assign dataGroup_hi_hi_1949 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1950;
  assign dataGroup_hi_hi_1950 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1951;
  assign dataGroup_hi_hi_1951 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1952;
  assign dataGroup_hi_hi_1952 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1953;
  assign dataGroup_hi_hi_1953 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1954;
  assign dataGroup_hi_hi_1954 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1955;
  assign dataGroup_hi_hi_1955 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1956;
  assign dataGroup_hi_hi_1956 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1957;
  assign dataGroup_hi_hi_1957 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1958;
  assign dataGroup_hi_hi_1958 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1959;
  assign dataGroup_hi_hi_1959 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1960;
  assign dataGroup_hi_hi_1960 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1961;
  assign dataGroup_hi_hi_1961 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1962;
  assign dataGroup_hi_hi_1962 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1963;
  assign dataGroup_hi_hi_1963 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1964;
  assign dataGroup_hi_hi_1964 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1965;
  assign dataGroup_hi_hi_1965 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1966;
  assign dataGroup_hi_hi_1966 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1967;
  assign dataGroup_hi_hi_1967 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1968;
  assign dataGroup_hi_hi_1968 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1969;
  assign dataGroup_hi_hi_1969 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1970;
  assign dataGroup_hi_hi_1970 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1971;
  assign dataGroup_hi_hi_1971 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1972;
  assign dataGroup_hi_hi_1972 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1973;
  assign dataGroup_hi_hi_1973 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1974;
  assign dataGroup_hi_hi_1974 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1975;
  assign dataGroup_hi_hi_1975 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1976;
  assign dataGroup_hi_hi_1976 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1977;
  assign dataGroup_hi_hi_1977 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1978;
  assign dataGroup_hi_hi_1978 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1979;
  assign dataGroup_hi_hi_1979 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1980;
  assign dataGroup_hi_hi_1980 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1981;
  assign dataGroup_hi_hi_1981 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1982;
  assign dataGroup_hi_hi_1982 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1983;
  assign dataGroup_hi_hi_1983 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1984;
  assign dataGroup_hi_hi_1984 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1985;
  assign dataGroup_hi_hi_1985 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1986;
  assign dataGroup_hi_hi_1986 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1987;
  assign dataGroup_hi_hi_1987 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1988;
  assign dataGroup_hi_hi_1988 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1989;
  assign dataGroup_hi_hi_1989 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1990;
  assign dataGroup_hi_hi_1990 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1991;
  assign dataGroup_hi_hi_1991 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1992;
  assign dataGroup_hi_hi_1992 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1993;
  assign dataGroup_hi_hi_1993 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1994;
  assign dataGroup_hi_hi_1994 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1995;
  assign dataGroup_hi_hi_1995 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1996;
  assign dataGroup_hi_hi_1996 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1997;
  assign dataGroup_hi_hi_1997 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1998;
  assign dataGroup_hi_hi_1998 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_1999;
  assign dataGroup_hi_hi_1999 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2000;
  assign dataGroup_hi_hi_2000 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2001;
  assign dataGroup_hi_hi_2001 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2002;
  assign dataGroup_hi_hi_2002 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2003;
  assign dataGroup_hi_hi_2003 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2004;
  assign dataGroup_hi_hi_2004 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2005;
  assign dataGroup_hi_hi_2005 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2006;
  assign dataGroup_hi_hi_2006 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2007;
  assign dataGroup_hi_hi_2007 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2008;
  assign dataGroup_hi_hi_2008 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2009;
  assign dataGroup_hi_hi_2009 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2010;
  assign dataGroup_hi_hi_2010 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2011;
  assign dataGroup_hi_hi_2011 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2012;
  assign dataGroup_hi_hi_2012 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2013;
  assign dataGroup_hi_hi_2013 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2014;
  assign dataGroup_hi_hi_2014 = _GEN_7;
  wire [511:0]  dataGroup_hi_hi_2015;
  assign dataGroup_hi_hi_2015 = _GEN_7;
  wire [1023:0] dataGroup_hi = {dataGroup_hi_hi, dataGroup_hi_lo};
  wire [7:0]    dataGroup_0 = dataGroup_lo[7:0];
  wire [1023:0] dataGroup_lo_1 = {dataGroup_lo_hi_1, dataGroup_lo_lo_1};
  wire [1023:0] dataGroup_hi_1 = {dataGroup_hi_hi_1, dataGroup_hi_lo_1};
  wire [7:0]    dataGroup_1 = dataGroup_lo_1[15:8];
  wire [1023:0] dataGroup_lo_2 = {dataGroup_lo_hi_2, dataGroup_lo_lo_2};
  wire [1023:0] dataGroup_hi_2 = {dataGroup_hi_hi_2, dataGroup_hi_lo_2};
  wire [7:0]    dataGroup_2 = dataGroup_lo_2[23:16];
  wire [1023:0] dataGroup_lo_3 = {dataGroup_lo_hi_3, dataGroup_lo_lo_3};
  wire [1023:0] dataGroup_hi_3 = {dataGroup_hi_hi_3, dataGroup_hi_lo_3};
  wire [7:0]    dataGroup_3 = dataGroup_lo_3[31:24];
  wire [1023:0] dataGroup_lo_4 = {dataGroup_lo_hi_4, dataGroup_lo_lo_4};
  wire [1023:0] dataGroup_hi_4 = {dataGroup_hi_hi_4, dataGroup_hi_lo_4};
  wire [7:0]    dataGroup_4 = dataGroup_lo_4[39:32];
  wire [1023:0] dataGroup_lo_5 = {dataGroup_lo_hi_5, dataGroup_lo_lo_5};
  wire [1023:0] dataGroup_hi_5 = {dataGroup_hi_hi_5, dataGroup_hi_lo_5};
  wire [7:0]    dataGroup_5 = dataGroup_lo_5[47:40];
  wire [1023:0] dataGroup_lo_6 = {dataGroup_lo_hi_6, dataGroup_lo_lo_6};
  wire [1023:0] dataGroup_hi_6 = {dataGroup_hi_hi_6, dataGroup_hi_lo_6};
  wire [7:0]    dataGroup_6 = dataGroup_lo_6[55:48];
  wire [1023:0] dataGroup_lo_7 = {dataGroup_lo_hi_7, dataGroup_lo_lo_7};
  wire [1023:0] dataGroup_hi_7 = {dataGroup_hi_hi_7, dataGroup_hi_lo_7};
  wire [7:0]    dataGroup_7 = dataGroup_lo_7[63:56];
  wire [1023:0] dataGroup_lo_8 = {dataGroup_lo_hi_8, dataGroup_lo_lo_8};
  wire [1023:0] dataGroup_hi_8 = {dataGroup_hi_hi_8, dataGroup_hi_lo_8};
  wire [7:0]    dataGroup_8 = dataGroup_lo_8[71:64];
  wire [1023:0] dataGroup_lo_9 = {dataGroup_lo_hi_9, dataGroup_lo_lo_9};
  wire [1023:0] dataGroup_hi_9 = {dataGroup_hi_hi_9, dataGroup_hi_lo_9};
  wire [7:0]    dataGroup_9 = dataGroup_lo_9[79:72];
  wire [1023:0] dataGroup_lo_10 = {dataGroup_lo_hi_10, dataGroup_lo_lo_10};
  wire [1023:0] dataGroup_hi_10 = {dataGroup_hi_hi_10, dataGroup_hi_lo_10};
  wire [7:0]    dataGroup_10 = dataGroup_lo_10[87:80];
  wire [1023:0] dataGroup_lo_11 = {dataGroup_lo_hi_11, dataGroup_lo_lo_11};
  wire [1023:0] dataGroup_hi_11 = {dataGroup_hi_hi_11, dataGroup_hi_lo_11};
  wire [7:0]    dataGroup_11 = dataGroup_lo_11[95:88];
  wire [1023:0] dataGroup_lo_12 = {dataGroup_lo_hi_12, dataGroup_lo_lo_12};
  wire [1023:0] dataGroup_hi_12 = {dataGroup_hi_hi_12, dataGroup_hi_lo_12};
  wire [7:0]    dataGroup_12 = dataGroup_lo_12[103:96];
  wire [1023:0] dataGroup_lo_13 = {dataGroup_lo_hi_13, dataGroup_lo_lo_13};
  wire [1023:0] dataGroup_hi_13 = {dataGroup_hi_hi_13, dataGroup_hi_lo_13};
  wire [7:0]    dataGroup_13 = dataGroup_lo_13[111:104];
  wire [1023:0] dataGroup_lo_14 = {dataGroup_lo_hi_14, dataGroup_lo_lo_14};
  wire [1023:0] dataGroup_hi_14 = {dataGroup_hi_hi_14, dataGroup_hi_lo_14};
  wire [7:0]    dataGroup_14 = dataGroup_lo_14[119:112];
  wire [1023:0] dataGroup_lo_15 = {dataGroup_lo_hi_15, dataGroup_lo_lo_15};
  wire [1023:0] dataGroup_hi_15 = {dataGroup_hi_hi_15, dataGroup_hi_lo_15};
  wire [7:0]    dataGroup_15 = dataGroup_lo_15[127:120];
  wire [1023:0] dataGroup_lo_16 = {dataGroup_lo_hi_16, dataGroup_lo_lo_16};
  wire [1023:0] dataGroup_hi_16 = {dataGroup_hi_hi_16, dataGroup_hi_lo_16};
  wire [7:0]    dataGroup_16 = dataGroup_lo_16[135:128];
  wire [1023:0] dataGroup_lo_17 = {dataGroup_lo_hi_17, dataGroup_lo_lo_17};
  wire [1023:0] dataGroup_hi_17 = {dataGroup_hi_hi_17, dataGroup_hi_lo_17};
  wire [7:0]    dataGroup_17 = dataGroup_lo_17[143:136];
  wire [1023:0] dataGroup_lo_18 = {dataGroup_lo_hi_18, dataGroup_lo_lo_18};
  wire [1023:0] dataGroup_hi_18 = {dataGroup_hi_hi_18, dataGroup_hi_lo_18};
  wire [7:0]    dataGroup_18 = dataGroup_lo_18[151:144];
  wire [1023:0] dataGroup_lo_19 = {dataGroup_lo_hi_19, dataGroup_lo_lo_19};
  wire [1023:0] dataGroup_hi_19 = {dataGroup_hi_hi_19, dataGroup_hi_lo_19};
  wire [7:0]    dataGroup_19 = dataGroup_lo_19[159:152];
  wire [1023:0] dataGroup_lo_20 = {dataGroup_lo_hi_20, dataGroup_lo_lo_20};
  wire [1023:0] dataGroup_hi_20 = {dataGroup_hi_hi_20, dataGroup_hi_lo_20};
  wire [7:0]    dataGroup_20 = dataGroup_lo_20[167:160];
  wire [1023:0] dataGroup_lo_21 = {dataGroup_lo_hi_21, dataGroup_lo_lo_21};
  wire [1023:0] dataGroup_hi_21 = {dataGroup_hi_hi_21, dataGroup_hi_lo_21};
  wire [7:0]    dataGroup_21 = dataGroup_lo_21[175:168];
  wire [1023:0] dataGroup_lo_22 = {dataGroup_lo_hi_22, dataGroup_lo_lo_22};
  wire [1023:0] dataGroup_hi_22 = {dataGroup_hi_hi_22, dataGroup_hi_lo_22};
  wire [7:0]    dataGroup_22 = dataGroup_lo_22[183:176];
  wire [1023:0] dataGroup_lo_23 = {dataGroup_lo_hi_23, dataGroup_lo_lo_23};
  wire [1023:0] dataGroup_hi_23 = {dataGroup_hi_hi_23, dataGroup_hi_lo_23};
  wire [7:0]    dataGroup_23 = dataGroup_lo_23[191:184];
  wire [1023:0] dataGroup_lo_24 = {dataGroup_lo_hi_24, dataGroup_lo_lo_24};
  wire [1023:0] dataGroup_hi_24 = {dataGroup_hi_hi_24, dataGroup_hi_lo_24};
  wire [7:0]    dataGroup_24 = dataGroup_lo_24[199:192];
  wire [1023:0] dataGroup_lo_25 = {dataGroup_lo_hi_25, dataGroup_lo_lo_25};
  wire [1023:0] dataGroup_hi_25 = {dataGroup_hi_hi_25, dataGroup_hi_lo_25};
  wire [7:0]    dataGroup_25 = dataGroup_lo_25[207:200];
  wire [1023:0] dataGroup_lo_26 = {dataGroup_lo_hi_26, dataGroup_lo_lo_26};
  wire [1023:0] dataGroup_hi_26 = {dataGroup_hi_hi_26, dataGroup_hi_lo_26};
  wire [7:0]    dataGroup_26 = dataGroup_lo_26[215:208];
  wire [1023:0] dataGroup_lo_27 = {dataGroup_lo_hi_27, dataGroup_lo_lo_27};
  wire [1023:0] dataGroup_hi_27 = {dataGroup_hi_hi_27, dataGroup_hi_lo_27};
  wire [7:0]    dataGroup_27 = dataGroup_lo_27[223:216];
  wire [1023:0] dataGroup_lo_28 = {dataGroup_lo_hi_28, dataGroup_lo_lo_28};
  wire [1023:0] dataGroup_hi_28 = {dataGroup_hi_hi_28, dataGroup_hi_lo_28};
  wire [7:0]    dataGroup_28 = dataGroup_lo_28[231:224];
  wire [1023:0] dataGroup_lo_29 = {dataGroup_lo_hi_29, dataGroup_lo_lo_29};
  wire [1023:0] dataGroup_hi_29 = {dataGroup_hi_hi_29, dataGroup_hi_lo_29};
  wire [7:0]    dataGroup_29 = dataGroup_lo_29[239:232];
  wire [1023:0] dataGroup_lo_30 = {dataGroup_lo_hi_30, dataGroup_lo_lo_30};
  wire [1023:0] dataGroup_hi_30 = {dataGroup_hi_hi_30, dataGroup_hi_lo_30};
  wire [7:0]    dataGroup_30 = dataGroup_lo_30[247:240];
  wire [1023:0] dataGroup_lo_31 = {dataGroup_lo_hi_31, dataGroup_lo_lo_31};
  wire [1023:0] dataGroup_hi_31 = {dataGroup_hi_hi_31, dataGroup_hi_lo_31};
  wire [7:0]    dataGroup_31 = dataGroup_lo_31[255:248];
  wire [15:0]   res_lo_lo_lo_lo = {dataGroup_1, dataGroup_0};
  wire [15:0]   res_lo_lo_lo_hi = {dataGroup_3, dataGroup_2};
  wire [31:0]   res_lo_lo_lo = {res_lo_lo_lo_hi, res_lo_lo_lo_lo};
  wire [15:0]   res_lo_lo_hi_lo = {dataGroup_5, dataGroup_4};
  wire [15:0]   res_lo_lo_hi_hi = {dataGroup_7, dataGroup_6};
  wire [31:0]   res_lo_lo_hi = {res_lo_lo_hi_hi, res_lo_lo_hi_lo};
  wire [63:0]   res_lo_lo = {res_lo_lo_hi, res_lo_lo_lo};
  wire [15:0]   res_lo_hi_lo_lo = {dataGroup_9, dataGroup_8};
  wire [15:0]   res_lo_hi_lo_hi = {dataGroup_11, dataGroup_10};
  wire [31:0]   res_lo_hi_lo = {res_lo_hi_lo_hi, res_lo_hi_lo_lo};
  wire [15:0]   res_lo_hi_hi_lo = {dataGroup_13, dataGroup_12};
  wire [15:0]   res_lo_hi_hi_hi = {dataGroup_15, dataGroup_14};
  wire [31:0]   res_lo_hi_hi = {res_lo_hi_hi_hi, res_lo_hi_hi_lo};
  wire [63:0]   res_lo_hi = {res_lo_hi_hi, res_lo_hi_lo};
  wire [127:0]  res_lo = {res_lo_hi, res_lo_lo};
  wire [15:0]   res_hi_lo_lo_lo = {dataGroup_17, dataGroup_16};
  wire [15:0]   res_hi_lo_lo_hi = {dataGroup_19, dataGroup_18};
  wire [31:0]   res_hi_lo_lo = {res_hi_lo_lo_hi, res_hi_lo_lo_lo};
  wire [15:0]   res_hi_lo_hi_lo = {dataGroup_21, dataGroup_20};
  wire [15:0]   res_hi_lo_hi_hi = {dataGroup_23, dataGroup_22};
  wire [31:0]   res_hi_lo_hi = {res_hi_lo_hi_hi, res_hi_lo_hi_lo};
  wire [63:0]   res_hi_lo = {res_hi_lo_hi, res_hi_lo_lo};
  wire [15:0]   res_hi_hi_lo_lo = {dataGroup_25, dataGroup_24};
  wire [15:0]   res_hi_hi_lo_hi = {dataGroup_27, dataGroup_26};
  wire [31:0]   res_hi_hi_lo = {res_hi_hi_lo_hi, res_hi_hi_lo_lo};
  wire [15:0]   res_hi_hi_hi_lo = {dataGroup_29, dataGroup_28};
  wire [15:0]   res_hi_hi_hi_hi = {dataGroup_31, dataGroup_30};
  wire [31:0]   res_hi_hi_hi = {res_hi_hi_hi_hi, res_hi_hi_hi_lo};
  wire [63:0]   res_hi_hi = {res_hi_hi_hi, res_hi_hi_lo};
  wire [127:0]  res_hi = {res_hi_hi, res_hi_lo};
  wire [255:0]  res = {res_hi, res_lo};
  wire [511:0]  lo_lo = {256'h0, res};
  wire [1023:0] lo = {512'h0, lo_lo};
  wire [2047:0] regroupLoadData_0_0 = {1024'h0, lo};
  wire [1023:0] dataGroup_lo_32 = {dataGroup_lo_hi_32, dataGroup_lo_lo_32};
  wire [1023:0] dataGroup_hi_32 = {dataGroup_hi_hi_32, dataGroup_hi_lo_32};
  wire [7:0]    dataGroup_0_1 = dataGroup_lo_32[7:0];
  wire [1023:0] dataGroup_lo_33 = {dataGroup_lo_hi_33, dataGroup_lo_lo_33};
  wire [1023:0] dataGroup_hi_33 = {dataGroup_hi_hi_33, dataGroup_hi_lo_33};
  wire [7:0]    dataGroup_1_1 = dataGroup_lo_33[23:16];
  wire [1023:0] dataGroup_lo_34 = {dataGroup_lo_hi_34, dataGroup_lo_lo_34};
  wire [1023:0] dataGroup_hi_34 = {dataGroup_hi_hi_34, dataGroup_hi_lo_34};
  wire [7:0]    dataGroup_2_1 = dataGroup_lo_34[39:32];
  wire [1023:0] dataGroup_lo_35 = {dataGroup_lo_hi_35, dataGroup_lo_lo_35};
  wire [1023:0] dataGroup_hi_35 = {dataGroup_hi_hi_35, dataGroup_hi_lo_35};
  wire [7:0]    dataGroup_3_1 = dataGroup_lo_35[55:48];
  wire [1023:0] dataGroup_lo_36 = {dataGroup_lo_hi_36, dataGroup_lo_lo_36};
  wire [1023:0] dataGroup_hi_36 = {dataGroup_hi_hi_36, dataGroup_hi_lo_36};
  wire [7:0]    dataGroup_4_1 = dataGroup_lo_36[71:64];
  wire [1023:0] dataGroup_lo_37 = {dataGroup_lo_hi_37, dataGroup_lo_lo_37};
  wire [1023:0] dataGroup_hi_37 = {dataGroup_hi_hi_37, dataGroup_hi_lo_37};
  wire [7:0]    dataGroup_5_1 = dataGroup_lo_37[87:80];
  wire [1023:0] dataGroup_lo_38 = {dataGroup_lo_hi_38, dataGroup_lo_lo_38};
  wire [1023:0] dataGroup_hi_38 = {dataGroup_hi_hi_38, dataGroup_hi_lo_38};
  wire [7:0]    dataGroup_6_1 = dataGroup_lo_38[103:96];
  wire [1023:0] dataGroup_lo_39 = {dataGroup_lo_hi_39, dataGroup_lo_lo_39};
  wire [1023:0] dataGroup_hi_39 = {dataGroup_hi_hi_39, dataGroup_hi_lo_39};
  wire [7:0]    dataGroup_7_1 = dataGroup_lo_39[119:112];
  wire [1023:0] dataGroup_lo_40 = {dataGroup_lo_hi_40, dataGroup_lo_lo_40};
  wire [1023:0] dataGroup_hi_40 = {dataGroup_hi_hi_40, dataGroup_hi_lo_40};
  wire [7:0]    dataGroup_8_1 = dataGroup_lo_40[135:128];
  wire [1023:0] dataGroup_lo_41 = {dataGroup_lo_hi_41, dataGroup_lo_lo_41};
  wire [1023:0] dataGroup_hi_41 = {dataGroup_hi_hi_41, dataGroup_hi_lo_41};
  wire [7:0]    dataGroup_9_1 = dataGroup_lo_41[151:144];
  wire [1023:0] dataGroup_lo_42 = {dataGroup_lo_hi_42, dataGroup_lo_lo_42};
  wire [1023:0] dataGroup_hi_42 = {dataGroup_hi_hi_42, dataGroup_hi_lo_42};
  wire [7:0]    dataGroup_10_1 = dataGroup_lo_42[167:160];
  wire [1023:0] dataGroup_lo_43 = {dataGroup_lo_hi_43, dataGroup_lo_lo_43};
  wire [1023:0] dataGroup_hi_43 = {dataGroup_hi_hi_43, dataGroup_hi_lo_43};
  wire [7:0]    dataGroup_11_1 = dataGroup_lo_43[183:176];
  wire [1023:0] dataGroup_lo_44 = {dataGroup_lo_hi_44, dataGroup_lo_lo_44};
  wire [1023:0] dataGroup_hi_44 = {dataGroup_hi_hi_44, dataGroup_hi_lo_44};
  wire [7:0]    dataGroup_12_1 = dataGroup_lo_44[199:192];
  wire [1023:0] dataGroup_lo_45 = {dataGroup_lo_hi_45, dataGroup_lo_lo_45};
  wire [1023:0] dataGroup_hi_45 = {dataGroup_hi_hi_45, dataGroup_hi_lo_45};
  wire [7:0]    dataGroup_13_1 = dataGroup_lo_45[215:208];
  wire [1023:0] dataGroup_lo_46 = {dataGroup_lo_hi_46, dataGroup_lo_lo_46};
  wire [1023:0] dataGroup_hi_46 = {dataGroup_hi_hi_46, dataGroup_hi_lo_46};
  wire [7:0]    dataGroup_14_1 = dataGroup_lo_46[231:224];
  wire [1023:0] dataGroup_lo_47 = {dataGroup_lo_hi_47, dataGroup_lo_lo_47};
  wire [1023:0] dataGroup_hi_47 = {dataGroup_hi_hi_47, dataGroup_hi_lo_47};
  wire [7:0]    dataGroup_15_1 = dataGroup_lo_47[247:240];
  wire [1023:0] dataGroup_lo_48 = {dataGroup_lo_hi_48, dataGroup_lo_lo_48};
  wire [1023:0] dataGroup_hi_48 = {dataGroup_hi_hi_48, dataGroup_hi_lo_48};
  wire [7:0]    dataGroup_16_1 = dataGroup_lo_48[263:256];
  wire [1023:0] dataGroup_lo_49 = {dataGroup_lo_hi_49, dataGroup_lo_lo_49};
  wire [1023:0] dataGroup_hi_49 = {dataGroup_hi_hi_49, dataGroup_hi_lo_49};
  wire [7:0]    dataGroup_17_1 = dataGroup_lo_49[279:272];
  wire [1023:0] dataGroup_lo_50 = {dataGroup_lo_hi_50, dataGroup_lo_lo_50};
  wire [1023:0] dataGroup_hi_50 = {dataGroup_hi_hi_50, dataGroup_hi_lo_50};
  wire [7:0]    dataGroup_18_1 = dataGroup_lo_50[295:288];
  wire [1023:0] dataGroup_lo_51 = {dataGroup_lo_hi_51, dataGroup_lo_lo_51};
  wire [1023:0] dataGroup_hi_51 = {dataGroup_hi_hi_51, dataGroup_hi_lo_51};
  wire [7:0]    dataGroup_19_1 = dataGroup_lo_51[311:304];
  wire [1023:0] dataGroup_lo_52 = {dataGroup_lo_hi_52, dataGroup_lo_lo_52};
  wire [1023:0] dataGroup_hi_52 = {dataGroup_hi_hi_52, dataGroup_hi_lo_52};
  wire [7:0]    dataGroup_20_1 = dataGroup_lo_52[327:320];
  wire [1023:0] dataGroup_lo_53 = {dataGroup_lo_hi_53, dataGroup_lo_lo_53};
  wire [1023:0] dataGroup_hi_53 = {dataGroup_hi_hi_53, dataGroup_hi_lo_53};
  wire [7:0]    dataGroup_21_1 = dataGroup_lo_53[343:336];
  wire [1023:0] dataGroup_lo_54 = {dataGroup_lo_hi_54, dataGroup_lo_lo_54};
  wire [1023:0] dataGroup_hi_54 = {dataGroup_hi_hi_54, dataGroup_hi_lo_54};
  wire [7:0]    dataGroup_22_1 = dataGroup_lo_54[359:352];
  wire [1023:0] dataGroup_lo_55 = {dataGroup_lo_hi_55, dataGroup_lo_lo_55};
  wire [1023:0] dataGroup_hi_55 = {dataGroup_hi_hi_55, dataGroup_hi_lo_55};
  wire [7:0]    dataGroup_23_1 = dataGroup_lo_55[375:368];
  wire [1023:0] dataGroup_lo_56 = {dataGroup_lo_hi_56, dataGroup_lo_lo_56};
  wire [1023:0] dataGroup_hi_56 = {dataGroup_hi_hi_56, dataGroup_hi_lo_56};
  wire [7:0]    dataGroup_24_1 = dataGroup_lo_56[391:384];
  wire [1023:0] dataGroup_lo_57 = {dataGroup_lo_hi_57, dataGroup_lo_lo_57};
  wire [1023:0] dataGroup_hi_57 = {dataGroup_hi_hi_57, dataGroup_hi_lo_57};
  wire [7:0]    dataGroup_25_1 = dataGroup_lo_57[407:400];
  wire [1023:0] dataGroup_lo_58 = {dataGroup_lo_hi_58, dataGroup_lo_lo_58};
  wire [1023:0] dataGroup_hi_58 = {dataGroup_hi_hi_58, dataGroup_hi_lo_58};
  wire [7:0]    dataGroup_26_1 = dataGroup_lo_58[423:416];
  wire [1023:0] dataGroup_lo_59 = {dataGroup_lo_hi_59, dataGroup_lo_lo_59};
  wire [1023:0] dataGroup_hi_59 = {dataGroup_hi_hi_59, dataGroup_hi_lo_59};
  wire [7:0]    dataGroup_27_1 = dataGroup_lo_59[439:432];
  wire [1023:0] dataGroup_lo_60 = {dataGroup_lo_hi_60, dataGroup_lo_lo_60};
  wire [1023:0] dataGroup_hi_60 = {dataGroup_hi_hi_60, dataGroup_hi_lo_60};
  wire [7:0]    dataGroup_28_1 = dataGroup_lo_60[455:448];
  wire [1023:0] dataGroup_lo_61 = {dataGroup_lo_hi_61, dataGroup_lo_lo_61};
  wire [1023:0] dataGroup_hi_61 = {dataGroup_hi_hi_61, dataGroup_hi_lo_61};
  wire [7:0]    dataGroup_29_1 = dataGroup_lo_61[471:464];
  wire [1023:0] dataGroup_lo_62 = {dataGroup_lo_hi_62, dataGroup_lo_lo_62};
  wire [1023:0] dataGroup_hi_62 = {dataGroup_hi_hi_62, dataGroup_hi_lo_62};
  wire [7:0]    dataGroup_30_1 = dataGroup_lo_62[487:480];
  wire [1023:0] dataGroup_lo_63 = {dataGroup_lo_hi_63, dataGroup_lo_lo_63};
  wire [1023:0] dataGroup_hi_63 = {dataGroup_hi_hi_63, dataGroup_hi_lo_63};
  wire [7:0]    dataGroup_31_1 = dataGroup_lo_63[503:496];
  wire [15:0]   res_lo_lo_lo_lo_1 = {dataGroup_1_1, dataGroup_0_1};
  wire [15:0]   res_lo_lo_lo_hi_1 = {dataGroup_3_1, dataGroup_2_1};
  wire [31:0]   res_lo_lo_lo_1 = {res_lo_lo_lo_hi_1, res_lo_lo_lo_lo_1};
  wire [15:0]   res_lo_lo_hi_lo_1 = {dataGroup_5_1, dataGroup_4_1};
  wire [15:0]   res_lo_lo_hi_hi_1 = {dataGroup_7_1, dataGroup_6_1};
  wire [31:0]   res_lo_lo_hi_1 = {res_lo_lo_hi_hi_1, res_lo_lo_hi_lo_1};
  wire [63:0]   res_lo_lo_1 = {res_lo_lo_hi_1, res_lo_lo_lo_1};
  wire [15:0]   res_lo_hi_lo_lo_1 = {dataGroup_9_1, dataGroup_8_1};
  wire [15:0]   res_lo_hi_lo_hi_1 = {dataGroup_11_1, dataGroup_10_1};
  wire [31:0]   res_lo_hi_lo_1 = {res_lo_hi_lo_hi_1, res_lo_hi_lo_lo_1};
  wire [15:0]   res_lo_hi_hi_lo_1 = {dataGroup_13_1, dataGroup_12_1};
  wire [15:0]   res_lo_hi_hi_hi_1 = {dataGroup_15_1, dataGroup_14_1};
  wire [31:0]   res_lo_hi_hi_1 = {res_lo_hi_hi_hi_1, res_lo_hi_hi_lo_1};
  wire [63:0]   res_lo_hi_1 = {res_lo_hi_hi_1, res_lo_hi_lo_1};
  wire [127:0]  res_lo_1 = {res_lo_hi_1, res_lo_lo_1};
  wire [15:0]   res_hi_lo_lo_lo_1 = {dataGroup_17_1, dataGroup_16_1};
  wire [15:0]   res_hi_lo_lo_hi_1 = {dataGroup_19_1, dataGroup_18_1};
  wire [31:0]   res_hi_lo_lo_1 = {res_hi_lo_lo_hi_1, res_hi_lo_lo_lo_1};
  wire [15:0]   res_hi_lo_hi_lo_1 = {dataGroup_21_1, dataGroup_20_1};
  wire [15:0]   res_hi_lo_hi_hi_1 = {dataGroup_23_1, dataGroup_22_1};
  wire [31:0]   res_hi_lo_hi_1 = {res_hi_lo_hi_hi_1, res_hi_lo_hi_lo_1};
  wire [63:0]   res_hi_lo_1 = {res_hi_lo_hi_1, res_hi_lo_lo_1};
  wire [15:0]   res_hi_hi_lo_lo_1 = {dataGroup_25_1, dataGroup_24_1};
  wire [15:0]   res_hi_hi_lo_hi_1 = {dataGroup_27_1, dataGroup_26_1};
  wire [31:0]   res_hi_hi_lo_1 = {res_hi_hi_lo_hi_1, res_hi_hi_lo_lo_1};
  wire [15:0]   res_hi_hi_hi_lo_1 = {dataGroup_29_1, dataGroup_28_1};
  wire [15:0]   res_hi_hi_hi_hi_1 = {dataGroup_31_1, dataGroup_30_1};
  wire [31:0]   res_hi_hi_hi_1 = {res_hi_hi_hi_hi_1, res_hi_hi_hi_lo_1};
  wire [63:0]   res_hi_hi_1 = {res_hi_hi_hi_1, res_hi_hi_lo_1};
  wire [127:0]  res_hi_1 = {res_hi_hi_1, res_hi_lo_1};
  wire [255:0]  res_8 = {res_hi_1, res_lo_1};
  wire [1023:0] dataGroup_lo_64 = {dataGroup_lo_hi_64, dataGroup_lo_lo_64};
  wire [1023:0] dataGroup_hi_64 = {dataGroup_hi_hi_64, dataGroup_hi_lo_64};
  wire [7:0]    dataGroup_0_2 = dataGroup_lo_64[15:8];
  wire [1023:0] dataGroup_lo_65 = {dataGroup_lo_hi_65, dataGroup_lo_lo_65};
  wire [1023:0] dataGroup_hi_65 = {dataGroup_hi_hi_65, dataGroup_hi_lo_65};
  wire [7:0]    dataGroup_1_2 = dataGroup_lo_65[31:24];
  wire [1023:0] dataGroup_lo_66 = {dataGroup_lo_hi_66, dataGroup_lo_lo_66};
  wire [1023:0] dataGroup_hi_66 = {dataGroup_hi_hi_66, dataGroup_hi_lo_66};
  wire [7:0]    dataGroup_2_2 = dataGroup_lo_66[47:40];
  wire [1023:0] dataGroup_lo_67 = {dataGroup_lo_hi_67, dataGroup_lo_lo_67};
  wire [1023:0] dataGroup_hi_67 = {dataGroup_hi_hi_67, dataGroup_hi_lo_67};
  wire [7:0]    dataGroup_3_2 = dataGroup_lo_67[63:56];
  wire [1023:0] dataGroup_lo_68 = {dataGroup_lo_hi_68, dataGroup_lo_lo_68};
  wire [1023:0] dataGroup_hi_68 = {dataGroup_hi_hi_68, dataGroup_hi_lo_68};
  wire [7:0]    dataGroup_4_2 = dataGroup_lo_68[79:72];
  wire [1023:0] dataGroup_lo_69 = {dataGroup_lo_hi_69, dataGroup_lo_lo_69};
  wire [1023:0] dataGroup_hi_69 = {dataGroup_hi_hi_69, dataGroup_hi_lo_69};
  wire [7:0]    dataGroup_5_2 = dataGroup_lo_69[95:88];
  wire [1023:0] dataGroup_lo_70 = {dataGroup_lo_hi_70, dataGroup_lo_lo_70};
  wire [1023:0] dataGroup_hi_70 = {dataGroup_hi_hi_70, dataGroup_hi_lo_70};
  wire [7:0]    dataGroup_6_2 = dataGroup_lo_70[111:104];
  wire [1023:0] dataGroup_lo_71 = {dataGroup_lo_hi_71, dataGroup_lo_lo_71};
  wire [1023:0] dataGroup_hi_71 = {dataGroup_hi_hi_71, dataGroup_hi_lo_71};
  wire [7:0]    dataGroup_7_2 = dataGroup_lo_71[127:120];
  wire [1023:0] dataGroup_lo_72 = {dataGroup_lo_hi_72, dataGroup_lo_lo_72};
  wire [1023:0] dataGroup_hi_72 = {dataGroup_hi_hi_72, dataGroup_hi_lo_72};
  wire [7:0]    dataGroup_8_2 = dataGroup_lo_72[143:136];
  wire [1023:0] dataGroup_lo_73 = {dataGroup_lo_hi_73, dataGroup_lo_lo_73};
  wire [1023:0] dataGroup_hi_73 = {dataGroup_hi_hi_73, dataGroup_hi_lo_73};
  wire [7:0]    dataGroup_9_2 = dataGroup_lo_73[159:152];
  wire [1023:0] dataGroup_lo_74 = {dataGroup_lo_hi_74, dataGroup_lo_lo_74};
  wire [1023:0] dataGroup_hi_74 = {dataGroup_hi_hi_74, dataGroup_hi_lo_74};
  wire [7:0]    dataGroup_10_2 = dataGroup_lo_74[175:168];
  wire [1023:0] dataGroup_lo_75 = {dataGroup_lo_hi_75, dataGroup_lo_lo_75};
  wire [1023:0] dataGroup_hi_75 = {dataGroup_hi_hi_75, dataGroup_hi_lo_75};
  wire [7:0]    dataGroup_11_2 = dataGroup_lo_75[191:184];
  wire [1023:0] dataGroup_lo_76 = {dataGroup_lo_hi_76, dataGroup_lo_lo_76};
  wire [1023:0] dataGroup_hi_76 = {dataGroup_hi_hi_76, dataGroup_hi_lo_76};
  wire [7:0]    dataGroup_12_2 = dataGroup_lo_76[207:200];
  wire [1023:0] dataGroup_lo_77 = {dataGroup_lo_hi_77, dataGroup_lo_lo_77};
  wire [1023:0] dataGroup_hi_77 = {dataGroup_hi_hi_77, dataGroup_hi_lo_77};
  wire [7:0]    dataGroup_13_2 = dataGroup_lo_77[223:216];
  wire [1023:0] dataGroup_lo_78 = {dataGroup_lo_hi_78, dataGroup_lo_lo_78};
  wire [1023:0] dataGroup_hi_78 = {dataGroup_hi_hi_78, dataGroup_hi_lo_78};
  wire [7:0]    dataGroup_14_2 = dataGroup_lo_78[239:232];
  wire [1023:0] dataGroup_lo_79 = {dataGroup_lo_hi_79, dataGroup_lo_lo_79};
  wire [1023:0] dataGroup_hi_79 = {dataGroup_hi_hi_79, dataGroup_hi_lo_79};
  wire [7:0]    dataGroup_15_2 = dataGroup_lo_79[255:248];
  wire [1023:0] dataGroup_lo_80 = {dataGroup_lo_hi_80, dataGroup_lo_lo_80};
  wire [1023:0] dataGroup_hi_80 = {dataGroup_hi_hi_80, dataGroup_hi_lo_80};
  wire [7:0]    dataGroup_16_2 = dataGroup_lo_80[271:264];
  wire [1023:0] dataGroup_lo_81 = {dataGroup_lo_hi_81, dataGroup_lo_lo_81};
  wire [1023:0] dataGroup_hi_81 = {dataGroup_hi_hi_81, dataGroup_hi_lo_81};
  wire [7:0]    dataGroup_17_2 = dataGroup_lo_81[287:280];
  wire [1023:0] dataGroup_lo_82 = {dataGroup_lo_hi_82, dataGroup_lo_lo_82};
  wire [1023:0] dataGroup_hi_82 = {dataGroup_hi_hi_82, dataGroup_hi_lo_82};
  wire [7:0]    dataGroup_18_2 = dataGroup_lo_82[303:296];
  wire [1023:0] dataGroup_lo_83 = {dataGroup_lo_hi_83, dataGroup_lo_lo_83};
  wire [1023:0] dataGroup_hi_83 = {dataGroup_hi_hi_83, dataGroup_hi_lo_83};
  wire [7:0]    dataGroup_19_2 = dataGroup_lo_83[319:312];
  wire [1023:0] dataGroup_lo_84 = {dataGroup_lo_hi_84, dataGroup_lo_lo_84};
  wire [1023:0] dataGroup_hi_84 = {dataGroup_hi_hi_84, dataGroup_hi_lo_84};
  wire [7:0]    dataGroup_20_2 = dataGroup_lo_84[335:328];
  wire [1023:0] dataGroup_lo_85 = {dataGroup_lo_hi_85, dataGroup_lo_lo_85};
  wire [1023:0] dataGroup_hi_85 = {dataGroup_hi_hi_85, dataGroup_hi_lo_85};
  wire [7:0]    dataGroup_21_2 = dataGroup_lo_85[351:344];
  wire [1023:0] dataGroup_lo_86 = {dataGroup_lo_hi_86, dataGroup_lo_lo_86};
  wire [1023:0] dataGroup_hi_86 = {dataGroup_hi_hi_86, dataGroup_hi_lo_86};
  wire [7:0]    dataGroup_22_2 = dataGroup_lo_86[367:360];
  wire [1023:0] dataGroup_lo_87 = {dataGroup_lo_hi_87, dataGroup_lo_lo_87};
  wire [1023:0] dataGroup_hi_87 = {dataGroup_hi_hi_87, dataGroup_hi_lo_87};
  wire [7:0]    dataGroup_23_2 = dataGroup_lo_87[383:376];
  wire [1023:0] dataGroup_lo_88 = {dataGroup_lo_hi_88, dataGroup_lo_lo_88};
  wire [1023:0] dataGroup_hi_88 = {dataGroup_hi_hi_88, dataGroup_hi_lo_88};
  wire [7:0]    dataGroup_24_2 = dataGroup_lo_88[399:392];
  wire [1023:0] dataGroup_lo_89 = {dataGroup_lo_hi_89, dataGroup_lo_lo_89};
  wire [1023:0] dataGroup_hi_89 = {dataGroup_hi_hi_89, dataGroup_hi_lo_89};
  wire [7:0]    dataGroup_25_2 = dataGroup_lo_89[415:408];
  wire [1023:0] dataGroup_lo_90 = {dataGroup_lo_hi_90, dataGroup_lo_lo_90};
  wire [1023:0] dataGroup_hi_90 = {dataGroup_hi_hi_90, dataGroup_hi_lo_90};
  wire [7:0]    dataGroup_26_2 = dataGroup_lo_90[431:424];
  wire [1023:0] dataGroup_lo_91 = {dataGroup_lo_hi_91, dataGroup_lo_lo_91};
  wire [1023:0] dataGroup_hi_91 = {dataGroup_hi_hi_91, dataGroup_hi_lo_91};
  wire [7:0]    dataGroup_27_2 = dataGroup_lo_91[447:440];
  wire [1023:0] dataGroup_lo_92 = {dataGroup_lo_hi_92, dataGroup_lo_lo_92};
  wire [1023:0] dataGroup_hi_92 = {dataGroup_hi_hi_92, dataGroup_hi_lo_92};
  wire [7:0]    dataGroup_28_2 = dataGroup_lo_92[463:456];
  wire [1023:0] dataGroup_lo_93 = {dataGroup_lo_hi_93, dataGroup_lo_lo_93};
  wire [1023:0] dataGroup_hi_93 = {dataGroup_hi_hi_93, dataGroup_hi_lo_93};
  wire [7:0]    dataGroup_29_2 = dataGroup_lo_93[479:472];
  wire [1023:0] dataGroup_lo_94 = {dataGroup_lo_hi_94, dataGroup_lo_lo_94};
  wire [1023:0] dataGroup_hi_94 = {dataGroup_hi_hi_94, dataGroup_hi_lo_94};
  wire [7:0]    dataGroup_30_2 = dataGroup_lo_94[495:488];
  wire [1023:0] dataGroup_lo_95 = {dataGroup_lo_hi_95, dataGroup_lo_lo_95};
  wire [1023:0] dataGroup_hi_95 = {dataGroup_hi_hi_95, dataGroup_hi_lo_95};
  wire [7:0]    dataGroup_31_2 = dataGroup_lo_95[511:504];
  wire [15:0]   res_lo_lo_lo_lo_2 = {dataGroup_1_2, dataGroup_0_2};
  wire [15:0]   res_lo_lo_lo_hi_2 = {dataGroup_3_2, dataGroup_2_2};
  wire [31:0]   res_lo_lo_lo_2 = {res_lo_lo_lo_hi_2, res_lo_lo_lo_lo_2};
  wire [15:0]   res_lo_lo_hi_lo_2 = {dataGroup_5_2, dataGroup_4_2};
  wire [15:0]   res_lo_lo_hi_hi_2 = {dataGroup_7_2, dataGroup_6_2};
  wire [31:0]   res_lo_lo_hi_2 = {res_lo_lo_hi_hi_2, res_lo_lo_hi_lo_2};
  wire [63:0]   res_lo_lo_2 = {res_lo_lo_hi_2, res_lo_lo_lo_2};
  wire [15:0]   res_lo_hi_lo_lo_2 = {dataGroup_9_2, dataGroup_8_2};
  wire [15:0]   res_lo_hi_lo_hi_2 = {dataGroup_11_2, dataGroup_10_2};
  wire [31:0]   res_lo_hi_lo_2 = {res_lo_hi_lo_hi_2, res_lo_hi_lo_lo_2};
  wire [15:0]   res_lo_hi_hi_lo_2 = {dataGroup_13_2, dataGroup_12_2};
  wire [15:0]   res_lo_hi_hi_hi_2 = {dataGroup_15_2, dataGroup_14_2};
  wire [31:0]   res_lo_hi_hi_2 = {res_lo_hi_hi_hi_2, res_lo_hi_hi_lo_2};
  wire [63:0]   res_lo_hi_2 = {res_lo_hi_hi_2, res_lo_hi_lo_2};
  wire [127:0]  res_lo_2 = {res_lo_hi_2, res_lo_lo_2};
  wire [15:0]   res_hi_lo_lo_lo_2 = {dataGroup_17_2, dataGroup_16_2};
  wire [15:0]   res_hi_lo_lo_hi_2 = {dataGroup_19_2, dataGroup_18_2};
  wire [31:0]   res_hi_lo_lo_2 = {res_hi_lo_lo_hi_2, res_hi_lo_lo_lo_2};
  wire [15:0]   res_hi_lo_hi_lo_2 = {dataGroup_21_2, dataGroup_20_2};
  wire [15:0]   res_hi_lo_hi_hi_2 = {dataGroup_23_2, dataGroup_22_2};
  wire [31:0]   res_hi_lo_hi_2 = {res_hi_lo_hi_hi_2, res_hi_lo_hi_lo_2};
  wire [63:0]   res_hi_lo_2 = {res_hi_lo_hi_2, res_hi_lo_lo_2};
  wire [15:0]   res_hi_hi_lo_lo_2 = {dataGroup_25_2, dataGroup_24_2};
  wire [15:0]   res_hi_hi_lo_hi_2 = {dataGroup_27_2, dataGroup_26_2};
  wire [31:0]   res_hi_hi_lo_2 = {res_hi_hi_lo_hi_2, res_hi_hi_lo_lo_2};
  wire [15:0]   res_hi_hi_hi_lo_2 = {dataGroup_29_2, dataGroup_28_2};
  wire [15:0]   res_hi_hi_hi_hi_2 = {dataGroup_31_2, dataGroup_30_2};
  wire [31:0]   res_hi_hi_hi_2 = {res_hi_hi_hi_hi_2, res_hi_hi_hi_lo_2};
  wire [63:0]   res_hi_hi_2 = {res_hi_hi_hi_2, res_hi_hi_lo_2};
  wire [127:0]  res_hi_2 = {res_hi_hi_2, res_hi_lo_2};
  wire [255:0]  res_9 = {res_hi_2, res_lo_2};
  wire [511:0]  lo_lo_1 = {res_9, res_8};
  wire [1023:0] lo_1 = {512'h0, lo_lo_1};
  wire [2047:0] regroupLoadData_0_1 = {1024'h0, lo_1};
  wire [1023:0] dataGroup_lo_96 = {dataGroup_lo_hi_96, dataGroup_lo_lo_96};
  wire [1023:0] dataGroup_hi_96 = {dataGroup_hi_hi_96, dataGroup_hi_lo_96};
  wire [7:0]    dataGroup_0_3 = dataGroup_lo_96[7:0];
  wire [1023:0] dataGroup_lo_97 = {dataGroup_lo_hi_97, dataGroup_lo_lo_97};
  wire [1023:0] dataGroup_hi_97 = {dataGroup_hi_hi_97, dataGroup_hi_lo_97};
  wire [7:0]    dataGroup_1_3 = dataGroup_lo_97[31:24];
  wire [1023:0] dataGroup_lo_98 = {dataGroup_lo_hi_98, dataGroup_lo_lo_98};
  wire [1023:0] dataGroup_hi_98 = {dataGroup_hi_hi_98, dataGroup_hi_lo_98};
  wire [7:0]    dataGroup_2_3 = dataGroup_lo_98[55:48];
  wire [1023:0] dataGroup_lo_99 = {dataGroup_lo_hi_99, dataGroup_lo_lo_99};
  wire [1023:0] dataGroup_hi_99 = {dataGroup_hi_hi_99, dataGroup_hi_lo_99};
  wire [7:0]    dataGroup_3_3 = dataGroup_lo_99[79:72];
  wire [1023:0] dataGroup_lo_100 = {dataGroup_lo_hi_100, dataGroup_lo_lo_100};
  wire [1023:0] dataGroup_hi_100 = {dataGroup_hi_hi_100, dataGroup_hi_lo_100};
  wire [7:0]    dataGroup_4_3 = dataGroup_lo_100[103:96];
  wire [1023:0] dataGroup_lo_101 = {dataGroup_lo_hi_101, dataGroup_lo_lo_101};
  wire [1023:0] dataGroup_hi_101 = {dataGroup_hi_hi_101, dataGroup_hi_lo_101};
  wire [7:0]    dataGroup_5_3 = dataGroup_lo_101[127:120];
  wire [1023:0] dataGroup_lo_102 = {dataGroup_lo_hi_102, dataGroup_lo_lo_102};
  wire [1023:0] dataGroup_hi_102 = {dataGroup_hi_hi_102, dataGroup_hi_lo_102};
  wire [7:0]    dataGroup_6_3 = dataGroup_lo_102[151:144];
  wire [1023:0] dataGroup_lo_103 = {dataGroup_lo_hi_103, dataGroup_lo_lo_103};
  wire [1023:0] dataGroup_hi_103 = {dataGroup_hi_hi_103, dataGroup_hi_lo_103};
  wire [7:0]    dataGroup_7_3 = dataGroup_lo_103[175:168];
  wire [1023:0] dataGroup_lo_104 = {dataGroup_lo_hi_104, dataGroup_lo_lo_104};
  wire [1023:0] dataGroup_hi_104 = {dataGroup_hi_hi_104, dataGroup_hi_lo_104};
  wire [7:0]    dataGroup_8_3 = dataGroup_lo_104[199:192];
  wire [1023:0] dataGroup_lo_105 = {dataGroup_lo_hi_105, dataGroup_lo_lo_105};
  wire [1023:0] dataGroup_hi_105 = {dataGroup_hi_hi_105, dataGroup_hi_lo_105};
  wire [7:0]    dataGroup_9_3 = dataGroup_lo_105[223:216];
  wire [1023:0] dataGroup_lo_106 = {dataGroup_lo_hi_106, dataGroup_lo_lo_106};
  wire [1023:0] dataGroup_hi_106 = {dataGroup_hi_hi_106, dataGroup_hi_lo_106};
  wire [7:0]    dataGroup_10_3 = dataGroup_lo_106[247:240];
  wire [1023:0] dataGroup_lo_107 = {dataGroup_lo_hi_107, dataGroup_lo_lo_107};
  wire [1023:0] dataGroup_hi_107 = {dataGroup_hi_hi_107, dataGroup_hi_lo_107};
  wire [7:0]    dataGroup_11_3 = dataGroup_lo_107[271:264];
  wire [1023:0] dataGroup_lo_108 = {dataGroup_lo_hi_108, dataGroup_lo_lo_108};
  wire [1023:0] dataGroup_hi_108 = {dataGroup_hi_hi_108, dataGroup_hi_lo_108};
  wire [7:0]    dataGroup_12_3 = dataGroup_lo_108[295:288];
  wire [1023:0] dataGroup_lo_109 = {dataGroup_lo_hi_109, dataGroup_lo_lo_109};
  wire [1023:0] dataGroup_hi_109 = {dataGroup_hi_hi_109, dataGroup_hi_lo_109};
  wire [7:0]    dataGroup_13_3 = dataGroup_lo_109[319:312];
  wire [1023:0] dataGroup_lo_110 = {dataGroup_lo_hi_110, dataGroup_lo_lo_110};
  wire [1023:0] dataGroup_hi_110 = {dataGroup_hi_hi_110, dataGroup_hi_lo_110};
  wire [7:0]    dataGroup_14_3 = dataGroup_lo_110[343:336];
  wire [1023:0] dataGroup_lo_111 = {dataGroup_lo_hi_111, dataGroup_lo_lo_111};
  wire [1023:0] dataGroup_hi_111 = {dataGroup_hi_hi_111, dataGroup_hi_lo_111};
  wire [7:0]    dataGroup_15_3 = dataGroup_lo_111[367:360];
  wire [1023:0] dataGroup_lo_112 = {dataGroup_lo_hi_112, dataGroup_lo_lo_112};
  wire [1023:0] dataGroup_hi_112 = {dataGroup_hi_hi_112, dataGroup_hi_lo_112};
  wire [7:0]    dataGroup_16_3 = dataGroup_lo_112[391:384];
  wire [1023:0] dataGroup_lo_113 = {dataGroup_lo_hi_113, dataGroup_lo_lo_113};
  wire [1023:0] dataGroup_hi_113 = {dataGroup_hi_hi_113, dataGroup_hi_lo_113};
  wire [7:0]    dataGroup_17_3 = dataGroup_lo_113[415:408];
  wire [1023:0] dataGroup_lo_114 = {dataGroup_lo_hi_114, dataGroup_lo_lo_114};
  wire [1023:0] dataGroup_hi_114 = {dataGroup_hi_hi_114, dataGroup_hi_lo_114};
  wire [7:0]    dataGroup_18_3 = dataGroup_lo_114[439:432];
  wire [1023:0] dataGroup_lo_115 = {dataGroup_lo_hi_115, dataGroup_lo_lo_115};
  wire [1023:0] dataGroup_hi_115 = {dataGroup_hi_hi_115, dataGroup_hi_lo_115};
  wire [7:0]    dataGroup_19_3 = dataGroup_lo_115[463:456];
  wire [1023:0] dataGroup_lo_116 = {dataGroup_lo_hi_116, dataGroup_lo_lo_116};
  wire [1023:0] dataGroup_hi_116 = {dataGroup_hi_hi_116, dataGroup_hi_lo_116};
  wire [7:0]    dataGroup_20_3 = dataGroup_lo_116[487:480];
  wire [1023:0] dataGroup_lo_117 = {dataGroup_lo_hi_117, dataGroup_lo_lo_117};
  wire [1023:0] dataGroup_hi_117 = {dataGroup_hi_hi_117, dataGroup_hi_lo_117};
  wire [7:0]    dataGroup_21_3 = dataGroup_lo_117[511:504];
  wire [1023:0] dataGroup_lo_118 = {dataGroup_lo_hi_118, dataGroup_lo_lo_118};
  wire [1023:0] dataGroup_hi_118 = {dataGroup_hi_hi_118, dataGroup_hi_lo_118};
  wire [7:0]    dataGroup_22_3 = dataGroup_lo_118[535:528];
  wire [1023:0] dataGroup_lo_119 = {dataGroup_lo_hi_119, dataGroup_lo_lo_119};
  wire [1023:0] dataGroup_hi_119 = {dataGroup_hi_hi_119, dataGroup_hi_lo_119};
  wire [7:0]    dataGroup_23_3 = dataGroup_lo_119[559:552];
  wire [1023:0] dataGroup_lo_120 = {dataGroup_lo_hi_120, dataGroup_lo_lo_120};
  wire [1023:0] dataGroup_hi_120 = {dataGroup_hi_hi_120, dataGroup_hi_lo_120};
  wire [7:0]    dataGroup_24_3 = dataGroup_lo_120[583:576];
  wire [1023:0] dataGroup_lo_121 = {dataGroup_lo_hi_121, dataGroup_lo_lo_121};
  wire [1023:0] dataGroup_hi_121 = {dataGroup_hi_hi_121, dataGroup_hi_lo_121};
  wire [7:0]    dataGroup_25_3 = dataGroup_lo_121[607:600];
  wire [1023:0] dataGroup_lo_122 = {dataGroup_lo_hi_122, dataGroup_lo_lo_122};
  wire [1023:0] dataGroup_hi_122 = {dataGroup_hi_hi_122, dataGroup_hi_lo_122};
  wire [7:0]    dataGroup_26_3 = dataGroup_lo_122[631:624];
  wire [1023:0] dataGroup_lo_123 = {dataGroup_lo_hi_123, dataGroup_lo_lo_123};
  wire [1023:0] dataGroup_hi_123 = {dataGroup_hi_hi_123, dataGroup_hi_lo_123};
  wire [7:0]    dataGroup_27_3 = dataGroup_lo_123[655:648];
  wire [1023:0] dataGroup_lo_124 = {dataGroup_lo_hi_124, dataGroup_lo_lo_124};
  wire [1023:0] dataGroup_hi_124 = {dataGroup_hi_hi_124, dataGroup_hi_lo_124};
  wire [7:0]    dataGroup_28_3 = dataGroup_lo_124[679:672];
  wire [1023:0] dataGroup_lo_125 = {dataGroup_lo_hi_125, dataGroup_lo_lo_125};
  wire [1023:0] dataGroup_hi_125 = {dataGroup_hi_hi_125, dataGroup_hi_lo_125};
  wire [7:0]    dataGroup_29_3 = dataGroup_lo_125[703:696];
  wire [1023:0] dataGroup_lo_126 = {dataGroup_lo_hi_126, dataGroup_lo_lo_126};
  wire [1023:0] dataGroup_hi_126 = {dataGroup_hi_hi_126, dataGroup_hi_lo_126};
  wire [7:0]    dataGroup_30_3 = dataGroup_lo_126[727:720];
  wire [1023:0] dataGroup_lo_127 = {dataGroup_lo_hi_127, dataGroup_lo_lo_127};
  wire [1023:0] dataGroup_hi_127 = {dataGroup_hi_hi_127, dataGroup_hi_lo_127};
  wire [7:0]    dataGroup_31_3 = dataGroup_lo_127[751:744];
  wire [15:0]   res_lo_lo_lo_lo_3 = {dataGroup_1_3, dataGroup_0_3};
  wire [15:0]   res_lo_lo_lo_hi_3 = {dataGroup_3_3, dataGroup_2_3};
  wire [31:0]   res_lo_lo_lo_3 = {res_lo_lo_lo_hi_3, res_lo_lo_lo_lo_3};
  wire [15:0]   res_lo_lo_hi_lo_3 = {dataGroup_5_3, dataGroup_4_3};
  wire [15:0]   res_lo_lo_hi_hi_3 = {dataGroup_7_3, dataGroup_6_3};
  wire [31:0]   res_lo_lo_hi_3 = {res_lo_lo_hi_hi_3, res_lo_lo_hi_lo_3};
  wire [63:0]   res_lo_lo_3 = {res_lo_lo_hi_3, res_lo_lo_lo_3};
  wire [15:0]   res_lo_hi_lo_lo_3 = {dataGroup_9_3, dataGroup_8_3};
  wire [15:0]   res_lo_hi_lo_hi_3 = {dataGroup_11_3, dataGroup_10_3};
  wire [31:0]   res_lo_hi_lo_3 = {res_lo_hi_lo_hi_3, res_lo_hi_lo_lo_3};
  wire [15:0]   res_lo_hi_hi_lo_3 = {dataGroup_13_3, dataGroup_12_3};
  wire [15:0]   res_lo_hi_hi_hi_3 = {dataGroup_15_3, dataGroup_14_3};
  wire [31:0]   res_lo_hi_hi_3 = {res_lo_hi_hi_hi_3, res_lo_hi_hi_lo_3};
  wire [63:0]   res_lo_hi_3 = {res_lo_hi_hi_3, res_lo_hi_lo_3};
  wire [127:0]  res_lo_3 = {res_lo_hi_3, res_lo_lo_3};
  wire [15:0]   res_hi_lo_lo_lo_3 = {dataGroup_17_3, dataGroup_16_3};
  wire [15:0]   res_hi_lo_lo_hi_3 = {dataGroup_19_3, dataGroup_18_3};
  wire [31:0]   res_hi_lo_lo_3 = {res_hi_lo_lo_hi_3, res_hi_lo_lo_lo_3};
  wire [15:0]   res_hi_lo_hi_lo_3 = {dataGroup_21_3, dataGroup_20_3};
  wire [15:0]   res_hi_lo_hi_hi_3 = {dataGroup_23_3, dataGroup_22_3};
  wire [31:0]   res_hi_lo_hi_3 = {res_hi_lo_hi_hi_3, res_hi_lo_hi_lo_3};
  wire [63:0]   res_hi_lo_3 = {res_hi_lo_hi_3, res_hi_lo_lo_3};
  wire [15:0]   res_hi_hi_lo_lo_3 = {dataGroup_25_3, dataGroup_24_3};
  wire [15:0]   res_hi_hi_lo_hi_3 = {dataGroup_27_3, dataGroup_26_3};
  wire [31:0]   res_hi_hi_lo_3 = {res_hi_hi_lo_hi_3, res_hi_hi_lo_lo_3};
  wire [15:0]   res_hi_hi_hi_lo_3 = {dataGroup_29_3, dataGroup_28_3};
  wire [15:0]   res_hi_hi_hi_hi_3 = {dataGroup_31_3, dataGroup_30_3};
  wire [31:0]   res_hi_hi_hi_3 = {res_hi_hi_hi_hi_3, res_hi_hi_hi_lo_3};
  wire [63:0]   res_hi_hi_3 = {res_hi_hi_hi_3, res_hi_hi_lo_3};
  wire [127:0]  res_hi_3 = {res_hi_hi_3, res_hi_lo_3};
  wire [255:0]  res_16 = {res_hi_3, res_lo_3};
  wire [1023:0] dataGroup_lo_128 = {dataGroup_lo_hi_128, dataGroup_lo_lo_128};
  wire [1023:0] dataGroup_hi_128 = {dataGroup_hi_hi_128, dataGroup_hi_lo_128};
  wire [7:0]    dataGroup_0_4 = dataGroup_lo_128[15:8];
  wire [1023:0] dataGroup_lo_129 = {dataGroup_lo_hi_129, dataGroup_lo_lo_129};
  wire [1023:0] dataGroup_hi_129 = {dataGroup_hi_hi_129, dataGroup_hi_lo_129};
  wire [7:0]    dataGroup_1_4 = dataGroup_lo_129[39:32];
  wire [1023:0] dataGroup_lo_130 = {dataGroup_lo_hi_130, dataGroup_lo_lo_130};
  wire [1023:0] dataGroup_hi_130 = {dataGroup_hi_hi_130, dataGroup_hi_lo_130};
  wire [7:0]    dataGroup_2_4 = dataGroup_lo_130[63:56];
  wire [1023:0] dataGroup_lo_131 = {dataGroup_lo_hi_131, dataGroup_lo_lo_131};
  wire [1023:0] dataGroup_hi_131 = {dataGroup_hi_hi_131, dataGroup_hi_lo_131};
  wire [7:0]    dataGroup_3_4 = dataGroup_lo_131[87:80];
  wire [1023:0] dataGroup_lo_132 = {dataGroup_lo_hi_132, dataGroup_lo_lo_132};
  wire [1023:0] dataGroup_hi_132 = {dataGroup_hi_hi_132, dataGroup_hi_lo_132};
  wire [7:0]    dataGroup_4_4 = dataGroup_lo_132[111:104];
  wire [1023:0] dataGroup_lo_133 = {dataGroup_lo_hi_133, dataGroup_lo_lo_133};
  wire [1023:0] dataGroup_hi_133 = {dataGroup_hi_hi_133, dataGroup_hi_lo_133};
  wire [7:0]    dataGroup_5_4 = dataGroup_lo_133[135:128];
  wire [1023:0] dataGroup_lo_134 = {dataGroup_lo_hi_134, dataGroup_lo_lo_134};
  wire [1023:0] dataGroup_hi_134 = {dataGroup_hi_hi_134, dataGroup_hi_lo_134};
  wire [7:0]    dataGroup_6_4 = dataGroup_lo_134[159:152];
  wire [1023:0] dataGroup_lo_135 = {dataGroup_lo_hi_135, dataGroup_lo_lo_135};
  wire [1023:0] dataGroup_hi_135 = {dataGroup_hi_hi_135, dataGroup_hi_lo_135};
  wire [7:0]    dataGroup_7_4 = dataGroup_lo_135[183:176];
  wire [1023:0] dataGroup_lo_136 = {dataGroup_lo_hi_136, dataGroup_lo_lo_136};
  wire [1023:0] dataGroup_hi_136 = {dataGroup_hi_hi_136, dataGroup_hi_lo_136};
  wire [7:0]    dataGroup_8_4 = dataGroup_lo_136[207:200];
  wire [1023:0] dataGroup_lo_137 = {dataGroup_lo_hi_137, dataGroup_lo_lo_137};
  wire [1023:0] dataGroup_hi_137 = {dataGroup_hi_hi_137, dataGroup_hi_lo_137};
  wire [7:0]    dataGroup_9_4 = dataGroup_lo_137[231:224];
  wire [1023:0] dataGroup_lo_138 = {dataGroup_lo_hi_138, dataGroup_lo_lo_138};
  wire [1023:0] dataGroup_hi_138 = {dataGroup_hi_hi_138, dataGroup_hi_lo_138};
  wire [7:0]    dataGroup_10_4 = dataGroup_lo_138[255:248];
  wire [1023:0] dataGroup_lo_139 = {dataGroup_lo_hi_139, dataGroup_lo_lo_139};
  wire [1023:0] dataGroup_hi_139 = {dataGroup_hi_hi_139, dataGroup_hi_lo_139};
  wire [7:0]    dataGroup_11_4 = dataGroup_lo_139[279:272];
  wire [1023:0] dataGroup_lo_140 = {dataGroup_lo_hi_140, dataGroup_lo_lo_140};
  wire [1023:0] dataGroup_hi_140 = {dataGroup_hi_hi_140, dataGroup_hi_lo_140};
  wire [7:0]    dataGroup_12_4 = dataGroup_lo_140[303:296];
  wire [1023:0] dataGroup_lo_141 = {dataGroup_lo_hi_141, dataGroup_lo_lo_141};
  wire [1023:0] dataGroup_hi_141 = {dataGroup_hi_hi_141, dataGroup_hi_lo_141};
  wire [7:0]    dataGroup_13_4 = dataGroup_lo_141[327:320];
  wire [1023:0] dataGroup_lo_142 = {dataGroup_lo_hi_142, dataGroup_lo_lo_142};
  wire [1023:0] dataGroup_hi_142 = {dataGroup_hi_hi_142, dataGroup_hi_lo_142};
  wire [7:0]    dataGroup_14_4 = dataGroup_lo_142[351:344];
  wire [1023:0] dataGroup_lo_143 = {dataGroup_lo_hi_143, dataGroup_lo_lo_143};
  wire [1023:0] dataGroup_hi_143 = {dataGroup_hi_hi_143, dataGroup_hi_lo_143};
  wire [7:0]    dataGroup_15_4 = dataGroup_lo_143[375:368];
  wire [1023:0] dataGroup_lo_144 = {dataGroup_lo_hi_144, dataGroup_lo_lo_144};
  wire [1023:0] dataGroup_hi_144 = {dataGroup_hi_hi_144, dataGroup_hi_lo_144};
  wire [7:0]    dataGroup_16_4 = dataGroup_lo_144[399:392];
  wire [1023:0] dataGroup_lo_145 = {dataGroup_lo_hi_145, dataGroup_lo_lo_145};
  wire [1023:0] dataGroup_hi_145 = {dataGroup_hi_hi_145, dataGroup_hi_lo_145};
  wire [7:0]    dataGroup_17_4 = dataGroup_lo_145[423:416];
  wire [1023:0] dataGroup_lo_146 = {dataGroup_lo_hi_146, dataGroup_lo_lo_146};
  wire [1023:0] dataGroup_hi_146 = {dataGroup_hi_hi_146, dataGroup_hi_lo_146};
  wire [7:0]    dataGroup_18_4 = dataGroup_lo_146[447:440];
  wire [1023:0] dataGroup_lo_147 = {dataGroup_lo_hi_147, dataGroup_lo_lo_147};
  wire [1023:0] dataGroup_hi_147 = {dataGroup_hi_hi_147, dataGroup_hi_lo_147};
  wire [7:0]    dataGroup_19_4 = dataGroup_lo_147[471:464];
  wire [1023:0] dataGroup_lo_148 = {dataGroup_lo_hi_148, dataGroup_lo_lo_148};
  wire [1023:0] dataGroup_hi_148 = {dataGroup_hi_hi_148, dataGroup_hi_lo_148};
  wire [7:0]    dataGroup_20_4 = dataGroup_lo_148[495:488];
  wire [1023:0] dataGroup_lo_149 = {dataGroup_lo_hi_149, dataGroup_lo_lo_149};
  wire [1023:0] dataGroup_hi_149 = {dataGroup_hi_hi_149, dataGroup_hi_lo_149};
  wire [7:0]    dataGroup_21_4 = dataGroup_lo_149[519:512];
  wire [1023:0] dataGroup_lo_150 = {dataGroup_lo_hi_150, dataGroup_lo_lo_150};
  wire [1023:0] dataGroup_hi_150 = {dataGroup_hi_hi_150, dataGroup_hi_lo_150};
  wire [7:0]    dataGroup_22_4 = dataGroup_lo_150[543:536];
  wire [1023:0] dataGroup_lo_151 = {dataGroup_lo_hi_151, dataGroup_lo_lo_151};
  wire [1023:0] dataGroup_hi_151 = {dataGroup_hi_hi_151, dataGroup_hi_lo_151};
  wire [7:0]    dataGroup_23_4 = dataGroup_lo_151[567:560];
  wire [1023:0] dataGroup_lo_152 = {dataGroup_lo_hi_152, dataGroup_lo_lo_152};
  wire [1023:0] dataGroup_hi_152 = {dataGroup_hi_hi_152, dataGroup_hi_lo_152};
  wire [7:0]    dataGroup_24_4 = dataGroup_lo_152[591:584];
  wire [1023:0] dataGroup_lo_153 = {dataGroup_lo_hi_153, dataGroup_lo_lo_153};
  wire [1023:0] dataGroup_hi_153 = {dataGroup_hi_hi_153, dataGroup_hi_lo_153};
  wire [7:0]    dataGroup_25_4 = dataGroup_lo_153[615:608];
  wire [1023:0] dataGroup_lo_154 = {dataGroup_lo_hi_154, dataGroup_lo_lo_154};
  wire [1023:0] dataGroup_hi_154 = {dataGroup_hi_hi_154, dataGroup_hi_lo_154};
  wire [7:0]    dataGroup_26_4 = dataGroup_lo_154[639:632];
  wire [1023:0] dataGroup_lo_155 = {dataGroup_lo_hi_155, dataGroup_lo_lo_155};
  wire [1023:0] dataGroup_hi_155 = {dataGroup_hi_hi_155, dataGroup_hi_lo_155};
  wire [7:0]    dataGroup_27_4 = dataGroup_lo_155[663:656];
  wire [1023:0] dataGroup_lo_156 = {dataGroup_lo_hi_156, dataGroup_lo_lo_156};
  wire [1023:0] dataGroup_hi_156 = {dataGroup_hi_hi_156, dataGroup_hi_lo_156};
  wire [7:0]    dataGroup_28_4 = dataGroup_lo_156[687:680];
  wire [1023:0] dataGroup_lo_157 = {dataGroup_lo_hi_157, dataGroup_lo_lo_157};
  wire [1023:0] dataGroup_hi_157 = {dataGroup_hi_hi_157, dataGroup_hi_lo_157};
  wire [7:0]    dataGroup_29_4 = dataGroup_lo_157[711:704];
  wire [1023:0] dataGroup_lo_158 = {dataGroup_lo_hi_158, dataGroup_lo_lo_158};
  wire [1023:0] dataGroup_hi_158 = {dataGroup_hi_hi_158, dataGroup_hi_lo_158};
  wire [7:0]    dataGroup_30_4 = dataGroup_lo_158[735:728];
  wire [1023:0] dataGroup_lo_159 = {dataGroup_lo_hi_159, dataGroup_lo_lo_159};
  wire [1023:0] dataGroup_hi_159 = {dataGroup_hi_hi_159, dataGroup_hi_lo_159};
  wire [7:0]    dataGroup_31_4 = dataGroup_lo_159[759:752];
  wire [15:0]   res_lo_lo_lo_lo_4 = {dataGroup_1_4, dataGroup_0_4};
  wire [15:0]   res_lo_lo_lo_hi_4 = {dataGroup_3_4, dataGroup_2_4};
  wire [31:0]   res_lo_lo_lo_4 = {res_lo_lo_lo_hi_4, res_lo_lo_lo_lo_4};
  wire [15:0]   res_lo_lo_hi_lo_4 = {dataGroup_5_4, dataGroup_4_4};
  wire [15:0]   res_lo_lo_hi_hi_4 = {dataGroup_7_4, dataGroup_6_4};
  wire [31:0]   res_lo_lo_hi_4 = {res_lo_lo_hi_hi_4, res_lo_lo_hi_lo_4};
  wire [63:0]   res_lo_lo_4 = {res_lo_lo_hi_4, res_lo_lo_lo_4};
  wire [15:0]   res_lo_hi_lo_lo_4 = {dataGroup_9_4, dataGroup_8_4};
  wire [15:0]   res_lo_hi_lo_hi_4 = {dataGroup_11_4, dataGroup_10_4};
  wire [31:0]   res_lo_hi_lo_4 = {res_lo_hi_lo_hi_4, res_lo_hi_lo_lo_4};
  wire [15:0]   res_lo_hi_hi_lo_4 = {dataGroup_13_4, dataGroup_12_4};
  wire [15:0]   res_lo_hi_hi_hi_4 = {dataGroup_15_4, dataGroup_14_4};
  wire [31:0]   res_lo_hi_hi_4 = {res_lo_hi_hi_hi_4, res_lo_hi_hi_lo_4};
  wire [63:0]   res_lo_hi_4 = {res_lo_hi_hi_4, res_lo_hi_lo_4};
  wire [127:0]  res_lo_4 = {res_lo_hi_4, res_lo_lo_4};
  wire [15:0]   res_hi_lo_lo_lo_4 = {dataGroup_17_4, dataGroup_16_4};
  wire [15:0]   res_hi_lo_lo_hi_4 = {dataGroup_19_4, dataGroup_18_4};
  wire [31:0]   res_hi_lo_lo_4 = {res_hi_lo_lo_hi_4, res_hi_lo_lo_lo_4};
  wire [15:0]   res_hi_lo_hi_lo_4 = {dataGroup_21_4, dataGroup_20_4};
  wire [15:0]   res_hi_lo_hi_hi_4 = {dataGroup_23_4, dataGroup_22_4};
  wire [31:0]   res_hi_lo_hi_4 = {res_hi_lo_hi_hi_4, res_hi_lo_hi_lo_4};
  wire [63:0]   res_hi_lo_4 = {res_hi_lo_hi_4, res_hi_lo_lo_4};
  wire [15:0]   res_hi_hi_lo_lo_4 = {dataGroup_25_4, dataGroup_24_4};
  wire [15:0]   res_hi_hi_lo_hi_4 = {dataGroup_27_4, dataGroup_26_4};
  wire [31:0]   res_hi_hi_lo_4 = {res_hi_hi_lo_hi_4, res_hi_hi_lo_lo_4};
  wire [15:0]   res_hi_hi_hi_lo_4 = {dataGroup_29_4, dataGroup_28_4};
  wire [15:0]   res_hi_hi_hi_hi_4 = {dataGroup_31_4, dataGroup_30_4};
  wire [31:0]   res_hi_hi_hi_4 = {res_hi_hi_hi_hi_4, res_hi_hi_hi_lo_4};
  wire [63:0]   res_hi_hi_4 = {res_hi_hi_hi_4, res_hi_hi_lo_4};
  wire [127:0]  res_hi_4 = {res_hi_hi_4, res_hi_lo_4};
  wire [255:0]  res_17 = {res_hi_4, res_lo_4};
  wire [1023:0] dataGroup_lo_160 = {dataGroup_lo_hi_160, dataGroup_lo_lo_160};
  wire [1023:0] dataGroup_hi_160 = {dataGroup_hi_hi_160, dataGroup_hi_lo_160};
  wire [7:0]    dataGroup_0_5 = dataGroup_lo_160[23:16];
  wire [1023:0] dataGroup_lo_161 = {dataGroup_lo_hi_161, dataGroup_lo_lo_161};
  wire [1023:0] dataGroup_hi_161 = {dataGroup_hi_hi_161, dataGroup_hi_lo_161};
  wire [7:0]    dataGroup_1_5 = dataGroup_lo_161[47:40];
  wire [1023:0] dataGroup_lo_162 = {dataGroup_lo_hi_162, dataGroup_lo_lo_162};
  wire [1023:0] dataGroup_hi_162 = {dataGroup_hi_hi_162, dataGroup_hi_lo_162};
  wire [7:0]    dataGroup_2_5 = dataGroup_lo_162[71:64];
  wire [1023:0] dataGroup_lo_163 = {dataGroup_lo_hi_163, dataGroup_lo_lo_163};
  wire [1023:0] dataGroup_hi_163 = {dataGroup_hi_hi_163, dataGroup_hi_lo_163};
  wire [7:0]    dataGroup_3_5 = dataGroup_lo_163[95:88];
  wire [1023:0] dataGroup_lo_164 = {dataGroup_lo_hi_164, dataGroup_lo_lo_164};
  wire [1023:0] dataGroup_hi_164 = {dataGroup_hi_hi_164, dataGroup_hi_lo_164};
  wire [7:0]    dataGroup_4_5 = dataGroup_lo_164[119:112];
  wire [1023:0] dataGroup_lo_165 = {dataGroup_lo_hi_165, dataGroup_lo_lo_165};
  wire [1023:0] dataGroup_hi_165 = {dataGroup_hi_hi_165, dataGroup_hi_lo_165};
  wire [7:0]    dataGroup_5_5 = dataGroup_lo_165[143:136];
  wire [1023:0] dataGroup_lo_166 = {dataGroup_lo_hi_166, dataGroup_lo_lo_166};
  wire [1023:0] dataGroup_hi_166 = {dataGroup_hi_hi_166, dataGroup_hi_lo_166};
  wire [7:0]    dataGroup_6_5 = dataGroup_lo_166[167:160];
  wire [1023:0] dataGroup_lo_167 = {dataGroup_lo_hi_167, dataGroup_lo_lo_167};
  wire [1023:0] dataGroup_hi_167 = {dataGroup_hi_hi_167, dataGroup_hi_lo_167};
  wire [7:0]    dataGroup_7_5 = dataGroup_lo_167[191:184];
  wire [1023:0] dataGroup_lo_168 = {dataGroup_lo_hi_168, dataGroup_lo_lo_168};
  wire [1023:0] dataGroup_hi_168 = {dataGroup_hi_hi_168, dataGroup_hi_lo_168};
  wire [7:0]    dataGroup_8_5 = dataGroup_lo_168[215:208];
  wire [1023:0] dataGroup_lo_169 = {dataGroup_lo_hi_169, dataGroup_lo_lo_169};
  wire [1023:0] dataGroup_hi_169 = {dataGroup_hi_hi_169, dataGroup_hi_lo_169};
  wire [7:0]    dataGroup_9_5 = dataGroup_lo_169[239:232];
  wire [1023:0] dataGroup_lo_170 = {dataGroup_lo_hi_170, dataGroup_lo_lo_170};
  wire [1023:0] dataGroup_hi_170 = {dataGroup_hi_hi_170, dataGroup_hi_lo_170};
  wire [7:0]    dataGroup_10_5 = dataGroup_lo_170[263:256];
  wire [1023:0] dataGroup_lo_171 = {dataGroup_lo_hi_171, dataGroup_lo_lo_171};
  wire [1023:0] dataGroup_hi_171 = {dataGroup_hi_hi_171, dataGroup_hi_lo_171};
  wire [7:0]    dataGroup_11_5 = dataGroup_lo_171[287:280];
  wire [1023:0] dataGroup_lo_172 = {dataGroup_lo_hi_172, dataGroup_lo_lo_172};
  wire [1023:0] dataGroup_hi_172 = {dataGroup_hi_hi_172, dataGroup_hi_lo_172};
  wire [7:0]    dataGroup_12_5 = dataGroup_lo_172[311:304];
  wire [1023:0] dataGroup_lo_173 = {dataGroup_lo_hi_173, dataGroup_lo_lo_173};
  wire [1023:0] dataGroup_hi_173 = {dataGroup_hi_hi_173, dataGroup_hi_lo_173};
  wire [7:0]    dataGroup_13_5 = dataGroup_lo_173[335:328];
  wire [1023:0] dataGroup_lo_174 = {dataGroup_lo_hi_174, dataGroup_lo_lo_174};
  wire [1023:0] dataGroup_hi_174 = {dataGroup_hi_hi_174, dataGroup_hi_lo_174};
  wire [7:0]    dataGroup_14_5 = dataGroup_lo_174[359:352];
  wire [1023:0] dataGroup_lo_175 = {dataGroup_lo_hi_175, dataGroup_lo_lo_175};
  wire [1023:0] dataGroup_hi_175 = {dataGroup_hi_hi_175, dataGroup_hi_lo_175};
  wire [7:0]    dataGroup_15_5 = dataGroup_lo_175[383:376];
  wire [1023:0] dataGroup_lo_176 = {dataGroup_lo_hi_176, dataGroup_lo_lo_176};
  wire [1023:0] dataGroup_hi_176 = {dataGroup_hi_hi_176, dataGroup_hi_lo_176};
  wire [7:0]    dataGroup_16_5 = dataGroup_lo_176[407:400];
  wire [1023:0] dataGroup_lo_177 = {dataGroup_lo_hi_177, dataGroup_lo_lo_177};
  wire [1023:0] dataGroup_hi_177 = {dataGroup_hi_hi_177, dataGroup_hi_lo_177};
  wire [7:0]    dataGroup_17_5 = dataGroup_lo_177[431:424];
  wire [1023:0] dataGroup_lo_178 = {dataGroup_lo_hi_178, dataGroup_lo_lo_178};
  wire [1023:0] dataGroup_hi_178 = {dataGroup_hi_hi_178, dataGroup_hi_lo_178};
  wire [7:0]    dataGroup_18_5 = dataGroup_lo_178[455:448];
  wire [1023:0] dataGroup_lo_179 = {dataGroup_lo_hi_179, dataGroup_lo_lo_179};
  wire [1023:0] dataGroup_hi_179 = {dataGroup_hi_hi_179, dataGroup_hi_lo_179};
  wire [7:0]    dataGroup_19_5 = dataGroup_lo_179[479:472];
  wire [1023:0] dataGroup_lo_180 = {dataGroup_lo_hi_180, dataGroup_lo_lo_180};
  wire [1023:0] dataGroup_hi_180 = {dataGroup_hi_hi_180, dataGroup_hi_lo_180};
  wire [7:0]    dataGroup_20_5 = dataGroup_lo_180[503:496];
  wire [1023:0] dataGroup_lo_181 = {dataGroup_lo_hi_181, dataGroup_lo_lo_181};
  wire [1023:0] dataGroup_hi_181 = {dataGroup_hi_hi_181, dataGroup_hi_lo_181};
  wire [7:0]    dataGroup_21_5 = dataGroup_lo_181[527:520];
  wire [1023:0] dataGroup_lo_182 = {dataGroup_lo_hi_182, dataGroup_lo_lo_182};
  wire [1023:0] dataGroup_hi_182 = {dataGroup_hi_hi_182, dataGroup_hi_lo_182};
  wire [7:0]    dataGroup_22_5 = dataGroup_lo_182[551:544];
  wire [1023:0] dataGroup_lo_183 = {dataGroup_lo_hi_183, dataGroup_lo_lo_183};
  wire [1023:0] dataGroup_hi_183 = {dataGroup_hi_hi_183, dataGroup_hi_lo_183};
  wire [7:0]    dataGroup_23_5 = dataGroup_lo_183[575:568];
  wire [1023:0] dataGroup_lo_184 = {dataGroup_lo_hi_184, dataGroup_lo_lo_184};
  wire [1023:0] dataGroup_hi_184 = {dataGroup_hi_hi_184, dataGroup_hi_lo_184};
  wire [7:0]    dataGroup_24_5 = dataGroup_lo_184[599:592];
  wire [1023:0] dataGroup_lo_185 = {dataGroup_lo_hi_185, dataGroup_lo_lo_185};
  wire [1023:0] dataGroup_hi_185 = {dataGroup_hi_hi_185, dataGroup_hi_lo_185};
  wire [7:0]    dataGroup_25_5 = dataGroup_lo_185[623:616];
  wire [1023:0] dataGroup_lo_186 = {dataGroup_lo_hi_186, dataGroup_lo_lo_186};
  wire [1023:0] dataGroup_hi_186 = {dataGroup_hi_hi_186, dataGroup_hi_lo_186};
  wire [7:0]    dataGroup_26_5 = dataGroup_lo_186[647:640];
  wire [1023:0] dataGroup_lo_187 = {dataGroup_lo_hi_187, dataGroup_lo_lo_187};
  wire [1023:0] dataGroup_hi_187 = {dataGroup_hi_hi_187, dataGroup_hi_lo_187};
  wire [7:0]    dataGroup_27_5 = dataGroup_lo_187[671:664];
  wire [1023:0] dataGroup_lo_188 = {dataGroup_lo_hi_188, dataGroup_lo_lo_188};
  wire [1023:0] dataGroup_hi_188 = {dataGroup_hi_hi_188, dataGroup_hi_lo_188};
  wire [7:0]    dataGroup_28_5 = dataGroup_lo_188[695:688];
  wire [1023:0] dataGroup_lo_189 = {dataGroup_lo_hi_189, dataGroup_lo_lo_189};
  wire [1023:0] dataGroup_hi_189 = {dataGroup_hi_hi_189, dataGroup_hi_lo_189};
  wire [7:0]    dataGroup_29_5 = dataGroup_lo_189[719:712];
  wire [1023:0] dataGroup_lo_190 = {dataGroup_lo_hi_190, dataGroup_lo_lo_190};
  wire [1023:0] dataGroup_hi_190 = {dataGroup_hi_hi_190, dataGroup_hi_lo_190};
  wire [7:0]    dataGroup_30_5 = dataGroup_lo_190[743:736];
  wire [1023:0] dataGroup_lo_191 = {dataGroup_lo_hi_191, dataGroup_lo_lo_191};
  wire [1023:0] dataGroup_hi_191 = {dataGroup_hi_hi_191, dataGroup_hi_lo_191};
  wire [7:0]    dataGroup_31_5 = dataGroup_lo_191[767:760];
  wire [15:0]   res_lo_lo_lo_lo_5 = {dataGroup_1_5, dataGroup_0_5};
  wire [15:0]   res_lo_lo_lo_hi_5 = {dataGroup_3_5, dataGroup_2_5};
  wire [31:0]   res_lo_lo_lo_5 = {res_lo_lo_lo_hi_5, res_lo_lo_lo_lo_5};
  wire [15:0]   res_lo_lo_hi_lo_5 = {dataGroup_5_5, dataGroup_4_5};
  wire [15:0]   res_lo_lo_hi_hi_5 = {dataGroup_7_5, dataGroup_6_5};
  wire [31:0]   res_lo_lo_hi_5 = {res_lo_lo_hi_hi_5, res_lo_lo_hi_lo_5};
  wire [63:0]   res_lo_lo_5 = {res_lo_lo_hi_5, res_lo_lo_lo_5};
  wire [15:0]   res_lo_hi_lo_lo_5 = {dataGroup_9_5, dataGroup_8_5};
  wire [15:0]   res_lo_hi_lo_hi_5 = {dataGroup_11_5, dataGroup_10_5};
  wire [31:0]   res_lo_hi_lo_5 = {res_lo_hi_lo_hi_5, res_lo_hi_lo_lo_5};
  wire [15:0]   res_lo_hi_hi_lo_5 = {dataGroup_13_5, dataGroup_12_5};
  wire [15:0]   res_lo_hi_hi_hi_5 = {dataGroup_15_5, dataGroup_14_5};
  wire [31:0]   res_lo_hi_hi_5 = {res_lo_hi_hi_hi_5, res_lo_hi_hi_lo_5};
  wire [63:0]   res_lo_hi_5 = {res_lo_hi_hi_5, res_lo_hi_lo_5};
  wire [127:0]  res_lo_5 = {res_lo_hi_5, res_lo_lo_5};
  wire [15:0]   res_hi_lo_lo_lo_5 = {dataGroup_17_5, dataGroup_16_5};
  wire [15:0]   res_hi_lo_lo_hi_5 = {dataGroup_19_5, dataGroup_18_5};
  wire [31:0]   res_hi_lo_lo_5 = {res_hi_lo_lo_hi_5, res_hi_lo_lo_lo_5};
  wire [15:0]   res_hi_lo_hi_lo_5 = {dataGroup_21_5, dataGroup_20_5};
  wire [15:0]   res_hi_lo_hi_hi_5 = {dataGroup_23_5, dataGroup_22_5};
  wire [31:0]   res_hi_lo_hi_5 = {res_hi_lo_hi_hi_5, res_hi_lo_hi_lo_5};
  wire [63:0]   res_hi_lo_5 = {res_hi_lo_hi_5, res_hi_lo_lo_5};
  wire [15:0]   res_hi_hi_lo_lo_5 = {dataGroup_25_5, dataGroup_24_5};
  wire [15:0]   res_hi_hi_lo_hi_5 = {dataGroup_27_5, dataGroup_26_5};
  wire [31:0]   res_hi_hi_lo_5 = {res_hi_hi_lo_hi_5, res_hi_hi_lo_lo_5};
  wire [15:0]   res_hi_hi_hi_lo_5 = {dataGroup_29_5, dataGroup_28_5};
  wire [15:0]   res_hi_hi_hi_hi_5 = {dataGroup_31_5, dataGroup_30_5};
  wire [31:0]   res_hi_hi_hi_5 = {res_hi_hi_hi_hi_5, res_hi_hi_hi_lo_5};
  wire [63:0]   res_hi_hi_5 = {res_hi_hi_hi_5, res_hi_hi_lo_5};
  wire [127:0]  res_hi_5 = {res_hi_hi_5, res_hi_lo_5};
  wire [255:0]  res_18 = {res_hi_5, res_lo_5};
  wire [511:0]  lo_lo_2 = {res_17, res_16};
  wire [511:0]  lo_hi_2 = {256'h0, res_18};
  wire [1023:0] lo_2 = {lo_hi_2, lo_lo_2};
  wire [2047:0] regroupLoadData_0_2 = {1024'h0, lo_2};
  wire [1023:0] dataGroup_lo_192 = {dataGroup_lo_hi_192, dataGroup_lo_lo_192};
  wire [1023:0] dataGroup_hi_192 = {dataGroup_hi_hi_192, dataGroup_hi_lo_192};
  wire [7:0]    dataGroup_0_6 = dataGroup_lo_192[7:0];
  wire [1023:0] dataGroup_lo_193 = {dataGroup_lo_hi_193, dataGroup_lo_lo_193};
  wire [1023:0] dataGroup_hi_193 = {dataGroup_hi_hi_193, dataGroup_hi_lo_193};
  wire [7:0]    dataGroup_1_6 = dataGroup_lo_193[39:32];
  wire [1023:0] dataGroup_lo_194 = {dataGroup_lo_hi_194, dataGroup_lo_lo_194};
  wire [1023:0] dataGroup_hi_194 = {dataGroup_hi_hi_194, dataGroup_hi_lo_194};
  wire [7:0]    dataGroup_2_6 = dataGroup_lo_194[71:64];
  wire [1023:0] dataGroup_lo_195 = {dataGroup_lo_hi_195, dataGroup_lo_lo_195};
  wire [1023:0] dataGroup_hi_195 = {dataGroup_hi_hi_195, dataGroup_hi_lo_195};
  wire [7:0]    dataGroup_3_6 = dataGroup_lo_195[103:96];
  wire [1023:0] dataGroup_lo_196 = {dataGroup_lo_hi_196, dataGroup_lo_lo_196};
  wire [1023:0] dataGroup_hi_196 = {dataGroup_hi_hi_196, dataGroup_hi_lo_196};
  wire [7:0]    dataGroup_4_6 = dataGroup_lo_196[135:128];
  wire [1023:0] dataGroup_lo_197 = {dataGroup_lo_hi_197, dataGroup_lo_lo_197};
  wire [1023:0] dataGroup_hi_197 = {dataGroup_hi_hi_197, dataGroup_hi_lo_197};
  wire [7:0]    dataGroup_5_6 = dataGroup_lo_197[167:160];
  wire [1023:0] dataGroup_lo_198 = {dataGroup_lo_hi_198, dataGroup_lo_lo_198};
  wire [1023:0] dataGroup_hi_198 = {dataGroup_hi_hi_198, dataGroup_hi_lo_198};
  wire [7:0]    dataGroup_6_6 = dataGroup_lo_198[199:192];
  wire [1023:0] dataGroup_lo_199 = {dataGroup_lo_hi_199, dataGroup_lo_lo_199};
  wire [1023:0] dataGroup_hi_199 = {dataGroup_hi_hi_199, dataGroup_hi_lo_199};
  wire [7:0]    dataGroup_7_6 = dataGroup_lo_199[231:224];
  wire [1023:0] dataGroup_lo_200 = {dataGroup_lo_hi_200, dataGroup_lo_lo_200};
  wire [1023:0] dataGroup_hi_200 = {dataGroup_hi_hi_200, dataGroup_hi_lo_200};
  wire [7:0]    dataGroup_8_6 = dataGroup_lo_200[263:256];
  wire [1023:0] dataGroup_lo_201 = {dataGroup_lo_hi_201, dataGroup_lo_lo_201};
  wire [1023:0] dataGroup_hi_201 = {dataGroup_hi_hi_201, dataGroup_hi_lo_201};
  wire [7:0]    dataGroup_9_6 = dataGroup_lo_201[295:288];
  wire [1023:0] dataGroup_lo_202 = {dataGroup_lo_hi_202, dataGroup_lo_lo_202};
  wire [1023:0] dataGroup_hi_202 = {dataGroup_hi_hi_202, dataGroup_hi_lo_202};
  wire [7:0]    dataGroup_10_6 = dataGroup_lo_202[327:320];
  wire [1023:0] dataGroup_lo_203 = {dataGroup_lo_hi_203, dataGroup_lo_lo_203};
  wire [1023:0] dataGroup_hi_203 = {dataGroup_hi_hi_203, dataGroup_hi_lo_203};
  wire [7:0]    dataGroup_11_6 = dataGroup_lo_203[359:352];
  wire [1023:0] dataGroup_lo_204 = {dataGroup_lo_hi_204, dataGroup_lo_lo_204};
  wire [1023:0] dataGroup_hi_204 = {dataGroup_hi_hi_204, dataGroup_hi_lo_204};
  wire [7:0]    dataGroup_12_6 = dataGroup_lo_204[391:384];
  wire [1023:0] dataGroup_lo_205 = {dataGroup_lo_hi_205, dataGroup_lo_lo_205};
  wire [1023:0] dataGroup_hi_205 = {dataGroup_hi_hi_205, dataGroup_hi_lo_205};
  wire [7:0]    dataGroup_13_6 = dataGroup_lo_205[423:416];
  wire [1023:0] dataGroup_lo_206 = {dataGroup_lo_hi_206, dataGroup_lo_lo_206};
  wire [1023:0] dataGroup_hi_206 = {dataGroup_hi_hi_206, dataGroup_hi_lo_206};
  wire [7:0]    dataGroup_14_6 = dataGroup_lo_206[455:448];
  wire [1023:0] dataGroup_lo_207 = {dataGroup_lo_hi_207, dataGroup_lo_lo_207};
  wire [1023:0] dataGroup_hi_207 = {dataGroup_hi_hi_207, dataGroup_hi_lo_207};
  wire [7:0]    dataGroup_15_6 = dataGroup_lo_207[487:480];
  wire [1023:0] dataGroup_lo_208 = {dataGroup_lo_hi_208, dataGroup_lo_lo_208};
  wire [1023:0] dataGroup_hi_208 = {dataGroup_hi_hi_208, dataGroup_hi_lo_208};
  wire [7:0]    dataGroup_16_6 = dataGroup_lo_208[519:512];
  wire [1023:0] dataGroup_lo_209 = {dataGroup_lo_hi_209, dataGroup_lo_lo_209};
  wire [1023:0] dataGroup_hi_209 = {dataGroup_hi_hi_209, dataGroup_hi_lo_209};
  wire [7:0]    dataGroup_17_6 = dataGroup_lo_209[551:544];
  wire [1023:0] dataGroup_lo_210 = {dataGroup_lo_hi_210, dataGroup_lo_lo_210};
  wire [1023:0] dataGroup_hi_210 = {dataGroup_hi_hi_210, dataGroup_hi_lo_210};
  wire [7:0]    dataGroup_18_6 = dataGroup_lo_210[583:576];
  wire [1023:0] dataGroup_lo_211 = {dataGroup_lo_hi_211, dataGroup_lo_lo_211};
  wire [1023:0] dataGroup_hi_211 = {dataGroup_hi_hi_211, dataGroup_hi_lo_211};
  wire [7:0]    dataGroup_19_6 = dataGroup_lo_211[615:608];
  wire [1023:0] dataGroup_lo_212 = {dataGroup_lo_hi_212, dataGroup_lo_lo_212};
  wire [1023:0] dataGroup_hi_212 = {dataGroup_hi_hi_212, dataGroup_hi_lo_212};
  wire [7:0]    dataGroup_20_6 = dataGroup_lo_212[647:640];
  wire [1023:0] dataGroup_lo_213 = {dataGroup_lo_hi_213, dataGroup_lo_lo_213};
  wire [1023:0] dataGroup_hi_213 = {dataGroup_hi_hi_213, dataGroup_hi_lo_213};
  wire [7:0]    dataGroup_21_6 = dataGroup_lo_213[679:672];
  wire [1023:0] dataGroup_lo_214 = {dataGroup_lo_hi_214, dataGroup_lo_lo_214};
  wire [1023:0] dataGroup_hi_214 = {dataGroup_hi_hi_214, dataGroup_hi_lo_214};
  wire [7:0]    dataGroup_22_6 = dataGroup_lo_214[711:704];
  wire [1023:0] dataGroup_lo_215 = {dataGroup_lo_hi_215, dataGroup_lo_lo_215};
  wire [1023:0] dataGroup_hi_215 = {dataGroup_hi_hi_215, dataGroup_hi_lo_215};
  wire [7:0]    dataGroup_23_6 = dataGroup_lo_215[743:736];
  wire [1023:0] dataGroup_lo_216 = {dataGroup_lo_hi_216, dataGroup_lo_lo_216};
  wire [1023:0] dataGroup_hi_216 = {dataGroup_hi_hi_216, dataGroup_hi_lo_216};
  wire [7:0]    dataGroup_24_6 = dataGroup_lo_216[775:768];
  wire [1023:0] dataGroup_lo_217 = {dataGroup_lo_hi_217, dataGroup_lo_lo_217};
  wire [1023:0] dataGroup_hi_217 = {dataGroup_hi_hi_217, dataGroup_hi_lo_217};
  wire [7:0]    dataGroup_25_6 = dataGroup_lo_217[807:800];
  wire [1023:0] dataGroup_lo_218 = {dataGroup_lo_hi_218, dataGroup_lo_lo_218};
  wire [1023:0] dataGroup_hi_218 = {dataGroup_hi_hi_218, dataGroup_hi_lo_218};
  wire [7:0]    dataGroup_26_6 = dataGroup_lo_218[839:832];
  wire [1023:0] dataGroup_lo_219 = {dataGroup_lo_hi_219, dataGroup_lo_lo_219};
  wire [1023:0] dataGroup_hi_219 = {dataGroup_hi_hi_219, dataGroup_hi_lo_219};
  wire [7:0]    dataGroup_27_6 = dataGroup_lo_219[871:864];
  wire [1023:0] dataGroup_lo_220 = {dataGroup_lo_hi_220, dataGroup_lo_lo_220};
  wire [1023:0] dataGroup_hi_220 = {dataGroup_hi_hi_220, dataGroup_hi_lo_220};
  wire [7:0]    dataGroup_28_6 = dataGroup_lo_220[903:896];
  wire [1023:0] dataGroup_lo_221 = {dataGroup_lo_hi_221, dataGroup_lo_lo_221};
  wire [1023:0] dataGroup_hi_221 = {dataGroup_hi_hi_221, dataGroup_hi_lo_221};
  wire [7:0]    dataGroup_29_6 = dataGroup_lo_221[935:928];
  wire [1023:0] dataGroup_lo_222 = {dataGroup_lo_hi_222, dataGroup_lo_lo_222};
  wire [1023:0] dataGroup_hi_222 = {dataGroup_hi_hi_222, dataGroup_hi_lo_222};
  wire [7:0]    dataGroup_30_6 = dataGroup_lo_222[967:960];
  wire [1023:0] dataGroup_lo_223 = {dataGroup_lo_hi_223, dataGroup_lo_lo_223};
  wire [1023:0] dataGroup_hi_223 = {dataGroup_hi_hi_223, dataGroup_hi_lo_223};
  wire [7:0]    dataGroup_31_6 = dataGroup_lo_223[999:992];
  wire [15:0]   res_lo_lo_lo_lo_6 = {dataGroup_1_6, dataGroup_0_6};
  wire [15:0]   res_lo_lo_lo_hi_6 = {dataGroup_3_6, dataGroup_2_6};
  wire [31:0]   res_lo_lo_lo_6 = {res_lo_lo_lo_hi_6, res_lo_lo_lo_lo_6};
  wire [15:0]   res_lo_lo_hi_lo_6 = {dataGroup_5_6, dataGroup_4_6};
  wire [15:0]   res_lo_lo_hi_hi_6 = {dataGroup_7_6, dataGroup_6_6};
  wire [31:0]   res_lo_lo_hi_6 = {res_lo_lo_hi_hi_6, res_lo_lo_hi_lo_6};
  wire [63:0]   res_lo_lo_6 = {res_lo_lo_hi_6, res_lo_lo_lo_6};
  wire [15:0]   res_lo_hi_lo_lo_6 = {dataGroup_9_6, dataGroup_8_6};
  wire [15:0]   res_lo_hi_lo_hi_6 = {dataGroup_11_6, dataGroup_10_6};
  wire [31:0]   res_lo_hi_lo_6 = {res_lo_hi_lo_hi_6, res_lo_hi_lo_lo_6};
  wire [15:0]   res_lo_hi_hi_lo_6 = {dataGroup_13_6, dataGroup_12_6};
  wire [15:0]   res_lo_hi_hi_hi_6 = {dataGroup_15_6, dataGroup_14_6};
  wire [31:0]   res_lo_hi_hi_6 = {res_lo_hi_hi_hi_6, res_lo_hi_hi_lo_6};
  wire [63:0]   res_lo_hi_6 = {res_lo_hi_hi_6, res_lo_hi_lo_6};
  wire [127:0]  res_lo_6 = {res_lo_hi_6, res_lo_lo_6};
  wire [15:0]   res_hi_lo_lo_lo_6 = {dataGroup_17_6, dataGroup_16_6};
  wire [15:0]   res_hi_lo_lo_hi_6 = {dataGroup_19_6, dataGroup_18_6};
  wire [31:0]   res_hi_lo_lo_6 = {res_hi_lo_lo_hi_6, res_hi_lo_lo_lo_6};
  wire [15:0]   res_hi_lo_hi_lo_6 = {dataGroup_21_6, dataGroup_20_6};
  wire [15:0]   res_hi_lo_hi_hi_6 = {dataGroup_23_6, dataGroup_22_6};
  wire [31:0]   res_hi_lo_hi_6 = {res_hi_lo_hi_hi_6, res_hi_lo_hi_lo_6};
  wire [63:0]   res_hi_lo_6 = {res_hi_lo_hi_6, res_hi_lo_lo_6};
  wire [15:0]   res_hi_hi_lo_lo_6 = {dataGroup_25_6, dataGroup_24_6};
  wire [15:0]   res_hi_hi_lo_hi_6 = {dataGroup_27_6, dataGroup_26_6};
  wire [31:0]   res_hi_hi_lo_6 = {res_hi_hi_lo_hi_6, res_hi_hi_lo_lo_6};
  wire [15:0]   res_hi_hi_hi_lo_6 = {dataGroup_29_6, dataGroup_28_6};
  wire [15:0]   res_hi_hi_hi_hi_6 = {dataGroup_31_6, dataGroup_30_6};
  wire [31:0]   res_hi_hi_hi_6 = {res_hi_hi_hi_hi_6, res_hi_hi_hi_lo_6};
  wire [63:0]   res_hi_hi_6 = {res_hi_hi_hi_6, res_hi_hi_lo_6};
  wire [127:0]  res_hi_6 = {res_hi_hi_6, res_hi_lo_6};
  wire [255:0]  res_24 = {res_hi_6, res_lo_6};
  wire [1023:0] dataGroup_lo_224 = {dataGroup_lo_hi_224, dataGroup_lo_lo_224};
  wire [1023:0] dataGroup_hi_224 = {dataGroup_hi_hi_224, dataGroup_hi_lo_224};
  wire [7:0]    dataGroup_0_7 = dataGroup_lo_224[15:8];
  wire [1023:0] dataGroup_lo_225 = {dataGroup_lo_hi_225, dataGroup_lo_lo_225};
  wire [1023:0] dataGroup_hi_225 = {dataGroup_hi_hi_225, dataGroup_hi_lo_225};
  wire [7:0]    dataGroup_1_7 = dataGroup_lo_225[47:40];
  wire [1023:0] dataGroup_lo_226 = {dataGroup_lo_hi_226, dataGroup_lo_lo_226};
  wire [1023:0] dataGroup_hi_226 = {dataGroup_hi_hi_226, dataGroup_hi_lo_226};
  wire [7:0]    dataGroup_2_7 = dataGroup_lo_226[79:72];
  wire [1023:0] dataGroup_lo_227 = {dataGroup_lo_hi_227, dataGroup_lo_lo_227};
  wire [1023:0] dataGroup_hi_227 = {dataGroup_hi_hi_227, dataGroup_hi_lo_227};
  wire [7:0]    dataGroup_3_7 = dataGroup_lo_227[111:104];
  wire [1023:0] dataGroup_lo_228 = {dataGroup_lo_hi_228, dataGroup_lo_lo_228};
  wire [1023:0] dataGroup_hi_228 = {dataGroup_hi_hi_228, dataGroup_hi_lo_228};
  wire [7:0]    dataGroup_4_7 = dataGroup_lo_228[143:136];
  wire [1023:0] dataGroup_lo_229 = {dataGroup_lo_hi_229, dataGroup_lo_lo_229};
  wire [1023:0] dataGroup_hi_229 = {dataGroup_hi_hi_229, dataGroup_hi_lo_229};
  wire [7:0]    dataGroup_5_7 = dataGroup_lo_229[175:168];
  wire [1023:0] dataGroup_lo_230 = {dataGroup_lo_hi_230, dataGroup_lo_lo_230};
  wire [1023:0] dataGroup_hi_230 = {dataGroup_hi_hi_230, dataGroup_hi_lo_230};
  wire [7:0]    dataGroup_6_7 = dataGroup_lo_230[207:200];
  wire [1023:0] dataGroup_lo_231 = {dataGroup_lo_hi_231, dataGroup_lo_lo_231};
  wire [1023:0] dataGroup_hi_231 = {dataGroup_hi_hi_231, dataGroup_hi_lo_231};
  wire [7:0]    dataGroup_7_7 = dataGroup_lo_231[239:232];
  wire [1023:0] dataGroup_lo_232 = {dataGroup_lo_hi_232, dataGroup_lo_lo_232};
  wire [1023:0] dataGroup_hi_232 = {dataGroup_hi_hi_232, dataGroup_hi_lo_232};
  wire [7:0]    dataGroup_8_7 = dataGroup_lo_232[271:264];
  wire [1023:0] dataGroup_lo_233 = {dataGroup_lo_hi_233, dataGroup_lo_lo_233};
  wire [1023:0] dataGroup_hi_233 = {dataGroup_hi_hi_233, dataGroup_hi_lo_233};
  wire [7:0]    dataGroup_9_7 = dataGroup_lo_233[303:296];
  wire [1023:0] dataGroup_lo_234 = {dataGroup_lo_hi_234, dataGroup_lo_lo_234};
  wire [1023:0] dataGroup_hi_234 = {dataGroup_hi_hi_234, dataGroup_hi_lo_234};
  wire [7:0]    dataGroup_10_7 = dataGroup_lo_234[335:328];
  wire [1023:0] dataGroup_lo_235 = {dataGroup_lo_hi_235, dataGroup_lo_lo_235};
  wire [1023:0] dataGroup_hi_235 = {dataGroup_hi_hi_235, dataGroup_hi_lo_235};
  wire [7:0]    dataGroup_11_7 = dataGroup_lo_235[367:360];
  wire [1023:0] dataGroup_lo_236 = {dataGroup_lo_hi_236, dataGroup_lo_lo_236};
  wire [1023:0] dataGroup_hi_236 = {dataGroup_hi_hi_236, dataGroup_hi_lo_236};
  wire [7:0]    dataGroup_12_7 = dataGroup_lo_236[399:392];
  wire [1023:0] dataGroup_lo_237 = {dataGroup_lo_hi_237, dataGroup_lo_lo_237};
  wire [1023:0] dataGroup_hi_237 = {dataGroup_hi_hi_237, dataGroup_hi_lo_237};
  wire [7:0]    dataGroup_13_7 = dataGroup_lo_237[431:424];
  wire [1023:0] dataGroup_lo_238 = {dataGroup_lo_hi_238, dataGroup_lo_lo_238};
  wire [1023:0] dataGroup_hi_238 = {dataGroup_hi_hi_238, dataGroup_hi_lo_238};
  wire [7:0]    dataGroup_14_7 = dataGroup_lo_238[463:456];
  wire [1023:0] dataGroup_lo_239 = {dataGroup_lo_hi_239, dataGroup_lo_lo_239};
  wire [1023:0] dataGroup_hi_239 = {dataGroup_hi_hi_239, dataGroup_hi_lo_239};
  wire [7:0]    dataGroup_15_7 = dataGroup_lo_239[495:488];
  wire [1023:0] dataGroup_lo_240 = {dataGroup_lo_hi_240, dataGroup_lo_lo_240};
  wire [1023:0] dataGroup_hi_240 = {dataGroup_hi_hi_240, dataGroup_hi_lo_240};
  wire [7:0]    dataGroup_16_7 = dataGroup_lo_240[527:520];
  wire [1023:0] dataGroup_lo_241 = {dataGroup_lo_hi_241, dataGroup_lo_lo_241};
  wire [1023:0] dataGroup_hi_241 = {dataGroup_hi_hi_241, dataGroup_hi_lo_241};
  wire [7:0]    dataGroup_17_7 = dataGroup_lo_241[559:552];
  wire [1023:0] dataGroup_lo_242 = {dataGroup_lo_hi_242, dataGroup_lo_lo_242};
  wire [1023:0] dataGroup_hi_242 = {dataGroup_hi_hi_242, dataGroup_hi_lo_242};
  wire [7:0]    dataGroup_18_7 = dataGroup_lo_242[591:584];
  wire [1023:0] dataGroup_lo_243 = {dataGroup_lo_hi_243, dataGroup_lo_lo_243};
  wire [1023:0] dataGroup_hi_243 = {dataGroup_hi_hi_243, dataGroup_hi_lo_243};
  wire [7:0]    dataGroup_19_7 = dataGroup_lo_243[623:616];
  wire [1023:0] dataGroup_lo_244 = {dataGroup_lo_hi_244, dataGroup_lo_lo_244};
  wire [1023:0] dataGroup_hi_244 = {dataGroup_hi_hi_244, dataGroup_hi_lo_244};
  wire [7:0]    dataGroup_20_7 = dataGroup_lo_244[655:648];
  wire [1023:0] dataGroup_lo_245 = {dataGroup_lo_hi_245, dataGroup_lo_lo_245};
  wire [1023:0] dataGroup_hi_245 = {dataGroup_hi_hi_245, dataGroup_hi_lo_245};
  wire [7:0]    dataGroup_21_7 = dataGroup_lo_245[687:680];
  wire [1023:0] dataGroup_lo_246 = {dataGroup_lo_hi_246, dataGroup_lo_lo_246};
  wire [1023:0] dataGroup_hi_246 = {dataGroup_hi_hi_246, dataGroup_hi_lo_246};
  wire [7:0]    dataGroup_22_7 = dataGroup_lo_246[719:712];
  wire [1023:0] dataGroup_lo_247 = {dataGroup_lo_hi_247, dataGroup_lo_lo_247};
  wire [1023:0] dataGroup_hi_247 = {dataGroup_hi_hi_247, dataGroup_hi_lo_247};
  wire [7:0]    dataGroup_23_7 = dataGroup_lo_247[751:744];
  wire [1023:0] dataGroup_lo_248 = {dataGroup_lo_hi_248, dataGroup_lo_lo_248};
  wire [1023:0] dataGroup_hi_248 = {dataGroup_hi_hi_248, dataGroup_hi_lo_248};
  wire [7:0]    dataGroup_24_7 = dataGroup_lo_248[783:776];
  wire [1023:0] dataGroup_lo_249 = {dataGroup_lo_hi_249, dataGroup_lo_lo_249};
  wire [1023:0] dataGroup_hi_249 = {dataGroup_hi_hi_249, dataGroup_hi_lo_249};
  wire [7:0]    dataGroup_25_7 = dataGroup_lo_249[815:808];
  wire [1023:0] dataGroup_lo_250 = {dataGroup_lo_hi_250, dataGroup_lo_lo_250};
  wire [1023:0] dataGroup_hi_250 = {dataGroup_hi_hi_250, dataGroup_hi_lo_250};
  wire [7:0]    dataGroup_26_7 = dataGroup_lo_250[847:840];
  wire [1023:0] dataGroup_lo_251 = {dataGroup_lo_hi_251, dataGroup_lo_lo_251};
  wire [1023:0] dataGroup_hi_251 = {dataGroup_hi_hi_251, dataGroup_hi_lo_251};
  wire [7:0]    dataGroup_27_7 = dataGroup_lo_251[879:872];
  wire [1023:0] dataGroup_lo_252 = {dataGroup_lo_hi_252, dataGroup_lo_lo_252};
  wire [1023:0] dataGroup_hi_252 = {dataGroup_hi_hi_252, dataGroup_hi_lo_252};
  wire [7:0]    dataGroup_28_7 = dataGroup_lo_252[911:904];
  wire [1023:0] dataGroup_lo_253 = {dataGroup_lo_hi_253, dataGroup_lo_lo_253};
  wire [1023:0] dataGroup_hi_253 = {dataGroup_hi_hi_253, dataGroup_hi_lo_253};
  wire [7:0]    dataGroup_29_7 = dataGroup_lo_253[943:936];
  wire [1023:0] dataGroup_lo_254 = {dataGroup_lo_hi_254, dataGroup_lo_lo_254};
  wire [1023:0] dataGroup_hi_254 = {dataGroup_hi_hi_254, dataGroup_hi_lo_254};
  wire [7:0]    dataGroup_30_7 = dataGroup_lo_254[975:968];
  wire [1023:0] dataGroup_lo_255 = {dataGroup_lo_hi_255, dataGroup_lo_lo_255};
  wire [1023:0] dataGroup_hi_255 = {dataGroup_hi_hi_255, dataGroup_hi_lo_255};
  wire [7:0]    dataGroup_31_7 = dataGroup_lo_255[1007:1000];
  wire [15:0]   res_lo_lo_lo_lo_7 = {dataGroup_1_7, dataGroup_0_7};
  wire [15:0]   res_lo_lo_lo_hi_7 = {dataGroup_3_7, dataGroup_2_7};
  wire [31:0]   res_lo_lo_lo_7 = {res_lo_lo_lo_hi_7, res_lo_lo_lo_lo_7};
  wire [15:0]   res_lo_lo_hi_lo_7 = {dataGroup_5_7, dataGroup_4_7};
  wire [15:0]   res_lo_lo_hi_hi_7 = {dataGroup_7_7, dataGroup_6_7};
  wire [31:0]   res_lo_lo_hi_7 = {res_lo_lo_hi_hi_7, res_lo_lo_hi_lo_7};
  wire [63:0]   res_lo_lo_7 = {res_lo_lo_hi_7, res_lo_lo_lo_7};
  wire [15:0]   res_lo_hi_lo_lo_7 = {dataGroup_9_7, dataGroup_8_7};
  wire [15:0]   res_lo_hi_lo_hi_7 = {dataGroup_11_7, dataGroup_10_7};
  wire [31:0]   res_lo_hi_lo_7 = {res_lo_hi_lo_hi_7, res_lo_hi_lo_lo_7};
  wire [15:0]   res_lo_hi_hi_lo_7 = {dataGroup_13_7, dataGroup_12_7};
  wire [15:0]   res_lo_hi_hi_hi_7 = {dataGroup_15_7, dataGroup_14_7};
  wire [31:0]   res_lo_hi_hi_7 = {res_lo_hi_hi_hi_7, res_lo_hi_hi_lo_7};
  wire [63:0]   res_lo_hi_7 = {res_lo_hi_hi_7, res_lo_hi_lo_7};
  wire [127:0]  res_lo_7 = {res_lo_hi_7, res_lo_lo_7};
  wire [15:0]   res_hi_lo_lo_lo_7 = {dataGroup_17_7, dataGroup_16_7};
  wire [15:0]   res_hi_lo_lo_hi_7 = {dataGroup_19_7, dataGroup_18_7};
  wire [31:0]   res_hi_lo_lo_7 = {res_hi_lo_lo_hi_7, res_hi_lo_lo_lo_7};
  wire [15:0]   res_hi_lo_hi_lo_7 = {dataGroup_21_7, dataGroup_20_7};
  wire [15:0]   res_hi_lo_hi_hi_7 = {dataGroup_23_7, dataGroup_22_7};
  wire [31:0]   res_hi_lo_hi_7 = {res_hi_lo_hi_hi_7, res_hi_lo_hi_lo_7};
  wire [63:0]   res_hi_lo_7 = {res_hi_lo_hi_7, res_hi_lo_lo_7};
  wire [15:0]   res_hi_hi_lo_lo_7 = {dataGroup_25_7, dataGroup_24_7};
  wire [15:0]   res_hi_hi_lo_hi_7 = {dataGroup_27_7, dataGroup_26_7};
  wire [31:0]   res_hi_hi_lo_7 = {res_hi_hi_lo_hi_7, res_hi_hi_lo_lo_7};
  wire [15:0]   res_hi_hi_hi_lo_7 = {dataGroup_29_7, dataGroup_28_7};
  wire [15:0]   res_hi_hi_hi_hi_7 = {dataGroup_31_7, dataGroup_30_7};
  wire [31:0]   res_hi_hi_hi_7 = {res_hi_hi_hi_hi_7, res_hi_hi_hi_lo_7};
  wire [63:0]   res_hi_hi_7 = {res_hi_hi_hi_7, res_hi_hi_lo_7};
  wire [127:0]  res_hi_7 = {res_hi_hi_7, res_hi_lo_7};
  wire [255:0]  res_25 = {res_hi_7, res_lo_7};
  wire [1023:0] dataGroup_lo_256 = {dataGroup_lo_hi_256, dataGroup_lo_lo_256};
  wire [1023:0] dataGroup_hi_256 = {dataGroup_hi_hi_256, dataGroup_hi_lo_256};
  wire [7:0]    dataGroup_0_8 = dataGroup_lo_256[23:16];
  wire [1023:0] dataGroup_lo_257 = {dataGroup_lo_hi_257, dataGroup_lo_lo_257};
  wire [1023:0] dataGroup_hi_257 = {dataGroup_hi_hi_257, dataGroup_hi_lo_257};
  wire [7:0]    dataGroup_1_8 = dataGroup_lo_257[55:48];
  wire [1023:0] dataGroup_lo_258 = {dataGroup_lo_hi_258, dataGroup_lo_lo_258};
  wire [1023:0] dataGroup_hi_258 = {dataGroup_hi_hi_258, dataGroup_hi_lo_258};
  wire [7:0]    dataGroup_2_8 = dataGroup_lo_258[87:80];
  wire [1023:0] dataGroup_lo_259 = {dataGroup_lo_hi_259, dataGroup_lo_lo_259};
  wire [1023:0] dataGroup_hi_259 = {dataGroup_hi_hi_259, dataGroup_hi_lo_259};
  wire [7:0]    dataGroup_3_8 = dataGroup_lo_259[119:112];
  wire [1023:0] dataGroup_lo_260 = {dataGroup_lo_hi_260, dataGroup_lo_lo_260};
  wire [1023:0] dataGroup_hi_260 = {dataGroup_hi_hi_260, dataGroup_hi_lo_260};
  wire [7:0]    dataGroup_4_8 = dataGroup_lo_260[151:144];
  wire [1023:0] dataGroup_lo_261 = {dataGroup_lo_hi_261, dataGroup_lo_lo_261};
  wire [1023:0] dataGroup_hi_261 = {dataGroup_hi_hi_261, dataGroup_hi_lo_261};
  wire [7:0]    dataGroup_5_8 = dataGroup_lo_261[183:176];
  wire [1023:0] dataGroup_lo_262 = {dataGroup_lo_hi_262, dataGroup_lo_lo_262};
  wire [1023:0] dataGroup_hi_262 = {dataGroup_hi_hi_262, dataGroup_hi_lo_262};
  wire [7:0]    dataGroup_6_8 = dataGroup_lo_262[215:208];
  wire [1023:0] dataGroup_lo_263 = {dataGroup_lo_hi_263, dataGroup_lo_lo_263};
  wire [1023:0] dataGroup_hi_263 = {dataGroup_hi_hi_263, dataGroup_hi_lo_263};
  wire [7:0]    dataGroup_7_8 = dataGroup_lo_263[247:240];
  wire [1023:0] dataGroup_lo_264 = {dataGroup_lo_hi_264, dataGroup_lo_lo_264};
  wire [1023:0] dataGroup_hi_264 = {dataGroup_hi_hi_264, dataGroup_hi_lo_264};
  wire [7:0]    dataGroup_8_8 = dataGroup_lo_264[279:272];
  wire [1023:0] dataGroup_lo_265 = {dataGroup_lo_hi_265, dataGroup_lo_lo_265};
  wire [1023:0] dataGroup_hi_265 = {dataGroup_hi_hi_265, dataGroup_hi_lo_265};
  wire [7:0]    dataGroup_9_8 = dataGroup_lo_265[311:304];
  wire [1023:0] dataGroup_lo_266 = {dataGroup_lo_hi_266, dataGroup_lo_lo_266};
  wire [1023:0] dataGroup_hi_266 = {dataGroup_hi_hi_266, dataGroup_hi_lo_266};
  wire [7:0]    dataGroup_10_8 = dataGroup_lo_266[343:336];
  wire [1023:0] dataGroup_lo_267 = {dataGroup_lo_hi_267, dataGroup_lo_lo_267};
  wire [1023:0] dataGroup_hi_267 = {dataGroup_hi_hi_267, dataGroup_hi_lo_267};
  wire [7:0]    dataGroup_11_8 = dataGroup_lo_267[375:368];
  wire [1023:0] dataGroup_lo_268 = {dataGroup_lo_hi_268, dataGroup_lo_lo_268};
  wire [1023:0] dataGroup_hi_268 = {dataGroup_hi_hi_268, dataGroup_hi_lo_268};
  wire [7:0]    dataGroup_12_8 = dataGroup_lo_268[407:400];
  wire [1023:0] dataGroup_lo_269 = {dataGroup_lo_hi_269, dataGroup_lo_lo_269};
  wire [1023:0] dataGroup_hi_269 = {dataGroup_hi_hi_269, dataGroup_hi_lo_269};
  wire [7:0]    dataGroup_13_8 = dataGroup_lo_269[439:432];
  wire [1023:0] dataGroup_lo_270 = {dataGroup_lo_hi_270, dataGroup_lo_lo_270};
  wire [1023:0] dataGroup_hi_270 = {dataGroup_hi_hi_270, dataGroup_hi_lo_270};
  wire [7:0]    dataGroup_14_8 = dataGroup_lo_270[471:464];
  wire [1023:0] dataGroup_lo_271 = {dataGroup_lo_hi_271, dataGroup_lo_lo_271};
  wire [1023:0] dataGroup_hi_271 = {dataGroup_hi_hi_271, dataGroup_hi_lo_271};
  wire [7:0]    dataGroup_15_8 = dataGroup_lo_271[503:496];
  wire [1023:0] dataGroup_lo_272 = {dataGroup_lo_hi_272, dataGroup_lo_lo_272};
  wire [1023:0] dataGroup_hi_272 = {dataGroup_hi_hi_272, dataGroup_hi_lo_272};
  wire [7:0]    dataGroup_16_8 = dataGroup_lo_272[535:528];
  wire [1023:0] dataGroup_lo_273 = {dataGroup_lo_hi_273, dataGroup_lo_lo_273};
  wire [1023:0] dataGroup_hi_273 = {dataGroup_hi_hi_273, dataGroup_hi_lo_273};
  wire [7:0]    dataGroup_17_8 = dataGroup_lo_273[567:560];
  wire [1023:0] dataGroup_lo_274 = {dataGroup_lo_hi_274, dataGroup_lo_lo_274};
  wire [1023:0] dataGroup_hi_274 = {dataGroup_hi_hi_274, dataGroup_hi_lo_274};
  wire [7:0]    dataGroup_18_8 = dataGroup_lo_274[599:592];
  wire [1023:0] dataGroup_lo_275 = {dataGroup_lo_hi_275, dataGroup_lo_lo_275};
  wire [1023:0] dataGroup_hi_275 = {dataGroup_hi_hi_275, dataGroup_hi_lo_275};
  wire [7:0]    dataGroup_19_8 = dataGroup_lo_275[631:624];
  wire [1023:0] dataGroup_lo_276 = {dataGroup_lo_hi_276, dataGroup_lo_lo_276};
  wire [1023:0] dataGroup_hi_276 = {dataGroup_hi_hi_276, dataGroup_hi_lo_276};
  wire [7:0]    dataGroup_20_8 = dataGroup_lo_276[663:656];
  wire [1023:0] dataGroup_lo_277 = {dataGroup_lo_hi_277, dataGroup_lo_lo_277};
  wire [1023:0] dataGroup_hi_277 = {dataGroup_hi_hi_277, dataGroup_hi_lo_277};
  wire [7:0]    dataGroup_21_8 = dataGroup_lo_277[695:688];
  wire [1023:0] dataGroup_lo_278 = {dataGroup_lo_hi_278, dataGroup_lo_lo_278};
  wire [1023:0] dataGroup_hi_278 = {dataGroup_hi_hi_278, dataGroup_hi_lo_278};
  wire [7:0]    dataGroup_22_8 = dataGroup_lo_278[727:720];
  wire [1023:0] dataGroup_lo_279 = {dataGroup_lo_hi_279, dataGroup_lo_lo_279};
  wire [1023:0] dataGroup_hi_279 = {dataGroup_hi_hi_279, dataGroup_hi_lo_279};
  wire [7:0]    dataGroup_23_8 = dataGroup_lo_279[759:752];
  wire [1023:0] dataGroup_lo_280 = {dataGroup_lo_hi_280, dataGroup_lo_lo_280};
  wire [1023:0] dataGroup_hi_280 = {dataGroup_hi_hi_280, dataGroup_hi_lo_280};
  wire [7:0]    dataGroup_24_8 = dataGroup_lo_280[791:784];
  wire [1023:0] dataGroup_lo_281 = {dataGroup_lo_hi_281, dataGroup_lo_lo_281};
  wire [1023:0] dataGroup_hi_281 = {dataGroup_hi_hi_281, dataGroup_hi_lo_281};
  wire [7:0]    dataGroup_25_8 = dataGroup_lo_281[823:816];
  wire [1023:0] dataGroup_lo_282 = {dataGroup_lo_hi_282, dataGroup_lo_lo_282};
  wire [1023:0] dataGroup_hi_282 = {dataGroup_hi_hi_282, dataGroup_hi_lo_282};
  wire [7:0]    dataGroup_26_8 = dataGroup_lo_282[855:848];
  wire [1023:0] dataGroup_lo_283 = {dataGroup_lo_hi_283, dataGroup_lo_lo_283};
  wire [1023:0] dataGroup_hi_283 = {dataGroup_hi_hi_283, dataGroup_hi_lo_283};
  wire [7:0]    dataGroup_27_8 = dataGroup_lo_283[887:880];
  wire [1023:0] dataGroup_lo_284 = {dataGroup_lo_hi_284, dataGroup_lo_lo_284};
  wire [1023:0] dataGroup_hi_284 = {dataGroup_hi_hi_284, dataGroup_hi_lo_284};
  wire [7:0]    dataGroup_28_8 = dataGroup_lo_284[919:912];
  wire [1023:0] dataGroup_lo_285 = {dataGroup_lo_hi_285, dataGroup_lo_lo_285};
  wire [1023:0] dataGroup_hi_285 = {dataGroup_hi_hi_285, dataGroup_hi_lo_285};
  wire [7:0]    dataGroup_29_8 = dataGroup_lo_285[951:944];
  wire [1023:0] dataGroup_lo_286 = {dataGroup_lo_hi_286, dataGroup_lo_lo_286};
  wire [1023:0] dataGroup_hi_286 = {dataGroup_hi_hi_286, dataGroup_hi_lo_286};
  wire [7:0]    dataGroup_30_8 = dataGroup_lo_286[983:976];
  wire [1023:0] dataGroup_lo_287 = {dataGroup_lo_hi_287, dataGroup_lo_lo_287};
  wire [1023:0] dataGroup_hi_287 = {dataGroup_hi_hi_287, dataGroup_hi_lo_287};
  wire [7:0]    dataGroup_31_8 = dataGroup_lo_287[1015:1008];
  wire [15:0]   res_lo_lo_lo_lo_8 = {dataGroup_1_8, dataGroup_0_8};
  wire [15:0]   res_lo_lo_lo_hi_8 = {dataGroup_3_8, dataGroup_2_8};
  wire [31:0]   res_lo_lo_lo_8 = {res_lo_lo_lo_hi_8, res_lo_lo_lo_lo_8};
  wire [15:0]   res_lo_lo_hi_lo_8 = {dataGroup_5_8, dataGroup_4_8};
  wire [15:0]   res_lo_lo_hi_hi_8 = {dataGroup_7_8, dataGroup_6_8};
  wire [31:0]   res_lo_lo_hi_8 = {res_lo_lo_hi_hi_8, res_lo_lo_hi_lo_8};
  wire [63:0]   res_lo_lo_8 = {res_lo_lo_hi_8, res_lo_lo_lo_8};
  wire [15:0]   res_lo_hi_lo_lo_8 = {dataGroup_9_8, dataGroup_8_8};
  wire [15:0]   res_lo_hi_lo_hi_8 = {dataGroup_11_8, dataGroup_10_8};
  wire [31:0]   res_lo_hi_lo_8 = {res_lo_hi_lo_hi_8, res_lo_hi_lo_lo_8};
  wire [15:0]   res_lo_hi_hi_lo_8 = {dataGroup_13_8, dataGroup_12_8};
  wire [15:0]   res_lo_hi_hi_hi_8 = {dataGroup_15_8, dataGroup_14_8};
  wire [31:0]   res_lo_hi_hi_8 = {res_lo_hi_hi_hi_8, res_lo_hi_hi_lo_8};
  wire [63:0]   res_lo_hi_8 = {res_lo_hi_hi_8, res_lo_hi_lo_8};
  wire [127:0]  res_lo_8 = {res_lo_hi_8, res_lo_lo_8};
  wire [15:0]   res_hi_lo_lo_lo_8 = {dataGroup_17_8, dataGroup_16_8};
  wire [15:0]   res_hi_lo_lo_hi_8 = {dataGroup_19_8, dataGroup_18_8};
  wire [31:0]   res_hi_lo_lo_8 = {res_hi_lo_lo_hi_8, res_hi_lo_lo_lo_8};
  wire [15:0]   res_hi_lo_hi_lo_8 = {dataGroup_21_8, dataGroup_20_8};
  wire [15:0]   res_hi_lo_hi_hi_8 = {dataGroup_23_8, dataGroup_22_8};
  wire [31:0]   res_hi_lo_hi_8 = {res_hi_lo_hi_hi_8, res_hi_lo_hi_lo_8};
  wire [63:0]   res_hi_lo_8 = {res_hi_lo_hi_8, res_hi_lo_lo_8};
  wire [15:0]   res_hi_hi_lo_lo_8 = {dataGroup_25_8, dataGroup_24_8};
  wire [15:0]   res_hi_hi_lo_hi_8 = {dataGroup_27_8, dataGroup_26_8};
  wire [31:0]   res_hi_hi_lo_8 = {res_hi_hi_lo_hi_8, res_hi_hi_lo_lo_8};
  wire [15:0]   res_hi_hi_hi_lo_8 = {dataGroup_29_8, dataGroup_28_8};
  wire [15:0]   res_hi_hi_hi_hi_8 = {dataGroup_31_8, dataGroup_30_8};
  wire [31:0]   res_hi_hi_hi_8 = {res_hi_hi_hi_hi_8, res_hi_hi_hi_lo_8};
  wire [63:0]   res_hi_hi_8 = {res_hi_hi_hi_8, res_hi_hi_lo_8};
  wire [127:0]  res_hi_8 = {res_hi_hi_8, res_hi_lo_8};
  wire [255:0]  res_26 = {res_hi_8, res_lo_8};
  wire [1023:0] dataGroup_lo_288 = {dataGroup_lo_hi_288, dataGroup_lo_lo_288};
  wire [1023:0] dataGroup_hi_288 = {dataGroup_hi_hi_288, dataGroup_hi_lo_288};
  wire [7:0]    dataGroup_0_9 = dataGroup_lo_288[31:24];
  wire [1023:0] dataGroup_lo_289 = {dataGroup_lo_hi_289, dataGroup_lo_lo_289};
  wire [1023:0] dataGroup_hi_289 = {dataGroup_hi_hi_289, dataGroup_hi_lo_289};
  wire [7:0]    dataGroup_1_9 = dataGroup_lo_289[63:56];
  wire [1023:0] dataGroup_lo_290 = {dataGroup_lo_hi_290, dataGroup_lo_lo_290};
  wire [1023:0] dataGroup_hi_290 = {dataGroup_hi_hi_290, dataGroup_hi_lo_290};
  wire [7:0]    dataGroup_2_9 = dataGroup_lo_290[95:88];
  wire [1023:0] dataGroup_lo_291 = {dataGroup_lo_hi_291, dataGroup_lo_lo_291};
  wire [1023:0] dataGroup_hi_291 = {dataGroup_hi_hi_291, dataGroup_hi_lo_291};
  wire [7:0]    dataGroup_3_9 = dataGroup_lo_291[127:120];
  wire [1023:0] dataGroup_lo_292 = {dataGroup_lo_hi_292, dataGroup_lo_lo_292};
  wire [1023:0] dataGroup_hi_292 = {dataGroup_hi_hi_292, dataGroup_hi_lo_292};
  wire [7:0]    dataGroup_4_9 = dataGroup_lo_292[159:152];
  wire [1023:0] dataGroup_lo_293 = {dataGroup_lo_hi_293, dataGroup_lo_lo_293};
  wire [1023:0] dataGroup_hi_293 = {dataGroup_hi_hi_293, dataGroup_hi_lo_293};
  wire [7:0]    dataGroup_5_9 = dataGroup_lo_293[191:184];
  wire [1023:0] dataGroup_lo_294 = {dataGroup_lo_hi_294, dataGroup_lo_lo_294};
  wire [1023:0] dataGroup_hi_294 = {dataGroup_hi_hi_294, dataGroup_hi_lo_294};
  wire [7:0]    dataGroup_6_9 = dataGroup_lo_294[223:216];
  wire [1023:0] dataGroup_lo_295 = {dataGroup_lo_hi_295, dataGroup_lo_lo_295};
  wire [1023:0] dataGroup_hi_295 = {dataGroup_hi_hi_295, dataGroup_hi_lo_295};
  wire [7:0]    dataGroup_7_9 = dataGroup_lo_295[255:248];
  wire [1023:0] dataGroup_lo_296 = {dataGroup_lo_hi_296, dataGroup_lo_lo_296};
  wire [1023:0] dataGroup_hi_296 = {dataGroup_hi_hi_296, dataGroup_hi_lo_296};
  wire [7:0]    dataGroup_8_9 = dataGroup_lo_296[287:280];
  wire [1023:0] dataGroup_lo_297 = {dataGroup_lo_hi_297, dataGroup_lo_lo_297};
  wire [1023:0] dataGroup_hi_297 = {dataGroup_hi_hi_297, dataGroup_hi_lo_297};
  wire [7:0]    dataGroup_9_9 = dataGroup_lo_297[319:312];
  wire [1023:0] dataGroup_lo_298 = {dataGroup_lo_hi_298, dataGroup_lo_lo_298};
  wire [1023:0] dataGroup_hi_298 = {dataGroup_hi_hi_298, dataGroup_hi_lo_298};
  wire [7:0]    dataGroup_10_9 = dataGroup_lo_298[351:344];
  wire [1023:0] dataGroup_lo_299 = {dataGroup_lo_hi_299, dataGroup_lo_lo_299};
  wire [1023:0] dataGroup_hi_299 = {dataGroup_hi_hi_299, dataGroup_hi_lo_299};
  wire [7:0]    dataGroup_11_9 = dataGroup_lo_299[383:376];
  wire [1023:0] dataGroup_lo_300 = {dataGroup_lo_hi_300, dataGroup_lo_lo_300};
  wire [1023:0] dataGroup_hi_300 = {dataGroup_hi_hi_300, dataGroup_hi_lo_300};
  wire [7:0]    dataGroup_12_9 = dataGroup_lo_300[415:408];
  wire [1023:0] dataGroup_lo_301 = {dataGroup_lo_hi_301, dataGroup_lo_lo_301};
  wire [1023:0] dataGroup_hi_301 = {dataGroup_hi_hi_301, dataGroup_hi_lo_301};
  wire [7:0]    dataGroup_13_9 = dataGroup_lo_301[447:440];
  wire [1023:0] dataGroup_lo_302 = {dataGroup_lo_hi_302, dataGroup_lo_lo_302};
  wire [1023:0] dataGroup_hi_302 = {dataGroup_hi_hi_302, dataGroup_hi_lo_302};
  wire [7:0]    dataGroup_14_9 = dataGroup_lo_302[479:472];
  wire [1023:0] dataGroup_lo_303 = {dataGroup_lo_hi_303, dataGroup_lo_lo_303};
  wire [1023:0] dataGroup_hi_303 = {dataGroup_hi_hi_303, dataGroup_hi_lo_303};
  wire [7:0]    dataGroup_15_9 = dataGroup_lo_303[511:504];
  wire [1023:0] dataGroup_lo_304 = {dataGroup_lo_hi_304, dataGroup_lo_lo_304};
  wire [1023:0] dataGroup_hi_304 = {dataGroup_hi_hi_304, dataGroup_hi_lo_304};
  wire [7:0]    dataGroup_16_9 = dataGroup_lo_304[543:536];
  wire [1023:0] dataGroup_lo_305 = {dataGroup_lo_hi_305, dataGroup_lo_lo_305};
  wire [1023:0] dataGroup_hi_305 = {dataGroup_hi_hi_305, dataGroup_hi_lo_305};
  wire [7:0]    dataGroup_17_9 = dataGroup_lo_305[575:568];
  wire [1023:0] dataGroup_lo_306 = {dataGroup_lo_hi_306, dataGroup_lo_lo_306};
  wire [1023:0] dataGroup_hi_306 = {dataGroup_hi_hi_306, dataGroup_hi_lo_306};
  wire [7:0]    dataGroup_18_9 = dataGroup_lo_306[607:600];
  wire [1023:0] dataGroup_lo_307 = {dataGroup_lo_hi_307, dataGroup_lo_lo_307};
  wire [1023:0] dataGroup_hi_307 = {dataGroup_hi_hi_307, dataGroup_hi_lo_307};
  wire [7:0]    dataGroup_19_9 = dataGroup_lo_307[639:632];
  wire [1023:0] dataGroup_lo_308 = {dataGroup_lo_hi_308, dataGroup_lo_lo_308};
  wire [1023:0] dataGroup_hi_308 = {dataGroup_hi_hi_308, dataGroup_hi_lo_308};
  wire [7:0]    dataGroup_20_9 = dataGroup_lo_308[671:664];
  wire [1023:0] dataGroup_lo_309 = {dataGroup_lo_hi_309, dataGroup_lo_lo_309};
  wire [1023:0] dataGroup_hi_309 = {dataGroup_hi_hi_309, dataGroup_hi_lo_309};
  wire [7:0]    dataGroup_21_9 = dataGroup_lo_309[703:696];
  wire [1023:0] dataGroup_lo_310 = {dataGroup_lo_hi_310, dataGroup_lo_lo_310};
  wire [1023:0] dataGroup_hi_310 = {dataGroup_hi_hi_310, dataGroup_hi_lo_310};
  wire [7:0]    dataGroup_22_9 = dataGroup_lo_310[735:728];
  wire [1023:0] dataGroup_lo_311 = {dataGroup_lo_hi_311, dataGroup_lo_lo_311};
  wire [1023:0] dataGroup_hi_311 = {dataGroup_hi_hi_311, dataGroup_hi_lo_311};
  wire [7:0]    dataGroup_23_9 = dataGroup_lo_311[767:760];
  wire [1023:0] dataGroup_lo_312 = {dataGroup_lo_hi_312, dataGroup_lo_lo_312};
  wire [1023:0] dataGroup_hi_312 = {dataGroup_hi_hi_312, dataGroup_hi_lo_312};
  wire [7:0]    dataGroup_24_9 = dataGroup_lo_312[799:792];
  wire [1023:0] dataGroup_lo_313 = {dataGroup_lo_hi_313, dataGroup_lo_lo_313};
  wire [1023:0] dataGroup_hi_313 = {dataGroup_hi_hi_313, dataGroup_hi_lo_313};
  wire [7:0]    dataGroup_25_9 = dataGroup_lo_313[831:824];
  wire [1023:0] dataGroup_lo_314 = {dataGroup_lo_hi_314, dataGroup_lo_lo_314};
  wire [1023:0] dataGroup_hi_314 = {dataGroup_hi_hi_314, dataGroup_hi_lo_314};
  wire [7:0]    dataGroup_26_9 = dataGroup_lo_314[863:856];
  wire [1023:0] dataGroup_lo_315 = {dataGroup_lo_hi_315, dataGroup_lo_lo_315};
  wire [1023:0] dataGroup_hi_315 = {dataGroup_hi_hi_315, dataGroup_hi_lo_315};
  wire [7:0]    dataGroup_27_9 = dataGroup_lo_315[895:888];
  wire [1023:0] dataGroup_lo_316 = {dataGroup_lo_hi_316, dataGroup_lo_lo_316};
  wire [1023:0] dataGroup_hi_316 = {dataGroup_hi_hi_316, dataGroup_hi_lo_316};
  wire [7:0]    dataGroup_28_9 = dataGroup_lo_316[927:920];
  wire [1023:0] dataGroup_lo_317 = {dataGroup_lo_hi_317, dataGroup_lo_lo_317};
  wire [1023:0] dataGroup_hi_317 = {dataGroup_hi_hi_317, dataGroup_hi_lo_317};
  wire [7:0]    dataGroup_29_9 = dataGroup_lo_317[959:952];
  wire [1023:0] dataGroup_lo_318 = {dataGroup_lo_hi_318, dataGroup_lo_lo_318};
  wire [1023:0] dataGroup_hi_318 = {dataGroup_hi_hi_318, dataGroup_hi_lo_318};
  wire [7:0]    dataGroup_30_9 = dataGroup_lo_318[991:984];
  wire [1023:0] dataGroup_lo_319 = {dataGroup_lo_hi_319, dataGroup_lo_lo_319};
  wire [1023:0] dataGroup_hi_319 = {dataGroup_hi_hi_319, dataGroup_hi_lo_319};
  wire [7:0]    dataGroup_31_9 = dataGroup_lo_319[1023:1016];
  wire [15:0]   res_lo_lo_lo_lo_9 = {dataGroup_1_9, dataGroup_0_9};
  wire [15:0]   res_lo_lo_lo_hi_9 = {dataGroup_3_9, dataGroup_2_9};
  wire [31:0]   res_lo_lo_lo_9 = {res_lo_lo_lo_hi_9, res_lo_lo_lo_lo_9};
  wire [15:0]   res_lo_lo_hi_lo_9 = {dataGroup_5_9, dataGroup_4_9};
  wire [15:0]   res_lo_lo_hi_hi_9 = {dataGroup_7_9, dataGroup_6_9};
  wire [31:0]   res_lo_lo_hi_9 = {res_lo_lo_hi_hi_9, res_lo_lo_hi_lo_9};
  wire [63:0]   res_lo_lo_9 = {res_lo_lo_hi_9, res_lo_lo_lo_9};
  wire [15:0]   res_lo_hi_lo_lo_9 = {dataGroup_9_9, dataGroup_8_9};
  wire [15:0]   res_lo_hi_lo_hi_9 = {dataGroup_11_9, dataGroup_10_9};
  wire [31:0]   res_lo_hi_lo_9 = {res_lo_hi_lo_hi_9, res_lo_hi_lo_lo_9};
  wire [15:0]   res_lo_hi_hi_lo_9 = {dataGroup_13_9, dataGroup_12_9};
  wire [15:0]   res_lo_hi_hi_hi_9 = {dataGroup_15_9, dataGroup_14_9};
  wire [31:0]   res_lo_hi_hi_9 = {res_lo_hi_hi_hi_9, res_lo_hi_hi_lo_9};
  wire [63:0]   res_lo_hi_9 = {res_lo_hi_hi_9, res_lo_hi_lo_9};
  wire [127:0]  res_lo_9 = {res_lo_hi_9, res_lo_lo_9};
  wire [15:0]   res_hi_lo_lo_lo_9 = {dataGroup_17_9, dataGroup_16_9};
  wire [15:0]   res_hi_lo_lo_hi_9 = {dataGroup_19_9, dataGroup_18_9};
  wire [31:0]   res_hi_lo_lo_9 = {res_hi_lo_lo_hi_9, res_hi_lo_lo_lo_9};
  wire [15:0]   res_hi_lo_hi_lo_9 = {dataGroup_21_9, dataGroup_20_9};
  wire [15:0]   res_hi_lo_hi_hi_9 = {dataGroup_23_9, dataGroup_22_9};
  wire [31:0]   res_hi_lo_hi_9 = {res_hi_lo_hi_hi_9, res_hi_lo_hi_lo_9};
  wire [63:0]   res_hi_lo_9 = {res_hi_lo_hi_9, res_hi_lo_lo_9};
  wire [15:0]   res_hi_hi_lo_lo_9 = {dataGroup_25_9, dataGroup_24_9};
  wire [15:0]   res_hi_hi_lo_hi_9 = {dataGroup_27_9, dataGroup_26_9};
  wire [31:0]   res_hi_hi_lo_9 = {res_hi_hi_lo_hi_9, res_hi_hi_lo_lo_9};
  wire [15:0]   res_hi_hi_hi_lo_9 = {dataGroup_29_9, dataGroup_28_9};
  wire [15:0]   res_hi_hi_hi_hi_9 = {dataGroup_31_9, dataGroup_30_9};
  wire [31:0]   res_hi_hi_hi_9 = {res_hi_hi_hi_hi_9, res_hi_hi_hi_lo_9};
  wire [63:0]   res_hi_hi_9 = {res_hi_hi_hi_9, res_hi_hi_lo_9};
  wire [127:0]  res_hi_9 = {res_hi_hi_9, res_hi_lo_9};
  wire [255:0]  res_27 = {res_hi_9, res_lo_9};
  wire [511:0]  lo_lo_3 = {res_25, res_24};
  wire [511:0]  lo_hi_3 = {res_27, res_26};
  wire [1023:0] lo_3 = {lo_hi_3, lo_lo_3};
  wire [2047:0] regroupLoadData_0_3 = {1024'h0, lo_3};
  wire [1023:0] dataGroup_lo_320 = {dataGroup_lo_hi_320, dataGroup_lo_lo_320};
  wire [1023:0] dataGroup_hi_320 = {dataGroup_hi_hi_320, dataGroup_hi_lo_320};
  wire [7:0]    dataGroup_0_10 = dataGroup_lo_320[7:0];
  wire [1023:0] dataGroup_lo_321 = {dataGroup_lo_hi_321, dataGroup_lo_lo_321};
  wire [1023:0] dataGroup_hi_321 = {dataGroup_hi_hi_321, dataGroup_hi_lo_321};
  wire [7:0]    dataGroup_1_10 = dataGroup_lo_321[47:40];
  wire [1023:0] dataGroup_lo_322 = {dataGroup_lo_hi_322, dataGroup_lo_lo_322};
  wire [1023:0] dataGroup_hi_322 = {dataGroup_hi_hi_322, dataGroup_hi_lo_322};
  wire [7:0]    dataGroup_2_10 = dataGroup_lo_322[87:80];
  wire [1023:0] dataGroup_lo_323 = {dataGroup_lo_hi_323, dataGroup_lo_lo_323};
  wire [1023:0] dataGroup_hi_323 = {dataGroup_hi_hi_323, dataGroup_hi_lo_323};
  wire [7:0]    dataGroup_3_10 = dataGroup_lo_323[127:120];
  wire [1023:0] dataGroup_lo_324 = {dataGroup_lo_hi_324, dataGroup_lo_lo_324};
  wire [1023:0] dataGroup_hi_324 = {dataGroup_hi_hi_324, dataGroup_hi_lo_324};
  wire [7:0]    dataGroup_4_10 = dataGroup_lo_324[167:160];
  wire [1023:0] dataGroup_lo_325 = {dataGroup_lo_hi_325, dataGroup_lo_lo_325};
  wire [1023:0] dataGroup_hi_325 = {dataGroup_hi_hi_325, dataGroup_hi_lo_325};
  wire [7:0]    dataGroup_5_10 = dataGroup_lo_325[207:200];
  wire [1023:0] dataGroup_lo_326 = {dataGroup_lo_hi_326, dataGroup_lo_lo_326};
  wire [1023:0] dataGroup_hi_326 = {dataGroup_hi_hi_326, dataGroup_hi_lo_326};
  wire [7:0]    dataGroup_6_10 = dataGroup_lo_326[247:240];
  wire [1023:0] dataGroup_lo_327 = {dataGroup_lo_hi_327, dataGroup_lo_lo_327};
  wire [1023:0] dataGroup_hi_327 = {dataGroup_hi_hi_327, dataGroup_hi_lo_327};
  wire [7:0]    dataGroup_7_10 = dataGroup_lo_327[287:280];
  wire [1023:0] dataGroup_lo_328 = {dataGroup_lo_hi_328, dataGroup_lo_lo_328};
  wire [1023:0] dataGroup_hi_328 = {dataGroup_hi_hi_328, dataGroup_hi_lo_328};
  wire [7:0]    dataGroup_8_10 = dataGroup_lo_328[327:320];
  wire [1023:0] dataGroup_lo_329 = {dataGroup_lo_hi_329, dataGroup_lo_lo_329};
  wire [1023:0] dataGroup_hi_329 = {dataGroup_hi_hi_329, dataGroup_hi_lo_329};
  wire [7:0]    dataGroup_9_10 = dataGroup_lo_329[367:360];
  wire [1023:0] dataGroup_lo_330 = {dataGroup_lo_hi_330, dataGroup_lo_lo_330};
  wire [1023:0] dataGroup_hi_330 = {dataGroup_hi_hi_330, dataGroup_hi_lo_330};
  wire [7:0]    dataGroup_10_10 = dataGroup_lo_330[407:400];
  wire [1023:0] dataGroup_lo_331 = {dataGroup_lo_hi_331, dataGroup_lo_lo_331};
  wire [1023:0] dataGroup_hi_331 = {dataGroup_hi_hi_331, dataGroup_hi_lo_331};
  wire [7:0]    dataGroup_11_10 = dataGroup_lo_331[447:440];
  wire [1023:0] dataGroup_lo_332 = {dataGroup_lo_hi_332, dataGroup_lo_lo_332};
  wire [1023:0] dataGroup_hi_332 = {dataGroup_hi_hi_332, dataGroup_hi_lo_332};
  wire [7:0]    dataGroup_12_10 = dataGroup_lo_332[487:480];
  wire [1023:0] dataGroup_lo_333 = {dataGroup_lo_hi_333, dataGroup_lo_lo_333};
  wire [1023:0] dataGroup_hi_333 = {dataGroup_hi_hi_333, dataGroup_hi_lo_333};
  wire [7:0]    dataGroup_13_10 = dataGroup_lo_333[527:520];
  wire [1023:0] dataGroup_lo_334 = {dataGroup_lo_hi_334, dataGroup_lo_lo_334};
  wire [1023:0] dataGroup_hi_334 = {dataGroup_hi_hi_334, dataGroup_hi_lo_334};
  wire [7:0]    dataGroup_14_10 = dataGroup_lo_334[567:560];
  wire [1023:0] dataGroup_lo_335 = {dataGroup_lo_hi_335, dataGroup_lo_lo_335};
  wire [1023:0] dataGroup_hi_335 = {dataGroup_hi_hi_335, dataGroup_hi_lo_335};
  wire [7:0]    dataGroup_15_10 = dataGroup_lo_335[607:600];
  wire [1023:0] dataGroup_lo_336 = {dataGroup_lo_hi_336, dataGroup_lo_lo_336};
  wire [1023:0] dataGroup_hi_336 = {dataGroup_hi_hi_336, dataGroup_hi_lo_336};
  wire [7:0]    dataGroup_16_10 = dataGroup_lo_336[647:640];
  wire [1023:0] dataGroup_lo_337 = {dataGroup_lo_hi_337, dataGroup_lo_lo_337};
  wire [1023:0] dataGroup_hi_337 = {dataGroup_hi_hi_337, dataGroup_hi_lo_337};
  wire [7:0]    dataGroup_17_10 = dataGroup_lo_337[687:680];
  wire [1023:0] dataGroup_lo_338 = {dataGroup_lo_hi_338, dataGroup_lo_lo_338};
  wire [1023:0] dataGroup_hi_338 = {dataGroup_hi_hi_338, dataGroup_hi_lo_338};
  wire [7:0]    dataGroup_18_10 = dataGroup_lo_338[727:720];
  wire [1023:0] dataGroup_lo_339 = {dataGroup_lo_hi_339, dataGroup_lo_lo_339};
  wire [1023:0] dataGroup_hi_339 = {dataGroup_hi_hi_339, dataGroup_hi_lo_339};
  wire [7:0]    dataGroup_19_10 = dataGroup_lo_339[767:760];
  wire [1023:0] dataGroup_lo_340 = {dataGroup_lo_hi_340, dataGroup_lo_lo_340};
  wire [1023:0] dataGroup_hi_340 = {dataGroup_hi_hi_340, dataGroup_hi_lo_340};
  wire [7:0]    dataGroup_20_10 = dataGroup_lo_340[807:800];
  wire [1023:0] dataGroup_lo_341 = {dataGroup_lo_hi_341, dataGroup_lo_lo_341};
  wire [1023:0] dataGroup_hi_341 = {dataGroup_hi_hi_341, dataGroup_hi_lo_341};
  wire [7:0]    dataGroup_21_10 = dataGroup_lo_341[847:840];
  wire [1023:0] dataGroup_lo_342 = {dataGroup_lo_hi_342, dataGroup_lo_lo_342};
  wire [1023:0] dataGroup_hi_342 = {dataGroup_hi_hi_342, dataGroup_hi_lo_342};
  wire [7:0]    dataGroup_22_10 = dataGroup_lo_342[887:880];
  wire [1023:0] dataGroup_lo_343 = {dataGroup_lo_hi_343, dataGroup_lo_lo_343};
  wire [1023:0] dataGroup_hi_343 = {dataGroup_hi_hi_343, dataGroup_hi_lo_343};
  wire [7:0]    dataGroup_23_10 = dataGroup_lo_343[927:920];
  wire [1023:0] dataGroup_lo_344 = {dataGroup_lo_hi_344, dataGroup_lo_lo_344};
  wire [1023:0] dataGroup_hi_344 = {dataGroup_hi_hi_344, dataGroup_hi_lo_344};
  wire [7:0]    dataGroup_24_10 = dataGroup_lo_344[967:960];
  wire [1023:0] dataGroup_lo_345 = {dataGroup_lo_hi_345, dataGroup_lo_lo_345};
  wire [1023:0] dataGroup_hi_345 = {dataGroup_hi_hi_345, dataGroup_hi_lo_345};
  wire [7:0]    dataGroup_25_10 = dataGroup_lo_345[1007:1000];
  wire [1023:0] dataGroup_lo_346 = {dataGroup_lo_hi_346, dataGroup_lo_lo_346};
  wire [1023:0] dataGroup_hi_346 = {dataGroup_hi_hi_346, dataGroup_hi_lo_346};
  wire [7:0]    dataGroup_26_10 = dataGroup_hi_346[23:16];
  wire [1023:0] dataGroup_lo_347 = {dataGroup_lo_hi_347, dataGroup_lo_lo_347};
  wire [1023:0] dataGroup_hi_347 = {dataGroup_hi_hi_347, dataGroup_hi_lo_347};
  wire [7:0]    dataGroup_27_10 = dataGroup_hi_347[63:56];
  wire [1023:0] dataGroup_lo_348 = {dataGroup_lo_hi_348, dataGroup_lo_lo_348};
  wire [1023:0] dataGroup_hi_348 = {dataGroup_hi_hi_348, dataGroup_hi_lo_348};
  wire [7:0]    dataGroup_28_10 = dataGroup_hi_348[103:96];
  wire [1023:0] dataGroup_lo_349 = {dataGroup_lo_hi_349, dataGroup_lo_lo_349};
  wire [1023:0] dataGroup_hi_349 = {dataGroup_hi_hi_349, dataGroup_hi_lo_349};
  wire [7:0]    dataGroup_29_10 = dataGroup_hi_349[143:136];
  wire [1023:0] dataGroup_lo_350 = {dataGroup_lo_hi_350, dataGroup_lo_lo_350};
  wire [1023:0] dataGroup_hi_350 = {dataGroup_hi_hi_350, dataGroup_hi_lo_350};
  wire [7:0]    dataGroup_30_10 = dataGroup_hi_350[183:176];
  wire [1023:0] dataGroup_lo_351 = {dataGroup_lo_hi_351, dataGroup_lo_lo_351};
  wire [1023:0] dataGroup_hi_351 = {dataGroup_hi_hi_351, dataGroup_hi_lo_351};
  wire [7:0]    dataGroup_31_10 = dataGroup_hi_351[223:216];
  wire [15:0]   res_lo_lo_lo_lo_10 = {dataGroup_1_10, dataGroup_0_10};
  wire [15:0]   res_lo_lo_lo_hi_10 = {dataGroup_3_10, dataGroup_2_10};
  wire [31:0]   res_lo_lo_lo_10 = {res_lo_lo_lo_hi_10, res_lo_lo_lo_lo_10};
  wire [15:0]   res_lo_lo_hi_lo_10 = {dataGroup_5_10, dataGroup_4_10};
  wire [15:0]   res_lo_lo_hi_hi_10 = {dataGroup_7_10, dataGroup_6_10};
  wire [31:0]   res_lo_lo_hi_10 = {res_lo_lo_hi_hi_10, res_lo_lo_hi_lo_10};
  wire [63:0]   res_lo_lo_10 = {res_lo_lo_hi_10, res_lo_lo_lo_10};
  wire [15:0]   res_lo_hi_lo_lo_10 = {dataGroup_9_10, dataGroup_8_10};
  wire [15:0]   res_lo_hi_lo_hi_10 = {dataGroup_11_10, dataGroup_10_10};
  wire [31:0]   res_lo_hi_lo_10 = {res_lo_hi_lo_hi_10, res_lo_hi_lo_lo_10};
  wire [15:0]   res_lo_hi_hi_lo_10 = {dataGroup_13_10, dataGroup_12_10};
  wire [15:0]   res_lo_hi_hi_hi_10 = {dataGroup_15_10, dataGroup_14_10};
  wire [31:0]   res_lo_hi_hi_10 = {res_lo_hi_hi_hi_10, res_lo_hi_hi_lo_10};
  wire [63:0]   res_lo_hi_10 = {res_lo_hi_hi_10, res_lo_hi_lo_10};
  wire [127:0]  res_lo_10 = {res_lo_hi_10, res_lo_lo_10};
  wire [15:0]   res_hi_lo_lo_lo_10 = {dataGroup_17_10, dataGroup_16_10};
  wire [15:0]   res_hi_lo_lo_hi_10 = {dataGroup_19_10, dataGroup_18_10};
  wire [31:0]   res_hi_lo_lo_10 = {res_hi_lo_lo_hi_10, res_hi_lo_lo_lo_10};
  wire [15:0]   res_hi_lo_hi_lo_10 = {dataGroup_21_10, dataGroup_20_10};
  wire [15:0]   res_hi_lo_hi_hi_10 = {dataGroup_23_10, dataGroup_22_10};
  wire [31:0]   res_hi_lo_hi_10 = {res_hi_lo_hi_hi_10, res_hi_lo_hi_lo_10};
  wire [63:0]   res_hi_lo_10 = {res_hi_lo_hi_10, res_hi_lo_lo_10};
  wire [15:0]   res_hi_hi_lo_lo_10 = {dataGroup_25_10, dataGroup_24_10};
  wire [15:0]   res_hi_hi_lo_hi_10 = {dataGroup_27_10, dataGroup_26_10};
  wire [31:0]   res_hi_hi_lo_10 = {res_hi_hi_lo_hi_10, res_hi_hi_lo_lo_10};
  wire [15:0]   res_hi_hi_hi_lo_10 = {dataGroup_29_10, dataGroup_28_10};
  wire [15:0]   res_hi_hi_hi_hi_10 = {dataGroup_31_10, dataGroup_30_10};
  wire [31:0]   res_hi_hi_hi_10 = {res_hi_hi_hi_hi_10, res_hi_hi_hi_lo_10};
  wire [63:0]   res_hi_hi_10 = {res_hi_hi_hi_10, res_hi_hi_lo_10};
  wire [127:0]  res_hi_10 = {res_hi_hi_10, res_hi_lo_10};
  wire [255:0]  res_32 = {res_hi_10, res_lo_10};
  wire [1023:0] dataGroup_lo_352 = {dataGroup_lo_hi_352, dataGroup_lo_lo_352};
  wire [1023:0] dataGroup_hi_352 = {dataGroup_hi_hi_352, dataGroup_hi_lo_352};
  wire [7:0]    dataGroup_0_11 = dataGroup_lo_352[15:8];
  wire [1023:0] dataGroup_lo_353 = {dataGroup_lo_hi_353, dataGroup_lo_lo_353};
  wire [1023:0] dataGroup_hi_353 = {dataGroup_hi_hi_353, dataGroup_hi_lo_353};
  wire [7:0]    dataGroup_1_11 = dataGroup_lo_353[55:48];
  wire [1023:0] dataGroup_lo_354 = {dataGroup_lo_hi_354, dataGroup_lo_lo_354};
  wire [1023:0] dataGroup_hi_354 = {dataGroup_hi_hi_354, dataGroup_hi_lo_354};
  wire [7:0]    dataGroup_2_11 = dataGroup_lo_354[95:88];
  wire [1023:0] dataGroup_lo_355 = {dataGroup_lo_hi_355, dataGroup_lo_lo_355};
  wire [1023:0] dataGroup_hi_355 = {dataGroup_hi_hi_355, dataGroup_hi_lo_355};
  wire [7:0]    dataGroup_3_11 = dataGroup_lo_355[135:128];
  wire [1023:0] dataGroup_lo_356 = {dataGroup_lo_hi_356, dataGroup_lo_lo_356};
  wire [1023:0] dataGroup_hi_356 = {dataGroup_hi_hi_356, dataGroup_hi_lo_356};
  wire [7:0]    dataGroup_4_11 = dataGroup_lo_356[175:168];
  wire [1023:0] dataGroup_lo_357 = {dataGroup_lo_hi_357, dataGroup_lo_lo_357};
  wire [1023:0] dataGroup_hi_357 = {dataGroup_hi_hi_357, dataGroup_hi_lo_357};
  wire [7:0]    dataGroup_5_11 = dataGroup_lo_357[215:208];
  wire [1023:0] dataGroup_lo_358 = {dataGroup_lo_hi_358, dataGroup_lo_lo_358};
  wire [1023:0] dataGroup_hi_358 = {dataGroup_hi_hi_358, dataGroup_hi_lo_358};
  wire [7:0]    dataGroup_6_11 = dataGroup_lo_358[255:248];
  wire [1023:0] dataGroup_lo_359 = {dataGroup_lo_hi_359, dataGroup_lo_lo_359};
  wire [1023:0] dataGroup_hi_359 = {dataGroup_hi_hi_359, dataGroup_hi_lo_359};
  wire [7:0]    dataGroup_7_11 = dataGroup_lo_359[295:288];
  wire [1023:0] dataGroup_lo_360 = {dataGroup_lo_hi_360, dataGroup_lo_lo_360};
  wire [1023:0] dataGroup_hi_360 = {dataGroup_hi_hi_360, dataGroup_hi_lo_360};
  wire [7:0]    dataGroup_8_11 = dataGroup_lo_360[335:328];
  wire [1023:0] dataGroup_lo_361 = {dataGroup_lo_hi_361, dataGroup_lo_lo_361};
  wire [1023:0] dataGroup_hi_361 = {dataGroup_hi_hi_361, dataGroup_hi_lo_361};
  wire [7:0]    dataGroup_9_11 = dataGroup_lo_361[375:368];
  wire [1023:0] dataGroup_lo_362 = {dataGroup_lo_hi_362, dataGroup_lo_lo_362};
  wire [1023:0] dataGroup_hi_362 = {dataGroup_hi_hi_362, dataGroup_hi_lo_362};
  wire [7:0]    dataGroup_10_11 = dataGroup_lo_362[415:408];
  wire [1023:0] dataGroup_lo_363 = {dataGroup_lo_hi_363, dataGroup_lo_lo_363};
  wire [1023:0] dataGroup_hi_363 = {dataGroup_hi_hi_363, dataGroup_hi_lo_363};
  wire [7:0]    dataGroup_11_11 = dataGroup_lo_363[455:448];
  wire [1023:0] dataGroup_lo_364 = {dataGroup_lo_hi_364, dataGroup_lo_lo_364};
  wire [1023:0] dataGroup_hi_364 = {dataGroup_hi_hi_364, dataGroup_hi_lo_364};
  wire [7:0]    dataGroup_12_11 = dataGroup_lo_364[495:488];
  wire [1023:0] dataGroup_lo_365 = {dataGroup_lo_hi_365, dataGroup_lo_lo_365};
  wire [1023:0] dataGroup_hi_365 = {dataGroup_hi_hi_365, dataGroup_hi_lo_365};
  wire [7:0]    dataGroup_13_11 = dataGroup_lo_365[535:528];
  wire [1023:0] dataGroup_lo_366 = {dataGroup_lo_hi_366, dataGroup_lo_lo_366};
  wire [1023:0] dataGroup_hi_366 = {dataGroup_hi_hi_366, dataGroup_hi_lo_366};
  wire [7:0]    dataGroup_14_11 = dataGroup_lo_366[575:568];
  wire [1023:0] dataGroup_lo_367 = {dataGroup_lo_hi_367, dataGroup_lo_lo_367};
  wire [1023:0] dataGroup_hi_367 = {dataGroup_hi_hi_367, dataGroup_hi_lo_367};
  wire [7:0]    dataGroup_15_11 = dataGroup_lo_367[615:608];
  wire [1023:0] dataGroup_lo_368 = {dataGroup_lo_hi_368, dataGroup_lo_lo_368};
  wire [1023:0] dataGroup_hi_368 = {dataGroup_hi_hi_368, dataGroup_hi_lo_368};
  wire [7:0]    dataGroup_16_11 = dataGroup_lo_368[655:648];
  wire [1023:0] dataGroup_lo_369 = {dataGroup_lo_hi_369, dataGroup_lo_lo_369};
  wire [1023:0] dataGroup_hi_369 = {dataGroup_hi_hi_369, dataGroup_hi_lo_369};
  wire [7:0]    dataGroup_17_11 = dataGroup_lo_369[695:688];
  wire [1023:0] dataGroup_lo_370 = {dataGroup_lo_hi_370, dataGroup_lo_lo_370};
  wire [1023:0] dataGroup_hi_370 = {dataGroup_hi_hi_370, dataGroup_hi_lo_370};
  wire [7:0]    dataGroup_18_11 = dataGroup_lo_370[735:728];
  wire [1023:0] dataGroup_lo_371 = {dataGroup_lo_hi_371, dataGroup_lo_lo_371};
  wire [1023:0] dataGroup_hi_371 = {dataGroup_hi_hi_371, dataGroup_hi_lo_371};
  wire [7:0]    dataGroup_19_11 = dataGroup_lo_371[775:768];
  wire [1023:0] dataGroup_lo_372 = {dataGroup_lo_hi_372, dataGroup_lo_lo_372};
  wire [1023:0] dataGroup_hi_372 = {dataGroup_hi_hi_372, dataGroup_hi_lo_372};
  wire [7:0]    dataGroup_20_11 = dataGroup_lo_372[815:808];
  wire [1023:0] dataGroup_lo_373 = {dataGroup_lo_hi_373, dataGroup_lo_lo_373};
  wire [1023:0] dataGroup_hi_373 = {dataGroup_hi_hi_373, dataGroup_hi_lo_373};
  wire [7:0]    dataGroup_21_11 = dataGroup_lo_373[855:848];
  wire [1023:0] dataGroup_lo_374 = {dataGroup_lo_hi_374, dataGroup_lo_lo_374};
  wire [1023:0] dataGroup_hi_374 = {dataGroup_hi_hi_374, dataGroup_hi_lo_374};
  wire [7:0]    dataGroup_22_11 = dataGroup_lo_374[895:888];
  wire [1023:0] dataGroup_lo_375 = {dataGroup_lo_hi_375, dataGroup_lo_lo_375};
  wire [1023:0] dataGroup_hi_375 = {dataGroup_hi_hi_375, dataGroup_hi_lo_375};
  wire [7:0]    dataGroup_23_11 = dataGroup_lo_375[935:928];
  wire [1023:0] dataGroup_lo_376 = {dataGroup_lo_hi_376, dataGroup_lo_lo_376};
  wire [1023:0] dataGroup_hi_376 = {dataGroup_hi_hi_376, dataGroup_hi_lo_376};
  wire [7:0]    dataGroup_24_11 = dataGroup_lo_376[975:968];
  wire [1023:0] dataGroup_lo_377 = {dataGroup_lo_hi_377, dataGroup_lo_lo_377};
  wire [1023:0] dataGroup_hi_377 = {dataGroup_hi_hi_377, dataGroup_hi_lo_377};
  wire [7:0]    dataGroup_25_11 = dataGroup_lo_377[1015:1008];
  wire [1023:0] dataGroup_lo_378 = {dataGroup_lo_hi_378, dataGroup_lo_lo_378};
  wire [1023:0] dataGroup_hi_378 = {dataGroup_hi_hi_378, dataGroup_hi_lo_378};
  wire [7:0]    dataGroup_26_11 = dataGroup_hi_378[31:24];
  wire [1023:0] dataGroup_lo_379 = {dataGroup_lo_hi_379, dataGroup_lo_lo_379};
  wire [1023:0] dataGroup_hi_379 = {dataGroup_hi_hi_379, dataGroup_hi_lo_379};
  wire [7:0]    dataGroup_27_11 = dataGroup_hi_379[71:64];
  wire [1023:0] dataGroup_lo_380 = {dataGroup_lo_hi_380, dataGroup_lo_lo_380};
  wire [1023:0] dataGroup_hi_380 = {dataGroup_hi_hi_380, dataGroup_hi_lo_380};
  wire [7:0]    dataGroup_28_11 = dataGroup_hi_380[111:104];
  wire [1023:0] dataGroup_lo_381 = {dataGroup_lo_hi_381, dataGroup_lo_lo_381};
  wire [1023:0] dataGroup_hi_381 = {dataGroup_hi_hi_381, dataGroup_hi_lo_381};
  wire [7:0]    dataGroup_29_11 = dataGroup_hi_381[151:144];
  wire [1023:0] dataGroup_lo_382 = {dataGroup_lo_hi_382, dataGroup_lo_lo_382};
  wire [1023:0] dataGroup_hi_382 = {dataGroup_hi_hi_382, dataGroup_hi_lo_382};
  wire [7:0]    dataGroup_30_11 = dataGroup_hi_382[191:184];
  wire [1023:0] dataGroup_lo_383 = {dataGroup_lo_hi_383, dataGroup_lo_lo_383};
  wire [1023:0] dataGroup_hi_383 = {dataGroup_hi_hi_383, dataGroup_hi_lo_383};
  wire [7:0]    dataGroup_31_11 = dataGroup_hi_383[231:224];
  wire [15:0]   res_lo_lo_lo_lo_11 = {dataGroup_1_11, dataGroup_0_11};
  wire [15:0]   res_lo_lo_lo_hi_11 = {dataGroup_3_11, dataGroup_2_11};
  wire [31:0]   res_lo_lo_lo_11 = {res_lo_lo_lo_hi_11, res_lo_lo_lo_lo_11};
  wire [15:0]   res_lo_lo_hi_lo_11 = {dataGroup_5_11, dataGroup_4_11};
  wire [15:0]   res_lo_lo_hi_hi_11 = {dataGroup_7_11, dataGroup_6_11};
  wire [31:0]   res_lo_lo_hi_11 = {res_lo_lo_hi_hi_11, res_lo_lo_hi_lo_11};
  wire [63:0]   res_lo_lo_11 = {res_lo_lo_hi_11, res_lo_lo_lo_11};
  wire [15:0]   res_lo_hi_lo_lo_11 = {dataGroup_9_11, dataGroup_8_11};
  wire [15:0]   res_lo_hi_lo_hi_11 = {dataGroup_11_11, dataGroup_10_11};
  wire [31:0]   res_lo_hi_lo_11 = {res_lo_hi_lo_hi_11, res_lo_hi_lo_lo_11};
  wire [15:0]   res_lo_hi_hi_lo_11 = {dataGroup_13_11, dataGroup_12_11};
  wire [15:0]   res_lo_hi_hi_hi_11 = {dataGroup_15_11, dataGroup_14_11};
  wire [31:0]   res_lo_hi_hi_11 = {res_lo_hi_hi_hi_11, res_lo_hi_hi_lo_11};
  wire [63:0]   res_lo_hi_11 = {res_lo_hi_hi_11, res_lo_hi_lo_11};
  wire [127:0]  res_lo_11 = {res_lo_hi_11, res_lo_lo_11};
  wire [15:0]   res_hi_lo_lo_lo_11 = {dataGroup_17_11, dataGroup_16_11};
  wire [15:0]   res_hi_lo_lo_hi_11 = {dataGroup_19_11, dataGroup_18_11};
  wire [31:0]   res_hi_lo_lo_11 = {res_hi_lo_lo_hi_11, res_hi_lo_lo_lo_11};
  wire [15:0]   res_hi_lo_hi_lo_11 = {dataGroup_21_11, dataGroup_20_11};
  wire [15:0]   res_hi_lo_hi_hi_11 = {dataGroup_23_11, dataGroup_22_11};
  wire [31:0]   res_hi_lo_hi_11 = {res_hi_lo_hi_hi_11, res_hi_lo_hi_lo_11};
  wire [63:0]   res_hi_lo_11 = {res_hi_lo_hi_11, res_hi_lo_lo_11};
  wire [15:0]   res_hi_hi_lo_lo_11 = {dataGroup_25_11, dataGroup_24_11};
  wire [15:0]   res_hi_hi_lo_hi_11 = {dataGroup_27_11, dataGroup_26_11};
  wire [31:0]   res_hi_hi_lo_11 = {res_hi_hi_lo_hi_11, res_hi_hi_lo_lo_11};
  wire [15:0]   res_hi_hi_hi_lo_11 = {dataGroup_29_11, dataGroup_28_11};
  wire [15:0]   res_hi_hi_hi_hi_11 = {dataGroup_31_11, dataGroup_30_11};
  wire [31:0]   res_hi_hi_hi_11 = {res_hi_hi_hi_hi_11, res_hi_hi_hi_lo_11};
  wire [63:0]   res_hi_hi_11 = {res_hi_hi_hi_11, res_hi_hi_lo_11};
  wire [127:0]  res_hi_11 = {res_hi_hi_11, res_hi_lo_11};
  wire [255:0]  res_33 = {res_hi_11, res_lo_11};
  wire [1023:0] dataGroup_lo_384 = {dataGroup_lo_hi_384, dataGroup_lo_lo_384};
  wire [1023:0] dataGroup_hi_384 = {dataGroup_hi_hi_384, dataGroup_hi_lo_384};
  wire [7:0]    dataGroup_0_12 = dataGroup_lo_384[23:16];
  wire [1023:0] dataGroup_lo_385 = {dataGroup_lo_hi_385, dataGroup_lo_lo_385};
  wire [1023:0] dataGroup_hi_385 = {dataGroup_hi_hi_385, dataGroup_hi_lo_385};
  wire [7:0]    dataGroup_1_12 = dataGroup_lo_385[63:56];
  wire [1023:0] dataGroup_lo_386 = {dataGroup_lo_hi_386, dataGroup_lo_lo_386};
  wire [1023:0] dataGroup_hi_386 = {dataGroup_hi_hi_386, dataGroup_hi_lo_386};
  wire [7:0]    dataGroup_2_12 = dataGroup_lo_386[103:96];
  wire [1023:0] dataGroup_lo_387 = {dataGroup_lo_hi_387, dataGroup_lo_lo_387};
  wire [1023:0] dataGroup_hi_387 = {dataGroup_hi_hi_387, dataGroup_hi_lo_387};
  wire [7:0]    dataGroup_3_12 = dataGroup_lo_387[143:136];
  wire [1023:0] dataGroup_lo_388 = {dataGroup_lo_hi_388, dataGroup_lo_lo_388};
  wire [1023:0] dataGroup_hi_388 = {dataGroup_hi_hi_388, dataGroup_hi_lo_388};
  wire [7:0]    dataGroup_4_12 = dataGroup_lo_388[183:176];
  wire [1023:0] dataGroup_lo_389 = {dataGroup_lo_hi_389, dataGroup_lo_lo_389};
  wire [1023:0] dataGroup_hi_389 = {dataGroup_hi_hi_389, dataGroup_hi_lo_389};
  wire [7:0]    dataGroup_5_12 = dataGroup_lo_389[223:216];
  wire [1023:0] dataGroup_lo_390 = {dataGroup_lo_hi_390, dataGroup_lo_lo_390};
  wire [1023:0] dataGroup_hi_390 = {dataGroup_hi_hi_390, dataGroup_hi_lo_390};
  wire [7:0]    dataGroup_6_12 = dataGroup_lo_390[263:256];
  wire [1023:0] dataGroup_lo_391 = {dataGroup_lo_hi_391, dataGroup_lo_lo_391};
  wire [1023:0] dataGroup_hi_391 = {dataGroup_hi_hi_391, dataGroup_hi_lo_391};
  wire [7:0]    dataGroup_7_12 = dataGroup_lo_391[303:296];
  wire [1023:0] dataGroup_lo_392 = {dataGroup_lo_hi_392, dataGroup_lo_lo_392};
  wire [1023:0] dataGroup_hi_392 = {dataGroup_hi_hi_392, dataGroup_hi_lo_392};
  wire [7:0]    dataGroup_8_12 = dataGroup_lo_392[343:336];
  wire [1023:0] dataGroup_lo_393 = {dataGroup_lo_hi_393, dataGroup_lo_lo_393};
  wire [1023:0] dataGroup_hi_393 = {dataGroup_hi_hi_393, dataGroup_hi_lo_393};
  wire [7:0]    dataGroup_9_12 = dataGroup_lo_393[383:376];
  wire [1023:0] dataGroup_lo_394 = {dataGroup_lo_hi_394, dataGroup_lo_lo_394};
  wire [1023:0] dataGroup_hi_394 = {dataGroup_hi_hi_394, dataGroup_hi_lo_394};
  wire [7:0]    dataGroup_10_12 = dataGroup_lo_394[423:416];
  wire [1023:0] dataGroup_lo_395 = {dataGroup_lo_hi_395, dataGroup_lo_lo_395};
  wire [1023:0] dataGroup_hi_395 = {dataGroup_hi_hi_395, dataGroup_hi_lo_395};
  wire [7:0]    dataGroup_11_12 = dataGroup_lo_395[463:456];
  wire [1023:0] dataGroup_lo_396 = {dataGroup_lo_hi_396, dataGroup_lo_lo_396};
  wire [1023:0] dataGroup_hi_396 = {dataGroup_hi_hi_396, dataGroup_hi_lo_396};
  wire [7:0]    dataGroup_12_12 = dataGroup_lo_396[503:496];
  wire [1023:0] dataGroup_lo_397 = {dataGroup_lo_hi_397, dataGroup_lo_lo_397};
  wire [1023:0] dataGroup_hi_397 = {dataGroup_hi_hi_397, dataGroup_hi_lo_397};
  wire [7:0]    dataGroup_13_12 = dataGroup_lo_397[543:536];
  wire [1023:0] dataGroup_lo_398 = {dataGroup_lo_hi_398, dataGroup_lo_lo_398};
  wire [1023:0] dataGroup_hi_398 = {dataGroup_hi_hi_398, dataGroup_hi_lo_398};
  wire [7:0]    dataGroup_14_12 = dataGroup_lo_398[583:576];
  wire [1023:0] dataGroup_lo_399 = {dataGroup_lo_hi_399, dataGroup_lo_lo_399};
  wire [1023:0] dataGroup_hi_399 = {dataGroup_hi_hi_399, dataGroup_hi_lo_399};
  wire [7:0]    dataGroup_15_12 = dataGroup_lo_399[623:616];
  wire [1023:0] dataGroup_lo_400 = {dataGroup_lo_hi_400, dataGroup_lo_lo_400};
  wire [1023:0] dataGroup_hi_400 = {dataGroup_hi_hi_400, dataGroup_hi_lo_400};
  wire [7:0]    dataGroup_16_12 = dataGroup_lo_400[663:656];
  wire [1023:0] dataGroup_lo_401 = {dataGroup_lo_hi_401, dataGroup_lo_lo_401};
  wire [1023:0] dataGroup_hi_401 = {dataGroup_hi_hi_401, dataGroup_hi_lo_401};
  wire [7:0]    dataGroup_17_12 = dataGroup_lo_401[703:696];
  wire [1023:0] dataGroup_lo_402 = {dataGroup_lo_hi_402, dataGroup_lo_lo_402};
  wire [1023:0] dataGroup_hi_402 = {dataGroup_hi_hi_402, dataGroup_hi_lo_402};
  wire [7:0]    dataGroup_18_12 = dataGroup_lo_402[743:736];
  wire [1023:0] dataGroup_lo_403 = {dataGroup_lo_hi_403, dataGroup_lo_lo_403};
  wire [1023:0] dataGroup_hi_403 = {dataGroup_hi_hi_403, dataGroup_hi_lo_403};
  wire [7:0]    dataGroup_19_12 = dataGroup_lo_403[783:776];
  wire [1023:0] dataGroup_lo_404 = {dataGroup_lo_hi_404, dataGroup_lo_lo_404};
  wire [1023:0] dataGroup_hi_404 = {dataGroup_hi_hi_404, dataGroup_hi_lo_404};
  wire [7:0]    dataGroup_20_12 = dataGroup_lo_404[823:816];
  wire [1023:0] dataGroup_lo_405 = {dataGroup_lo_hi_405, dataGroup_lo_lo_405};
  wire [1023:0] dataGroup_hi_405 = {dataGroup_hi_hi_405, dataGroup_hi_lo_405};
  wire [7:0]    dataGroup_21_12 = dataGroup_lo_405[863:856];
  wire [1023:0] dataGroup_lo_406 = {dataGroup_lo_hi_406, dataGroup_lo_lo_406};
  wire [1023:0] dataGroup_hi_406 = {dataGroup_hi_hi_406, dataGroup_hi_lo_406};
  wire [7:0]    dataGroup_22_12 = dataGroup_lo_406[903:896];
  wire [1023:0] dataGroup_lo_407 = {dataGroup_lo_hi_407, dataGroup_lo_lo_407};
  wire [1023:0] dataGroup_hi_407 = {dataGroup_hi_hi_407, dataGroup_hi_lo_407};
  wire [7:0]    dataGroup_23_12 = dataGroup_lo_407[943:936];
  wire [1023:0] dataGroup_lo_408 = {dataGroup_lo_hi_408, dataGroup_lo_lo_408};
  wire [1023:0] dataGroup_hi_408 = {dataGroup_hi_hi_408, dataGroup_hi_lo_408};
  wire [7:0]    dataGroup_24_12 = dataGroup_lo_408[983:976];
  wire [1023:0] dataGroup_lo_409 = {dataGroup_lo_hi_409, dataGroup_lo_lo_409};
  wire [1023:0] dataGroup_hi_409 = {dataGroup_hi_hi_409, dataGroup_hi_lo_409};
  wire [7:0]    dataGroup_25_12 = dataGroup_lo_409[1023:1016];
  wire [1023:0] dataGroup_lo_410 = {dataGroup_lo_hi_410, dataGroup_lo_lo_410};
  wire [1023:0] dataGroup_hi_410 = {dataGroup_hi_hi_410, dataGroup_hi_lo_410};
  wire [7:0]    dataGroup_26_12 = dataGroup_hi_410[39:32];
  wire [1023:0] dataGroup_lo_411 = {dataGroup_lo_hi_411, dataGroup_lo_lo_411};
  wire [1023:0] dataGroup_hi_411 = {dataGroup_hi_hi_411, dataGroup_hi_lo_411};
  wire [7:0]    dataGroup_27_12 = dataGroup_hi_411[79:72];
  wire [1023:0] dataGroup_lo_412 = {dataGroup_lo_hi_412, dataGroup_lo_lo_412};
  wire [1023:0] dataGroup_hi_412 = {dataGroup_hi_hi_412, dataGroup_hi_lo_412};
  wire [7:0]    dataGroup_28_12 = dataGroup_hi_412[119:112];
  wire [1023:0] dataGroup_lo_413 = {dataGroup_lo_hi_413, dataGroup_lo_lo_413};
  wire [1023:0] dataGroup_hi_413 = {dataGroup_hi_hi_413, dataGroup_hi_lo_413};
  wire [7:0]    dataGroup_29_12 = dataGroup_hi_413[159:152];
  wire [1023:0] dataGroup_lo_414 = {dataGroup_lo_hi_414, dataGroup_lo_lo_414};
  wire [1023:0] dataGroup_hi_414 = {dataGroup_hi_hi_414, dataGroup_hi_lo_414};
  wire [7:0]    dataGroup_30_12 = dataGroup_hi_414[199:192];
  wire [1023:0] dataGroup_lo_415 = {dataGroup_lo_hi_415, dataGroup_lo_lo_415};
  wire [1023:0] dataGroup_hi_415 = {dataGroup_hi_hi_415, dataGroup_hi_lo_415};
  wire [7:0]    dataGroup_31_12 = dataGroup_hi_415[239:232];
  wire [15:0]   res_lo_lo_lo_lo_12 = {dataGroup_1_12, dataGroup_0_12};
  wire [15:0]   res_lo_lo_lo_hi_12 = {dataGroup_3_12, dataGroup_2_12};
  wire [31:0]   res_lo_lo_lo_12 = {res_lo_lo_lo_hi_12, res_lo_lo_lo_lo_12};
  wire [15:0]   res_lo_lo_hi_lo_12 = {dataGroup_5_12, dataGroup_4_12};
  wire [15:0]   res_lo_lo_hi_hi_12 = {dataGroup_7_12, dataGroup_6_12};
  wire [31:0]   res_lo_lo_hi_12 = {res_lo_lo_hi_hi_12, res_lo_lo_hi_lo_12};
  wire [63:0]   res_lo_lo_12 = {res_lo_lo_hi_12, res_lo_lo_lo_12};
  wire [15:0]   res_lo_hi_lo_lo_12 = {dataGroup_9_12, dataGroup_8_12};
  wire [15:0]   res_lo_hi_lo_hi_12 = {dataGroup_11_12, dataGroup_10_12};
  wire [31:0]   res_lo_hi_lo_12 = {res_lo_hi_lo_hi_12, res_lo_hi_lo_lo_12};
  wire [15:0]   res_lo_hi_hi_lo_12 = {dataGroup_13_12, dataGroup_12_12};
  wire [15:0]   res_lo_hi_hi_hi_12 = {dataGroup_15_12, dataGroup_14_12};
  wire [31:0]   res_lo_hi_hi_12 = {res_lo_hi_hi_hi_12, res_lo_hi_hi_lo_12};
  wire [63:0]   res_lo_hi_12 = {res_lo_hi_hi_12, res_lo_hi_lo_12};
  wire [127:0]  res_lo_12 = {res_lo_hi_12, res_lo_lo_12};
  wire [15:0]   res_hi_lo_lo_lo_12 = {dataGroup_17_12, dataGroup_16_12};
  wire [15:0]   res_hi_lo_lo_hi_12 = {dataGroup_19_12, dataGroup_18_12};
  wire [31:0]   res_hi_lo_lo_12 = {res_hi_lo_lo_hi_12, res_hi_lo_lo_lo_12};
  wire [15:0]   res_hi_lo_hi_lo_12 = {dataGroup_21_12, dataGroup_20_12};
  wire [15:0]   res_hi_lo_hi_hi_12 = {dataGroup_23_12, dataGroup_22_12};
  wire [31:0]   res_hi_lo_hi_12 = {res_hi_lo_hi_hi_12, res_hi_lo_hi_lo_12};
  wire [63:0]   res_hi_lo_12 = {res_hi_lo_hi_12, res_hi_lo_lo_12};
  wire [15:0]   res_hi_hi_lo_lo_12 = {dataGroup_25_12, dataGroup_24_12};
  wire [15:0]   res_hi_hi_lo_hi_12 = {dataGroup_27_12, dataGroup_26_12};
  wire [31:0]   res_hi_hi_lo_12 = {res_hi_hi_lo_hi_12, res_hi_hi_lo_lo_12};
  wire [15:0]   res_hi_hi_hi_lo_12 = {dataGroup_29_12, dataGroup_28_12};
  wire [15:0]   res_hi_hi_hi_hi_12 = {dataGroup_31_12, dataGroup_30_12};
  wire [31:0]   res_hi_hi_hi_12 = {res_hi_hi_hi_hi_12, res_hi_hi_hi_lo_12};
  wire [63:0]   res_hi_hi_12 = {res_hi_hi_hi_12, res_hi_hi_lo_12};
  wire [127:0]  res_hi_12 = {res_hi_hi_12, res_hi_lo_12};
  wire [255:0]  res_34 = {res_hi_12, res_lo_12};
  wire [1023:0] dataGroup_lo_416 = {dataGroup_lo_hi_416, dataGroup_lo_lo_416};
  wire [1023:0] dataGroup_hi_416 = {dataGroup_hi_hi_416, dataGroup_hi_lo_416};
  wire [7:0]    dataGroup_0_13 = dataGroup_lo_416[31:24];
  wire [1023:0] dataGroup_lo_417 = {dataGroup_lo_hi_417, dataGroup_lo_lo_417};
  wire [1023:0] dataGroup_hi_417 = {dataGroup_hi_hi_417, dataGroup_hi_lo_417};
  wire [7:0]    dataGroup_1_13 = dataGroup_lo_417[71:64];
  wire [1023:0] dataGroup_lo_418 = {dataGroup_lo_hi_418, dataGroup_lo_lo_418};
  wire [1023:0] dataGroup_hi_418 = {dataGroup_hi_hi_418, dataGroup_hi_lo_418};
  wire [7:0]    dataGroup_2_13 = dataGroup_lo_418[111:104];
  wire [1023:0] dataGroup_lo_419 = {dataGroup_lo_hi_419, dataGroup_lo_lo_419};
  wire [1023:0] dataGroup_hi_419 = {dataGroup_hi_hi_419, dataGroup_hi_lo_419};
  wire [7:0]    dataGroup_3_13 = dataGroup_lo_419[151:144];
  wire [1023:0] dataGroup_lo_420 = {dataGroup_lo_hi_420, dataGroup_lo_lo_420};
  wire [1023:0] dataGroup_hi_420 = {dataGroup_hi_hi_420, dataGroup_hi_lo_420};
  wire [7:0]    dataGroup_4_13 = dataGroup_lo_420[191:184];
  wire [1023:0] dataGroup_lo_421 = {dataGroup_lo_hi_421, dataGroup_lo_lo_421};
  wire [1023:0] dataGroup_hi_421 = {dataGroup_hi_hi_421, dataGroup_hi_lo_421};
  wire [7:0]    dataGroup_5_13 = dataGroup_lo_421[231:224];
  wire [1023:0] dataGroup_lo_422 = {dataGroup_lo_hi_422, dataGroup_lo_lo_422};
  wire [1023:0] dataGroup_hi_422 = {dataGroup_hi_hi_422, dataGroup_hi_lo_422};
  wire [7:0]    dataGroup_6_13 = dataGroup_lo_422[271:264];
  wire [1023:0] dataGroup_lo_423 = {dataGroup_lo_hi_423, dataGroup_lo_lo_423};
  wire [1023:0] dataGroup_hi_423 = {dataGroup_hi_hi_423, dataGroup_hi_lo_423};
  wire [7:0]    dataGroup_7_13 = dataGroup_lo_423[311:304];
  wire [1023:0] dataGroup_lo_424 = {dataGroup_lo_hi_424, dataGroup_lo_lo_424};
  wire [1023:0] dataGroup_hi_424 = {dataGroup_hi_hi_424, dataGroup_hi_lo_424};
  wire [7:0]    dataGroup_8_13 = dataGroup_lo_424[351:344];
  wire [1023:0] dataGroup_lo_425 = {dataGroup_lo_hi_425, dataGroup_lo_lo_425};
  wire [1023:0] dataGroup_hi_425 = {dataGroup_hi_hi_425, dataGroup_hi_lo_425};
  wire [7:0]    dataGroup_9_13 = dataGroup_lo_425[391:384];
  wire [1023:0] dataGroup_lo_426 = {dataGroup_lo_hi_426, dataGroup_lo_lo_426};
  wire [1023:0] dataGroup_hi_426 = {dataGroup_hi_hi_426, dataGroup_hi_lo_426};
  wire [7:0]    dataGroup_10_13 = dataGroup_lo_426[431:424];
  wire [1023:0] dataGroup_lo_427 = {dataGroup_lo_hi_427, dataGroup_lo_lo_427};
  wire [1023:0] dataGroup_hi_427 = {dataGroup_hi_hi_427, dataGroup_hi_lo_427};
  wire [7:0]    dataGroup_11_13 = dataGroup_lo_427[471:464];
  wire [1023:0] dataGroup_lo_428 = {dataGroup_lo_hi_428, dataGroup_lo_lo_428};
  wire [1023:0] dataGroup_hi_428 = {dataGroup_hi_hi_428, dataGroup_hi_lo_428};
  wire [7:0]    dataGroup_12_13 = dataGroup_lo_428[511:504];
  wire [1023:0] dataGroup_lo_429 = {dataGroup_lo_hi_429, dataGroup_lo_lo_429};
  wire [1023:0] dataGroup_hi_429 = {dataGroup_hi_hi_429, dataGroup_hi_lo_429};
  wire [7:0]    dataGroup_13_13 = dataGroup_lo_429[551:544];
  wire [1023:0] dataGroup_lo_430 = {dataGroup_lo_hi_430, dataGroup_lo_lo_430};
  wire [1023:0] dataGroup_hi_430 = {dataGroup_hi_hi_430, dataGroup_hi_lo_430};
  wire [7:0]    dataGroup_14_13 = dataGroup_lo_430[591:584];
  wire [1023:0] dataGroup_lo_431 = {dataGroup_lo_hi_431, dataGroup_lo_lo_431};
  wire [1023:0] dataGroup_hi_431 = {dataGroup_hi_hi_431, dataGroup_hi_lo_431};
  wire [7:0]    dataGroup_15_13 = dataGroup_lo_431[631:624];
  wire [1023:0] dataGroup_lo_432 = {dataGroup_lo_hi_432, dataGroup_lo_lo_432};
  wire [1023:0] dataGroup_hi_432 = {dataGroup_hi_hi_432, dataGroup_hi_lo_432};
  wire [7:0]    dataGroup_16_13 = dataGroup_lo_432[671:664];
  wire [1023:0] dataGroup_lo_433 = {dataGroup_lo_hi_433, dataGroup_lo_lo_433};
  wire [1023:0] dataGroup_hi_433 = {dataGroup_hi_hi_433, dataGroup_hi_lo_433};
  wire [7:0]    dataGroup_17_13 = dataGroup_lo_433[711:704];
  wire [1023:0] dataGroup_lo_434 = {dataGroup_lo_hi_434, dataGroup_lo_lo_434};
  wire [1023:0] dataGroup_hi_434 = {dataGroup_hi_hi_434, dataGroup_hi_lo_434};
  wire [7:0]    dataGroup_18_13 = dataGroup_lo_434[751:744];
  wire [1023:0] dataGroup_lo_435 = {dataGroup_lo_hi_435, dataGroup_lo_lo_435};
  wire [1023:0] dataGroup_hi_435 = {dataGroup_hi_hi_435, dataGroup_hi_lo_435};
  wire [7:0]    dataGroup_19_13 = dataGroup_lo_435[791:784];
  wire [1023:0] dataGroup_lo_436 = {dataGroup_lo_hi_436, dataGroup_lo_lo_436};
  wire [1023:0] dataGroup_hi_436 = {dataGroup_hi_hi_436, dataGroup_hi_lo_436};
  wire [7:0]    dataGroup_20_13 = dataGroup_lo_436[831:824];
  wire [1023:0] dataGroup_lo_437 = {dataGroup_lo_hi_437, dataGroup_lo_lo_437};
  wire [1023:0] dataGroup_hi_437 = {dataGroup_hi_hi_437, dataGroup_hi_lo_437};
  wire [7:0]    dataGroup_21_13 = dataGroup_lo_437[871:864];
  wire [1023:0] dataGroup_lo_438 = {dataGroup_lo_hi_438, dataGroup_lo_lo_438};
  wire [1023:0] dataGroup_hi_438 = {dataGroup_hi_hi_438, dataGroup_hi_lo_438};
  wire [7:0]    dataGroup_22_13 = dataGroup_lo_438[911:904];
  wire [1023:0] dataGroup_lo_439 = {dataGroup_lo_hi_439, dataGroup_lo_lo_439};
  wire [1023:0] dataGroup_hi_439 = {dataGroup_hi_hi_439, dataGroup_hi_lo_439};
  wire [7:0]    dataGroup_23_13 = dataGroup_lo_439[951:944];
  wire [1023:0] dataGroup_lo_440 = {dataGroup_lo_hi_440, dataGroup_lo_lo_440};
  wire [1023:0] dataGroup_hi_440 = {dataGroup_hi_hi_440, dataGroup_hi_lo_440};
  wire [7:0]    dataGroup_24_13 = dataGroup_lo_440[991:984];
  wire [1023:0] dataGroup_lo_441 = {dataGroup_lo_hi_441, dataGroup_lo_lo_441};
  wire [1023:0] dataGroup_hi_441 = {dataGroup_hi_hi_441, dataGroup_hi_lo_441};
  wire [7:0]    dataGroup_25_13 = dataGroup_hi_441[7:0];
  wire [1023:0] dataGroup_lo_442 = {dataGroup_lo_hi_442, dataGroup_lo_lo_442};
  wire [1023:0] dataGroup_hi_442 = {dataGroup_hi_hi_442, dataGroup_hi_lo_442};
  wire [7:0]    dataGroup_26_13 = dataGroup_hi_442[47:40];
  wire [1023:0] dataGroup_lo_443 = {dataGroup_lo_hi_443, dataGroup_lo_lo_443};
  wire [1023:0] dataGroup_hi_443 = {dataGroup_hi_hi_443, dataGroup_hi_lo_443};
  wire [7:0]    dataGroup_27_13 = dataGroup_hi_443[87:80];
  wire [1023:0] dataGroup_lo_444 = {dataGroup_lo_hi_444, dataGroup_lo_lo_444};
  wire [1023:0] dataGroup_hi_444 = {dataGroup_hi_hi_444, dataGroup_hi_lo_444};
  wire [7:0]    dataGroup_28_13 = dataGroup_hi_444[127:120];
  wire [1023:0] dataGroup_lo_445 = {dataGroup_lo_hi_445, dataGroup_lo_lo_445};
  wire [1023:0] dataGroup_hi_445 = {dataGroup_hi_hi_445, dataGroup_hi_lo_445};
  wire [7:0]    dataGroup_29_13 = dataGroup_hi_445[167:160];
  wire [1023:0] dataGroup_lo_446 = {dataGroup_lo_hi_446, dataGroup_lo_lo_446};
  wire [1023:0] dataGroup_hi_446 = {dataGroup_hi_hi_446, dataGroup_hi_lo_446};
  wire [7:0]    dataGroup_30_13 = dataGroup_hi_446[207:200];
  wire [1023:0] dataGroup_lo_447 = {dataGroup_lo_hi_447, dataGroup_lo_lo_447};
  wire [1023:0] dataGroup_hi_447 = {dataGroup_hi_hi_447, dataGroup_hi_lo_447};
  wire [7:0]    dataGroup_31_13 = dataGroup_hi_447[247:240];
  wire [15:0]   res_lo_lo_lo_lo_13 = {dataGroup_1_13, dataGroup_0_13};
  wire [15:0]   res_lo_lo_lo_hi_13 = {dataGroup_3_13, dataGroup_2_13};
  wire [31:0]   res_lo_lo_lo_13 = {res_lo_lo_lo_hi_13, res_lo_lo_lo_lo_13};
  wire [15:0]   res_lo_lo_hi_lo_13 = {dataGroup_5_13, dataGroup_4_13};
  wire [15:0]   res_lo_lo_hi_hi_13 = {dataGroup_7_13, dataGroup_6_13};
  wire [31:0]   res_lo_lo_hi_13 = {res_lo_lo_hi_hi_13, res_lo_lo_hi_lo_13};
  wire [63:0]   res_lo_lo_13 = {res_lo_lo_hi_13, res_lo_lo_lo_13};
  wire [15:0]   res_lo_hi_lo_lo_13 = {dataGroup_9_13, dataGroup_8_13};
  wire [15:0]   res_lo_hi_lo_hi_13 = {dataGroup_11_13, dataGroup_10_13};
  wire [31:0]   res_lo_hi_lo_13 = {res_lo_hi_lo_hi_13, res_lo_hi_lo_lo_13};
  wire [15:0]   res_lo_hi_hi_lo_13 = {dataGroup_13_13, dataGroup_12_13};
  wire [15:0]   res_lo_hi_hi_hi_13 = {dataGroup_15_13, dataGroup_14_13};
  wire [31:0]   res_lo_hi_hi_13 = {res_lo_hi_hi_hi_13, res_lo_hi_hi_lo_13};
  wire [63:0]   res_lo_hi_13 = {res_lo_hi_hi_13, res_lo_hi_lo_13};
  wire [127:0]  res_lo_13 = {res_lo_hi_13, res_lo_lo_13};
  wire [15:0]   res_hi_lo_lo_lo_13 = {dataGroup_17_13, dataGroup_16_13};
  wire [15:0]   res_hi_lo_lo_hi_13 = {dataGroup_19_13, dataGroup_18_13};
  wire [31:0]   res_hi_lo_lo_13 = {res_hi_lo_lo_hi_13, res_hi_lo_lo_lo_13};
  wire [15:0]   res_hi_lo_hi_lo_13 = {dataGroup_21_13, dataGroup_20_13};
  wire [15:0]   res_hi_lo_hi_hi_13 = {dataGroup_23_13, dataGroup_22_13};
  wire [31:0]   res_hi_lo_hi_13 = {res_hi_lo_hi_hi_13, res_hi_lo_hi_lo_13};
  wire [63:0]   res_hi_lo_13 = {res_hi_lo_hi_13, res_hi_lo_lo_13};
  wire [15:0]   res_hi_hi_lo_lo_13 = {dataGroup_25_13, dataGroup_24_13};
  wire [15:0]   res_hi_hi_lo_hi_13 = {dataGroup_27_13, dataGroup_26_13};
  wire [31:0]   res_hi_hi_lo_13 = {res_hi_hi_lo_hi_13, res_hi_hi_lo_lo_13};
  wire [15:0]   res_hi_hi_hi_lo_13 = {dataGroup_29_13, dataGroup_28_13};
  wire [15:0]   res_hi_hi_hi_hi_13 = {dataGroup_31_13, dataGroup_30_13};
  wire [31:0]   res_hi_hi_hi_13 = {res_hi_hi_hi_hi_13, res_hi_hi_hi_lo_13};
  wire [63:0]   res_hi_hi_13 = {res_hi_hi_hi_13, res_hi_hi_lo_13};
  wire [127:0]  res_hi_13 = {res_hi_hi_13, res_hi_lo_13};
  wire [255:0]  res_35 = {res_hi_13, res_lo_13};
  wire [1023:0] dataGroup_lo_448 = {dataGroup_lo_hi_448, dataGroup_lo_lo_448};
  wire [1023:0] dataGroup_hi_448 = {dataGroup_hi_hi_448, dataGroup_hi_lo_448};
  wire [7:0]    dataGroup_0_14 = dataGroup_lo_448[39:32];
  wire [1023:0] dataGroup_lo_449 = {dataGroup_lo_hi_449, dataGroup_lo_lo_449};
  wire [1023:0] dataGroup_hi_449 = {dataGroup_hi_hi_449, dataGroup_hi_lo_449};
  wire [7:0]    dataGroup_1_14 = dataGroup_lo_449[79:72];
  wire [1023:0] dataGroup_lo_450 = {dataGroup_lo_hi_450, dataGroup_lo_lo_450};
  wire [1023:0] dataGroup_hi_450 = {dataGroup_hi_hi_450, dataGroup_hi_lo_450};
  wire [7:0]    dataGroup_2_14 = dataGroup_lo_450[119:112];
  wire [1023:0] dataGroup_lo_451 = {dataGroup_lo_hi_451, dataGroup_lo_lo_451};
  wire [1023:0] dataGroup_hi_451 = {dataGroup_hi_hi_451, dataGroup_hi_lo_451};
  wire [7:0]    dataGroup_3_14 = dataGroup_lo_451[159:152];
  wire [1023:0] dataGroup_lo_452 = {dataGroup_lo_hi_452, dataGroup_lo_lo_452};
  wire [1023:0] dataGroup_hi_452 = {dataGroup_hi_hi_452, dataGroup_hi_lo_452};
  wire [7:0]    dataGroup_4_14 = dataGroup_lo_452[199:192];
  wire [1023:0] dataGroup_lo_453 = {dataGroup_lo_hi_453, dataGroup_lo_lo_453};
  wire [1023:0] dataGroup_hi_453 = {dataGroup_hi_hi_453, dataGroup_hi_lo_453};
  wire [7:0]    dataGroup_5_14 = dataGroup_lo_453[239:232];
  wire [1023:0] dataGroup_lo_454 = {dataGroup_lo_hi_454, dataGroup_lo_lo_454};
  wire [1023:0] dataGroup_hi_454 = {dataGroup_hi_hi_454, dataGroup_hi_lo_454};
  wire [7:0]    dataGroup_6_14 = dataGroup_lo_454[279:272];
  wire [1023:0] dataGroup_lo_455 = {dataGroup_lo_hi_455, dataGroup_lo_lo_455};
  wire [1023:0] dataGroup_hi_455 = {dataGroup_hi_hi_455, dataGroup_hi_lo_455};
  wire [7:0]    dataGroup_7_14 = dataGroup_lo_455[319:312];
  wire [1023:0] dataGroup_lo_456 = {dataGroup_lo_hi_456, dataGroup_lo_lo_456};
  wire [1023:0] dataGroup_hi_456 = {dataGroup_hi_hi_456, dataGroup_hi_lo_456};
  wire [7:0]    dataGroup_8_14 = dataGroup_lo_456[359:352];
  wire [1023:0] dataGroup_lo_457 = {dataGroup_lo_hi_457, dataGroup_lo_lo_457};
  wire [1023:0] dataGroup_hi_457 = {dataGroup_hi_hi_457, dataGroup_hi_lo_457};
  wire [7:0]    dataGroup_9_14 = dataGroup_lo_457[399:392];
  wire [1023:0] dataGroup_lo_458 = {dataGroup_lo_hi_458, dataGroup_lo_lo_458};
  wire [1023:0] dataGroup_hi_458 = {dataGroup_hi_hi_458, dataGroup_hi_lo_458};
  wire [7:0]    dataGroup_10_14 = dataGroup_lo_458[439:432];
  wire [1023:0] dataGroup_lo_459 = {dataGroup_lo_hi_459, dataGroup_lo_lo_459};
  wire [1023:0] dataGroup_hi_459 = {dataGroup_hi_hi_459, dataGroup_hi_lo_459};
  wire [7:0]    dataGroup_11_14 = dataGroup_lo_459[479:472];
  wire [1023:0] dataGroup_lo_460 = {dataGroup_lo_hi_460, dataGroup_lo_lo_460};
  wire [1023:0] dataGroup_hi_460 = {dataGroup_hi_hi_460, dataGroup_hi_lo_460};
  wire [7:0]    dataGroup_12_14 = dataGroup_lo_460[519:512];
  wire [1023:0] dataGroup_lo_461 = {dataGroup_lo_hi_461, dataGroup_lo_lo_461};
  wire [1023:0] dataGroup_hi_461 = {dataGroup_hi_hi_461, dataGroup_hi_lo_461};
  wire [7:0]    dataGroup_13_14 = dataGroup_lo_461[559:552];
  wire [1023:0] dataGroup_lo_462 = {dataGroup_lo_hi_462, dataGroup_lo_lo_462};
  wire [1023:0] dataGroup_hi_462 = {dataGroup_hi_hi_462, dataGroup_hi_lo_462};
  wire [7:0]    dataGroup_14_14 = dataGroup_lo_462[599:592];
  wire [1023:0] dataGroup_lo_463 = {dataGroup_lo_hi_463, dataGroup_lo_lo_463};
  wire [1023:0] dataGroup_hi_463 = {dataGroup_hi_hi_463, dataGroup_hi_lo_463};
  wire [7:0]    dataGroup_15_14 = dataGroup_lo_463[639:632];
  wire [1023:0] dataGroup_lo_464 = {dataGroup_lo_hi_464, dataGroup_lo_lo_464};
  wire [1023:0] dataGroup_hi_464 = {dataGroup_hi_hi_464, dataGroup_hi_lo_464};
  wire [7:0]    dataGroup_16_14 = dataGroup_lo_464[679:672];
  wire [1023:0] dataGroup_lo_465 = {dataGroup_lo_hi_465, dataGroup_lo_lo_465};
  wire [1023:0] dataGroup_hi_465 = {dataGroup_hi_hi_465, dataGroup_hi_lo_465};
  wire [7:0]    dataGroup_17_14 = dataGroup_lo_465[719:712];
  wire [1023:0] dataGroup_lo_466 = {dataGroup_lo_hi_466, dataGroup_lo_lo_466};
  wire [1023:0] dataGroup_hi_466 = {dataGroup_hi_hi_466, dataGroup_hi_lo_466};
  wire [7:0]    dataGroup_18_14 = dataGroup_lo_466[759:752];
  wire [1023:0] dataGroup_lo_467 = {dataGroup_lo_hi_467, dataGroup_lo_lo_467};
  wire [1023:0] dataGroup_hi_467 = {dataGroup_hi_hi_467, dataGroup_hi_lo_467};
  wire [7:0]    dataGroup_19_14 = dataGroup_lo_467[799:792];
  wire [1023:0] dataGroup_lo_468 = {dataGroup_lo_hi_468, dataGroup_lo_lo_468};
  wire [1023:0] dataGroup_hi_468 = {dataGroup_hi_hi_468, dataGroup_hi_lo_468};
  wire [7:0]    dataGroup_20_14 = dataGroup_lo_468[839:832];
  wire [1023:0] dataGroup_lo_469 = {dataGroup_lo_hi_469, dataGroup_lo_lo_469};
  wire [1023:0] dataGroup_hi_469 = {dataGroup_hi_hi_469, dataGroup_hi_lo_469};
  wire [7:0]    dataGroup_21_14 = dataGroup_lo_469[879:872];
  wire [1023:0] dataGroup_lo_470 = {dataGroup_lo_hi_470, dataGroup_lo_lo_470};
  wire [1023:0] dataGroup_hi_470 = {dataGroup_hi_hi_470, dataGroup_hi_lo_470};
  wire [7:0]    dataGroup_22_14 = dataGroup_lo_470[919:912];
  wire [1023:0] dataGroup_lo_471 = {dataGroup_lo_hi_471, dataGroup_lo_lo_471};
  wire [1023:0] dataGroup_hi_471 = {dataGroup_hi_hi_471, dataGroup_hi_lo_471};
  wire [7:0]    dataGroup_23_14 = dataGroup_lo_471[959:952];
  wire [1023:0] dataGroup_lo_472 = {dataGroup_lo_hi_472, dataGroup_lo_lo_472};
  wire [1023:0] dataGroup_hi_472 = {dataGroup_hi_hi_472, dataGroup_hi_lo_472};
  wire [7:0]    dataGroup_24_14 = dataGroup_lo_472[999:992];
  wire [1023:0] dataGroup_lo_473 = {dataGroup_lo_hi_473, dataGroup_lo_lo_473};
  wire [1023:0] dataGroup_hi_473 = {dataGroup_hi_hi_473, dataGroup_hi_lo_473};
  wire [7:0]    dataGroup_25_14 = dataGroup_hi_473[15:8];
  wire [1023:0] dataGroup_lo_474 = {dataGroup_lo_hi_474, dataGroup_lo_lo_474};
  wire [1023:0] dataGroup_hi_474 = {dataGroup_hi_hi_474, dataGroup_hi_lo_474};
  wire [7:0]    dataGroup_26_14 = dataGroup_hi_474[55:48];
  wire [1023:0] dataGroup_lo_475 = {dataGroup_lo_hi_475, dataGroup_lo_lo_475};
  wire [1023:0] dataGroup_hi_475 = {dataGroup_hi_hi_475, dataGroup_hi_lo_475};
  wire [7:0]    dataGroup_27_14 = dataGroup_hi_475[95:88];
  wire [1023:0] dataGroup_lo_476 = {dataGroup_lo_hi_476, dataGroup_lo_lo_476};
  wire [1023:0] dataGroup_hi_476 = {dataGroup_hi_hi_476, dataGroup_hi_lo_476};
  wire [7:0]    dataGroup_28_14 = dataGroup_hi_476[135:128];
  wire [1023:0] dataGroup_lo_477 = {dataGroup_lo_hi_477, dataGroup_lo_lo_477};
  wire [1023:0] dataGroup_hi_477 = {dataGroup_hi_hi_477, dataGroup_hi_lo_477};
  wire [7:0]    dataGroup_29_14 = dataGroup_hi_477[175:168];
  wire [1023:0] dataGroup_lo_478 = {dataGroup_lo_hi_478, dataGroup_lo_lo_478};
  wire [1023:0] dataGroup_hi_478 = {dataGroup_hi_hi_478, dataGroup_hi_lo_478};
  wire [7:0]    dataGroup_30_14 = dataGroup_hi_478[215:208];
  wire [1023:0] dataGroup_lo_479 = {dataGroup_lo_hi_479, dataGroup_lo_lo_479};
  wire [1023:0] dataGroup_hi_479 = {dataGroup_hi_hi_479, dataGroup_hi_lo_479};
  wire [7:0]    dataGroup_31_14 = dataGroup_hi_479[255:248];
  wire [15:0]   res_lo_lo_lo_lo_14 = {dataGroup_1_14, dataGroup_0_14};
  wire [15:0]   res_lo_lo_lo_hi_14 = {dataGroup_3_14, dataGroup_2_14};
  wire [31:0]   res_lo_lo_lo_14 = {res_lo_lo_lo_hi_14, res_lo_lo_lo_lo_14};
  wire [15:0]   res_lo_lo_hi_lo_14 = {dataGroup_5_14, dataGroup_4_14};
  wire [15:0]   res_lo_lo_hi_hi_14 = {dataGroup_7_14, dataGroup_6_14};
  wire [31:0]   res_lo_lo_hi_14 = {res_lo_lo_hi_hi_14, res_lo_lo_hi_lo_14};
  wire [63:0]   res_lo_lo_14 = {res_lo_lo_hi_14, res_lo_lo_lo_14};
  wire [15:0]   res_lo_hi_lo_lo_14 = {dataGroup_9_14, dataGroup_8_14};
  wire [15:0]   res_lo_hi_lo_hi_14 = {dataGroup_11_14, dataGroup_10_14};
  wire [31:0]   res_lo_hi_lo_14 = {res_lo_hi_lo_hi_14, res_lo_hi_lo_lo_14};
  wire [15:0]   res_lo_hi_hi_lo_14 = {dataGroup_13_14, dataGroup_12_14};
  wire [15:0]   res_lo_hi_hi_hi_14 = {dataGroup_15_14, dataGroup_14_14};
  wire [31:0]   res_lo_hi_hi_14 = {res_lo_hi_hi_hi_14, res_lo_hi_hi_lo_14};
  wire [63:0]   res_lo_hi_14 = {res_lo_hi_hi_14, res_lo_hi_lo_14};
  wire [127:0]  res_lo_14 = {res_lo_hi_14, res_lo_lo_14};
  wire [15:0]   res_hi_lo_lo_lo_14 = {dataGroup_17_14, dataGroup_16_14};
  wire [15:0]   res_hi_lo_lo_hi_14 = {dataGroup_19_14, dataGroup_18_14};
  wire [31:0]   res_hi_lo_lo_14 = {res_hi_lo_lo_hi_14, res_hi_lo_lo_lo_14};
  wire [15:0]   res_hi_lo_hi_lo_14 = {dataGroup_21_14, dataGroup_20_14};
  wire [15:0]   res_hi_lo_hi_hi_14 = {dataGroup_23_14, dataGroup_22_14};
  wire [31:0]   res_hi_lo_hi_14 = {res_hi_lo_hi_hi_14, res_hi_lo_hi_lo_14};
  wire [63:0]   res_hi_lo_14 = {res_hi_lo_hi_14, res_hi_lo_lo_14};
  wire [15:0]   res_hi_hi_lo_lo_14 = {dataGroup_25_14, dataGroup_24_14};
  wire [15:0]   res_hi_hi_lo_hi_14 = {dataGroup_27_14, dataGroup_26_14};
  wire [31:0]   res_hi_hi_lo_14 = {res_hi_hi_lo_hi_14, res_hi_hi_lo_lo_14};
  wire [15:0]   res_hi_hi_hi_lo_14 = {dataGroup_29_14, dataGroup_28_14};
  wire [15:0]   res_hi_hi_hi_hi_14 = {dataGroup_31_14, dataGroup_30_14};
  wire [31:0]   res_hi_hi_hi_14 = {res_hi_hi_hi_hi_14, res_hi_hi_hi_lo_14};
  wire [63:0]   res_hi_hi_14 = {res_hi_hi_hi_14, res_hi_hi_lo_14};
  wire [127:0]  res_hi_14 = {res_hi_hi_14, res_hi_lo_14};
  wire [255:0]  res_36 = {res_hi_14, res_lo_14};
  wire [511:0]  lo_lo_4 = {res_33, res_32};
  wire [511:0]  lo_hi_4 = {res_35, res_34};
  wire [1023:0] lo_4 = {lo_hi_4, lo_lo_4};
  wire [511:0]  hi_lo_4 = {256'h0, res_36};
  wire [1023:0] hi_4 = {512'h0, hi_lo_4};
  wire [2047:0] regroupLoadData_0_4 = {hi_4, lo_4};
  wire [1023:0] dataGroup_lo_480 = {dataGroup_lo_hi_480, dataGroup_lo_lo_480};
  wire [1023:0] dataGroup_hi_480 = {dataGroup_hi_hi_480, dataGroup_hi_lo_480};
  wire [7:0]    dataGroup_0_15 = dataGroup_lo_480[7:0];
  wire [1023:0] dataGroup_lo_481 = {dataGroup_lo_hi_481, dataGroup_lo_lo_481};
  wire [1023:0] dataGroup_hi_481 = {dataGroup_hi_hi_481, dataGroup_hi_lo_481};
  wire [7:0]    dataGroup_1_15 = dataGroup_lo_481[55:48];
  wire [1023:0] dataGroup_lo_482 = {dataGroup_lo_hi_482, dataGroup_lo_lo_482};
  wire [1023:0] dataGroup_hi_482 = {dataGroup_hi_hi_482, dataGroup_hi_lo_482};
  wire [7:0]    dataGroup_2_15 = dataGroup_lo_482[103:96];
  wire [1023:0] dataGroup_lo_483 = {dataGroup_lo_hi_483, dataGroup_lo_lo_483};
  wire [1023:0] dataGroup_hi_483 = {dataGroup_hi_hi_483, dataGroup_hi_lo_483};
  wire [7:0]    dataGroup_3_15 = dataGroup_lo_483[151:144];
  wire [1023:0] dataGroup_lo_484 = {dataGroup_lo_hi_484, dataGroup_lo_lo_484};
  wire [1023:0] dataGroup_hi_484 = {dataGroup_hi_hi_484, dataGroup_hi_lo_484};
  wire [7:0]    dataGroup_4_15 = dataGroup_lo_484[199:192];
  wire [1023:0] dataGroup_lo_485 = {dataGroup_lo_hi_485, dataGroup_lo_lo_485};
  wire [1023:0] dataGroup_hi_485 = {dataGroup_hi_hi_485, dataGroup_hi_lo_485};
  wire [7:0]    dataGroup_5_15 = dataGroup_lo_485[247:240];
  wire [1023:0] dataGroup_lo_486 = {dataGroup_lo_hi_486, dataGroup_lo_lo_486};
  wire [1023:0] dataGroup_hi_486 = {dataGroup_hi_hi_486, dataGroup_hi_lo_486};
  wire [7:0]    dataGroup_6_15 = dataGroup_lo_486[295:288];
  wire [1023:0] dataGroup_lo_487 = {dataGroup_lo_hi_487, dataGroup_lo_lo_487};
  wire [1023:0] dataGroup_hi_487 = {dataGroup_hi_hi_487, dataGroup_hi_lo_487};
  wire [7:0]    dataGroup_7_15 = dataGroup_lo_487[343:336];
  wire [1023:0] dataGroup_lo_488 = {dataGroup_lo_hi_488, dataGroup_lo_lo_488};
  wire [1023:0] dataGroup_hi_488 = {dataGroup_hi_hi_488, dataGroup_hi_lo_488};
  wire [7:0]    dataGroup_8_15 = dataGroup_lo_488[391:384];
  wire [1023:0] dataGroup_lo_489 = {dataGroup_lo_hi_489, dataGroup_lo_lo_489};
  wire [1023:0] dataGroup_hi_489 = {dataGroup_hi_hi_489, dataGroup_hi_lo_489};
  wire [7:0]    dataGroup_9_15 = dataGroup_lo_489[439:432];
  wire [1023:0] dataGroup_lo_490 = {dataGroup_lo_hi_490, dataGroup_lo_lo_490};
  wire [1023:0] dataGroup_hi_490 = {dataGroup_hi_hi_490, dataGroup_hi_lo_490};
  wire [7:0]    dataGroup_10_15 = dataGroup_lo_490[487:480];
  wire [1023:0] dataGroup_lo_491 = {dataGroup_lo_hi_491, dataGroup_lo_lo_491};
  wire [1023:0] dataGroup_hi_491 = {dataGroup_hi_hi_491, dataGroup_hi_lo_491};
  wire [7:0]    dataGroup_11_15 = dataGroup_lo_491[535:528];
  wire [1023:0] dataGroup_lo_492 = {dataGroup_lo_hi_492, dataGroup_lo_lo_492};
  wire [1023:0] dataGroup_hi_492 = {dataGroup_hi_hi_492, dataGroup_hi_lo_492};
  wire [7:0]    dataGroup_12_15 = dataGroup_lo_492[583:576];
  wire [1023:0] dataGroup_lo_493 = {dataGroup_lo_hi_493, dataGroup_lo_lo_493};
  wire [1023:0] dataGroup_hi_493 = {dataGroup_hi_hi_493, dataGroup_hi_lo_493};
  wire [7:0]    dataGroup_13_15 = dataGroup_lo_493[631:624];
  wire [1023:0] dataGroup_lo_494 = {dataGroup_lo_hi_494, dataGroup_lo_lo_494};
  wire [1023:0] dataGroup_hi_494 = {dataGroup_hi_hi_494, dataGroup_hi_lo_494};
  wire [7:0]    dataGroup_14_15 = dataGroup_lo_494[679:672];
  wire [1023:0] dataGroup_lo_495 = {dataGroup_lo_hi_495, dataGroup_lo_lo_495};
  wire [1023:0] dataGroup_hi_495 = {dataGroup_hi_hi_495, dataGroup_hi_lo_495};
  wire [7:0]    dataGroup_15_15 = dataGroup_lo_495[727:720];
  wire [1023:0] dataGroup_lo_496 = {dataGroup_lo_hi_496, dataGroup_lo_lo_496};
  wire [1023:0] dataGroup_hi_496 = {dataGroup_hi_hi_496, dataGroup_hi_lo_496};
  wire [7:0]    dataGroup_16_15 = dataGroup_lo_496[775:768];
  wire [1023:0] dataGroup_lo_497 = {dataGroup_lo_hi_497, dataGroup_lo_lo_497};
  wire [1023:0] dataGroup_hi_497 = {dataGroup_hi_hi_497, dataGroup_hi_lo_497};
  wire [7:0]    dataGroup_17_15 = dataGroup_lo_497[823:816];
  wire [1023:0] dataGroup_lo_498 = {dataGroup_lo_hi_498, dataGroup_lo_lo_498};
  wire [1023:0] dataGroup_hi_498 = {dataGroup_hi_hi_498, dataGroup_hi_lo_498};
  wire [7:0]    dataGroup_18_15 = dataGroup_lo_498[871:864];
  wire [1023:0] dataGroup_lo_499 = {dataGroup_lo_hi_499, dataGroup_lo_lo_499};
  wire [1023:0] dataGroup_hi_499 = {dataGroup_hi_hi_499, dataGroup_hi_lo_499};
  wire [7:0]    dataGroup_19_15 = dataGroup_lo_499[919:912];
  wire [1023:0] dataGroup_lo_500 = {dataGroup_lo_hi_500, dataGroup_lo_lo_500};
  wire [1023:0] dataGroup_hi_500 = {dataGroup_hi_hi_500, dataGroup_hi_lo_500};
  wire [7:0]    dataGroup_20_15 = dataGroup_lo_500[967:960];
  wire [1023:0] dataGroup_lo_501 = {dataGroup_lo_hi_501, dataGroup_lo_lo_501};
  wire [1023:0] dataGroup_hi_501 = {dataGroup_hi_hi_501, dataGroup_hi_lo_501};
  wire [7:0]    dataGroup_21_15 = dataGroup_lo_501[1015:1008];
  wire [1023:0] dataGroup_lo_502 = {dataGroup_lo_hi_502, dataGroup_lo_lo_502};
  wire [1023:0] dataGroup_hi_502 = {dataGroup_hi_hi_502, dataGroup_hi_lo_502};
  wire [7:0]    dataGroup_22_15 = dataGroup_hi_502[39:32];
  wire [1023:0] dataGroup_lo_503 = {dataGroup_lo_hi_503, dataGroup_lo_lo_503};
  wire [1023:0] dataGroup_hi_503 = {dataGroup_hi_hi_503, dataGroup_hi_lo_503};
  wire [7:0]    dataGroup_23_15 = dataGroup_hi_503[87:80];
  wire [1023:0] dataGroup_lo_504 = {dataGroup_lo_hi_504, dataGroup_lo_lo_504};
  wire [1023:0] dataGroup_hi_504 = {dataGroup_hi_hi_504, dataGroup_hi_lo_504};
  wire [7:0]    dataGroup_24_15 = dataGroup_hi_504[135:128];
  wire [1023:0] dataGroup_lo_505 = {dataGroup_lo_hi_505, dataGroup_lo_lo_505};
  wire [1023:0] dataGroup_hi_505 = {dataGroup_hi_hi_505, dataGroup_hi_lo_505};
  wire [7:0]    dataGroup_25_15 = dataGroup_hi_505[183:176];
  wire [1023:0] dataGroup_lo_506 = {dataGroup_lo_hi_506, dataGroup_lo_lo_506};
  wire [1023:0] dataGroup_hi_506 = {dataGroup_hi_hi_506, dataGroup_hi_lo_506};
  wire [7:0]    dataGroup_26_15 = dataGroup_hi_506[231:224];
  wire [1023:0] dataGroup_lo_507 = {dataGroup_lo_hi_507, dataGroup_lo_lo_507};
  wire [1023:0] dataGroup_hi_507 = {dataGroup_hi_hi_507, dataGroup_hi_lo_507};
  wire [7:0]    dataGroup_27_15 = dataGroup_hi_507[279:272];
  wire [1023:0] dataGroup_lo_508 = {dataGroup_lo_hi_508, dataGroup_lo_lo_508};
  wire [1023:0] dataGroup_hi_508 = {dataGroup_hi_hi_508, dataGroup_hi_lo_508};
  wire [7:0]    dataGroup_28_15 = dataGroup_hi_508[327:320];
  wire [1023:0] dataGroup_lo_509 = {dataGroup_lo_hi_509, dataGroup_lo_lo_509};
  wire [1023:0] dataGroup_hi_509 = {dataGroup_hi_hi_509, dataGroup_hi_lo_509};
  wire [7:0]    dataGroup_29_15 = dataGroup_hi_509[375:368];
  wire [1023:0] dataGroup_lo_510 = {dataGroup_lo_hi_510, dataGroup_lo_lo_510};
  wire [1023:0] dataGroup_hi_510 = {dataGroup_hi_hi_510, dataGroup_hi_lo_510};
  wire [7:0]    dataGroup_30_15 = dataGroup_hi_510[423:416];
  wire [1023:0] dataGroup_lo_511 = {dataGroup_lo_hi_511, dataGroup_lo_lo_511};
  wire [1023:0] dataGroup_hi_511 = {dataGroup_hi_hi_511, dataGroup_hi_lo_511};
  wire [7:0]    dataGroup_31_15 = dataGroup_hi_511[471:464];
  wire [15:0]   res_lo_lo_lo_lo_15 = {dataGroup_1_15, dataGroup_0_15};
  wire [15:0]   res_lo_lo_lo_hi_15 = {dataGroup_3_15, dataGroup_2_15};
  wire [31:0]   res_lo_lo_lo_15 = {res_lo_lo_lo_hi_15, res_lo_lo_lo_lo_15};
  wire [15:0]   res_lo_lo_hi_lo_15 = {dataGroup_5_15, dataGroup_4_15};
  wire [15:0]   res_lo_lo_hi_hi_15 = {dataGroup_7_15, dataGroup_6_15};
  wire [31:0]   res_lo_lo_hi_15 = {res_lo_lo_hi_hi_15, res_lo_lo_hi_lo_15};
  wire [63:0]   res_lo_lo_15 = {res_lo_lo_hi_15, res_lo_lo_lo_15};
  wire [15:0]   res_lo_hi_lo_lo_15 = {dataGroup_9_15, dataGroup_8_15};
  wire [15:0]   res_lo_hi_lo_hi_15 = {dataGroup_11_15, dataGroup_10_15};
  wire [31:0]   res_lo_hi_lo_15 = {res_lo_hi_lo_hi_15, res_lo_hi_lo_lo_15};
  wire [15:0]   res_lo_hi_hi_lo_15 = {dataGroup_13_15, dataGroup_12_15};
  wire [15:0]   res_lo_hi_hi_hi_15 = {dataGroup_15_15, dataGroup_14_15};
  wire [31:0]   res_lo_hi_hi_15 = {res_lo_hi_hi_hi_15, res_lo_hi_hi_lo_15};
  wire [63:0]   res_lo_hi_15 = {res_lo_hi_hi_15, res_lo_hi_lo_15};
  wire [127:0]  res_lo_15 = {res_lo_hi_15, res_lo_lo_15};
  wire [15:0]   res_hi_lo_lo_lo_15 = {dataGroup_17_15, dataGroup_16_15};
  wire [15:0]   res_hi_lo_lo_hi_15 = {dataGroup_19_15, dataGroup_18_15};
  wire [31:0]   res_hi_lo_lo_15 = {res_hi_lo_lo_hi_15, res_hi_lo_lo_lo_15};
  wire [15:0]   res_hi_lo_hi_lo_15 = {dataGroup_21_15, dataGroup_20_15};
  wire [15:0]   res_hi_lo_hi_hi_15 = {dataGroup_23_15, dataGroup_22_15};
  wire [31:0]   res_hi_lo_hi_15 = {res_hi_lo_hi_hi_15, res_hi_lo_hi_lo_15};
  wire [63:0]   res_hi_lo_15 = {res_hi_lo_hi_15, res_hi_lo_lo_15};
  wire [15:0]   res_hi_hi_lo_lo_15 = {dataGroup_25_15, dataGroup_24_15};
  wire [15:0]   res_hi_hi_lo_hi_15 = {dataGroup_27_15, dataGroup_26_15};
  wire [31:0]   res_hi_hi_lo_15 = {res_hi_hi_lo_hi_15, res_hi_hi_lo_lo_15};
  wire [15:0]   res_hi_hi_hi_lo_15 = {dataGroup_29_15, dataGroup_28_15};
  wire [15:0]   res_hi_hi_hi_hi_15 = {dataGroup_31_15, dataGroup_30_15};
  wire [31:0]   res_hi_hi_hi_15 = {res_hi_hi_hi_hi_15, res_hi_hi_hi_lo_15};
  wire [63:0]   res_hi_hi_15 = {res_hi_hi_hi_15, res_hi_hi_lo_15};
  wire [127:0]  res_hi_15 = {res_hi_hi_15, res_hi_lo_15};
  wire [255:0]  res_40 = {res_hi_15, res_lo_15};
  wire [1023:0] dataGroup_lo_512 = {dataGroup_lo_hi_512, dataGroup_lo_lo_512};
  wire [1023:0] dataGroup_hi_512 = {dataGroup_hi_hi_512, dataGroup_hi_lo_512};
  wire [7:0]    dataGroup_0_16 = dataGroup_lo_512[15:8];
  wire [1023:0] dataGroup_lo_513 = {dataGroup_lo_hi_513, dataGroup_lo_lo_513};
  wire [1023:0] dataGroup_hi_513 = {dataGroup_hi_hi_513, dataGroup_hi_lo_513};
  wire [7:0]    dataGroup_1_16 = dataGroup_lo_513[63:56];
  wire [1023:0] dataGroup_lo_514 = {dataGroup_lo_hi_514, dataGroup_lo_lo_514};
  wire [1023:0] dataGroup_hi_514 = {dataGroup_hi_hi_514, dataGroup_hi_lo_514};
  wire [7:0]    dataGroup_2_16 = dataGroup_lo_514[111:104];
  wire [1023:0] dataGroup_lo_515 = {dataGroup_lo_hi_515, dataGroup_lo_lo_515};
  wire [1023:0] dataGroup_hi_515 = {dataGroup_hi_hi_515, dataGroup_hi_lo_515};
  wire [7:0]    dataGroup_3_16 = dataGroup_lo_515[159:152];
  wire [1023:0] dataGroup_lo_516 = {dataGroup_lo_hi_516, dataGroup_lo_lo_516};
  wire [1023:0] dataGroup_hi_516 = {dataGroup_hi_hi_516, dataGroup_hi_lo_516};
  wire [7:0]    dataGroup_4_16 = dataGroup_lo_516[207:200];
  wire [1023:0] dataGroup_lo_517 = {dataGroup_lo_hi_517, dataGroup_lo_lo_517};
  wire [1023:0] dataGroup_hi_517 = {dataGroup_hi_hi_517, dataGroup_hi_lo_517};
  wire [7:0]    dataGroup_5_16 = dataGroup_lo_517[255:248];
  wire [1023:0] dataGroup_lo_518 = {dataGroup_lo_hi_518, dataGroup_lo_lo_518};
  wire [1023:0] dataGroup_hi_518 = {dataGroup_hi_hi_518, dataGroup_hi_lo_518};
  wire [7:0]    dataGroup_6_16 = dataGroup_lo_518[303:296];
  wire [1023:0] dataGroup_lo_519 = {dataGroup_lo_hi_519, dataGroup_lo_lo_519};
  wire [1023:0] dataGroup_hi_519 = {dataGroup_hi_hi_519, dataGroup_hi_lo_519};
  wire [7:0]    dataGroup_7_16 = dataGroup_lo_519[351:344];
  wire [1023:0] dataGroup_lo_520 = {dataGroup_lo_hi_520, dataGroup_lo_lo_520};
  wire [1023:0] dataGroup_hi_520 = {dataGroup_hi_hi_520, dataGroup_hi_lo_520};
  wire [7:0]    dataGroup_8_16 = dataGroup_lo_520[399:392];
  wire [1023:0] dataGroup_lo_521 = {dataGroup_lo_hi_521, dataGroup_lo_lo_521};
  wire [1023:0] dataGroup_hi_521 = {dataGroup_hi_hi_521, dataGroup_hi_lo_521};
  wire [7:0]    dataGroup_9_16 = dataGroup_lo_521[447:440];
  wire [1023:0] dataGroup_lo_522 = {dataGroup_lo_hi_522, dataGroup_lo_lo_522};
  wire [1023:0] dataGroup_hi_522 = {dataGroup_hi_hi_522, dataGroup_hi_lo_522};
  wire [7:0]    dataGroup_10_16 = dataGroup_lo_522[495:488];
  wire [1023:0] dataGroup_lo_523 = {dataGroup_lo_hi_523, dataGroup_lo_lo_523};
  wire [1023:0] dataGroup_hi_523 = {dataGroup_hi_hi_523, dataGroup_hi_lo_523};
  wire [7:0]    dataGroup_11_16 = dataGroup_lo_523[543:536];
  wire [1023:0] dataGroup_lo_524 = {dataGroup_lo_hi_524, dataGroup_lo_lo_524};
  wire [1023:0] dataGroup_hi_524 = {dataGroup_hi_hi_524, dataGroup_hi_lo_524};
  wire [7:0]    dataGroup_12_16 = dataGroup_lo_524[591:584];
  wire [1023:0] dataGroup_lo_525 = {dataGroup_lo_hi_525, dataGroup_lo_lo_525};
  wire [1023:0] dataGroup_hi_525 = {dataGroup_hi_hi_525, dataGroup_hi_lo_525};
  wire [7:0]    dataGroup_13_16 = dataGroup_lo_525[639:632];
  wire [1023:0] dataGroup_lo_526 = {dataGroup_lo_hi_526, dataGroup_lo_lo_526};
  wire [1023:0] dataGroup_hi_526 = {dataGroup_hi_hi_526, dataGroup_hi_lo_526};
  wire [7:0]    dataGroup_14_16 = dataGroup_lo_526[687:680];
  wire [1023:0] dataGroup_lo_527 = {dataGroup_lo_hi_527, dataGroup_lo_lo_527};
  wire [1023:0] dataGroup_hi_527 = {dataGroup_hi_hi_527, dataGroup_hi_lo_527};
  wire [7:0]    dataGroup_15_16 = dataGroup_lo_527[735:728];
  wire [1023:0] dataGroup_lo_528 = {dataGroup_lo_hi_528, dataGroup_lo_lo_528};
  wire [1023:0] dataGroup_hi_528 = {dataGroup_hi_hi_528, dataGroup_hi_lo_528};
  wire [7:0]    dataGroup_16_16 = dataGroup_lo_528[783:776];
  wire [1023:0] dataGroup_lo_529 = {dataGroup_lo_hi_529, dataGroup_lo_lo_529};
  wire [1023:0] dataGroup_hi_529 = {dataGroup_hi_hi_529, dataGroup_hi_lo_529};
  wire [7:0]    dataGroup_17_16 = dataGroup_lo_529[831:824];
  wire [1023:0] dataGroup_lo_530 = {dataGroup_lo_hi_530, dataGroup_lo_lo_530};
  wire [1023:0] dataGroup_hi_530 = {dataGroup_hi_hi_530, dataGroup_hi_lo_530};
  wire [7:0]    dataGroup_18_16 = dataGroup_lo_530[879:872];
  wire [1023:0] dataGroup_lo_531 = {dataGroup_lo_hi_531, dataGroup_lo_lo_531};
  wire [1023:0] dataGroup_hi_531 = {dataGroup_hi_hi_531, dataGroup_hi_lo_531};
  wire [7:0]    dataGroup_19_16 = dataGroup_lo_531[927:920];
  wire [1023:0] dataGroup_lo_532 = {dataGroup_lo_hi_532, dataGroup_lo_lo_532};
  wire [1023:0] dataGroup_hi_532 = {dataGroup_hi_hi_532, dataGroup_hi_lo_532};
  wire [7:0]    dataGroup_20_16 = dataGroup_lo_532[975:968];
  wire [1023:0] dataGroup_lo_533 = {dataGroup_lo_hi_533, dataGroup_lo_lo_533};
  wire [1023:0] dataGroup_hi_533 = {dataGroup_hi_hi_533, dataGroup_hi_lo_533};
  wire [7:0]    dataGroup_21_16 = dataGroup_lo_533[1023:1016];
  wire [1023:0] dataGroup_lo_534 = {dataGroup_lo_hi_534, dataGroup_lo_lo_534};
  wire [1023:0] dataGroup_hi_534 = {dataGroup_hi_hi_534, dataGroup_hi_lo_534};
  wire [7:0]    dataGroup_22_16 = dataGroup_hi_534[47:40];
  wire [1023:0] dataGroup_lo_535 = {dataGroup_lo_hi_535, dataGroup_lo_lo_535};
  wire [1023:0] dataGroup_hi_535 = {dataGroup_hi_hi_535, dataGroup_hi_lo_535};
  wire [7:0]    dataGroup_23_16 = dataGroup_hi_535[95:88];
  wire [1023:0] dataGroup_lo_536 = {dataGroup_lo_hi_536, dataGroup_lo_lo_536};
  wire [1023:0] dataGroup_hi_536 = {dataGroup_hi_hi_536, dataGroup_hi_lo_536};
  wire [7:0]    dataGroup_24_16 = dataGroup_hi_536[143:136];
  wire [1023:0] dataGroup_lo_537 = {dataGroup_lo_hi_537, dataGroup_lo_lo_537};
  wire [1023:0] dataGroup_hi_537 = {dataGroup_hi_hi_537, dataGroup_hi_lo_537};
  wire [7:0]    dataGroup_25_16 = dataGroup_hi_537[191:184];
  wire [1023:0] dataGroup_lo_538 = {dataGroup_lo_hi_538, dataGroup_lo_lo_538};
  wire [1023:0] dataGroup_hi_538 = {dataGroup_hi_hi_538, dataGroup_hi_lo_538};
  wire [7:0]    dataGroup_26_16 = dataGroup_hi_538[239:232];
  wire [1023:0] dataGroup_lo_539 = {dataGroup_lo_hi_539, dataGroup_lo_lo_539};
  wire [1023:0] dataGroup_hi_539 = {dataGroup_hi_hi_539, dataGroup_hi_lo_539};
  wire [7:0]    dataGroup_27_16 = dataGroup_hi_539[287:280];
  wire [1023:0] dataGroup_lo_540 = {dataGroup_lo_hi_540, dataGroup_lo_lo_540};
  wire [1023:0] dataGroup_hi_540 = {dataGroup_hi_hi_540, dataGroup_hi_lo_540};
  wire [7:0]    dataGroup_28_16 = dataGroup_hi_540[335:328];
  wire [1023:0] dataGroup_lo_541 = {dataGroup_lo_hi_541, dataGroup_lo_lo_541};
  wire [1023:0] dataGroup_hi_541 = {dataGroup_hi_hi_541, dataGroup_hi_lo_541};
  wire [7:0]    dataGroup_29_16 = dataGroup_hi_541[383:376];
  wire [1023:0] dataGroup_lo_542 = {dataGroup_lo_hi_542, dataGroup_lo_lo_542};
  wire [1023:0] dataGroup_hi_542 = {dataGroup_hi_hi_542, dataGroup_hi_lo_542};
  wire [7:0]    dataGroup_30_16 = dataGroup_hi_542[431:424];
  wire [1023:0] dataGroup_lo_543 = {dataGroup_lo_hi_543, dataGroup_lo_lo_543};
  wire [1023:0] dataGroup_hi_543 = {dataGroup_hi_hi_543, dataGroup_hi_lo_543};
  wire [7:0]    dataGroup_31_16 = dataGroup_hi_543[479:472];
  wire [15:0]   res_lo_lo_lo_lo_16 = {dataGroup_1_16, dataGroup_0_16};
  wire [15:0]   res_lo_lo_lo_hi_16 = {dataGroup_3_16, dataGroup_2_16};
  wire [31:0]   res_lo_lo_lo_16 = {res_lo_lo_lo_hi_16, res_lo_lo_lo_lo_16};
  wire [15:0]   res_lo_lo_hi_lo_16 = {dataGroup_5_16, dataGroup_4_16};
  wire [15:0]   res_lo_lo_hi_hi_16 = {dataGroup_7_16, dataGroup_6_16};
  wire [31:0]   res_lo_lo_hi_16 = {res_lo_lo_hi_hi_16, res_lo_lo_hi_lo_16};
  wire [63:0]   res_lo_lo_16 = {res_lo_lo_hi_16, res_lo_lo_lo_16};
  wire [15:0]   res_lo_hi_lo_lo_16 = {dataGroup_9_16, dataGroup_8_16};
  wire [15:0]   res_lo_hi_lo_hi_16 = {dataGroup_11_16, dataGroup_10_16};
  wire [31:0]   res_lo_hi_lo_16 = {res_lo_hi_lo_hi_16, res_lo_hi_lo_lo_16};
  wire [15:0]   res_lo_hi_hi_lo_16 = {dataGroup_13_16, dataGroup_12_16};
  wire [15:0]   res_lo_hi_hi_hi_16 = {dataGroup_15_16, dataGroup_14_16};
  wire [31:0]   res_lo_hi_hi_16 = {res_lo_hi_hi_hi_16, res_lo_hi_hi_lo_16};
  wire [63:0]   res_lo_hi_16 = {res_lo_hi_hi_16, res_lo_hi_lo_16};
  wire [127:0]  res_lo_16 = {res_lo_hi_16, res_lo_lo_16};
  wire [15:0]   res_hi_lo_lo_lo_16 = {dataGroup_17_16, dataGroup_16_16};
  wire [15:0]   res_hi_lo_lo_hi_16 = {dataGroup_19_16, dataGroup_18_16};
  wire [31:0]   res_hi_lo_lo_16 = {res_hi_lo_lo_hi_16, res_hi_lo_lo_lo_16};
  wire [15:0]   res_hi_lo_hi_lo_16 = {dataGroup_21_16, dataGroup_20_16};
  wire [15:0]   res_hi_lo_hi_hi_16 = {dataGroup_23_16, dataGroup_22_16};
  wire [31:0]   res_hi_lo_hi_16 = {res_hi_lo_hi_hi_16, res_hi_lo_hi_lo_16};
  wire [63:0]   res_hi_lo_16 = {res_hi_lo_hi_16, res_hi_lo_lo_16};
  wire [15:0]   res_hi_hi_lo_lo_16 = {dataGroup_25_16, dataGroup_24_16};
  wire [15:0]   res_hi_hi_lo_hi_16 = {dataGroup_27_16, dataGroup_26_16};
  wire [31:0]   res_hi_hi_lo_16 = {res_hi_hi_lo_hi_16, res_hi_hi_lo_lo_16};
  wire [15:0]   res_hi_hi_hi_lo_16 = {dataGroup_29_16, dataGroup_28_16};
  wire [15:0]   res_hi_hi_hi_hi_16 = {dataGroup_31_16, dataGroup_30_16};
  wire [31:0]   res_hi_hi_hi_16 = {res_hi_hi_hi_hi_16, res_hi_hi_hi_lo_16};
  wire [63:0]   res_hi_hi_16 = {res_hi_hi_hi_16, res_hi_hi_lo_16};
  wire [127:0]  res_hi_16 = {res_hi_hi_16, res_hi_lo_16};
  wire [255:0]  res_41 = {res_hi_16, res_lo_16};
  wire [1023:0] dataGroup_lo_544 = {dataGroup_lo_hi_544, dataGroup_lo_lo_544};
  wire [1023:0] dataGroup_hi_544 = {dataGroup_hi_hi_544, dataGroup_hi_lo_544};
  wire [7:0]    dataGroup_0_17 = dataGroup_lo_544[23:16];
  wire [1023:0] dataGroup_lo_545 = {dataGroup_lo_hi_545, dataGroup_lo_lo_545};
  wire [1023:0] dataGroup_hi_545 = {dataGroup_hi_hi_545, dataGroup_hi_lo_545};
  wire [7:0]    dataGroup_1_17 = dataGroup_lo_545[71:64];
  wire [1023:0] dataGroup_lo_546 = {dataGroup_lo_hi_546, dataGroup_lo_lo_546};
  wire [1023:0] dataGroup_hi_546 = {dataGroup_hi_hi_546, dataGroup_hi_lo_546};
  wire [7:0]    dataGroup_2_17 = dataGroup_lo_546[119:112];
  wire [1023:0] dataGroup_lo_547 = {dataGroup_lo_hi_547, dataGroup_lo_lo_547};
  wire [1023:0] dataGroup_hi_547 = {dataGroup_hi_hi_547, dataGroup_hi_lo_547};
  wire [7:0]    dataGroup_3_17 = dataGroup_lo_547[167:160];
  wire [1023:0] dataGroup_lo_548 = {dataGroup_lo_hi_548, dataGroup_lo_lo_548};
  wire [1023:0] dataGroup_hi_548 = {dataGroup_hi_hi_548, dataGroup_hi_lo_548};
  wire [7:0]    dataGroup_4_17 = dataGroup_lo_548[215:208];
  wire [1023:0] dataGroup_lo_549 = {dataGroup_lo_hi_549, dataGroup_lo_lo_549};
  wire [1023:0] dataGroup_hi_549 = {dataGroup_hi_hi_549, dataGroup_hi_lo_549};
  wire [7:0]    dataGroup_5_17 = dataGroup_lo_549[263:256];
  wire [1023:0] dataGroup_lo_550 = {dataGroup_lo_hi_550, dataGroup_lo_lo_550};
  wire [1023:0] dataGroup_hi_550 = {dataGroup_hi_hi_550, dataGroup_hi_lo_550};
  wire [7:0]    dataGroup_6_17 = dataGroup_lo_550[311:304];
  wire [1023:0] dataGroup_lo_551 = {dataGroup_lo_hi_551, dataGroup_lo_lo_551};
  wire [1023:0] dataGroup_hi_551 = {dataGroup_hi_hi_551, dataGroup_hi_lo_551};
  wire [7:0]    dataGroup_7_17 = dataGroup_lo_551[359:352];
  wire [1023:0] dataGroup_lo_552 = {dataGroup_lo_hi_552, dataGroup_lo_lo_552};
  wire [1023:0] dataGroup_hi_552 = {dataGroup_hi_hi_552, dataGroup_hi_lo_552};
  wire [7:0]    dataGroup_8_17 = dataGroup_lo_552[407:400];
  wire [1023:0] dataGroup_lo_553 = {dataGroup_lo_hi_553, dataGroup_lo_lo_553};
  wire [1023:0] dataGroup_hi_553 = {dataGroup_hi_hi_553, dataGroup_hi_lo_553};
  wire [7:0]    dataGroup_9_17 = dataGroup_lo_553[455:448];
  wire [1023:0] dataGroup_lo_554 = {dataGroup_lo_hi_554, dataGroup_lo_lo_554};
  wire [1023:0] dataGroup_hi_554 = {dataGroup_hi_hi_554, dataGroup_hi_lo_554};
  wire [7:0]    dataGroup_10_17 = dataGroup_lo_554[503:496];
  wire [1023:0] dataGroup_lo_555 = {dataGroup_lo_hi_555, dataGroup_lo_lo_555};
  wire [1023:0] dataGroup_hi_555 = {dataGroup_hi_hi_555, dataGroup_hi_lo_555};
  wire [7:0]    dataGroup_11_17 = dataGroup_lo_555[551:544];
  wire [1023:0] dataGroup_lo_556 = {dataGroup_lo_hi_556, dataGroup_lo_lo_556};
  wire [1023:0] dataGroup_hi_556 = {dataGroup_hi_hi_556, dataGroup_hi_lo_556};
  wire [7:0]    dataGroup_12_17 = dataGroup_lo_556[599:592];
  wire [1023:0] dataGroup_lo_557 = {dataGroup_lo_hi_557, dataGroup_lo_lo_557};
  wire [1023:0] dataGroup_hi_557 = {dataGroup_hi_hi_557, dataGroup_hi_lo_557};
  wire [7:0]    dataGroup_13_17 = dataGroup_lo_557[647:640];
  wire [1023:0] dataGroup_lo_558 = {dataGroup_lo_hi_558, dataGroup_lo_lo_558};
  wire [1023:0] dataGroup_hi_558 = {dataGroup_hi_hi_558, dataGroup_hi_lo_558};
  wire [7:0]    dataGroup_14_17 = dataGroup_lo_558[695:688];
  wire [1023:0] dataGroup_lo_559 = {dataGroup_lo_hi_559, dataGroup_lo_lo_559};
  wire [1023:0] dataGroup_hi_559 = {dataGroup_hi_hi_559, dataGroup_hi_lo_559};
  wire [7:0]    dataGroup_15_17 = dataGroup_lo_559[743:736];
  wire [1023:0] dataGroup_lo_560 = {dataGroup_lo_hi_560, dataGroup_lo_lo_560};
  wire [1023:0] dataGroup_hi_560 = {dataGroup_hi_hi_560, dataGroup_hi_lo_560};
  wire [7:0]    dataGroup_16_17 = dataGroup_lo_560[791:784];
  wire [1023:0] dataGroup_lo_561 = {dataGroup_lo_hi_561, dataGroup_lo_lo_561};
  wire [1023:0] dataGroup_hi_561 = {dataGroup_hi_hi_561, dataGroup_hi_lo_561};
  wire [7:0]    dataGroup_17_17 = dataGroup_lo_561[839:832];
  wire [1023:0] dataGroup_lo_562 = {dataGroup_lo_hi_562, dataGroup_lo_lo_562};
  wire [1023:0] dataGroup_hi_562 = {dataGroup_hi_hi_562, dataGroup_hi_lo_562};
  wire [7:0]    dataGroup_18_17 = dataGroup_lo_562[887:880];
  wire [1023:0] dataGroup_lo_563 = {dataGroup_lo_hi_563, dataGroup_lo_lo_563};
  wire [1023:0] dataGroup_hi_563 = {dataGroup_hi_hi_563, dataGroup_hi_lo_563};
  wire [7:0]    dataGroup_19_17 = dataGroup_lo_563[935:928];
  wire [1023:0] dataGroup_lo_564 = {dataGroup_lo_hi_564, dataGroup_lo_lo_564};
  wire [1023:0] dataGroup_hi_564 = {dataGroup_hi_hi_564, dataGroup_hi_lo_564};
  wire [7:0]    dataGroup_20_17 = dataGroup_lo_564[983:976];
  wire [1023:0] dataGroup_lo_565 = {dataGroup_lo_hi_565, dataGroup_lo_lo_565};
  wire [1023:0] dataGroup_hi_565 = {dataGroup_hi_hi_565, dataGroup_hi_lo_565};
  wire [7:0]    dataGroup_21_17 = dataGroup_hi_565[7:0];
  wire [1023:0] dataGroup_lo_566 = {dataGroup_lo_hi_566, dataGroup_lo_lo_566};
  wire [1023:0] dataGroup_hi_566 = {dataGroup_hi_hi_566, dataGroup_hi_lo_566};
  wire [7:0]    dataGroup_22_17 = dataGroup_hi_566[55:48];
  wire [1023:0] dataGroup_lo_567 = {dataGroup_lo_hi_567, dataGroup_lo_lo_567};
  wire [1023:0] dataGroup_hi_567 = {dataGroup_hi_hi_567, dataGroup_hi_lo_567};
  wire [7:0]    dataGroup_23_17 = dataGroup_hi_567[103:96];
  wire [1023:0] dataGroup_lo_568 = {dataGroup_lo_hi_568, dataGroup_lo_lo_568};
  wire [1023:0] dataGroup_hi_568 = {dataGroup_hi_hi_568, dataGroup_hi_lo_568};
  wire [7:0]    dataGroup_24_17 = dataGroup_hi_568[151:144];
  wire [1023:0] dataGroup_lo_569 = {dataGroup_lo_hi_569, dataGroup_lo_lo_569};
  wire [1023:0] dataGroup_hi_569 = {dataGroup_hi_hi_569, dataGroup_hi_lo_569};
  wire [7:0]    dataGroup_25_17 = dataGroup_hi_569[199:192];
  wire [1023:0] dataGroup_lo_570 = {dataGroup_lo_hi_570, dataGroup_lo_lo_570};
  wire [1023:0] dataGroup_hi_570 = {dataGroup_hi_hi_570, dataGroup_hi_lo_570};
  wire [7:0]    dataGroup_26_17 = dataGroup_hi_570[247:240];
  wire [1023:0] dataGroup_lo_571 = {dataGroup_lo_hi_571, dataGroup_lo_lo_571};
  wire [1023:0] dataGroup_hi_571 = {dataGroup_hi_hi_571, dataGroup_hi_lo_571};
  wire [7:0]    dataGroup_27_17 = dataGroup_hi_571[295:288];
  wire [1023:0] dataGroup_lo_572 = {dataGroup_lo_hi_572, dataGroup_lo_lo_572};
  wire [1023:0] dataGroup_hi_572 = {dataGroup_hi_hi_572, dataGroup_hi_lo_572};
  wire [7:0]    dataGroup_28_17 = dataGroup_hi_572[343:336];
  wire [1023:0] dataGroup_lo_573 = {dataGroup_lo_hi_573, dataGroup_lo_lo_573};
  wire [1023:0] dataGroup_hi_573 = {dataGroup_hi_hi_573, dataGroup_hi_lo_573};
  wire [7:0]    dataGroup_29_17 = dataGroup_hi_573[391:384];
  wire [1023:0] dataGroup_lo_574 = {dataGroup_lo_hi_574, dataGroup_lo_lo_574};
  wire [1023:0] dataGroup_hi_574 = {dataGroup_hi_hi_574, dataGroup_hi_lo_574};
  wire [7:0]    dataGroup_30_17 = dataGroup_hi_574[439:432];
  wire [1023:0] dataGroup_lo_575 = {dataGroup_lo_hi_575, dataGroup_lo_lo_575};
  wire [1023:0] dataGroup_hi_575 = {dataGroup_hi_hi_575, dataGroup_hi_lo_575};
  wire [7:0]    dataGroup_31_17 = dataGroup_hi_575[487:480];
  wire [15:0]   res_lo_lo_lo_lo_17 = {dataGroup_1_17, dataGroup_0_17};
  wire [15:0]   res_lo_lo_lo_hi_17 = {dataGroup_3_17, dataGroup_2_17};
  wire [31:0]   res_lo_lo_lo_17 = {res_lo_lo_lo_hi_17, res_lo_lo_lo_lo_17};
  wire [15:0]   res_lo_lo_hi_lo_17 = {dataGroup_5_17, dataGroup_4_17};
  wire [15:0]   res_lo_lo_hi_hi_17 = {dataGroup_7_17, dataGroup_6_17};
  wire [31:0]   res_lo_lo_hi_17 = {res_lo_lo_hi_hi_17, res_lo_lo_hi_lo_17};
  wire [63:0]   res_lo_lo_17 = {res_lo_lo_hi_17, res_lo_lo_lo_17};
  wire [15:0]   res_lo_hi_lo_lo_17 = {dataGroup_9_17, dataGroup_8_17};
  wire [15:0]   res_lo_hi_lo_hi_17 = {dataGroup_11_17, dataGroup_10_17};
  wire [31:0]   res_lo_hi_lo_17 = {res_lo_hi_lo_hi_17, res_lo_hi_lo_lo_17};
  wire [15:0]   res_lo_hi_hi_lo_17 = {dataGroup_13_17, dataGroup_12_17};
  wire [15:0]   res_lo_hi_hi_hi_17 = {dataGroup_15_17, dataGroup_14_17};
  wire [31:0]   res_lo_hi_hi_17 = {res_lo_hi_hi_hi_17, res_lo_hi_hi_lo_17};
  wire [63:0]   res_lo_hi_17 = {res_lo_hi_hi_17, res_lo_hi_lo_17};
  wire [127:0]  res_lo_17 = {res_lo_hi_17, res_lo_lo_17};
  wire [15:0]   res_hi_lo_lo_lo_17 = {dataGroup_17_17, dataGroup_16_17};
  wire [15:0]   res_hi_lo_lo_hi_17 = {dataGroup_19_17, dataGroup_18_17};
  wire [31:0]   res_hi_lo_lo_17 = {res_hi_lo_lo_hi_17, res_hi_lo_lo_lo_17};
  wire [15:0]   res_hi_lo_hi_lo_17 = {dataGroup_21_17, dataGroup_20_17};
  wire [15:0]   res_hi_lo_hi_hi_17 = {dataGroup_23_17, dataGroup_22_17};
  wire [31:0]   res_hi_lo_hi_17 = {res_hi_lo_hi_hi_17, res_hi_lo_hi_lo_17};
  wire [63:0]   res_hi_lo_17 = {res_hi_lo_hi_17, res_hi_lo_lo_17};
  wire [15:0]   res_hi_hi_lo_lo_17 = {dataGroup_25_17, dataGroup_24_17};
  wire [15:0]   res_hi_hi_lo_hi_17 = {dataGroup_27_17, dataGroup_26_17};
  wire [31:0]   res_hi_hi_lo_17 = {res_hi_hi_lo_hi_17, res_hi_hi_lo_lo_17};
  wire [15:0]   res_hi_hi_hi_lo_17 = {dataGroup_29_17, dataGroup_28_17};
  wire [15:0]   res_hi_hi_hi_hi_17 = {dataGroup_31_17, dataGroup_30_17};
  wire [31:0]   res_hi_hi_hi_17 = {res_hi_hi_hi_hi_17, res_hi_hi_hi_lo_17};
  wire [63:0]   res_hi_hi_17 = {res_hi_hi_hi_17, res_hi_hi_lo_17};
  wire [127:0]  res_hi_17 = {res_hi_hi_17, res_hi_lo_17};
  wire [255:0]  res_42 = {res_hi_17, res_lo_17};
  wire [1023:0] dataGroup_lo_576 = {dataGroup_lo_hi_576, dataGroup_lo_lo_576};
  wire [1023:0] dataGroup_hi_576 = {dataGroup_hi_hi_576, dataGroup_hi_lo_576};
  wire [7:0]    dataGroup_0_18 = dataGroup_lo_576[31:24];
  wire [1023:0] dataGroup_lo_577 = {dataGroup_lo_hi_577, dataGroup_lo_lo_577};
  wire [1023:0] dataGroup_hi_577 = {dataGroup_hi_hi_577, dataGroup_hi_lo_577};
  wire [7:0]    dataGroup_1_18 = dataGroup_lo_577[79:72];
  wire [1023:0] dataGroup_lo_578 = {dataGroup_lo_hi_578, dataGroup_lo_lo_578};
  wire [1023:0] dataGroup_hi_578 = {dataGroup_hi_hi_578, dataGroup_hi_lo_578};
  wire [7:0]    dataGroup_2_18 = dataGroup_lo_578[127:120];
  wire [1023:0] dataGroup_lo_579 = {dataGroup_lo_hi_579, dataGroup_lo_lo_579};
  wire [1023:0] dataGroup_hi_579 = {dataGroup_hi_hi_579, dataGroup_hi_lo_579};
  wire [7:0]    dataGroup_3_18 = dataGroup_lo_579[175:168];
  wire [1023:0] dataGroup_lo_580 = {dataGroup_lo_hi_580, dataGroup_lo_lo_580};
  wire [1023:0] dataGroup_hi_580 = {dataGroup_hi_hi_580, dataGroup_hi_lo_580};
  wire [7:0]    dataGroup_4_18 = dataGroup_lo_580[223:216];
  wire [1023:0] dataGroup_lo_581 = {dataGroup_lo_hi_581, dataGroup_lo_lo_581};
  wire [1023:0] dataGroup_hi_581 = {dataGroup_hi_hi_581, dataGroup_hi_lo_581};
  wire [7:0]    dataGroup_5_18 = dataGroup_lo_581[271:264];
  wire [1023:0] dataGroup_lo_582 = {dataGroup_lo_hi_582, dataGroup_lo_lo_582};
  wire [1023:0] dataGroup_hi_582 = {dataGroup_hi_hi_582, dataGroup_hi_lo_582};
  wire [7:0]    dataGroup_6_18 = dataGroup_lo_582[319:312];
  wire [1023:0] dataGroup_lo_583 = {dataGroup_lo_hi_583, dataGroup_lo_lo_583};
  wire [1023:0] dataGroup_hi_583 = {dataGroup_hi_hi_583, dataGroup_hi_lo_583};
  wire [7:0]    dataGroup_7_18 = dataGroup_lo_583[367:360];
  wire [1023:0] dataGroup_lo_584 = {dataGroup_lo_hi_584, dataGroup_lo_lo_584};
  wire [1023:0] dataGroup_hi_584 = {dataGroup_hi_hi_584, dataGroup_hi_lo_584};
  wire [7:0]    dataGroup_8_18 = dataGroup_lo_584[415:408];
  wire [1023:0] dataGroup_lo_585 = {dataGroup_lo_hi_585, dataGroup_lo_lo_585};
  wire [1023:0] dataGroup_hi_585 = {dataGroup_hi_hi_585, dataGroup_hi_lo_585};
  wire [7:0]    dataGroup_9_18 = dataGroup_lo_585[463:456];
  wire [1023:0] dataGroup_lo_586 = {dataGroup_lo_hi_586, dataGroup_lo_lo_586};
  wire [1023:0] dataGroup_hi_586 = {dataGroup_hi_hi_586, dataGroup_hi_lo_586};
  wire [7:0]    dataGroup_10_18 = dataGroup_lo_586[511:504];
  wire [1023:0] dataGroup_lo_587 = {dataGroup_lo_hi_587, dataGroup_lo_lo_587};
  wire [1023:0] dataGroup_hi_587 = {dataGroup_hi_hi_587, dataGroup_hi_lo_587};
  wire [7:0]    dataGroup_11_18 = dataGroup_lo_587[559:552];
  wire [1023:0] dataGroup_lo_588 = {dataGroup_lo_hi_588, dataGroup_lo_lo_588};
  wire [1023:0] dataGroup_hi_588 = {dataGroup_hi_hi_588, dataGroup_hi_lo_588};
  wire [7:0]    dataGroup_12_18 = dataGroup_lo_588[607:600];
  wire [1023:0] dataGroup_lo_589 = {dataGroup_lo_hi_589, dataGroup_lo_lo_589};
  wire [1023:0] dataGroup_hi_589 = {dataGroup_hi_hi_589, dataGroup_hi_lo_589};
  wire [7:0]    dataGroup_13_18 = dataGroup_lo_589[655:648];
  wire [1023:0] dataGroup_lo_590 = {dataGroup_lo_hi_590, dataGroup_lo_lo_590};
  wire [1023:0] dataGroup_hi_590 = {dataGroup_hi_hi_590, dataGroup_hi_lo_590};
  wire [7:0]    dataGroup_14_18 = dataGroup_lo_590[703:696];
  wire [1023:0] dataGroup_lo_591 = {dataGroup_lo_hi_591, dataGroup_lo_lo_591};
  wire [1023:0] dataGroup_hi_591 = {dataGroup_hi_hi_591, dataGroup_hi_lo_591};
  wire [7:0]    dataGroup_15_18 = dataGroup_lo_591[751:744];
  wire [1023:0] dataGroup_lo_592 = {dataGroup_lo_hi_592, dataGroup_lo_lo_592};
  wire [1023:0] dataGroup_hi_592 = {dataGroup_hi_hi_592, dataGroup_hi_lo_592};
  wire [7:0]    dataGroup_16_18 = dataGroup_lo_592[799:792];
  wire [1023:0] dataGroup_lo_593 = {dataGroup_lo_hi_593, dataGroup_lo_lo_593};
  wire [1023:0] dataGroup_hi_593 = {dataGroup_hi_hi_593, dataGroup_hi_lo_593};
  wire [7:0]    dataGroup_17_18 = dataGroup_lo_593[847:840];
  wire [1023:0] dataGroup_lo_594 = {dataGroup_lo_hi_594, dataGroup_lo_lo_594};
  wire [1023:0] dataGroup_hi_594 = {dataGroup_hi_hi_594, dataGroup_hi_lo_594};
  wire [7:0]    dataGroup_18_18 = dataGroup_lo_594[895:888];
  wire [1023:0] dataGroup_lo_595 = {dataGroup_lo_hi_595, dataGroup_lo_lo_595};
  wire [1023:0] dataGroup_hi_595 = {dataGroup_hi_hi_595, dataGroup_hi_lo_595};
  wire [7:0]    dataGroup_19_18 = dataGroup_lo_595[943:936];
  wire [1023:0] dataGroup_lo_596 = {dataGroup_lo_hi_596, dataGroup_lo_lo_596};
  wire [1023:0] dataGroup_hi_596 = {dataGroup_hi_hi_596, dataGroup_hi_lo_596};
  wire [7:0]    dataGroup_20_18 = dataGroup_lo_596[991:984];
  wire [1023:0] dataGroup_lo_597 = {dataGroup_lo_hi_597, dataGroup_lo_lo_597};
  wire [1023:0] dataGroup_hi_597 = {dataGroup_hi_hi_597, dataGroup_hi_lo_597};
  wire [7:0]    dataGroup_21_18 = dataGroup_hi_597[15:8];
  wire [1023:0] dataGroup_lo_598 = {dataGroup_lo_hi_598, dataGroup_lo_lo_598};
  wire [1023:0] dataGroup_hi_598 = {dataGroup_hi_hi_598, dataGroup_hi_lo_598};
  wire [7:0]    dataGroup_22_18 = dataGroup_hi_598[63:56];
  wire [1023:0] dataGroup_lo_599 = {dataGroup_lo_hi_599, dataGroup_lo_lo_599};
  wire [1023:0] dataGroup_hi_599 = {dataGroup_hi_hi_599, dataGroup_hi_lo_599};
  wire [7:0]    dataGroup_23_18 = dataGroup_hi_599[111:104];
  wire [1023:0] dataGroup_lo_600 = {dataGroup_lo_hi_600, dataGroup_lo_lo_600};
  wire [1023:0] dataGroup_hi_600 = {dataGroup_hi_hi_600, dataGroup_hi_lo_600};
  wire [7:0]    dataGroup_24_18 = dataGroup_hi_600[159:152];
  wire [1023:0] dataGroup_lo_601 = {dataGroup_lo_hi_601, dataGroup_lo_lo_601};
  wire [1023:0] dataGroup_hi_601 = {dataGroup_hi_hi_601, dataGroup_hi_lo_601};
  wire [7:0]    dataGroup_25_18 = dataGroup_hi_601[207:200];
  wire [1023:0] dataGroup_lo_602 = {dataGroup_lo_hi_602, dataGroup_lo_lo_602};
  wire [1023:0] dataGroup_hi_602 = {dataGroup_hi_hi_602, dataGroup_hi_lo_602};
  wire [7:0]    dataGroup_26_18 = dataGroup_hi_602[255:248];
  wire [1023:0] dataGroup_lo_603 = {dataGroup_lo_hi_603, dataGroup_lo_lo_603};
  wire [1023:0] dataGroup_hi_603 = {dataGroup_hi_hi_603, dataGroup_hi_lo_603};
  wire [7:0]    dataGroup_27_18 = dataGroup_hi_603[303:296];
  wire [1023:0] dataGroup_lo_604 = {dataGroup_lo_hi_604, dataGroup_lo_lo_604};
  wire [1023:0] dataGroup_hi_604 = {dataGroup_hi_hi_604, dataGroup_hi_lo_604};
  wire [7:0]    dataGroup_28_18 = dataGroup_hi_604[351:344];
  wire [1023:0] dataGroup_lo_605 = {dataGroup_lo_hi_605, dataGroup_lo_lo_605};
  wire [1023:0] dataGroup_hi_605 = {dataGroup_hi_hi_605, dataGroup_hi_lo_605};
  wire [7:0]    dataGroup_29_18 = dataGroup_hi_605[399:392];
  wire [1023:0] dataGroup_lo_606 = {dataGroup_lo_hi_606, dataGroup_lo_lo_606};
  wire [1023:0] dataGroup_hi_606 = {dataGroup_hi_hi_606, dataGroup_hi_lo_606};
  wire [7:0]    dataGroup_30_18 = dataGroup_hi_606[447:440];
  wire [1023:0] dataGroup_lo_607 = {dataGroup_lo_hi_607, dataGroup_lo_lo_607};
  wire [1023:0] dataGroup_hi_607 = {dataGroup_hi_hi_607, dataGroup_hi_lo_607};
  wire [7:0]    dataGroup_31_18 = dataGroup_hi_607[495:488];
  wire [15:0]   res_lo_lo_lo_lo_18 = {dataGroup_1_18, dataGroup_0_18};
  wire [15:0]   res_lo_lo_lo_hi_18 = {dataGroup_3_18, dataGroup_2_18};
  wire [31:0]   res_lo_lo_lo_18 = {res_lo_lo_lo_hi_18, res_lo_lo_lo_lo_18};
  wire [15:0]   res_lo_lo_hi_lo_18 = {dataGroup_5_18, dataGroup_4_18};
  wire [15:0]   res_lo_lo_hi_hi_18 = {dataGroup_7_18, dataGroup_6_18};
  wire [31:0]   res_lo_lo_hi_18 = {res_lo_lo_hi_hi_18, res_lo_lo_hi_lo_18};
  wire [63:0]   res_lo_lo_18 = {res_lo_lo_hi_18, res_lo_lo_lo_18};
  wire [15:0]   res_lo_hi_lo_lo_18 = {dataGroup_9_18, dataGroup_8_18};
  wire [15:0]   res_lo_hi_lo_hi_18 = {dataGroup_11_18, dataGroup_10_18};
  wire [31:0]   res_lo_hi_lo_18 = {res_lo_hi_lo_hi_18, res_lo_hi_lo_lo_18};
  wire [15:0]   res_lo_hi_hi_lo_18 = {dataGroup_13_18, dataGroup_12_18};
  wire [15:0]   res_lo_hi_hi_hi_18 = {dataGroup_15_18, dataGroup_14_18};
  wire [31:0]   res_lo_hi_hi_18 = {res_lo_hi_hi_hi_18, res_lo_hi_hi_lo_18};
  wire [63:0]   res_lo_hi_18 = {res_lo_hi_hi_18, res_lo_hi_lo_18};
  wire [127:0]  res_lo_18 = {res_lo_hi_18, res_lo_lo_18};
  wire [15:0]   res_hi_lo_lo_lo_18 = {dataGroup_17_18, dataGroup_16_18};
  wire [15:0]   res_hi_lo_lo_hi_18 = {dataGroup_19_18, dataGroup_18_18};
  wire [31:0]   res_hi_lo_lo_18 = {res_hi_lo_lo_hi_18, res_hi_lo_lo_lo_18};
  wire [15:0]   res_hi_lo_hi_lo_18 = {dataGroup_21_18, dataGroup_20_18};
  wire [15:0]   res_hi_lo_hi_hi_18 = {dataGroup_23_18, dataGroup_22_18};
  wire [31:0]   res_hi_lo_hi_18 = {res_hi_lo_hi_hi_18, res_hi_lo_hi_lo_18};
  wire [63:0]   res_hi_lo_18 = {res_hi_lo_hi_18, res_hi_lo_lo_18};
  wire [15:0]   res_hi_hi_lo_lo_18 = {dataGroup_25_18, dataGroup_24_18};
  wire [15:0]   res_hi_hi_lo_hi_18 = {dataGroup_27_18, dataGroup_26_18};
  wire [31:0]   res_hi_hi_lo_18 = {res_hi_hi_lo_hi_18, res_hi_hi_lo_lo_18};
  wire [15:0]   res_hi_hi_hi_lo_18 = {dataGroup_29_18, dataGroup_28_18};
  wire [15:0]   res_hi_hi_hi_hi_18 = {dataGroup_31_18, dataGroup_30_18};
  wire [31:0]   res_hi_hi_hi_18 = {res_hi_hi_hi_hi_18, res_hi_hi_hi_lo_18};
  wire [63:0]   res_hi_hi_18 = {res_hi_hi_hi_18, res_hi_hi_lo_18};
  wire [127:0]  res_hi_18 = {res_hi_hi_18, res_hi_lo_18};
  wire [255:0]  res_43 = {res_hi_18, res_lo_18};
  wire [1023:0] dataGroup_lo_608 = {dataGroup_lo_hi_608, dataGroup_lo_lo_608};
  wire [1023:0] dataGroup_hi_608 = {dataGroup_hi_hi_608, dataGroup_hi_lo_608};
  wire [7:0]    dataGroup_0_19 = dataGroup_lo_608[39:32];
  wire [1023:0] dataGroup_lo_609 = {dataGroup_lo_hi_609, dataGroup_lo_lo_609};
  wire [1023:0] dataGroup_hi_609 = {dataGroup_hi_hi_609, dataGroup_hi_lo_609};
  wire [7:0]    dataGroup_1_19 = dataGroup_lo_609[87:80];
  wire [1023:0] dataGroup_lo_610 = {dataGroup_lo_hi_610, dataGroup_lo_lo_610};
  wire [1023:0] dataGroup_hi_610 = {dataGroup_hi_hi_610, dataGroup_hi_lo_610};
  wire [7:0]    dataGroup_2_19 = dataGroup_lo_610[135:128];
  wire [1023:0] dataGroup_lo_611 = {dataGroup_lo_hi_611, dataGroup_lo_lo_611};
  wire [1023:0] dataGroup_hi_611 = {dataGroup_hi_hi_611, dataGroup_hi_lo_611};
  wire [7:0]    dataGroup_3_19 = dataGroup_lo_611[183:176];
  wire [1023:0] dataGroup_lo_612 = {dataGroup_lo_hi_612, dataGroup_lo_lo_612};
  wire [1023:0] dataGroup_hi_612 = {dataGroup_hi_hi_612, dataGroup_hi_lo_612};
  wire [7:0]    dataGroup_4_19 = dataGroup_lo_612[231:224];
  wire [1023:0] dataGroup_lo_613 = {dataGroup_lo_hi_613, dataGroup_lo_lo_613};
  wire [1023:0] dataGroup_hi_613 = {dataGroup_hi_hi_613, dataGroup_hi_lo_613};
  wire [7:0]    dataGroup_5_19 = dataGroup_lo_613[279:272];
  wire [1023:0] dataGroup_lo_614 = {dataGroup_lo_hi_614, dataGroup_lo_lo_614};
  wire [1023:0] dataGroup_hi_614 = {dataGroup_hi_hi_614, dataGroup_hi_lo_614};
  wire [7:0]    dataGroup_6_19 = dataGroup_lo_614[327:320];
  wire [1023:0] dataGroup_lo_615 = {dataGroup_lo_hi_615, dataGroup_lo_lo_615};
  wire [1023:0] dataGroup_hi_615 = {dataGroup_hi_hi_615, dataGroup_hi_lo_615};
  wire [7:0]    dataGroup_7_19 = dataGroup_lo_615[375:368];
  wire [1023:0] dataGroup_lo_616 = {dataGroup_lo_hi_616, dataGroup_lo_lo_616};
  wire [1023:0] dataGroup_hi_616 = {dataGroup_hi_hi_616, dataGroup_hi_lo_616};
  wire [7:0]    dataGroup_8_19 = dataGroup_lo_616[423:416];
  wire [1023:0] dataGroup_lo_617 = {dataGroup_lo_hi_617, dataGroup_lo_lo_617};
  wire [1023:0] dataGroup_hi_617 = {dataGroup_hi_hi_617, dataGroup_hi_lo_617};
  wire [7:0]    dataGroup_9_19 = dataGroup_lo_617[471:464];
  wire [1023:0] dataGroup_lo_618 = {dataGroup_lo_hi_618, dataGroup_lo_lo_618};
  wire [1023:0] dataGroup_hi_618 = {dataGroup_hi_hi_618, dataGroup_hi_lo_618};
  wire [7:0]    dataGroup_10_19 = dataGroup_lo_618[519:512];
  wire [1023:0] dataGroup_lo_619 = {dataGroup_lo_hi_619, dataGroup_lo_lo_619};
  wire [1023:0] dataGroup_hi_619 = {dataGroup_hi_hi_619, dataGroup_hi_lo_619};
  wire [7:0]    dataGroup_11_19 = dataGroup_lo_619[567:560];
  wire [1023:0] dataGroup_lo_620 = {dataGroup_lo_hi_620, dataGroup_lo_lo_620};
  wire [1023:0] dataGroup_hi_620 = {dataGroup_hi_hi_620, dataGroup_hi_lo_620};
  wire [7:0]    dataGroup_12_19 = dataGroup_lo_620[615:608];
  wire [1023:0] dataGroup_lo_621 = {dataGroup_lo_hi_621, dataGroup_lo_lo_621};
  wire [1023:0] dataGroup_hi_621 = {dataGroup_hi_hi_621, dataGroup_hi_lo_621};
  wire [7:0]    dataGroup_13_19 = dataGroup_lo_621[663:656];
  wire [1023:0] dataGroup_lo_622 = {dataGroup_lo_hi_622, dataGroup_lo_lo_622};
  wire [1023:0] dataGroup_hi_622 = {dataGroup_hi_hi_622, dataGroup_hi_lo_622};
  wire [7:0]    dataGroup_14_19 = dataGroup_lo_622[711:704];
  wire [1023:0] dataGroup_lo_623 = {dataGroup_lo_hi_623, dataGroup_lo_lo_623};
  wire [1023:0] dataGroup_hi_623 = {dataGroup_hi_hi_623, dataGroup_hi_lo_623};
  wire [7:0]    dataGroup_15_19 = dataGroup_lo_623[759:752];
  wire [1023:0] dataGroup_lo_624 = {dataGroup_lo_hi_624, dataGroup_lo_lo_624};
  wire [1023:0] dataGroup_hi_624 = {dataGroup_hi_hi_624, dataGroup_hi_lo_624};
  wire [7:0]    dataGroup_16_19 = dataGroup_lo_624[807:800];
  wire [1023:0] dataGroup_lo_625 = {dataGroup_lo_hi_625, dataGroup_lo_lo_625};
  wire [1023:0] dataGroup_hi_625 = {dataGroup_hi_hi_625, dataGroup_hi_lo_625};
  wire [7:0]    dataGroup_17_19 = dataGroup_lo_625[855:848];
  wire [1023:0] dataGroup_lo_626 = {dataGroup_lo_hi_626, dataGroup_lo_lo_626};
  wire [1023:0] dataGroup_hi_626 = {dataGroup_hi_hi_626, dataGroup_hi_lo_626};
  wire [7:0]    dataGroup_18_19 = dataGroup_lo_626[903:896];
  wire [1023:0] dataGroup_lo_627 = {dataGroup_lo_hi_627, dataGroup_lo_lo_627};
  wire [1023:0] dataGroup_hi_627 = {dataGroup_hi_hi_627, dataGroup_hi_lo_627};
  wire [7:0]    dataGroup_19_19 = dataGroup_lo_627[951:944];
  wire [1023:0] dataGroup_lo_628 = {dataGroup_lo_hi_628, dataGroup_lo_lo_628};
  wire [1023:0] dataGroup_hi_628 = {dataGroup_hi_hi_628, dataGroup_hi_lo_628};
  wire [7:0]    dataGroup_20_19 = dataGroup_lo_628[999:992];
  wire [1023:0] dataGroup_lo_629 = {dataGroup_lo_hi_629, dataGroup_lo_lo_629};
  wire [1023:0] dataGroup_hi_629 = {dataGroup_hi_hi_629, dataGroup_hi_lo_629};
  wire [7:0]    dataGroup_21_19 = dataGroup_hi_629[23:16];
  wire [1023:0] dataGroup_lo_630 = {dataGroup_lo_hi_630, dataGroup_lo_lo_630};
  wire [1023:0] dataGroup_hi_630 = {dataGroup_hi_hi_630, dataGroup_hi_lo_630};
  wire [7:0]    dataGroup_22_19 = dataGroup_hi_630[71:64];
  wire [1023:0] dataGroup_lo_631 = {dataGroup_lo_hi_631, dataGroup_lo_lo_631};
  wire [1023:0] dataGroup_hi_631 = {dataGroup_hi_hi_631, dataGroup_hi_lo_631};
  wire [7:0]    dataGroup_23_19 = dataGroup_hi_631[119:112];
  wire [1023:0] dataGroup_lo_632 = {dataGroup_lo_hi_632, dataGroup_lo_lo_632};
  wire [1023:0] dataGroup_hi_632 = {dataGroup_hi_hi_632, dataGroup_hi_lo_632};
  wire [7:0]    dataGroup_24_19 = dataGroup_hi_632[167:160];
  wire [1023:0] dataGroup_lo_633 = {dataGroup_lo_hi_633, dataGroup_lo_lo_633};
  wire [1023:0] dataGroup_hi_633 = {dataGroup_hi_hi_633, dataGroup_hi_lo_633};
  wire [7:0]    dataGroup_25_19 = dataGroup_hi_633[215:208];
  wire [1023:0] dataGroup_lo_634 = {dataGroup_lo_hi_634, dataGroup_lo_lo_634};
  wire [1023:0] dataGroup_hi_634 = {dataGroup_hi_hi_634, dataGroup_hi_lo_634};
  wire [7:0]    dataGroup_26_19 = dataGroup_hi_634[263:256];
  wire [1023:0] dataGroup_lo_635 = {dataGroup_lo_hi_635, dataGroup_lo_lo_635};
  wire [1023:0] dataGroup_hi_635 = {dataGroup_hi_hi_635, dataGroup_hi_lo_635};
  wire [7:0]    dataGroup_27_19 = dataGroup_hi_635[311:304];
  wire [1023:0] dataGroup_lo_636 = {dataGroup_lo_hi_636, dataGroup_lo_lo_636};
  wire [1023:0] dataGroup_hi_636 = {dataGroup_hi_hi_636, dataGroup_hi_lo_636};
  wire [7:0]    dataGroup_28_19 = dataGroup_hi_636[359:352];
  wire [1023:0] dataGroup_lo_637 = {dataGroup_lo_hi_637, dataGroup_lo_lo_637};
  wire [1023:0] dataGroup_hi_637 = {dataGroup_hi_hi_637, dataGroup_hi_lo_637};
  wire [7:0]    dataGroup_29_19 = dataGroup_hi_637[407:400];
  wire [1023:0] dataGroup_lo_638 = {dataGroup_lo_hi_638, dataGroup_lo_lo_638};
  wire [1023:0] dataGroup_hi_638 = {dataGroup_hi_hi_638, dataGroup_hi_lo_638};
  wire [7:0]    dataGroup_30_19 = dataGroup_hi_638[455:448];
  wire [1023:0] dataGroup_lo_639 = {dataGroup_lo_hi_639, dataGroup_lo_lo_639};
  wire [1023:0] dataGroup_hi_639 = {dataGroup_hi_hi_639, dataGroup_hi_lo_639};
  wire [7:0]    dataGroup_31_19 = dataGroup_hi_639[503:496];
  wire [15:0]   res_lo_lo_lo_lo_19 = {dataGroup_1_19, dataGroup_0_19};
  wire [15:0]   res_lo_lo_lo_hi_19 = {dataGroup_3_19, dataGroup_2_19};
  wire [31:0]   res_lo_lo_lo_19 = {res_lo_lo_lo_hi_19, res_lo_lo_lo_lo_19};
  wire [15:0]   res_lo_lo_hi_lo_19 = {dataGroup_5_19, dataGroup_4_19};
  wire [15:0]   res_lo_lo_hi_hi_19 = {dataGroup_7_19, dataGroup_6_19};
  wire [31:0]   res_lo_lo_hi_19 = {res_lo_lo_hi_hi_19, res_lo_lo_hi_lo_19};
  wire [63:0]   res_lo_lo_19 = {res_lo_lo_hi_19, res_lo_lo_lo_19};
  wire [15:0]   res_lo_hi_lo_lo_19 = {dataGroup_9_19, dataGroup_8_19};
  wire [15:0]   res_lo_hi_lo_hi_19 = {dataGroup_11_19, dataGroup_10_19};
  wire [31:0]   res_lo_hi_lo_19 = {res_lo_hi_lo_hi_19, res_lo_hi_lo_lo_19};
  wire [15:0]   res_lo_hi_hi_lo_19 = {dataGroup_13_19, dataGroup_12_19};
  wire [15:0]   res_lo_hi_hi_hi_19 = {dataGroup_15_19, dataGroup_14_19};
  wire [31:0]   res_lo_hi_hi_19 = {res_lo_hi_hi_hi_19, res_lo_hi_hi_lo_19};
  wire [63:0]   res_lo_hi_19 = {res_lo_hi_hi_19, res_lo_hi_lo_19};
  wire [127:0]  res_lo_19 = {res_lo_hi_19, res_lo_lo_19};
  wire [15:0]   res_hi_lo_lo_lo_19 = {dataGroup_17_19, dataGroup_16_19};
  wire [15:0]   res_hi_lo_lo_hi_19 = {dataGroup_19_19, dataGroup_18_19};
  wire [31:0]   res_hi_lo_lo_19 = {res_hi_lo_lo_hi_19, res_hi_lo_lo_lo_19};
  wire [15:0]   res_hi_lo_hi_lo_19 = {dataGroup_21_19, dataGroup_20_19};
  wire [15:0]   res_hi_lo_hi_hi_19 = {dataGroup_23_19, dataGroup_22_19};
  wire [31:0]   res_hi_lo_hi_19 = {res_hi_lo_hi_hi_19, res_hi_lo_hi_lo_19};
  wire [63:0]   res_hi_lo_19 = {res_hi_lo_hi_19, res_hi_lo_lo_19};
  wire [15:0]   res_hi_hi_lo_lo_19 = {dataGroup_25_19, dataGroup_24_19};
  wire [15:0]   res_hi_hi_lo_hi_19 = {dataGroup_27_19, dataGroup_26_19};
  wire [31:0]   res_hi_hi_lo_19 = {res_hi_hi_lo_hi_19, res_hi_hi_lo_lo_19};
  wire [15:0]   res_hi_hi_hi_lo_19 = {dataGroup_29_19, dataGroup_28_19};
  wire [15:0]   res_hi_hi_hi_hi_19 = {dataGroup_31_19, dataGroup_30_19};
  wire [31:0]   res_hi_hi_hi_19 = {res_hi_hi_hi_hi_19, res_hi_hi_hi_lo_19};
  wire [63:0]   res_hi_hi_19 = {res_hi_hi_hi_19, res_hi_hi_lo_19};
  wire [127:0]  res_hi_19 = {res_hi_hi_19, res_hi_lo_19};
  wire [255:0]  res_44 = {res_hi_19, res_lo_19};
  wire [1023:0] dataGroup_lo_640 = {dataGroup_lo_hi_640, dataGroup_lo_lo_640};
  wire [1023:0] dataGroup_hi_640 = {dataGroup_hi_hi_640, dataGroup_hi_lo_640};
  wire [7:0]    dataGroup_0_20 = dataGroup_lo_640[47:40];
  wire [1023:0] dataGroup_lo_641 = {dataGroup_lo_hi_641, dataGroup_lo_lo_641};
  wire [1023:0] dataGroup_hi_641 = {dataGroup_hi_hi_641, dataGroup_hi_lo_641};
  wire [7:0]    dataGroup_1_20 = dataGroup_lo_641[95:88];
  wire [1023:0] dataGroup_lo_642 = {dataGroup_lo_hi_642, dataGroup_lo_lo_642};
  wire [1023:0] dataGroup_hi_642 = {dataGroup_hi_hi_642, dataGroup_hi_lo_642};
  wire [7:0]    dataGroup_2_20 = dataGroup_lo_642[143:136];
  wire [1023:0] dataGroup_lo_643 = {dataGroup_lo_hi_643, dataGroup_lo_lo_643};
  wire [1023:0] dataGroup_hi_643 = {dataGroup_hi_hi_643, dataGroup_hi_lo_643};
  wire [7:0]    dataGroup_3_20 = dataGroup_lo_643[191:184];
  wire [1023:0] dataGroup_lo_644 = {dataGroup_lo_hi_644, dataGroup_lo_lo_644};
  wire [1023:0] dataGroup_hi_644 = {dataGroup_hi_hi_644, dataGroup_hi_lo_644};
  wire [7:0]    dataGroup_4_20 = dataGroup_lo_644[239:232];
  wire [1023:0] dataGroup_lo_645 = {dataGroup_lo_hi_645, dataGroup_lo_lo_645};
  wire [1023:0] dataGroup_hi_645 = {dataGroup_hi_hi_645, dataGroup_hi_lo_645};
  wire [7:0]    dataGroup_5_20 = dataGroup_lo_645[287:280];
  wire [1023:0] dataGroup_lo_646 = {dataGroup_lo_hi_646, dataGroup_lo_lo_646};
  wire [1023:0] dataGroup_hi_646 = {dataGroup_hi_hi_646, dataGroup_hi_lo_646};
  wire [7:0]    dataGroup_6_20 = dataGroup_lo_646[335:328];
  wire [1023:0] dataGroup_lo_647 = {dataGroup_lo_hi_647, dataGroup_lo_lo_647};
  wire [1023:0] dataGroup_hi_647 = {dataGroup_hi_hi_647, dataGroup_hi_lo_647};
  wire [7:0]    dataGroup_7_20 = dataGroup_lo_647[383:376];
  wire [1023:0] dataGroup_lo_648 = {dataGroup_lo_hi_648, dataGroup_lo_lo_648};
  wire [1023:0] dataGroup_hi_648 = {dataGroup_hi_hi_648, dataGroup_hi_lo_648};
  wire [7:0]    dataGroup_8_20 = dataGroup_lo_648[431:424];
  wire [1023:0] dataGroup_lo_649 = {dataGroup_lo_hi_649, dataGroup_lo_lo_649};
  wire [1023:0] dataGroup_hi_649 = {dataGroup_hi_hi_649, dataGroup_hi_lo_649};
  wire [7:0]    dataGroup_9_20 = dataGroup_lo_649[479:472];
  wire [1023:0] dataGroup_lo_650 = {dataGroup_lo_hi_650, dataGroup_lo_lo_650};
  wire [1023:0] dataGroup_hi_650 = {dataGroup_hi_hi_650, dataGroup_hi_lo_650};
  wire [7:0]    dataGroup_10_20 = dataGroup_lo_650[527:520];
  wire [1023:0] dataGroup_lo_651 = {dataGroup_lo_hi_651, dataGroup_lo_lo_651};
  wire [1023:0] dataGroup_hi_651 = {dataGroup_hi_hi_651, dataGroup_hi_lo_651};
  wire [7:0]    dataGroup_11_20 = dataGroup_lo_651[575:568];
  wire [1023:0] dataGroup_lo_652 = {dataGroup_lo_hi_652, dataGroup_lo_lo_652};
  wire [1023:0] dataGroup_hi_652 = {dataGroup_hi_hi_652, dataGroup_hi_lo_652};
  wire [7:0]    dataGroup_12_20 = dataGroup_lo_652[623:616];
  wire [1023:0] dataGroup_lo_653 = {dataGroup_lo_hi_653, dataGroup_lo_lo_653};
  wire [1023:0] dataGroup_hi_653 = {dataGroup_hi_hi_653, dataGroup_hi_lo_653};
  wire [7:0]    dataGroup_13_20 = dataGroup_lo_653[671:664];
  wire [1023:0] dataGroup_lo_654 = {dataGroup_lo_hi_654, dataGroup_lo_lo_654};
  wire [1023:0] dataGroup_hi_654 = {dataGroup_hi_hi_654, dataGroup_hi_lo_654};
  wire [7:0]    dataGroup_14_20 = dataGroup_lo_654[719:712];
  wire [1023:0] dataGroup_lo_655 = {dataGroup_lo_hi_655, dataGroup_lo_lo_655};
  wire [1023:0] dataGroup_hi_655 = {dataGroup_hi_hi_655, dataGroup_hi_lo_655};
  wire [7:0]    dataGroup_15_20 = dataGroup_lo_655[767:760];
  wire [1023:0] dataGroup_lo_656 = {dataGroup_lo_hi_656, dataGroup_lo_lo_656};
  wire [1023:0] dataGroup_hi_656 = {dataGroup_hi_hi_656, dataGroup_hi_lo_656};
  wire [7:0]    dataGroup_16_20 = dataGroup_lo_656[815:808];
  wire [1023:0] dataGroup_lo_657 = {dataGroup_lo_hi_657, dataGroup_lo_lo_657};
  wire [1023:0] dataGroup_hi_657 = {dataGroup_hi_hi_657, dataGroup_hi_lo_657};
  wire [7:0]    dataGroup_17_20 = dataGroup_lo_657[863:856];
  wire [1023:0] dataGroup_lo_658 = {dataGroup_lo_hi_658, dataGroup_lo_lo_658};
  wire [1023:0] dataGroup_hi_658 = {dataGroup_hi_hi_658, dataGroup_hi_lo_658};
  wire [7:0]    dataGroup_18_20 = dataGroup_lo_658[911:904];
  wire [1023:0] dataGroup_lo_659 = {dataGroup_lo_hi_659, dataGroup_lo_lo_659};
  wire [1023:0] dataGroup_hi_659 = {dataGroup_hi_hi_659, dataGroup_hi_lo_659};
  wire [7:0]    dataGroup_19_20 = dataGroup_lo_659[959:952];
  wire [1023:0] dataGroup_lo_660 = {dataGroup_lo_hi_660, dataGroup_lo_lo_660};
  wire [1023:0] dataGroup_hi_660 = {dataGroup_hi_hi_660, dataGroup_hi_lo_660};
  wire [7:0]    dataGroup_20_20 = dataGroup_lo_660[1007:1000];
  wire [1023:0] dataGroup_lo_661 = {dataGroup_lo_hi_661, dataGroup_lo_lo_661};
  wire [1023:0] dataGroup_hi_661 = {dataGroup_hi_hi_661, dataGroup_hi_lo_661};
  wire [7:0]    dataGroup_21_20 = dataGroup_hi_661[31:24];
  wire [1023:0] dataGroup_lo_662 = {dataGroup_lo_hi_662, dataGroup_lo_lo_662};
  wire [1023:0] dataGroup_hi_662 = {dataGroup_hi_hi_662, dataGroup_hi_lo_662};
  wire [7:0]    dataGroup_22_20 = dataGroup_hi_662[79:72];
  wire [1023:0] dataGroup_lo_663 = {dataGroup_lo_hi_663, dataGroup_lo_lo_663};
  wire [1023:0] dataGroup_hi_663 = {dataGroup_hi_hi_663, dataGroup_hi_lo_663};
  wire [7:0]    dataGroup_23_20 = dataGroup_hi_663[127:120];
  wire [1023:0] dataGroup_lo_664 = {dataGroup_lo_hi_664, dataGroup_lo_lo_664};
  wire [1023:0] dataGroup_hi_664 = {dataGroup_hi_hi_664, dataGroup_hi_lo_664};
  wire [7:0]    dataGroup_24_20 = dataGroup_hi_664[175:168];
  wire [1023:0] dataGroup_lo_665 = {dataGroup_lo_hi_665, dataGroup_lo_lo_665};
  wire [1023:0] dataGroup_hi_665 = {dataGroup_hi_hi_665, dataGroup_hi_lo_665};
  wire [7:0]    dataGroup_25_20 = dataGroup_hi_665[223:216];
  wire [1023:0] dataGroup_lo_666 = {dataGroup_lo_hi_666, dataGroup_lo_lo_666};
  wire [1023:0] dataGroup_hi_666 = {dataGroup_hi_hi_666, dataGroup_hi_lo_666};
  wire [7:0]    dataGroup_26_20 = dataGroup_hi_666[271:264];
  wire [1023:0] dataGroup_lo_667 = {dataGroup_lo_hi_667, dataGroup_lo_lo_667};
  wire [1023:0] dataGroup_hi_667 = {dataGroup_hi_hi_667, dataGroup_hi_lo_667};
  wire [7:0]    dataGroup_27_20 = dataGroup_hi_667[319:312];
  wire [1023:0] dataGroup_lo_668 = {dataGroup_lo_hi_668, dataGroup_lo_lo_668};
  wire [1023:0] dataGroup_hi_668 = {dataGroup_hi_hi_668, dataGroup_hi_lo_668};
  wire [7:0]    dataGroup_28_20 = dataGroup_hi_668[367:360];
  wire [1023:0] dataGroup_lo_669 = {dataGroup_lo_hi_669, dataGroup_lo_lo_669};
  wire [1023:0] dataGroup_hi_669 = {dataGroup_hi_hi_669, dataGroup_hi_lo_669};
  wire [7:0]    dataGroup_29_20 = dataGroup_hi_669[415:408];
  wire [1023:0] dataGroup_lo_670 = {dataGroup_lo_hi_670, dataGroup_lo_lo_670};
  wire [1023:0] dataGroup_hi_670 = {dataGroup_hi_hi_670, dataGroup_hi_lo_670};
  wire [7:0]    dataGroup_30_20 = dataGroup_hi_670[463:456];
  wire [1023:0] dataGroup_lo_671 = {dataGroup_lo_hi_671, dataGroup_lo_lo_671};
  wire [1023:0] dataGroup_hi_671 = {dataGroup_hi_hi_671, dataGroup_hi_lo_671};
  wire [7:0]    dataGroup_31_20 = dataGroup_hi_671[511:504];
  wire [15:0]   res_lo_lo_lo_lo_20 = {dataGroup_1_20, dataGroup_0_20};
  wire [15:0]   res_lo_lo_lo_hi_20 = {dataGroup_3_20, dataGroup_2_20};
  wire [31:0]   res_lo_lo_lo_20 = {res_lo_lo_lo_hi_20, res_lo_lo_lo_lo_20};
  wire [15:0]   res_lo_lo_hi_lo_20 = {dataGroup_5_20, dataGroup_4_20};
  wire [15:0]   res_lo_lo_hi_hi_20 = {dataGroup_7_20, dataGroup_6_20};
  wire [31:0]   res_lo_lo_hi_20 = {res_lo_lo_hi_hi_20, res_lo_lo_hi_lo_20};
  wire [63:0]   res_lo_lo_20 = {res_lo_lo_hi_20, res_lo_lo_lo_20};
  wire [15:0]   res_lo_hi_lo_lo_20 = {dataGroup_9_20, dataGroup_8_20};
  wire [15:0]   res_lo_hi_lo_hi_20 = {dataGroup_11_20, dataGroup_10_20};
  wire [31:0]   res_lo_hi_lo_20 = {res_lo_hi_lo_hi_20, res_lo_hi_lo_lo_20};
  wire [15:0]   res_lo_hi_hi_lo_20 = {dataGroup_13_20, dataGroup_12_20};
  wire [15:0]   res_lo_hi_hi_hi_20 = {dataGroup_15_20, dataGroup_14_20};
  wire [31:0]   res_lo_hi_hi_20 = {res_lo_hi_hi_hi_20, res_lo_hi_hi_lo_20};
  wire [63:0]   res_lo_hi_20 = {res_lo_hi_hi_20, res_lo_hi_lo_20};
  wire [127:0]  res_lo_20 = {res_lo_hi_20, res_lo_lo_20};
  wire [15:0]   res_hi_lo_lo_lo_20 = {dataGroup_17_20, dataGroup_16_20};
  wire [15:0]   res_hi_lo_lo_hi_20 = {dataGroup_19_20, dataGroup_18_20};
  wire [31:0]   res_hi_lo_lo_20 = {res_hi_lo_lo_hi_20, res_hi_lo_lo_lo_20};
  wire [15:0]   res_hi_lo_hi_lo_20 = {dataGroup_21_20, dataGroup_20_20};
  wire [15:0]   res_hi_lo_hi_hi_20 = {dataGroup_23_20, dataGroup_22_20};
  wire [31:0]   res_hi_lo_hi_20 = {res_hi_lo_hi_hi_20, res_hi_lo_hi_lo_20};
  wire [63:0]   res_hi_lo_20 = {res_hi_lo_hi_20, res_hi_lo_lo_20};
  wire [15:0]   res_hi_hi_lo_lo_20 = {dataGroup_25_20, dataGroup_24_20};
  wire [15:0]   res_hi_hi_lo_hi_20 = {dataGroup_27_20, dataGroup_26_20};
  wire [31:0]   res_hi_hi_lo_20 = {res_hi_hi_lo_hi_20, res_hi_hi_lo_lo_20};
  wire [15:0]   res_hi_hi_hi_lo_20 = {dataGroup_29_20, dataGroup_28_20};
  wire [15:0]   res_hi_hi_hi_hi_20 = {dataGroup_31_20, dataGroup_30_20};
  wire [31:0]   res_hi_hi_hi_20 = {res_hi_hi_hi_hi_20, res_hi_hi_hi_lo_20};
  wire [63:0]   res_hi_hi_20 = {res_hi_hi_hi_20, res_hi_hi_lo_20};
  wire [127:0]  res_hi_20 = {res_hi_hi_20, res_hi_lo_20};
  wire [255:0]  res_45 = {res_hi_20, res_lo_20};
  wire [511:0]  lo_lo_5 = {res_41, res_40};
  wire [511:0]  lo_hi_5 = {res_43, res_42};
  wire [1023:0] lo_5 = {lo_hi_5, lo_lo_5};
  wire [511:0]  hi_lo_5 = {res_45, res_44};
  wire [1023:0] hi_5 = {512'h0, hi_lo_5};
  wire [2047:0] regroupLoadData_0_5 = {hi_5, lo_5};
  wire [1023:0] dataGroup_lo_672 = {dataGroup_lo_hi_672, dataGroup_lo_lo_672};
  wire [1023:0] dataGroup_hi_672 = {dataGroup_hi_hi_672, dataGroup_hi_lo_672};
  wire [7:0]    dataGroup_0_21 = dataGroup_lo_672[7:0];
  wire [1023:0] dataGroup_lo_673 = {dataGroup_lo_hi_673, dataGroup_lo_lo_673};
  wire [1023:0] dataGroup_hi_673 = {dataGroup_hi_hi_673, dataGroup_hi_lo_673};
  wire [7:0]    dataGroup_1_21 = dataGroup_lo_673[63:56];
  wire [1023:0] dataGroup_lo_674 = {dataGroup_lo_hi_674, dataGroup_lo_lo_674};
  wire [1023:0] dataGroup_hi_674 = {dataGroup_hi_hi_674, dataGroup_hi_lo_674};
  wire [7:0]    dataGroup_2_21 = dataGroup_lo_674[119:112];
  wire [1023:0] dataGroup_lo_675 = {dataGroup_lo_hi_675, dataGroup_lo_lo_675};
  wire [1023:0] dataGroup_hi_675 = {dataGroup_hi_hi_675, dataGroup_hi_lo_675};
  wire [7:0]    dataGroup_3_21 = dataGroup_lo_675[175:168];
  wire [1023:0] dataGroup_lo_676 = {dataGroup_lo_hi_676, dataGroup_lo_lo_676};
  wire [1023:0] dataGroup_hi_676 = {dataGroup_hi_hi_676, dataGroup_hi_lo_676};
  wire [7:0]    dataGroup_4_21 = dataGroup_lo_676[231:224];
  wire [1023:0] dataGroup_lo_677 = {dataGroup_lo_hi_677, dataGroup_lo_lo_677};
  wire [1023:0] dataGroup_hi_677 = {dataGroup_hi_hi_677, dataGroup_hi_lo_677};
  wire [7:0]    dataGroup_5_21 = dataGroup_lo_677[287:280];
  wire [1023:0] dataGroup_lo_678 = {dataGroup_lo_hi_678, dataGroup_lo_lo_678};
  wire [1023:0] dataGroup_hi_678 = {dataGroup_hi_hi_678, dataGroup_hi_lo_678};
  wire [7:0]    dataGroup_6_21 = dataGroup_lo_678[343:336];
  wire [1023:0] dataGroup_lo_679 = {dataGroup_lo_hi_679, dataGroup_lo_lo_679};
  wire [1023:0] dataGroup_hi_679 = {dataGroup_hi_hi_679, dataGroup_hi_lo_679};
  wire [7:0]    dataGroup_7_21 = dataGroup_lo_679[399:392];
  wire [1023:0] dataGroup_lo_680 = {dataGroup_lo_hi_680, dataGroup_lo_lo_680};
  wire [1023:0] dataGroup_hi_680 = {dataGroup_hi_hi_680, dataGroup_hi_lo_680};
  wire [7:0]    dataGroup_8_21 = dataGroup_lo_680[455:448];
  wire [1023:0] dataGroup_lo_681 = {dataGroup_lo_hi_681, dataGroup_lo_lo_681};
  wire [1023:0] dataGroup_hi_681 = {dataGroup_hi_hi_681, dataGroup_hi_lo_681};
  wire [7:0]    dataGroup_9_21 = dataGroup_lo_681[511:504];
  wire [1023:0] dataGroup_lo_682 = {dataGroup_lo_hi_682, dataGroup_lo_lo_682};
  wire [1023:0] dataGroup_hi_682 = {dataGroup_hi_hi_682, dataGroup_hi_lo_682};
  wire [7:0]    dataGroup_10_21 = dataGroup_lo_682[567:560];
  wire [1023:0] dataGroup_lo_683 = {dataGroup_lo_hi_683, dataGroup_lo_lo_683};
  wire [1023:0] dataGroup_hi_683 = {dataGroup_hi_hi_683, dataGroup_hi_lo_683};
  wire [7:0]    dataGroup_11_21 = dataGroup_lo_683[623:616];
  wire [1023:0] dataGroup_lo_684 = {dataGroup_lo_hi_684, dataGroup_lo_lo_684};
  wire [1023:0] dataGroup_hi_684 = {dataGroup_hi_hi_684, dataGroup_hi_lo_684};
  wire [7:0]    dataGroup_12_21 = dataGroup_lo_684[679:672];
  wire [1023:0] dataGroup_lo_685 = {dataGroup_lo_hi_685, dataGroup_lo_lo_685};
  wire [1023:0] dataGroup_hi_685 = {dataGroup_hi_hi_685, dataGroup_hi_lo_685};
  wire [7:0]    dataGroup_13_21 = dataGroup_lo_685[735:728];
  wire [1023:0] dataGroup_lo_686 = {dataGroup_lo_hi_686, dataGroup_lo_lo_686};
  wire [1023:0] dataGroup_hi_686 = {dataGroup_hi_hi_686, dataGroup_hi_lo_686};
  wire [7:0]    dataGroup_14_21 = dataGroup_lo_686[791:784];
  wire [1023:0] dataGroup_lo_687 = {dataGroup_lo_hi_687, dataGroup_lo_lo_687};
  wire [1023:0] dataGroup_hi_687 = {dataGroup_hi_hi_687, dataGroup_hi_lo_687};
  wire [7:0]    dataGroup_15_21 = dataGroup_lo_687[847:840];
  wire [1023:0] dataGroup_lo_688 = {dataGroup_lo_hi_688, dataGroup_lo_lo_688};
  wire [1023:0] dataGroup_hi_688 = {dataGroup_hi_hi_688, dataGroup_hi_lo_688};
  wire [7:0]    dataGroup_16_21 = dataGroup_lo_688[903:896];
  wire [1023:0] dataGroup_lo_689 = {dataGroup_lo_hi_689, dataGroup_lo_lo_689};
  wire [1023:0] dataGroup_hi_689 = {dataGroup_hi_hi_689, dataGroup_hi_lo_689};
  wire [7:0]    dataGroup_17_21 = dataGroup_lo_689[959:952];
  wire [1023:0] dataGroup_lo_690 = {dataGroup_lo_hi_690, dataGroup_lo_lo_690};
  wire [1023:0] dataGroup_hi_690 = {dataGroup_hi_hi_690, dataGroup_hi_lo_690};
  wire [7:0]    dataGroup_18_21 = dataGroup_lo_690[1015:1008];
  wire [1023:0] dataGroup_lo_691 = {dataGroup_lo_hi_691, dataGroup_lo_lo_691};
  wire [1023:0] dataGroup_hi_691 = {dataGroup_hi_hi_691, dataGroup_hi_lo_691};
  wire [7:0]    dataGroup_19_21 = dataGroup_hi_691[47:40];
  wire [1023:0] dataGroup_lo_692 = {dataGroup_lo_hi_692, dataGroup_lo_lo_692};
  wire [1023:0] dataGroup_hi_692 = {dataGroup_hi_hi_692, dataGroup_hi_lo_692};
  wire [7:0]    dataGroup_20_21 = dataGroup_hi_692[103:96];
  wire [1023:0] dataGroup_lo_693 = {dataGroup_lo_hi_693, dataGroup_lo_lo_693};
  wire [1023:0] dataGroup_hi_693 = {dataGroup_hi_hi_693, dataGroup_hi_lo_693};
  wire [7:0]    dataGroup_21_21 = dataGroup_hi_693[159:152];
  wire [1023:0] dataGroup_lo_694 = {dataGroup_lo_hi_694, dataGroup_lo_lo_694};
  wire [1023:0] dataGroup_hi_694 = {dataGroup_hi_hi_694, dataGroup_hi_lo_694};
  wire [7:0]    dataGroup_22_21 = dataGroup_hi_694[215:208];
  wire [1023:0] dataGroup_lo_695 = {dataGroup_lo_hi_695, dataGroup_lo_lo_695};
  wire [1023:0] dataGroup_hi_695 = {dataGroup_hi_hi_695, dataGroup_hi_lo_695};
  wire [7:0]    dataGroup_23_21 = dataGroup_hi_695[271:264];
  wire [1023:0] dataGroup_lo_696 = {dataGroup_lo_hi_696, dataGroup_lo_lo_696};
  wire [1023:0] dataGroup_hi_696 = {dataGroup_hi_hi_696, dataGroup_hi_lo_696};
  wire [7:0]    dataGroup_24_21 = dataGroup_hi_696[327:320];
  wire [1023:0] dataGroup_lo_697 = {dataGroup_lo_hi_697, dataGroup_lo_lo_697};
  wire [1023:0] dataGroup_hi_697 = {dataGroup_hi_hi_697, dataGroup_hi_lo_697};
  wire [7:0]    dataGroup_25_21 = dataGroup_hi_697[383:376];
  wire [1023:0] dataGroup_lo_698 = {dataGroup_lo_hi_698, dataGroup_lo_lo_698};
  wire [1023:0] dataGroup_hi_698 = {dataGroup_hi_hi_698, dataGroup_hi_lo_698};
  wire [7:0]    dataGroup_26_21 = dataGroup_hi_698[439:432];
  wire [1023:0] dataGroup_lo_699 = {dataGroup_lo_hi_699, dataGroup_lo_lo_699};
  wire [1023:0] dataGroup_hi_699 = {dataGroup_hi_hi_699, dataGroup_hi_lo_699};
  wire [7:0]    dataGroup_27_21 = dataGroup_hi_699[495:488];
  wire [1023:0] dataGroup_lo_700 = {dataGroup_lo_hi_700, dataGroup_lo_lo_700};
  wire [1023:0] dataGroup_hi_700 = {dataGroup_hi_hi_700, dataGroup_hi_lo_700};
  wire [7:0]    dataGroup_28_21 = dataGroup_hi_700[551:544];
  wire [1023:0] dataGroup_lo_701 = {dataGroup_lo_hi_701, dataGroup_lo_lo_701};
  wire [1023:0] dataGroup_hi_701 = {dataGroup_hi_hi_701, dataGroup_hi_lo_701};
  wire [7:0]    dataGroup_29_21 = dataGroup_hi_701[607:600];
  wire [1023:0] dataGroup_lo_702 = {dataGroup_lo_hi_702, dataGroup_lo_lo_702};
  wire [1023:0] dataGroup_hi_702 = {dataGroup_hi_hi_702, dataGroup_hi_lo_702};
  wire [7:0]    dataGroup_30_21 = dataGroup_hi_702[663:656];
  wire [1023:0] dataGroup_lo_703 = {dataGroup_lo_hi_703, dataGroup_lo_lo_703};
  wire [1023:0] dataGroup_hi_703 = {dataGroup_hi_hi_703, dataGroup_hi_lo_703};
  wire [7:0]    dataGroup_31_21 = dataGroup_hi_703[719:712];
  wire [15:0]   res_lo_lo_lo_lo_21 = {dataGroup_1_21, dataGroup_0_21};
  wire [15:0]   res_lo_lo_lo_hi_21 = {dataGroup_3_21, dataGroup_2_21};
  wire [31:0]   res_lo_lo_lo_21 = {res_lo_lo_lo_hi_21, res_lo_lo_lo_lo_21};
  wire [15:0]   res_lo_lo_hi_lo_21 = {dataGroup_5_21, dataGroup_4_21};
  wire [15:0]   res_lo_lo_hi_hi_21 = {dataGroup_7_21, dataGroup_6_21};
  wire [31:0]   res_lo_lo_hi_21 = {res_lo_lo_hi_hi_21, res_lo_lo_hi_lo_21};
  wire [63:0]   res_lo_lo_21 = {res_lo_lo_hi_21, res_lo_lo_lo_21};
  wire [15:0]   res_lo_hi_lo_lo_21 = {dataGroup_9_21, dataGroup_8_21};
  wire [15:0]   res_lo_hi_lo_hi_21 = {dataGroup_11_21, dataGroup_10_21};
  wire [31:0]   res_lo_hi_lo_21 = {res_lo_hi_lo_hi_21, res_lo_hi_lo_lo_21};
  wire [15:0]   res_lo_hi_hi_lo_21 = {dataGroup_13_21, dataGroup_12_21};
  wire [15:0]   res_lo_hi_hi_hi_21 = {dataGroup_15_21, dataGroup_14_21};
  wire [31:0]   res_lo_hi_hi_21 = {res_lo_hi_hi_hi_21, res_lo_hi_hi_lo_21};
  wire [63:0]   res_lo_hi_21 = {res_lo_hi_hi_21, res_lo_hi_lo_21};
  wire [127:0]  res_lo_21 = {res_lo_hi_21, res_lo_lo_21};
  wire [15:0]   res_hi_lo_lo_lo_21 = {dataGroup_17_21, dataGroup_16_21};
  wire [15:0]   res_hi_lo_lo_hi_21 = {dataGroup_19_21, dataGroup_18_21};
  wire [31:0]   res_hi_lo_lo_21 = {res_hi_lo_lo_hi_21, res_hi_lo_lo_lo_21};
  wire [15:0]   res_hi_lo_hi_lo_21 = {dataGroup_21_21, dataGroup_20_21};
  wire [15:0]   res_hi_lo_hi_hi_21 = {dataGroup_23_21, dataGroup_22_21};
  wire [31:0]   res_hi_lo_hi_21 = {res_hi_lo_hi_hi_21, res_hi_lo_hi_lo_21};
  wire [63:0]   res_hi_lo_21 = {res_hi_lo_hi_21, res_hi_lo_lo_21};
  wire [15:0]   res_hi_hi_lo_lo_21 = {dataGroup_25_21, dataGroup_24_21};
  wire [15:0]   res_hi_hi_lo_hi_21 = {dataGroup_27_21, dataGroup_26_21};
  wire [31:0]   res_hi_hi_lo_21 = {res_hi_hi_lo_hi_21, res_hi_hi_lo_lo_21};
  wire [15:0]   res_hi_hi_hi_lo_21 = {dataGroup_29_21, dataGroup_28_21};
  wire [15:0]   res_hi_hi_hi_hi_21 = {dataGroup_31_21, dataGroup_30_21};
  wire [31:0]   res_hi_hi_hi_21 = {res_hi_hi_hi_hi_21, res_hi_hi_hi_lo_21};
  wire [63:0]   res_hi_hi_21 = {res_hi_hi_hi_21, res_hi_hi_lo_21};
  wire [127:0]  res_hi_21 = {res_hi_hi_21, res_hi_lo_21};
  wire [255:0]  res_48 = {res_hi_21, res_lo_21};
  wire [1023:0] dataGroup_lo_704 = {dataGroup_lo_hi_704, dataGroup_lo_lo_704};
  wire [1023:0] dataGroup_hi_704 = {dataGroup_hi_hi_704, dataGroup_hi_lo_704};
  wire [7:0]    dataGroup_0_22 = dataGroup_lo_704[15:8];
  wire [1023:0] dataGroup_lo_705 = {dataGroup_lo_hi_705, dataGroup_lo_lo_705};
  wire [1023:0] dataGroup_hi_705 = {dataGroup_hi_hi_705, dataGroup_hi_lo_705};
  wire [7:0]    dataGroup_1_22 = dataGroup_lo_705[71:64];
  wire [1023:0] dataGroup_lo_706 = {dataGroup_lo_hi_706, dataGroup_lo_lo_706};
  wire [1023:0] dataGroup_hi_706 = {dataGroup_hi_hi_706, dataGroup_hi_lo_706};
  wire [7:0]    dataGroup_2_22 = dataGroup_lo_706[127:120];
  wire [1023:0] dataGroup_lo_707 = {dataGroup_lo_hi_707, dataGroup_lo_lo_707};
  wire [1023:0] dataGroup_hi_707 = {dataGroup_hi_hi_707, dataGroup_hi_lo_707};
  wire [7:0]    dataGroup_3_22 = dataGroup_lo_707[183:176];
  wire [1023:0] dataGroup_lo_708 = {dataGroup_lo_hi_708, dataGroup_lo_lo_708};
  wire [1023:0] dataGroup_hi_708 = {dataGroup_hi_hi_708, dataGroup_hi_lo_708};
  wire [7:0]    dataGroup_4_22 = dataGroup_lo_708[239:232];
  wire [1023:0] dataGroup_lo_709 = {dataGroup_lo_hi_709, dataGroup_lo_lo_709};
  wire [1023:0] dataGroup_hi_709 = {dataGroup_hi_hi_709, dataGroup_hi_lo_709};
  wire [7:0]    dataGroup_5_22 = dataGroup_lo_709[295:288];
  wire [1023:0] dataGroup_lo_710 = {dataGroup_lo_hi_710, dataGroup_lo_lo_710};
  wire [1023:0] dataGroup_hi_710 = {dataGroup_hi_hi_710, dataGroup_hi_lo_710};
  wire [7:0]    dataGroup_6_22 = dataGroup_lo_710[351:344];
  wire [1023:0] dataGroup_lo_711 = {dataGroup_lo_hi_711, dataGroup_lo_lo_711};
  wire [1023:0] dataGroup_hi_711 = {dataGroup_hi_hi_711, dataGroup_hi_lo_711};
  wire [7:0]    dataGroup_7_22 = dataGroup_lo_711[407:400];
  wire [1023:0] dataGroup_lo_712 = {dataGroup_lo_hi_712, dataGroup_lo_lo_712};
  wire [1023:0] dataGroup_hi_712 = {dataGroup_hi_hi_712, dataGroup_hi_lo_712};
  wire [7:0]    dataGroup_8_22 = dataGroup_lo_712[463:456];
  wire [1023:0] dataGroup_lo_713 = {dataGroup_lo_hi_713, dataGroup_lo_lo_713};
  wire [1023:0] dataGroup_hi_713 = {dataGroup_hi_hi_713, dataGroup_hi_lo_713};
  wire [7:0]    dataGroup_9_22 = dataGroup_lo_713[519:512];
  wire [1023:0] dataGroup_lo_714 = {dataGroup_lo_hi_714, dataGroup_lo_lo_714};
  wire [1023:0] dataGroup_hi_714 = {dataGroup_hi_hi_714, dataGroup_hi_lo_714};
  wire [7:0]    dataGroup_10_22 = dataGroup_lo_714[575:568];
  wire [1023:0] dataGroup_lo_715 = {dataGroup_lo_hi_715, dataGroup_lo_lo_715};
  wire [1023:0] dataGroup_hi_715 = {dataGroup_hi_hi_715, dataGroup_hi_lo_715};
  wire [7:0]    dataGroup_11_22 = dataGroup_lo_715[631:624];
  wire [1023:0] dataGroup_lo_716 = {dataGroup_lo_hi_716, dataGroup_lo_lo_716};
  wire [1023:0] dataGroup_hi_716 = {dataGroup_hi_hi_716, dataGroup_hi_lo_716};
  wire [7:0]    dataGroup_12_22 = dataGroup_lo_716[687:680];
  wire [1023:0] dataGroup_lo_717 = {dataGroup_lo_hi_717, dataGroup_lo_lo_717};
  wire [1023:0] dataGroup_hi_717 = {dataGroup_hi_hi_717, dataGroup_hi_lo_717};
  wire [7:0]    dataGroup_13_22 = dataGroup_lo_717[743:736];
  wire [1023:0] dataGroup_lo_718 = {dataGroup_lo_hi_718, dataGroup_lo_lo_718};
  wire [1023:0] dataGroup_hi_718 = {dataGroup_hi_hi_718, dataGroup_hi_lo_718};
  wire [7:0]    dataGroup_14_22 = dataGroup_lo_718[799:792];
  wire [1023:0] dataGroup_lo_719 = {dataGroup_lo_hi_719, dataGroup_lo_lo_719};
  wire [1023:0] dataGroup_hi_719 = {dataGroup_hi_hi_719, dataGroup_hi_lo_719};
  wire [7:0]    dataGroup_15_22 = dataGroup_lo_719[855:848];
  wire [1023:0] dataGroup_lo_720 = {dataGroup_lo_hi_720, dataGroup_lo_lo_720};
  wire [1023:0] dataGroup_hi_720 = {dataGroup_hi_hi_720, dataGroup_hi_lo_720};
  wire [7:0]    dataGroup_16_22 = dataGroup_lo_720[911:904];
  wire [1023:0] dataGroup_lo_721 = {dataGroup_lo_hi_721, dataGroup_lo_lo_721};
  wire [1023:0] dataGroup_hi_721 = {dataGroup_hi_hi_721, dataGroup_hi_lo_721};
  wire [7:0]    dataGroup_17_22 = dataGroup_lo_721[967:960];
  wire [1023:0] dataGroup_lo_722 = {dataGroup_lo_hi_722, dataGroup_lo_lo_722};
  wire [1023:0] dataGroup_hi_722 = {dataGroup_hi_hi_722, dataGroup_hi_lo_722};
  wire [7:0]    dataGroup_18_22 = dataGroup_lo_722[1023:1016];
  wire [1023:0] dataGroup_lo_723 = {dataGroup_lo_hi_723, dataGroup_lo_lo_723};
  wire [1023:0] dataGroup_hi_723 = {dataGroup_hi_hi_723, dataGroup_hi_lo_723};
  wire [7:0]    dataGroup_19_22 = dataGroup_hi_723[55:48];
  wire [1023:0] dataGroup_lo_724 = {dataGroup_lo_hi_724, dataGroup_lo_lo_724};
  wire [1023:0] dataGroup_hi_724 = {dataGroup_hi_hi_724, dataGroup_hi_lo_724};
  wire [7:0]    dataGroup_20_22 = dataGroup_hi_724[111:104];
  wire [1023:0] dataGroup_lo_725 = {dataGroup_lo_hi_725, dataGroup_lo_lo_725};
  wire [1023:0] dataGroup_hi_725 = {dataGroup_hi_hi_725, dataGroup_hi_lo_725};
  wire [7:0]    dataGroup_21_22 = dataGroup_hi_725[167:160];
  wire [1023:0] dataGroup_lo_726 = {dataGroup_lo_hi_726, dataGroup_lo_lo_726};
  wire [1023:0] dataGroup_hi_726 = {dataGroup_hi_hi_726, dataGroup_hi_lo_726};
  wire [7:0]    dataGroup_22_22 = dataGroup_hi_726[223:216];
  wire [1023:0] dataGroup_lo_727 = {dataGroup_lo_hi_727, dataGroup_lo_lo_727};
  wire [1023:0] dataGroup_hi_727 = {dataGroup_hi_hi_727, dataGroup_hi_lo_727};
  wire [7:0]    dataGroup_23_22 = dataGroup_hi_727[279:272];
  wire [1023:0] dataGroup_lo_728 = {dataGroup_lo_hi_728, dataGroup_lo_lo_728};
  wire [1023:0] dataGroup_hi_728 = {dataGroup_hi_hi_728, dataGroup_hi_lo_728};
  wire [7:0]    dataGroup_24_22 = dataGroup_hi_728[335:328];
  wire [1023:0] dataGroup_lo_729 = {dataGroup_lo_hi_729, dataGroup_lo_lo_729};
  wire [1023:0] dataGroup_hi_729 = {dataGroup_hi_hi_729, dataGroup_hi_lo_729};
  wire [7:0]    dataGroup_25_22 = dataGroup_hi_729[391:384];
  wire [1023:0] dataGroup_lo_730 = {dataGroup_lo_hi_730, dataGroup_lo_lo_730};
  wire [1023:0] dataGroup_hi_730 = {dataGroup_hi_hi_730, dataGroup_hi_lo_730};
  wire [7:0]    dataGroup_26_22 = dataGroup_hi_730[447:440];
  wire [1023:0] dataGroup_lo_731 = {dataGroup_lo_hi_731, dataGroup_lo_lo_731};
  wire [1023:0] dataGroup_hi_731 = {dataGroup_hi_hi_731, dataGroup_hi_lo_731};
  wire [7:0]    dataGroup_27_22 = dataGroup_hi_731[503:496];
  wire [1023:0] dataGroup_lo_732 = {dataGroup_lo_hi_732, dataGroup_lo_lo_732};
  wire [1023:0] dataGroup_hi_732 = {dataGroup_hi_hi_732, dataGroup_hi_lo_732};
  wire [7:0]    dataGroup_28_22 = dataGroup_hi_732[559:552];
  wire [1023:0] dataGroup_lo_733 = {dataGroup_lo_hi_733, dataGroup_lo_lo_733};
  wire [1023:0] dataGroup_hi_733 = {dataGroup_hi_hi_733, dataGroup_hi_lo_733};
  wire [7:0]    dataGroup_29_22 = dataGroup_hi_733[615:608];
  wire [1023:0] dataGroup_lo_734 = {dataGroup_lo_hi_734, dataGroup_lo_lo_734};
  wire [1023:0] dataGroup_hi_734 = {dataGroup_hi_hi_734, dataGroup_hi_lo_734};
  wire [7:0]    dataGroup_30_22 = dataGroup_hi_734[671:664];
  wire [1023:0] dataGroup_lo_735 = {dataGroup_lo_hi_735, dataGroup_lo_lo_735};
  wire [1023:0] dataGroup_hi_735 = {dataGroup_hi_hi_735, dataGroup_hi_lo_735};
  wire [7:0]    dataGroup_31_22 = dataGroup_hi_735[727:720];
  wire [15:0]   res_lo_lo_lo_lo_22 = {dataGroup_1_22, dataGroup_0_22};
  wire [15:0]   res_lo_lo_lo_hi_22 = {dataGroup_3_22, dataGroup_2_22};
  wire [31:0]   res_lo_lo_lo_22 = {res_lo_lo_lo_hi_22, res_lo_lo_lo_lo_22};
  wire [15:0]   res_lo_lo_hi_lo_22 = {dataGroup_5_22, dataGroup_4_22};
  wire [15:0]   res_lo_lo_hi_hi_22 = {dataGroup_7_22, dataGroup_6_22};
  wire [31:0]   res_lo_lo_hi_22 = {res_lo_lo_hi_hi_22, res_lo_lo_hi_lo_22};
  wire [63:0]   res_lo_lo_22 = {res_lo_lo_hi_22, res_lo_lo_lo_22};
  wire [15:0]   res_lo_hi_lo_lo_22 = {dataGroup_9_22, dataGroup_8_22};
  wire [15:0]   res_lo_hi_lo_hi_22 = {dataGroup_11_22, dataGroup_10_22};
  wire [31:0]   res_lo_hi_lo_22 = {res_lo_hi_lo_hi_22, res_lo_hi_lo_lo_22};
  wire [15:0]   res_lo_hi_hi_lo_22 = {dataGroup_13_22, dataGroup_12_22};
  wire [15:0]   res_lo_hi_hi_hi_22 = {dataGroup_15_22, dataGroup_14_22};
  wire [31:0]   res_lo_hi_hi_22 = {res_lo_hi_hi_hi_22, res_lo_hi_hi_lo_22};
  wire [63:0]   res_lo_hi_22 = {res_lo_hi_hi_22, res_lo_hi_lo_22};
  wire [127:0]  res_lo_22 = {res_lo_hi_22, res_lo_lo_22};
  wire [15:0]   res_hi_lo_lo_lo_22 = {dataGroup_17_22, dataGroup_16_22};
  wire [15:0]   res_hi_lo_lo_hi_22 = {dataGroup_19_22, dataGroup_18_22};
  wire [31:0]   res_hi_lo_lo_22 = {res_hi_lo_lo_hi_22, res_hi_lo_lo_lo_22};
  wire [15:0]   res_hi_lo_hi_lo_22 = {dataGroup_21_22, dataGroup_20_22};
  wire [15:0]   res_hi_lo_hi_hi_22 = {dataGroup_23_22, dataGroup_22_22};
  wire [31:0]   res_hi_lo_hi_22 = {res_hi_lo_hi_hi_22, res_hi_lo_hi_lo_22};
  wire [63:0]   res_hi_lo_22 = {res_hi_lo_hi_22, res_hi_lo_lo_22};
  wire [15:0]   res_hi_hi_lo_lo_22 = {dataGroup_25_22, dataGroup_24_22};
  wire [15:0]   res_hi_hi_lo_hi_22 = {dataGroup_27_22, dataGroup_26_22};
  wire [31:0]   res_hi_hi_lo_22 = {res_hi_hi_lo_hi_22, res_hi_hi_lo_lo_22};
  wire [15:0]   res_hi_hi_hi_lo_22 = {dataGroup_29_22, dataGroup_28_22};
  wire [15:0]   res_hi_hi_hi_hi_22 = {dataGroup_31_22, dataGroup_30_22};
  wire [31:0]   res_hi_hi_hi_22 = {res_hi_hi_hi_hi_22, res_hi_hi_hi_lo_22};
  wire [63:0]   res_hi_hi_22 = {res_hi_hi_hi_22, res_hi_hi_lo_22};
  wire [127:0]  res_hi_22 = {res_hi_hi_22, res_hi_lo_22};
  wire [255:0]  res_49 = {res_hi_22, res_lo_22};
  wire [1023:0] dataGroup_lo_736 = {dataGroup_lo_hi_736, dataGroup_lo_lo_736};
  wire [1023:0] dataGroup_hi_736 = {dataGroup_hi_hi_736, dataGroup_hi_lo_736};
  wire [7:0]    dataGroup_0_23 = dataGroup_lo_736[23:16];
  wire [1023:0] dataGroup_lo_737 = {dataGroup_lo_hi_737, dataGroup_lo_lo_737};
  wire [1023:0] dataGroup_hi_737 = {dataGroup_hi_hi_737, dataGroup_hi_lo_737};
  wire [7:0]    dataGroup_1_23 = dataGroup_lo_737[79:72];
  wire [1023:0] dataGroup_lo_738 = {dataGroup_lo_hi_738, dataGroup_lo_lo_738};
  wire [1023:0] dataGroup_hi_738 = {dataGroup_hi_hi_738, dataGroup_hi_lo_738};
  wire [7:0]    dataGroup_2_23 = dataGroup_lo_738[135:128];
  wire [1023:0] dataGroup_lo_739 = {dataGroup_lo_hi_739, dataGroup_lo_lo_739};
  wire [1023:0] dataGroup_hi_739 = {dataGroup_hi_hi_739, dataGroup_hi_lo_739};
  wire [7:0]    dataGroup_3_23 = dataGroup_lo_739[191:184];
  wire [1023:0] dataGroup_lo_740 = {dataGroup_lo_hi_740, dataGroup_lo_lo_740};
  wire [1023:0] dataGroup_hi_740 = {dataGroup_hi_hi_740, dataGroup_hi_lo_740};
  wire [7:0]    dataGroup_4_23 = dataGroup_lo_740[247:240];
  wire [1023:0] dataGroup_lo_741 = {dataGroup_lo_hi_741, dataGroup_lo_lo_741};
  wire [1023:0] dataGroup_hi_741 = {dataGroup_hi_hi_741, dataGroup_hi_lo_741};
  wire [7:0]    dataGroup_5_23 = dataGroup_lo_741[303:296];
  wire [1023:0] dataGroup_lo_742 = {dataGroup_lo_hi_742, dataGroup_lo_lo_742};
  wire [1023:0] dataGroup_hi_742 = {dataGroup_hi_hi_742, dataGroup_hi_lo_742};
  wire [7:0]    dataGroup_6_23 = dataGroup_lo_742[359:352];
  wire [1023:0] dataGroup_lo_743 = {dataGroup_lo_hi_743, dataGroup_lo_lo_743};
  wire [1023:0] dataGroup_hi_743 = {dataGroup_hi_hi_743, dataGroup_hi_lo_743};
  wire [7:0]    dataGroup_7_23 = dataGroup_lo_743[415:408];
  wire [1023:0] dataGroup_lo_744 = {dataGroup_lo_hi_744, dataGroup_lo_lo_744};
  wire [1023:0] dataGroup_hi_744 = {dataGroup_hi_hi_744, dataGroup_hi_lo_744};
  wire [7:0]    dataGroup_8_23 = dataGroup_lo_744[471:464];
  wire [1023:0] dataGroup_lo_745 = {dataGroup_lo_hi_745, dataGroup_lo_lo_745};
  wire [1023:0] dataGroup_hi_745 = {dataGroup_hi_hi_745, dataGroup_hi_lo_745};
  wire [7:0]    dataGroup_9_23 = dataGroup_lo_745[527:520];
  wire [1023:0] dataGroup_lo_746 = {dataGroup_lo_hi_746, dataGroup_lo_lo_746};
  wire [1023:0] dataGroup_hi_746 = {dataGroup_hi_hi_746, dataGroup_hi_lo_746};
  wire [7:0]    dataGroup_10_23 = dataGroup_lo_746[583:576];
  wire [1023:0] dataGroup_lo_747 = {dataGroup_lo_hi_747, dataGroup_lo_lo_747};
  wire [1023:0] dataGroup_hi_747 = {dataGroup_hi_hi_747, dataGroup_hi_lo_747};
  wire [7:0]    dataGroup_11_23 = dataGroup_lo_747[639:632];
  wire [1023:0] dataGroup_lo_748 = {dataGroup_lo_hi_748, dataGroup_lo_lo_748};
  wire [1023:0] dataGroup_hi_748 = {dataGroup_hi_hi_748, dataGroup_hi_lo_748};
  wire [7:0]    dataGroup_12_23 = dataGroup_lo_748[695:688];
  wire [1023:0] dataGroup_lo_749 = {dataGroup_lo_hi_749, dataGroup_lo_lo_749};
  wire [1023:0] dataGroup_hi_749 = {dataGroup_hi_hi_749, dataGroup_hi_lo_749};
  wire [7:0]    dataGroup_13_23 = dataGroup_lo_749[751:744];
  wire [1023:0] dataGroup_lo_750 = {dataGroup_lo_hi_750, dataGroup_lo_lo_750};
  wire [1023:0] dataGroup_hi_750 = {dataGroup_hi_hi_750, dataGroup_hi_lo_750};
  wire [7:0]    dataGroup_14_23 = dataGroup_lo_750[807:800];
  wire [1023:0] dataGroup_lo_751 = {dataGroup_lo_hi_751, dataGroup_lo_lo_751};
  wire [1023:0] dataGroup_hi_751 = {dataGroup_hi_hi_751, dataGroup_hi_lo_751};
  wire [7:0]    dataGroup_15_23 = dataGroup_lo_751[863:856];
  wire [1023:0] dataGroup_lo_752 = {dataGroup_lo_hi_752, dataGroup_lo_lo_752};
  wire [1023:0] dataGroup_hi_752 = {dataGroup_hi_hi_752, dataGroup_hi_lo_752};
  wire [7:0]    dataGroup_16_23 = dataGroup_lo_752[919:912];
  wire [1023:0] dataGroup_lo_753 = {dataGroup_lo_hi_753, dataGroup_lo_lo_753};
  wire [1023:0] dataGroup_hi_753 = {dataGroup_hi_hi_753, dataGroup_hi_lo_753};
  wire [7:0]    dataGroup_17_23 = dataGroup_lo_753[975:968];
  wire [1023:0] dataGroup_lo_754 = {dataGroup_lo_hi_754, dataGroup_lo_lo_754};
  wire [1023:0] dataGroup_hi_754 = {dataGroup_hi_hi_754, dataGroup_hi_lo_754};
  wire [7:0]    dataGroup_18_23 = dataGroup_hi_754[7:0];
  wire [1023:0] dataGroup_lo_755 = {dataGroup_lo_hi_755, dataGroup_lo_lo_755};
  wire [1023:0] dataGroup_hi_755 = {dataGroup_hi_hi_755, dataGroup_hi_lo_755};
  wire [7:0]    dataGroup_19_23 = dataGroup_hi_755[63:56];
  wire [1023:0] dataGroup_lo_756 = {dataGroup_lo_hi_756, dataGroup_lo_lo_756};
  wire [1023:0] dataGroup_hi_756 = {dataGroup_hi_hi_756, dataGroup_hi_lo_756};
  wire [7:0]    dataGroup_20_23 = dataGroup_hi_756[119:112];
  wire [1023:0] dataGroup_lo_757 = {dataGroup_lo_hi_757, dataGroup_lo_lo_757};
  wire [1023:0] dataGroup_hi_757 = {dataGroup_hi_hi_757, dataGroup_hi_lo_757};
  wire [7:0]    dataGroup_21_23 = dataGroup_hi_757[175:168];
  wire [1023:0] dataGroup_lo_758 = {dataGroup_lo_hi_758, dataGroup_lo_lo_758};
  wire [1023:0] dataGroup_hi_758 = {dataGroup_hi_hi_758, dataGroup_hi_lo_758};
  wire [7:0]    dataGroup_22_23 = dataGroup_hi_758[231:224];
  wire [1023:0] dataGroup_lo_759 = {dataGroup_lo_hi_759, dataGroup_lo_lo_759};
  wire [1023:0] dataGroup_hi_759 = {dataGroup_hi_hi_759, dataGroup_hi_lo_759};
  wire [7:0]    dataGroup_23_23 = dataGroup_hi_759[287:280];
  wire [1023:0] dataGroup_lo_760 = {dataGroup_lo_hi_760, dataGroup_lo_lo_760};
  wire [1023:0] dataGroup_hi_760 = {dataGroup_hi_hi_760, dataGroup_hi_lo_760};
  wire [7:0]    dataGroup_24_23 = dataGroup_hi_760[343:336];
  wire [1023:0] dataGroup_lo_761 = {dataGroup_lo_hi_761, dataGroup_lo_lo_761};
  wire [1023:0] dataGroup_hi_761 = {dataGroup_hi_hi_761, dataGroup_hi_lo_761};
  wire [7:0]    dataGroup_25_23 = dataGroup_hi_761[399:392];
  wire [1023:0] dataGroup_lo_762 = {dataGroup_lo_hi_762, dataGroup_lo_lo_762};
  wire [1023:0] dataGroup_hi_762 = {dataGroup_hi_hi_762, dataGroup_hi_lo_762};
  wire [7:0]    dataGroup_26_23 = dataGroup_hi_762[455:448];
  wire [1023:0] dataGroup_lo_763 = {dataGroup_lo_hi_763, dataGroup_lo_lo_763};
  wire [1023:0] dataGroup_hi_763 = {dataGroup_hi_hi_763, dataGroup_hi_lo_763};
  wire [7:0]    dataGroup_27_23 = dataGroup_hi_763[511:504];
  wire [1023:0] dataGroup_lo_764 = {dataGroup_lo_hi_764, dataGroup_lo_lo_764};
  wire [1023:0] dataGroup_hi_764 = {dataGroup_hi_hi_764, dataGroup_hi_lo_764};
  wire [7:0]    dataGroup_28_23 = dataGroup_hi_764[567:560];
  wire [1023:0] dataGroup_lo_765 = {dataGroup_lo_hi_765, dataGroup_lo_lo_765};
  wire [1023:0] dataGroup_hi_765 = {dataGroup_hi_hi_765, dataGroup_hi_lo_765};
  wire [7:0]    dataGroup_29_23 = dataGroup_hi_765[623:616];
  wire [1023:0] dataGroup_lo_766 = {dataGroup_lo_hi_766, dataGroup_lo_lo_766};
  wire [1023:0] dataGroup_hi_766 = {dataGroup_hi_hi_766, dataGroup_hi_lo_766};
  wire [7:0]    dataGroup_30_23 = dataGroup_hi_766[679:672];
  wire [1023:0] dataGroup_lo_767 = {dataGroup_lo_hi_767, dataGroup_lo_lo_767};
  wire [1023:0] dataGroup_hi_767 = {dataGroup_hi_hi_767, dataGroup_hi_lo_767};
  wire [7:0]    dataGroup_31_23 = dataGroup_hi_767[735:728];
  wire [15:0]   res_lo_lo_lo_lo_23 = {dataGroup_1_23, dataGroup_0_23};
  wire [15:0]   res_lo_lo_lo_hi_23 = {dataGroup_3_23, dataGroup_2_23};
  wire [31:0]   res_lo_lo_lo_23 = {res_lo_lo_lo_hi_23, res_lo_lo_lo_lo_23};
  wire [15:0]   res_lo_lo_hi_lo_23 = {dataGroup_5_23, dataGroup_4_23};
  wire [15:0]   res_lo_lo_hi_hi_23 = {dataGroup_7_23, dataGroup_6_23};
  wire [31:0]   res_lo_lo_hi_23 = {res_lo_lo_hi_hi_23, res_lo_lo_hi_lo_23};
  wire [63:0]   res_lo_lo_23 = {res_lo_lo_hi_23, res_lo_lo_lo_23};
  wire [15:0]   res_lo_hi_lo_lo_23 = {dataGroup_9_23, dataGroup_8_23};
  wire [15:0]   res_lo_hi_lo_hi_23 = {dataGroup_11_23, dataGroup_10_23};
  wire [31:0]   res_lo_hi_lo_23 = {res_lo_hi_lo_hi_23, res_lo_hi_lo_lo_23};
  wire [15:0]   res_lo_hi_hi_lo_23 = {dataGroup_13_23, dataGroup_12_23};
  wire [15:0]   res_lo_hi_hi_hi_23 = {dataGroup_15_23, dataGroup_14_23};
  wire [31:0]   res_lo_hi_hi_23 = {res_lo_hi_hi_hi_23, res_lo_hi_hi_lo_23};
  wire [63:0]   res_lo_hi_23 = {res_lo_hi_hi_23, res_lo_hi_lo_23};
  wire [127:0]  res_lo_23 = {res_lo_hi_23, res_lo_lo_23};
  wire [15:0]   res_hi_lo_lo_lo_23 = {dataGroup_17_23, dataGroup_16_23};
  wire [15:0]   res_hi_lo_lo_hi_23 = {dataGroup_19_23, dataGroup_18_23};
  wire [31:0]   res_hi_lo_lo_23 = {res_hi_lo_lo_hi_23, res_hi_lo_lo_lo_23};
  wire [15:0]   res_hi_lo_hi_lo_23 = {dataGroup_21_23, dataGroup_20_23};
  wire [15:0]   res_hi_lo_hi_hi_23 = {dataGroup_23_23, dataGroup_22_23};
  wire [31:0]   res_hi_lo_hi_23 = {res_hi_lo_hi_hi_23, res_hi_lo_hi_lo_23};
  wire [63:0]   res_hi_lo_23 = {res_hi_lo_hi_23, res_hi_lo_lo_23};
  wire [15:0]   res_hi_hi_lo_lo_23 = {dataGroup_25_23, dataGroup_24_23};
  wire [15:0]   res_hi_hi_lo_hi_23 = {dataGroup_27_23, dataGroup_26_23};
  wire [31:0]   res_hi_hi_lo_23 = {res_hi_hi_lo_hi_23, res_hi_hi_lo_lo_23};
  wire [15:0]   res_hi_hi_hi_lo_23 = {dataGroup_29_23, dataGroup_28_23};
  wire [15:0]   res_hi_hi_hi_hi_23 = {dataGroup_31_23, dataGroup_30_23};
  wire [31:0]   res_hi_hi_hi_23 = {res_hi_hi_hi_hi_23, res_hi_hi_hi_lo_23};
  wire [63:0]   res_hi_hi_23 = {res_hi_hi_hi_23, res_hi_hi_lo_23};
  wire [127:0]  res_hi_23 = {res_hi_hi_23, res_hi_lo_23};
  wire [255:0]  res_50 = {res_hi_23, res_lo_23};
  wire [1023:0] dataGroup_lo_768 = {dataGroup_lo_hi_768, dataGroup_lo_lo_768};
  wire [1023:0] dataGroup_hi_768 = {dataGroup_hi_hi_768, dataGroup_hi_lo_768};
  wire [7:0]    dataGroup_0_24 = dataGroup_lo_768[31:24];
  wire [1023:0] dataGroup_lo_769 = {dataGroup_lo_hi_769, dataGroup_lo_lo_769};
  wire [1023:0] dataGroup_hi_769 = {dataGroup_hi_hi_769, dataGroup_hi_lo_769};
  wire [7:0]    dataGroup_1_24 = dataGroup_lo_769[87:80];
  wire [1023:0] dataGroup_lo_770 = {dataGroup_lo_hi_770, dataGroup_lo_lo_770};
  wire [1023:0] dataGroup_hi_770 = {dataGroup_hi_hi_770, dataGroup_hi_lo_770};
  wire [7:0]    dataGroup_2_24 = dataGroup_lo_770[143:136];
  wire [1023:0] dataGroup_lo_771 = {dataGroup_lo_hi_771, dataGroup_lo_lo_771};
  wire [1023:0] dataGroup_hi_771 = {dataGroup_hi_hi_771, dataGroup_hi_lo_771};
  wire [7:0]    dataGroup_3_24 = dataGroup_lo_771[199:192];
  wire [1023:0] dataGroup_lo_772 = {dataGroup_lo_hi_772, dataGroup_lo_lo_772};
  wire [1023:0] dataGroup_hi_772 = {dataGroup_hi_hi_772, dataGroup_hi_lo_772};
  wire [7:0]    dataGroup_4_24 = dataGroup_lo_772[255:248];
  wire [1023:0] dataGroup_lo_773 = {dataGroup_lo_hi_773, dataGroup_lo_lo_773};
  wire [1023:0] dataGroup_hi_773 = {dataGroup_hi_hi_773, dataGroup_hi_lo_773};
  wire [7:0]    dataGroup_5_24 = dataGroup_lo_773[311:304];
  wire [1023:0] dataGroup_lo_774 = {dataGroup_lo_hi_774, dataGroup_lo_lo_774};
  wire [1023:0] dataGroup_hi_774 = {dataGroup_hi_hi_774, dataGroup_hi_lo_774};
  wire [7:0]    dataGroup_6_24 = dataGroup_lo_774[367:360];
  wire [1023:0] dataGroup_lo_775 = {dataGroup_lo_hi_775, dataGroup_lo_lo_775};
  wire [1023:0] dataGroup_hi_775 = {dataGroup_hi_hi_775, dataGroup_hi_lo_775};
  wire [7:0]    dataGroup_7_24 = dataGroup_lo_775[423:416];
  wire [1023:0] dataGroup_lo_776 = {dataGroup_lo_hi_776, dataGroup_lo_lo_776};
  wire [1023:0] dataGroup_hi_776 = {dataGroup_hi_hi_776, dataGroup_hi_lo_776};
  wire [7:0]    dataGroup_8_24 = dataGroup_lo_776[479:472];
  wire [1023:0] dataGroup_lo_777 = {dataGroup_lo_hi_777, dataGroup_lo_lo_777};
  wire [1023:0] dataGroup_hi_777 = {dataGroup_hi_hi_777, dataGroup_hi_lo_777};
  wire [7:0]    dataGroup_9_24 = dataGroup_lo_777[535:528];
  wire [1023:0] dataGroup_lo_778 = {dataGroup_lo_hi_778, dataGroup_lo_lo_778};
  wire [1023:0] dataGroup_hi_778 = {dataGroup_hi_hi_778, dataGroup_hi_lo_778};
  wire [7:0]    dataGroup_10_24 = dataGroup_lo_778[591:584];
  wire [1023:0] dataGroup_lo_779 = {dataGroup_lo_hi_779, dataGroup_lo_lo_779};
  wire [1023:0] dataGroup_hi_779 = {dataGroup_hi_hi_779, dataGroup_hi_lo_779};
  wire [7:0]    dataGroup_11_24 = dataGroup_lo_779[647:640];
  wire [1023:0] dataGroup_lo_780 = {dataGroup_lo_hi_780, dataGroup_lo_lo_780};
  wire [1023:0] dataGroup_hi_780 = {dataGroup_hi_hi_780, dataGroup_hi_lo_780};
  wire [7:0]    dataGroup_12_24 = dataGroup_lo_780[703:696];
  wire [1023:0] dataGroup_lo_781 = {dataGroup_lo_hi_781, dataGroup_lo_lo_781};
  wire [1023:0] dataGroup_hi_781 = {dataGroup_hi_hi_781, dataGroup_hi_lo_781};
  wire [7:0]    dataGroup_13_24 = dataGroup_lo_781[759:752];
  wire [1023:0] dataGroup_lo_782 = {dataGroup_lo_hi_782, dataGroup_lo_lo_782};
  wire [1023:0] dataGroup_hi_782 = {dataGroup_hi_hi_782, dataGroup_hi_lo_782};
  wire [7:0]    dataGroup_14_24 = dataGroup_lo_782[815:808];
  wire [1023:0] dataGroup_lo_783 = {dataGroup_lo_hi_783, dataGroup_lo_lo_783};
  wire [1023:0] dataGroup_hi_783 = {dataGroup_hi_hi_783, dataGroup_hi_lo_783};
  wire [7:0]    dataGroup_15_24 = dataGroup_lo_783[871:864];
  wire [1023:0] dataGroup_lo_784 = {dataGroup_lo_hi_784, dataGroup_lo_lo_784};
  wire [1023:0] dataGroup_hi_784 = {dataGroup_hi_hi_784, dataGroup_hi_lo_784};
  wire [7:0]    dataGroup_16_24 = dataGroup_lo_784[927:920];
  wire [1023:0] dataGroup_lo_785 = {dataGroup_lo_hi_785, dataGroup_lo_lo_785};
  wire [1023:0] dataGroup_hi_785 = {dataGroup_hi_hi_785, dataGroup_hi_lo_785};
  wire [7:0]    dataGroup_17_24 = dataGroup_lo_785[983:976];
  wire [1023:0] dataGroup_lo_786 = {dataGroup_lo_hi_786, dataGroup_lo_lo_786};
  wire [1023:0] dataGroup_hi_786 = {dataGroup_hi_hi_786, dataGroup_hi_lo_786};
  wire [7:0]    dataGroup_18_24 = dataGroup_hi_786[15:8];
  wire [1023:0] dataGroup_lo_787 = {dataGroup_lo_hi_787, dataGroup_lo_lo_787};
  wire [1023:0] dataGroup_hi_787 = {dataGroup_hi_hi_787, dataGroup_hi_lo_787};
  wire [7:0]    dataGroup_19_24 = dataGroup_hi_787[71:64];
  wire [1023:0] dataGroup_lo_788 = {dataGroup_lo_hi_788, dataGroup_lo_lo_788};
  wire [1023:0] dataGroup_hi_788 = {dataGroup_hi_hi_788, dataGroup_hi_lo_788};
  wire [7:0]    dataGroup_20_24 = dataGroup_hi_788[127:120];
  wire [1023:0] dataGroup_lo_789 = {dataGroup_lo_hi_789, dataGroup_lo_lo_789};
  wire [1023:0] dataGroup_hi_789 = {dataGroup_hi_hi_789, dataGroup_hi_lo_789};
  wire [7:0]    dataGroup_21_24 = dataGroup_hi_789[183:176];
  wire [1023:0] dataGroup_lo_790 = {dataGroup_lo_hi_790, dataGroup_lo_lo_790};
  wire [1023:0] dataGroup_hi_790 = {dataGroup_hi_hi_790, dataGroup_hi_lo_790};
  wire [7:0]    dataGroup_22_24 = dataGroup_hi_790[239:232];
  wire [1023:0] dataGroup_lo_791 = {dataGroup_lo_hi_791, dataGroup_lo_lo_791};
  wire [1023:0] dataGroup_hi_791 = {dataGroup_hi_hi_791, dataGroup_hi_lo_791};
  wire [7:0]    dataGroup_23_24 = dataGroup_hi_791[295:288];
  wire [1023:0] dataGroup_lo_792 = {dataGroup_lo_hi_792, dataGroup_lo_lo_792};
  wire [1023:0] dataGroup_hi_792 = {dataGroup_hi_hi_792, dataGroup_hi_lo_792};
  wire [7:0]    dataGroup_24_24 = dataGroup_hi_792[351:344];
  wire [1023:0] dataGroup_lo_793 = {dataGroup_lo_hi_793, dataGroup_lo_lo_793};
  wire [1023:0] dataGroup_hi_793 = {dataGroup_hi_hi_793, dataGroup_hi_lo_793};
  wire [7:0]    dataGroup_25_24 = dataGroup_hi_793[407:400];
  wire [1023:0] dataGroup_lo_794 = {dataGroup_lo_hi_794, dataGroup_lo_lo_794};
  wire [1023:0] dataGroup_hi_794 = {dataGroup_hi_hi_794, dataGroup_hi_lo_794};
  wire [7:0]    dataGroup_26_24 = dataGroup_hi_794[463:456];
  wire [1023:0] dataGroup_lo_795 = {dataGroup_lo_hi_795, dataGroup_lo_lo_795};
  wire [1023:0] dataGroup_hi_795 = {dataGroup_hi_hi_795, dataGroup_hi_lo_795};
  wire [7:0]    dataGroup_27_24 = dataGroup_hi_795[519:512];
  wire [1023:0] dataGroup_lo_796 = {dataGroup_lo_hi_796, dataGroup_lo_lo_796};
  wire [1023:0] dataGroup_hi_796 = {dataGroup_hi_hi_796, dataGroup_hi_lo_796};
  wire [7:0]    dataGroup_28_24 = dataGroup_hi_796[575:568];
  wire [1023:0] dataGroup_lo_797 = {dataGroup_lo_hi_797, dataGroup_lo_lo_797};
  wire [1023:0] dataGroup_hi_797 = {dataGroup_hi_hi_797, dataGroup_hi_lo_797};
  wire [7:0]    dataGroup_29_24 = dataGroup_hi_797[631:624];
  wire [1023:0] dataGroup_lo_798 = {dataGroup_lo_hi_798, dataGroup_lo_lo_798};
  wire [1023:0] dataGroup_hi_798 = {dataGroup_hi_hi_798, dataGroup_hi_lo_798};
  wire [7:0]    dataGroup_30_24 = dataGroup_hi_798[687:680];
  wire [1023:0] dataGroup_lo_799 = {dataGroup_lo_hi_799, dataGroup_lo_lo_799};
  wire [1023:0] dataGroup_hi_799 = {dataGroup_hi_hi_799, dataGroup_hi_lo_799};
  wire [7:0]    dataGroup_31_24 = dataGroup_hi_799[743:736];
  wire [15:0]   res_lo_lo_lo_lo_24 = {dataGroup_1_24, dataGroup_0_24};
  wire [15:0]   res_lo_lo_lo_hi_24 = {dataGroup_3_24, dataGroup_2_24};
  wire [31:0]   res_lo_lo_lo_24 = {res_lo_lo_lo_hi_24, res_lo_lo_lo_lo_24};
  wire [15:0]   res_lo_lo_hi_lo_24 = {dataGroup_5_24, dataGroup_4_24};
  wire [15:0]   res_lo_lo_hi_hi_24 = {dataGroup_7_24, dataGroup_6_24};
  wire [31:0]   res_lo_lo_hi_24 = {res_lo_lo_hi_hi_24, res_lo_lo_hi_lo_24};
  wire [63:0]   res_lo_lo_24 = {res_lo_lo_hi_24, res_lo_lo_lo_24};
  wire [15:0]   res_lo_hi_lo_lo_24 = {dataGroup_9_24, dataGroup_8_24};
  wire [15:0]   res_lo_hi_lo_hi_24 = {dataGroup_11_24, dataGroup_10_24};
  wire [31:0]   res_lo_hi_lo_24 = {res_lo_hi_lo_hi_24, res_lo_hi_lo_lo_24};
  wire [15:0]   res_lo_hi_hi_lo_24 = {dataGroup_13_24, dataGroup_12_24};
  wire [15:0]   res_lo_hi_hi_hi_24 = {dataGroup_15_24, dataGroup_14_24};
  wire [31:0]   res_lo_hi_hi_24 = {res_lo_hi_hi_hi_24, res_lo_hi_hi_lo_24};
  wire [63:0]   res_lo_hi_24 = {res_lo_hi_hi_24, res_lo_hi_lo_24};
  wire [127:0]  res_lo_24 = {res_lo_hi_24, res_lo_lo_24};
  wire [15:0]   res_hi_lo_lo_lo_24 = {dataGroup_17_24, dataGroup_16_24};
  wire [15:0]   res_hi_lo_lo_hi_24 = {dataGroup_19_24, dataGroup_18_24};
  wire [31:0]   res_hi_lo_lo_24 = {res_hi_lo_lo_hi_24, res_hi_lo_lo_lo_24};
  wire [15:0]   res_hi_lo_hi_lo_24 = {dataGroup_21_24, dataGroup_20_24};
  wire [15:0]   res_hi_lo_hi_hi_24 = {dataGroup_23_24, dataGroup_22_24};
  wire [31:0]   res_hi_lo_hi_24 = {res_hi_lo_hi_hi_24, res_hi_lo_hi_lo_24};
  wire [63:0]   res_hi_lo_24 = {res_hi_lo_hi_24, res_hi_lo_lo_24};
  wire [15:0]   res_hi_hi_lo_lo_24 = {dataGroup_25_24, dataGroup_24_24};
  wire [15:0]   res_hi_hi_lo_hi_24 = {dataGroup_27_24, dataGroup_26_24};
  wire [31:0]   res_hi_hi_lo_24 = {res_hi_hi_lo_hi_24, res_hi_hi_lo_lo_24};
  wire [15:0]   res_hi_hi_hi_lo_24 = {dataGroup_29_24, dataGroup_28_24};
  wire [15:0]   res_hi_hi_hi_hi_24 = {dataGroup_31_24, dataGroup_30_24};
  wire [31:0]   res_hi_hi_hi_24 = {res_hi_hi_hi_hi_24, res_hi_hi_hi_lo_24};
  wire [63:0]   res_hi_hi_24 = {res_hi_hi_hi_24, res_hi_hi_lo_24};
  wire [127:0]  res_hi_24 = {res_hi_hi_24, res_hi_lo_24};
  wire [255:0]  res_51 = {res_hi_24, res_lo_24};
  wire [1023:0] dataGroup_lo_800 = {dataGroup_lo_hi_800, dataGroup_lo_lo_800};
  wire [1023:0] dataGroup_hi_800 = {dataGroup_hi_hi_800, dataGroup_hi_lo_800};
  wire [7:0]    dataGroup_0_25 = dataGroup_lo_800[39:32];
  wire [1023:0] dataGroup_lo_801 = {dataGroup_lo_hi_801, dataGroup_lo_lo_801};
  wire [1023:0] dataGroup_hi_801 = {dataGroup_hi_hi_801, dataGroup_hi_lo_801};
  wire [7:0]    dataGroup_1_25 = dataGroup_lo_801[95:88];
  wire [1023:0] dataGroup_lo_802 = {dataGroup_lo_hi_802, dataGroup_lo_lo_802};
  wire [1023:0] dataGroup_hi_802 = {dataGroup_hi_hi_802, dataGroup_hi_lo_802};
  wire [7:0]    dataGroup_2_25 = dataGroup_lo_802[151:144];
  wire [1023:0] dataGroup_lo_803 = {dataGroup_lo_hi_803, dataGroup_lo_lo_803};
  wire [1023:0] dataGroup_hi_803 = {dataGroup_hi_hi_803, dataGroup_hi_lo_803};
  wire [7:0]    dataGroup_3_25 = dataGroup_lo_803[207:200];
  wire [1023:0] dataGroup_lo_804 = {dataGroup_lo_hi_804, dataGroup_lo_lo_804};
  wire [1023:0] dataGroup_hi_804 = {dataGroup_hi_hi_804, dataGroup_hi_lo_804};
  wire [7:0]    dataGroup_4_25 = dataGroup_lo_804[263:256];
  wire [1023:0] dataGroup_lo_805 = {dataGroup_lo_hi_805, dataGroup_lo_lo_805};
  wire [1023:0] dataGroup_hi_805 = {dataGroup_hi_hi_805, dataGroup_hi_lo_805};
  wire [7:0]    dataGroup_5_25 = dataGroup_lo_805[319:312];
  wire [1023:0] dataGroup_lo_806 = {dataGroup_lo_hi_806, dataGroup_lo_lo_806};
  wire [1023:0] dataGroup_hi_806 = {dataGroup_hi_hi_806, dataGroup_hi_lo_806};
  wire [7:0]    dataGroup_6_25 = dataGroup_lo_806[375:368];
  wire [1023:0] dataGroup_lo_807 = {dataGroup_lo_hi_807, dataGroup_lo_lo_807};
  wire [1023:0] dataGroup_hi_807 = {dataGroup_hi_hi_807, dataGroup_hi_lo_807};
  wire [7:0]    dataGroup_7_25 = dataGroup_lo_807[431:424];
  wire [1023:0] dataGroup_lo_808 = {dataGroup_lo_hi_808, dataGroup_lo_lo_808};
  wire [1023:0] dataGroup_hi_808 = {dataGroup_hi_hi_808, dataGroup_hi_lo_808};
  wire [7:0]    dataGroup_8_25 = dataGroup_lo_808[487:480];
  wire [1023:0] dataGroup_lo_809 = {dataGroup_lo_hi_809, dataGroup_lo_lo_809};
  wire [1023:0] dataGroup_hi_809 = {dataGroup_hi_hi_809, dataGroup_hi_lo_809};
  wire [7:0]    dataGroup_9_25 = dataGroup_lo_809[543:536];
  wire [1023:0] dataGroup_lo_810 = {dataGroup_lo_hi_810, dataGroup_lo_lo_810};
  wire [1023:0] dataGroup_hi_810 = {dataGroup_hi_hi_810, dataGroup_hi_lo_810};
  wire [7:0]    dataGroup_10_25 = dataGroup_lo_810[599:592];
  wire [1023:0] dataGroup_lo_811 = {dataGroup_lo_hi_811, dataGroup_lo_lo_811};
  wire [1023:0] dataGroup_hi_811 = {dataGroup_hi_hi_811, dataGroup_hi_lo_811};
  wire [7:0]    dataGroup_11_25 = dataGroup_lo_811[655:648];
  wire [1023:0] dataGroup_lo_812 = {dataGroup_lo_hi_812, dataGroup_lo_lo_812};
  wire [1023:0] dataGroup_hi_812 = {dataGroup_hi_hi_812, dataGroup_hi_lo_812};
  wire [7:0]    dataGroup_12_25 = dataGroup_lo_812[711:704];
  wire [1023:0] dataGroup_lo_813 = {dataGroup_lo_hi_813, dataGroup_lo_lo_813};
  wire [1023:0] dataGroup_hi_813 = {dataGroup_hi_hi_813, dataGroup_hi_lo_813};
  wire [7:0]    dataGroup_13_25 = dataGroup_lo_813[767:760];
  wire [1023:0] dataGroup_lo_814 = {dataGroup_lo_hi_814, dataGroup_lo_lo_814};
  wire [1023:0] dataGroup_hi_814 = {dataGroup_hi_hi_814, dataGroup_hi_lo_814};
  wire [7:0]    dataGroup_14_25 = dataGroup_lo_814[823:816];
  wire [1023:0] dataGroup_lo_815 = {dataGroup_lo_hi_815, dataGroup_lo_lo_815};
  wire [1023:0] dataGroup_hi_815 = {dataGroup_hi_hi_815, dataGroup_hi_lo_815};
  wire [7:0]    dataGroup_15_25 = dataGroup_lo_815[879:872];
  wire [1023:0] dataGroup_lo_816 = {dataGroup_lo_hi_816, dataGroup_lo_lo_816};
  wire [1023:0] dataGroup_hi_816 = {dataGroup_hi_hi_816, dataGroup_hi_lo_816};
  wire [7:0]    dataGroup_16_25 = dataGroup_lo_816[935:928];
  wire [1023:0] dataGroup_lo_817 = {dataGroup_lo_hi_817, dataGroup_lo_lo_817};
  wire [1023:0] dataGroup_hi_817 = {dataGroup_hi_hi_817, dataGroup_hi_lo_817};
  wire [7:0]    dataGroup_17_25 = dataGroup_lo_817[991:984];
  wire [1023:0] dataGroup_lo_818 = {dataGroup_lo_hi_818, dataGroup_lo_lo_818};
  wire [1023:0] dataGroup_hi_818 = {dataGroup_hi_hi_818, dataGroup_hi_lo_818};
  wire [7:0]    dataGroup_18_25 = dataGroup_hi_818[23:16];
  wire [1023:0] dataGroup_lo_819 = {dataGroup_lo_hi_819, dataGroup_lo_lo_819};
  wire [1023:0] dataGroup_hi_819 = {dataGroup_hi_hi_819, dataGroup_hi_lo_819};
  wire [7:0]    dataGroup_19_25 = dataGroup_hi_819[79:72];
  wire [1023:0] dataGroup_lo_820 = {dataGroup_lo_hi_820, dataGroup_lo_lo_820};
  wire [1023:0] dataGroup_hi_820 = {dataGroup_hi_hi_820, dataGroup_hi_lo_820};
  wire [7:0]    dataGroup_20_25 = dataGroup_hi_820[135:128];
  wire [1023:0] dataGroup_lo_821 = {dataGroup_lo_hi_821, dataGroup_lo_lo_821};
  wire [1023:0] dataGroup_hi_821 = {dataGroup_hi_hi_821, dataGroup_hi_lo_821};
  wire [7:0]    dataGroup_21_25 = dataGroup_hi_821[191:184];
  wire [1023:0] dataGroup_lo_822 = {dataGroup_lo_hi_822, dataGroup_lo_lo_822};
  wire [1023:0] dataGroup_hi_822 = {dataGroup_hi_hi_822, dataGroup_hi_lo_822};
  wire [7:0]    dataGroup_22_25 = dataGroup_hi_822[247:240];
  wire [1023:0] dataGroup_lo_823 = {dataGroup_lo_hi_823, dataGroup_lo_lo_823};
  wire [1023:0] dataGroup_hi_823 = {dataGroup_hi_hi_823, dataGroup_hi_lo_823};
  wire [7:0]    dataGroup_23_25 = dataGroup_hi_823[303:296];
  wire [1023:0] dataGroup_lo_824 = {dataGroup_lo_hi_824, dataGroup_lo_lo_824};
  wire [1023:0] dataGroup_hi_824 = {dataGroup_hi_hi_824, dataGroup_hi_lo_824};
  wire [7:0]    dataGroup_24_25 = dataGroup_hi_824[359:352];
  wire [1023:0] dataGroup_lo_825 = {dataGroup_lo_hi_825, dataGroup_lo_lo_825};
  wire [1023:0] dataGroup_hi_825 = {dataGroup_hi_hi_825, dataGroup_hi_lo_825};
  wire [7:0]    dataGroup_25_25 = dataGroup_hi_825[415:408];
  wire [1023:0] dataGroup_lo_826 = {dataGroup_lo_hi_826, dataGroup_lo_lo_826};
  wire [1023:0] dataGroup_hi_826 = {dataGroup_hi_hi_826, dataGroup_hi_lo_826};
  wire [7:0]    dataGroup_26_25 = dataGroup_hi_826[471:464];
  wire [1023:0] dataGroup_lo_827 = {dataGroup_lo_hi_827, dataGroup_lo_lo_827};
  wire [1023:0] dataGroup_hi_827 = {dataGroup_hi_hi_827, dataGroup_hi_lo_827};
  wire [7:0]    dataGroup_27_25 = dataGroup_hi_827[527:520];
  wire [1023:0] dataGroup_lo_828 = {dataGroup_lo_hi_828, dataGroup_lo_lo_828};
  wire [1023:0] dataGroup_hi_828 = {dataGroup_hi_hi_828, dataGroup_hi_lo_828};
  wire [7:0]    dataGroup_28_25 = dataGroup_hi_828[583:576];
  wire [1023:0] dataGroup_lo_829 = {dataGroup_lo_hi_829, dataGroup_lo_lo_829};
  wire [1023:0] dataGroup_hi_829 = {dataGroup_hi_hi_829, dataGroup_hi_lo_829};
  wire [7:0]    dataGroup_29_25 = dataGroup_hi_829[639:632];
  wire [1023:0] dataGroup_lo_830 = {dataGroup_lo_hi_830, dataGroup_lo_lo_830};
  wire [1023:0] dataGroup_hi_830 = {dataGroup_hi_hi_830, dataGroup_hi_lo_830};
  wire [7:0]    dataGroup_30_25 = dataGroup_hi_830[695:688];
  wire [1023:0] dataGroup_lo_831 = {dataGroup_lo_hi_831, dataGroup_lo_lo_831};
  wire [1023:0] dataGroup_hi_831 = {dataGroup_hi_hi_831, dataGroup_hi_lo_831};
  wire [7:0]    dataGroup_31_25 = dataGroup_hi_831[751:744];
  wire [15:0]   res_lo_lo_lo_lo_25 = {dataGroup_1_25, dataGroup_0_25};
  wire [15:0]   res_lo_lo_lo_hi_25 = {dataGroup_3_25, dataGroup_2_25};
  wire [31:0]   res_lo_lo_lo_25 = {res_lo_lo_lo_hi_25, res_lo_lo_lo_lo_25};
  wire [15:0]   res_lo_lo_hi_lo_25 = {dataGroup_5_25, dataGroup_4_25};
  wire [15:0]   res_lo_lo_hi_hi_25 = {dataGroup_7_25, dataGroup_6_25};
  wire [31:0]   res_lo_lo_hi_25 = {res_lo_lo_hi_hi_25, res_lo_lo_hi_lo_25};
  wire [63:0]   res_lo_lo_25 = {res_lo_lo_hi_25, res_lo_lo_lo_25};
  wire [15:0]   res_lo_hi_lo_lo_25 = {dataGroup_9_25, dataGroup_8_25};
  wire [15:0]   res_lo_hi_lo_hi_25 = {dataGroup_11_25, dataGroup_10_25};
  wire [31:0]   res_lo_hi_lo_25 = {res_lo_hi_lo_hi_25, res_lo_hi_lo_lo_25};
  wire [15:0]   res_lo_hi_hi_lo_25 = {dataGroup_13_25, dataGroup_12_25};
  wire [15:0]   res_lo_hi_hi_hi_25 = {dataGroup_15_25, dataGroup_14_25};
  wire [31:0]   res_lo_hi_hi_25 = {res_lo_hi_hi_hi_25, res_lo_hi_hi_lo_25};
  wire [63:0]   res_lo_hi_25 = {res_lo_hi_hi_25, res_lo_hi_lo_25};
  wire [127:0]  res_lo_25 = {res_lo_hi_25, res_lo_lo_25};
  wire [15:0]   res_hi_lo_lo_lo_25 = {dataGroup_17_25, dataGroup_16_25};
  wire [15:0]   res_hi_lo_lo_hi_25 = {dataGroup_19_25, dataGroup_18_25};
  wire [31:0]   res_hi_lo_lo_25 = {res_hi_lo_lo_hi_25, res_hi_lo_lo_lo_25};
  wire [15:0]   res_hi_lo_hi_lo_25 = {dataGroup_21_25, dataGroup_20_25};
  wire [15:0]   res_hi_lo_hi_hi_25 = {dataGroup_23_25, dataGroup_22_25};
  wire [31:0]   res_hi_lo_hi_25 = {res_hi_lo_hi_hi_25, res_hi_lo_hi_lo_25};
  wire [63:0]   res_hi_lo_25 = {res_hi_lo_hi_25, res_hi_lo_lo_25};
  wire [15:0]   res_hi_hi_lo_lo_25 = {dataGroup_25_25, dataGroup_24_25};
  wire [15:0]   res_hi_hi_lo_hi_25 = {dataGroup_27_25, dataGroup_26_25};
  wire [31:0]   res_hi_hi_lo_25 = {res_hi_hi_lo_hi_25, res_hi_hi_lo_lo_25};
  wire [15:0]   res_hi_hi_hi_lo_25 = {dataGroup_29_25, dataGroup_28_25};
  wire [15:0]   res_hi_hi_hi_hi_25 = {dataGroup_31_25, dataGroup_30_25};
  wire [31:0]   res_hi_hi_hi_25 = {res_hi_hi_hi_hi_25, res_hi_hi_hi_lo_25};
  wire [63:0]   res_hi_hi_25 = {res_hi_hi_hi_25, res_hi_hi_lo_25};
  wire [127:0]  res_hi_25 = {res_hi_hi_25, res_hi_lo_25};
  wire [255:0]  res_52 = {res_hi_25, res_lo_25};
  wire [1023:0] dataGroup_lo_832 = {dataGroup_lo_hi_832, dataGroup_lo_lo_832};
  wire [1023:0] dataGroup_hi_832 = {dataGroup_hi_hi_832, dataGroup_hi_lo_832};
  wire [7:0]    dataGroup_0_26 = dataGroup_lo_832[47:40];
  wire [1023:0] dataGroup_lo_833 = {dataGroup_lo_hi_833, dataGroup_lo_lo_833};
  wire [1023:0] dataGroup_hi_833 = {dataGroup_hi_hi_833, dataGroup_hi_lo_833};
  wire [7:0]    dataGroup_1_26 = dataGroup_lo_833[103:96];
  wire [1023:0] dataGroup_lo_834 = {dataGroup_lo_hi_834, dataGroup_lo_lo_834};
  wire [1023:0] dataGroup_hi_834 = {dataGroup_hi_hi_834, dataGroup_hi_lo_834};
  wire [7:0]    dataGroup_2_26 = dataGroup_lo_834[159:152];
  wire [1023:0] dataGroup_lo_835 = {dataGroup_lo_hi_835, dataGroup_lo_lo_835};
  wire [1023:0] dataGroup_hi_835 = {dataGroup_hi_hi_835, dataGroup_hi_lo_835};
  wire [7:0]    dataGroup_3_26 = dataGroup_lo_835[215:208];
  wire [1023:0] dataGroup_lo_836 = {dataGroup_lo_hi_836, dataGroup_lo_lo_836};
  wire [1023:0] dataGroup_hi_836 = {dataGroup_hi_hi_836, dataGroup_hi_lo_836};
  wire [7:0]    dataGroup_4_26 = dataGroup_lo_836[271:264];
  wire [1023:0] dataGroup_lo_837 = {dataGroup_lo_hi_837, dataGroup_lo_lo_837};
  wire [1023:0] dataGroup_hi_837 = {dataGroup_hi_hi_837, dataGroup_hi_lo_837};
  wire [7:0]    dataGroup_5_26 = dataGroup_lo_837[327:320];
  wire [1023:0] dataGroup_lo_838 = {dataGroup_lo_hi_838, dataGroup_lo_lo_838};
  wire [1023:0] dataGroup_hi_838 = {dataGroup_hi_hi_838, dataGroup_hi_lo_838};
  wire [7:0]    dataGroup_6_26 = dataGroup_lo_838[383:376];
  wire [1023:0] dataGroup_lo_839 = {dataGroup_lo_hi_839, dataGroup_lo_lo_839};
  wire [1023:0] dataGroup_hi_839 = {dataGroup_hi_hi_839, dataGroup_hi_lo_839};
  wire [7:0]    dataGroup_7_26 = dataGroup_lo_839[439:432];
  wire [1023:0] dataGroup_lo_840 = {dataGroup_lo_hi_840, dataGroup_lo_lo_840};
  wire [1023:0] dataGroup_hi_840 = {dataGroup_hi_hi_840, dataGroup_hi_lo_840};
  wire [7:0]    dataGroup_8_26 = dataGroup_lo_840[495:488];
  wire [1023:0] dataGroup_lo_841 = {dataGroup_lo_hi_841, dataGroup_lo_lo_841};
  wire [1023:0] dataGroup_hi_841 = {dataGroup_hi_hi_841, dataGroup_hi_lo_841};
  wire [7:0]    dataGroup_9_26 = dataGroup_lo_841[551:544];
  wire [1023:0] dataGroup_lo_842 = {dataGroup_lo_hi_842, dataGroup_lo_lo_842};
  wire [1023:0] dataGroup_hi_842 = {dataGroup_hi_hi_842, dataGroup_hi_lo_842};
  wire [7:0]    dataGroup_10_26 = dataGroup_lo_842[607:600];
  wire [1023:0] dataGroup_lo_843 = {dataGroup_lo_hi_843, dataGroup_lo_lo_843};
  wire [1023:0] dataGroup_hi_843 = {dataGroup_hi_hi_843, dataGroup_hi_lo_843};
  wire [7:0]    dataGroup_11_26 = dataGroup_lo_843[663:656];
  wire [1023:0] dataGroup_lo_844 = {dataGroup_lo_hi_844, dataGroup_lo_lo_844};
  wire [1023:0] dataGroup_hi_844 = {dataGroup_hi_hi_844, dataGroup_hi_lo_844};
  wire [7:0]    dataGroup_12_26 = dataGroup_lo_844[719:712];
  wire [1023:0] dataGroup_lo_845 = {dataGroup_lo_hi_845, dataGroup_lo_lo_845};
  wire [1023:0] dataGroup_hi_845 = {dataGroup_hi_hi_845, dataGroup_hi_lo_845};
  wire [7:0]    dataGroup_13_26 = dataGroup_lo_845[775:768];
  wire [1023:0] dataGroup_lo_846 = {dataGroup_lo_hi_846, dataGroup_lo_lo_846};
  wire [1023:0] dataGroup_hi_846 = {dataGroup_hi_hi_846, dataGroup_hi_lo_846};
  wire [7:0]    dataGroup_14_26 = dataGroup_lo_846[831:824];
  wire [1023:0] dataGroup_lo_847 = {dataGroup_lo_hi_847, dataGroup_lo_lo_847};
  wire [1023:0] dataGroup_hi_847 = {dataGroup_hi_hi_847, dataGroup_hi_lo_847};
  wire [7:0]    dataGroup_15_26 = dataGroup_lo_847[887:880];
  wire [1023:0] dataGroup_lo_848 = {dataGroup_lo_hi_848, dataGroup_lo_lo_848};
  wire [1023:0] dataGroup_hi_848 = {dataGroup_hi_hi_848, dataGroup_hi_lo_848};
  wire [7:0]    dataGroup_16_26 = dataGroup_lo_848[943:936];
  wire [1023:0] dataGroup_lo_849 = {dataGroup_lo_hi_849, dataGroup_lo_lo_849};
  wire [1023:0] dataGroup_hi_849 = {dataGroup_hi_hi_849, dataGroup_hi_lo_849};
  wire [7:0]    dataGroup_17_26 = dataGroup_lo_849[999:992];
  wire [1023:0] dataGroup_lo_850 = {dataGroup_lo_hi_850, dataGroup_lo_lo_850};
  wire [1023:0] dataGroup_hi_850 = {dataGroup_hi_hi_850, dataGroup_hi_lo_850};
  wire [7:0]    dataGroup_18_26 = dataGroup_hi_850[31:24];
  wire [1023:0] dataGroup_lo_851 = {dataGroup_lo_hi_851, dataGroup_lo_lo_851};
  wire [1023:0] dataGroup_hi_851 = {dataGroup_hi_hi_851, dataGroup_hi_lo_851};
  wire [7:0]    dataGroup_19_26 = dataGroup_hi_851[87:80];
  wire [1023:0] dataGroup_lo_852 = {dataGroup_lo_hi_852, dataGroup_lo_lo_852};
  wire [1023:0] dataGroup_hi_852 = {dataGroup_hi_hi_852, dataGroup_hi_lo_852};
  wire [7:0]    dataGroup_20_26 = dataGroup_hi_852[143:136];
  wire [1023:0] dataGroup_lo_853 = {dataGroup_lo_hi_853, dataGroup_lo_lo_853};
  wire [1023:0] dataGroup_hi_853 = {dataGroup_hi_hi_853, dataGroup_hi_lo_853};
  wire [7:0]    dataGroup_21_26 = dataGroup_hi_853[199:192];
  wire [1023:0] dataGroup_lo_854 = {dataGroup_lo_hi_854, dataGroup_lo_lo_854};
  wire [1023:0] dataGroup_hi_854 = {dataGroup_hi_hi_854, dataGroup_hi_lo_854};
  wire [7:0]    dataGroup_22_26 = dataGroup_hi_854[255:248];
  wire [1023:0] dataGroup_lo_855 = {dataGroup_lo_hi_855, dataGroup_lo_lo_855};
  wire [1023:0] dataGroup_hi_855 = {dataGroup_hi_hi_855, dataGroup_hi_lo_855};
  wire [7:0]    dataGroup_23_26 = dataGroup_hi_855[311:304];
  wire [1023:0] dataGroup_lo_856 = {dataGroup_lo_hi_856, dataGroup_lo_lo_856};
  wire [1023:0] dataGroup_hi_856 = {dataGroup_hi_hi_856, dataGroup_hi_lo_856};
  wire [7:0]    dataGroup_24_26 = dataGroup_hi_856[367:360];
  wire [1023:0] dataGroup_lo_857 = {dataGroup_lo_hi_857, dataGroup_lo_lo_857};
  wire [1023:0] dataGroup_hi_857 = {dataGroup_hi_hi_857, dataGroup_hi_lo_857};
  wire [7:0]    dataGroup_25_26 = dataGroup_hi_857[423:416];
  wire [1023:0] dataGroup_lo_858 = {dataGroup_lo_hi_858, dataGroup_lo_lo_858};
  wire [1023:0] dataGroup_hi_858 = {dataGroup_hi_hi_858, dataGroup_hi_lo_858};
  wire [7:0]    dataGroup_26_26 = dataGroup_hi_858[479:472];
  wire [1023:0] dataGroup_lo_859 = {dataGroup_lo_hi_859, dataGroup_lo_lo_859};
  wire [1023:0] dataGroup_hi_859 = {dataGroup_hi_hi_859, dataGroup_hi_lo_859};
  wire [7:0]    dataGroup_27_26 = dataGroup_hi_859[535:528];
  wire [1023:0] dataGroup_lo_860 = {dataGroup_lo_hi_860, dataGroup_lo_lo_860};
  wire [1023:0] dataGroup_hi_860 = {dataGroup_hi_hi_860, dataGroup_hi_lo_860};
  wire [7:0]    dataGroup_28_26 = dataGroup_hi_860[591:584];
  wire [1023:0] dataGroup_lo_861 = {dataGroup_lo_hi_861, dataGroup_lo_lo_861};
  wire [1023:0] dataGroup_hi_861 = {dataGroup_hi_hi_861, dataGroup_hi_lo_861};
  wire [7:0]    dataGroup_29_26 = dataGroup_hi_861[647:640];
  wire [1023:0] dataGroup_lo_862 = {dataGroup_lo_hi_862, dataGroup_lo_lo_862};
  wire [1023:0] dataGroup_hi_862 = {dataGroup_hi_hi_862, dataGroup_hi_lo_862};
  wire [7:0]    dataGroup_30_26 = dataGroup_hi_862[703:696];
  wire [1023:0] dataGroup_lo_863 = {dataGroup_lo_hi_863, dataGroup_lo_lo_863};
  wire [1023:0] dataGroup_hi_863 = {dataGroup_hi_hi_863, dataGroup_hi_lo_863};
  wire [7:0]    dataGroup_31_26 = dataGroup_hi_863[759:752];
  wire [15:0]   res_lo_lo_lo_lo_26 = {dataGroup_1_26, dataGroup_0_26};
  wire [15:0]   res_lo_lo_lo_hi_26 = {dataGroup_3_26, dataGroup_2_26};
  wire [31:0]   res_lo_lo_lo_26 = {res_lo_lo_lo_hi_26, res_lo_lo_lo_lo_26};
  wire [15:0]   res_lo_lo_hi_lo_26 = {dataGroup_5_26, dataGroup_4_26};
  wire [15:0]   res_lo_lo_hi_hi_26 = {dataGroup_7_26, dataGroup_6_26};
  wire [31:0]   res_lo_lo_hi_26 = {res_lo_lo_hi_hi_26, res_lo_lo_hi_lo_26};
  wire [63:0]   res_lo_lo_26 = {res_lo_lo_hi_26, res_lo_lo_lo_26};
  wire [15:0]   res_lo_hi_lo_lo_26 = {dataGroup_9_26, dataGroup_8_26};
  wire [15:0]   res_lo_hi_lo_hi_26 = {dataGroup_11_26, dataGroup_10_26};
  wire [31:0]   res_lo_hi_lo_26 = {res_lo_hi_lo_hi_26, res_lo_hi_lo_lo_26};
  wire [15:0]   res_lo_hi_hi_lo_26 = {dataGroup_13_26, dataGroup_12_26};
  wire [15:0]   res_lo_hi_hi_hi_26 = {dataGroup_15_26, dataGroup_14_26};
  wire [31:0]   res_lo_hi_hi_26 = {res_lo_hi_hi_hi_26, res_lo_hi_hi_lo_26};
  wire [63:0]   res_lo_hi_26 = {res_lo_hi_hi_26, res_lo_hi_lo_26};
  wire [127:0]  res_lo_26 = {res_lo_hi_26, res_lo_lo_26};
  wire [15:0]   res_hi_lo_lo_lo_26 = {dataGroup_17_26, dataGroup_16_26};
  wire [15:0]   res_hi_lo_lo_hi_26 = {dataGroup_19_26, dataGroup_18_26};
  wire [31:0]   res_hi_lo_lo_26 = {res_hi_lo_lo_hi_26, res_hi_lo_lo_lo_26};
  wire [15:0]   res_hi_lo_hi_lo_26 = {dataGroup_21_26, dataGroup_20_26};
  wire [15:0]   res_hi_lo_hi_hi_26 = {dataGroup_23_26, dataGroup_22_26};
  wire [31:0]   res_hi_lo_hi_26 = {res_hi_lo_hi_hi_26, res_hi_lo_hi_lo_26};
  wire [63:0]   res_hi_lo_26 = {res_hi_lo_hi_26, res_hi_lo_lo_26};
  wire [15:0]   res_hi_hi_lo_lo_26 = {dataGroup_25_26, dataGroup_24_26};
  wire [15:0]   res_hi_hi_lo_hi_26 = {dataGroup_27_26, dataGroup_26_26};
  wire [31:0]   res_hi_hi_lo_26 = {res_hi_hi_lo_hi_26, res_hi_hi_lo_lo_26};
  wire [15:0]   res_hi_hi_hi_lo_26 = {dataGroup_29_26, dataGroup_28_26};
  wire [15:0]   res_hi_hi_hi_hi_26 = {dataGroup_31_26, dataGroup_30_26};
  wire [31:0]   res_hi_hi_hi_26 = {res_hi_hi_hi_hi_26, res_hi_hi_hi_lo_26};
  wire [63:0]   res_hi_hi_26 = {res_hi_hi_hi_26, res_hi_hi_lo_26};
  wire [127:0]  res_hi_26 = {res_hi_hi_26, res_hi_lo_26};
  wire [255:0]  res_53 = {res_hi_26, res_lo_26};
  wire [1023:0] dataGroup_lo_864 = {dataGroup_lo_hi_864, dataGroup_lo_lo_864};
  wire [1023:0] dataGroup_hi_864 = {dataGroup_hi_hi_864, dataGroup_hi_lo_864};
  wire [7:0]    dataGroup_0_27 = dataGroup_lo_864[55:48];
  wire [1023:0] dataGroup_lo_865 = {dataGroup_lo_hi_865, dataGroup_lo_lo_865};
  wire [1023:0] dataGroup_hi_865 = {dataGroup_hi_hi_865, dataGroup_hi_lo_865};
  wire [7:0]    dataGroup_1_27 = dataGroup_lo_865[111:104];
  wire [1023:0] dataGroup_lo_866 = {dataGroup_lo_hi_866, dataGroup_lo_lo_866};
  wire [1023:0] dataGroup_hi_866 = {dataGroup_hi_hi_866, dataGroup_hi_lo_866};
  wire [7:0]    dataGroup_2_27 = dataGroup_lo_866[167:160];
  wire [1023:0] dataGroup_lo_867 = {dataGroup_lo_hi_867, dataGroup_lo_lo_867};
  wire [1023:0] dataGroup_hi_867 = {dataGroup_hi_hi_867, dataGroup_hi_lo_867};
  wire [7:0]    dataGroup_3_27 = dataGroup_lo_867[223:216];
  wire [1023:0] dataGroup_lo_868 = {dataGroup_lo_hi_868, dataGroup_lo_lo_868};
  wire [1023:0] dataGroup_hi_868 = {dataGroup_hi_hi_868, dataGroup_hi_lo_868};
  wire [7:0]    dataGroup_4_27 = dataGroup_lo_868[279:272];
  wire [1023:0] dataGroup_lo_869 = {dataGroup_lo_hi_869, dataGroup_lo_lo_869};
  wire [1023:0] dataGroup_hi_869 = {dataGroup_hi_hi_869, dataGroup_hi_lo_869};
  wire [7:0]    dataGroup_5_27 = dataGroup_lo_869[335:328];
  wire [1023:0] dataGroup_lo_870 = {dataGroup_lo_hi_870, dataGroup_lo_lo_870};
  wire [1023:0] dataGroup_hi_870 = {dataGroup_hi_hi_870, dataGroup_hi_lo_870};
  wire [7:0]    dataGroup_6_27 = dataGroup_lo_870[391:384];
  wire [1023:0] dataGroup_lo_871 = {dataGroup_lo_hi_871, dataGroup_lo_lo_871};
  wire [1023:0] dataGroup_hi_871 = {dataGroup_hi_hi_871, dataGroup_hi_lo_871};
  wire [7:0]    dataGroup_7_27 = dataGroup_lo_871[447:440];
  wire [1023:0] dataGroup_lo_872 = {dataGroup_lo_hi_872, dataGroup_lo_lo_872};
  wire [1023:0] dataGroup_hi_872 = {dataGroup_hi_hi_872, dataGroup_hi_lo_872};
  wire [7:0]    dataGroup_8_27 = dataGroup_lo_872[503:496];
  wire [1023:0] dataGroup_lo_873 = {dataGroup_lo_hi_873, dataGroup_lo_lo_873};
  wire [1023:0] dataGroup_hi_873 = {dataGroup_hi_hi_873, dataGroup_hi_lo_873};
  wire [7:0]    dataGroup_9_27 = dataGroup_lo_873[559:552];
  wire [1023:0] dataGroup_lo_874 = {dataGroup_lo_hi_874, dataGroup_lo_lo_874};
  wire [1023:0] dataGroup_hi_874 = {dataGroup_hi_hi_874, dataGroup_hi_lo_874};
  wire [7:0]    dataGroup_10_27 = dataGroup_lo_874[615:608];
  wire [1023:0] dataGroup_lo_875 = {dataGroup_lo_hi_875, dataGroup_lo_lo_875};
  wire [1023:0] dataGroup_hi_875 = {dataGroup_hi_hi_875, dataGroup_hi_lo_875};
  wire [7:0]    dataGroup_11_27 = dataGroup_lo_875[671:664];
  wire [1023:0] dataGroup_lo_876 = {dataGroup_lo_hi_876, dataGroup_lo_lo_876};
  wire [1023:0] dataGroup_hi_876 = {dataGroup_hi_hi_876, dataGroup_hi_lo_876};
  wire [7:0]    dataGroup_12_27 = dataGroup_lo_876[727:720];
  wire [1023:0] dataGroup_lo_877 = {dataGroup_lo_hi_877, dataGroup_lo_lo_877};
  wire [1023:0] dataGroup_hi_877 = {dataGroup_hi_hi_877, dataGroup_hi_lo_877};
  wire [7:0]    dataGroup_13_27 = dataGroup_lo_877[783:776];
  wire [1023:0] dataGroup_lo_878 = {dataGroup_lo_hi_878, dataGroup_lo_lo_878};
  wire [1023:0] dataGroup_hi_878 = {dataGroup_hi_hi_878, dataGroup_hi_lo_878};
  wire [7:0]    dataGroup_14_27 = dataGroup_lo_878[839:832];
  wire [1023:0] dataGroup_lo_879 = {dataGroup_lo_hi_879, dataGroup_lo_lo_879};
  wire [1023:0] dataGroup_hi_879 = {dataGroup_hi_hi_879, dataGroup_hi_lo_879};
  wire [7:0]    dataGroup_15_27 = dataGroup_lo_879[895:888];
  wire [1023:0] dataGroup_lo_880 = {dataGroup_lo_hi_880, dataGroup_lo_lo_880};
  wire [1023:0] dataGroup_hi_880 = {dataGroup_hi_hi_880, dataGroup_hi_lo_880};
  wire [7:0]    dataGroup_16_27 = dataGroup_lo_880[951:944];
  wire [1023:0] dataGroup_lo_881 = {dataGroup_lo_hi_881, dataGroup_lo_lo_881};
  wire [1023:0] dataGroup_hi_881 = {dataGroup_hi_hi_881, dataGroup_hi_lo_881};
  wire [7:0]    dataGroup_17_27 = dataGroup_lo_881[1007:1000];
  wire [1023:0] dataGroup_lo_882 = {dataGroup_lo_hi_882, dataGroup_lo_lo_882};
  wire [1023:0] dataGroup_hi_882 = {dataGroup_hi_hi_882, dataGroup_hi_lo_882};
  wire [7:0]    dataGroup_18_27 = dataGroup_hi_882[39:32];
  wire [1023:0] dataGroup_lo_883 = {dataGroup_lo_hi_883, dataGroup_lo_lo_883};
  wire [1023:0] dataGroup_hi_883 = {dataGroup_hi_hi_883, dataGroup_hi_lo_883};
  wire [7:0]    dataGroup_19_27 = dataGroup_hi_883[95:88];
  wire [1023:0] dataGroup_lo_884 = {dataGroup_lo_hi_884, dataGroup_lo_lo_884};
  wire [1023:0] dataGroup_hi_884 = {dataGroup_hi_hi_884, dataGroup_hi_lo_884};
  wire [7:0]    dataGroup_20_27 = dataGroup_hi_884[151:144];
  wire [1023:0] dataGroup_lo_885 = {dataGroup_lo_hi_885, dataGroup_lo_lo_885};
  wire [1023:0] dataGroup_hi_885 = {dataGroup_hi_hi_885, dataGroup_hi_lo_885};
  wire [7:0]    dataGroup_21_27 = dataGroup_hi_885[207:200];
  wire [1023:0] dataGroup_lo_886 = {dataGroup_lo_hi_886, dataGroup_lo_lo_886};
  wire [1023:0] dataGroup_hi_886 = {dataGroup_hi_hi_886, dataGroup_hi_lo_886};
  wire [7:0]    dataGroup_22_27 = dataGroup_hi_886[263:256];
  wire [1023:0] dataGroup_lo_887 = {dataGroup_lo_hi_887, dataGroup_lo_lo_887};
  wire [1023:0] dataGroup_hi_887 = {dataGroup_hi_hi_887, dataGroup_hi_lo_887};
  wire [7:0]    dataGroup_23_27 = dataGroup_hi_887[319:312];
  wire [1023:0] dataGroup_lo_888 = {dataGroup_lo_hi_888, dataGroup_lo_lo_888};
  wire [1023:0] dataGroup_hi_888 = {dataGroup_hi_hi_888, dataGroup_hi_lo_888};
  wire [7:0]    dataGroup_24_27 = dataGroup_hi_888[375:368];
  wire [1023:0] dataGroup_lo_889 = {dataGroup_lo_hi_889, dataGroup_lo_lo_889};
  wire [1023:0] dataGroup_hi_889 = {dataGroup_hi_hi_889, dataGroup_hi_lo_889};
  wire [7:0]    dataGroup_25_27 = dataGroup_hi_889[431:424];
  wire [1023:0] dataGroup_lo_890 = {dataGroup_lo_hi_890, dataGroup_lo_lo_890};
  wire [1023:0] dataGroup_hi_890 = {dataGroup_hi_hi_890, dataGroup_hi_lo_890};
  wire [7:0]    dataGroup_26_27 = dataGroup_hi_890[487:480];
  wire [1023:0] dataGroup_lo_891 = {dataGroup_lo_hi_891, dataGroup_lo_lo_891};
  wire [1023:0] dataGroup_hi_891 = {dataGroup_hi_hi_891, dataGroup_hi_lo_891};
  wire [7:0]    dataGroup_27_27 = dataGroup_hi_891[543:536];
  wire [1023:0] dataGroup_lo_892 = {dataGroup_lo_hi_892, dataGroup_lo_lo_892};
  wire [1023:0] dataGroup_hi_892 = {dataGroup_hi_hi_892, dataGroup_hi_lo_892};
  wire [7:0]    dataGroup_28_27 = dataGroup_hi_892[599:592];
  wire [1023:0] dataGroup_lo_893 = {dataGroup_lo_hi_893, dataGroup_lo_lo_893};
  wire [1023:0] dataGroup_hi_893 = {dataGroup_hi_hi_893, dataGroup_hi_lo_893};
  wire [7:0]    dataGroup_29_27 = dataGroup_hi_893[655:648];
  wire [1023:0] dataGroup_lo_894 = {dataGroup_lo_hi_894, dataGroup_lo_lo_894};
  wire [1023:0] dataGroup_hi_894 = {dataGroup_hi_hi_894, dataGroup_hi_lo_894};
  wire [7:0]    dataGroup_30_27 = dataGroup_hi_894[711:704];
  wire [1023:0] dataGroup_lo_895 = {dataGroup_lo_hi_895, dataGroup_lo_lo_895};
  wire [1023:0] dataGroup_hi_895 = {dataGroup_hi_hi_895, dataGroup_hi_lo_895};
  wire [7:0]    dataGroup_31_27 = dataGroup_hi_895[767:760];
  wire [15:0]   res_lo_lo_lo_lo_27 = {dataGroup_1_27, dataGroup_0_27};
  wire [15:0]   res_lo_lo_lo_hi_27 = {dataGroup_3_27, dataGroup_2_27};
  wire [31:0]   res_lo_lo_lo_27 = {res_lo_lo_lo_hi_27, res_lo_lo_lo_lo_27};
  wire [15:0]   res_lo_lo_hi_lo_27 = {dataGroup_5_27, dataGroup_4_27};
  wire [15:0]   res_lo_lo_hi_hi_27 = {dataGroup_7_27, dataGroup_6_27};
  wire [31:0]   res_lo_lo_hi_27 = {res_lo_lo_hi_hi_27, res_lo_lo_hi_lo_27};
  wire [63:0]   res_lo_lo_27 = {res_lo_lo_hi_27, res_lo_lo_lo_27};
  wire [15:0]   res_lo_hi_lo_lo_27 = {dataGroup_9_27, dataGroup_8_27};
  wire [15:0]   res_lo_hi_lo_hi_27 = {dataGroup_11_27, dataGroup_10_27};
  wire [31:0]   res_lo_hi_lo_27 = {res_lo_hi_lo_hi_27, res_lo_hi_lo_lo_27};
  wire [15:0]   res_lo_hi_hi_lo_27 = {dataGroup_13_27, dataGroup_12_27};
  wire [15:0]   res_lo_hi_hi_hi_27 = {dataGroup_15_27, dataGroup_14_27};
  wire [31:0]   res_lo_hi_hi_27 = {res_lo_hi_hi_hi_27, res_lo_hi_hi_lo_27};
  wire [63:0]   res_lo_hi_27 = {res_lo_hi_hi_27, res_lo_hi_lo_27};
  wire [127:0]  res_lo_27 = {res_lo_hi_27, res_lo_lo_27};
  wire [15:0]   res_hi_lo_lo_lo_27 = {dataGroup_17_27, dataGroup_16_27};
  wire [15:0]   res_hi_lo_lo_hi_27 = {dataGroup_19_27, dataGroup_18_27};
  wire [31:0]   res_hi_lo_lo_27 = {res_hi_lo_lo_hi_27, res_hi_lo_lo_lo_27};
  wire [15:0]   res_hi_lo_hi_lo_27 = {dataGroup_21_27, dataGroup_20_27};
  wire [15:0]   res_hi_lo_hi_hi_27 = {dataGroup_23_27, dataGroup_22_27};
  wire [31:0]   res_hi_lo_hi_27 = {res_hi_lo_hi_hi_27, res_hi_lo_hi_lo_27};
  wire [63:0]   res_hi_lo_27 = {res_hi_lo_hi_27, res_hi_lo_lo_27};
  wire [15:0]   res_hi_hi_lo_lo_27 = {dataGroup_25_27, dataGroup_24_27};
  wire [15:0]   res_hi_hi_lo_hi_27 = {dataGroup_27_27, dataGroup_26_27};
  wire [31:0]   res_hi_hi_lo_27 = {res_hi_hi_lo_hi_27, res_hi_hi_lo_lo_27};
  wire [15:0]   res_hi_hi_hi_lo_27 = {dataGroup_29_27, dataGroup_28_27};
  wire [15:0]   res_hi_hi_hi_hi_27 = {dataGroup_31_27, dataGroup_30_27};
  wire [31:0]   res_hi_hi_hi_27 = {res_hi_hi_hi_hi_27, res_hi_hi_hi_lo_27};
  wire [63:0]   res_hi_hi_27 = {res_hi_hi_hi_27, res_hi_hi_lo_27};
  wire [127:0]  res_hi_27 = {res_hi_hi_27, res_hi_lo_27};
  wire [255:0]  res_54 = {res_hi_27, res_lo_27};
  wire [511:0]  lo_lo_6 = {res_49, res_48};
  wire [511:0]  lo_hi_6 = {res_51, res_50};
  wire [1023:0] lo_6 = {lo_hi_6, lo_lo_6};
  wire [511:0]  hi_lo_6 = {res_53, res_52};
  wire [511:0]  hi_hi_6 = {256'h0, res_54};
  wire [1023:0] hi_6 = {hi_hi_6, hi_lo_6};
  wire [2047:0] regroupLoadData_0_6 = {hi_6, lo_6};
  wire [1023:0] dataGroup_lo_896 = {dataGroup_lo_hi_896, dataGroup_lo_lo_896};
  wire [1023:0] dataGroup_hi_896 = {dataGroup_hi_hi_896, dataGroup_hi_lo_896};
  wire [7:0]    dataGroup_0_28 = dataGroup_lo_896[7:0];
  wire [1023:0] dataGroup_lo_897 = {dataGroup_lo_hi_897, dataGroup_lo_lo_897};
  wire [1023:0] dataGroup_hi_897 = {dataGroup_hi_hi_897, dataGroup_hi_lo_897};
  wire [7:0]    dataGroup_1_28 = dataGroup_lo_897[71:64];
  wire [1023:0] dataGroup_lo_898 = {dataGroup_lo_hi_898, dataGroup_lo_lo_898};
  wire [1023:0] dataGroup_hi_898 = {dataGroup_hi_hi_898, dataGroup_hi_lo_898};
  wire [7:0]    dataGroup_2_28 = dataGroup_lo_898[135:128];
  wire [1023:0] dataGroup_lo_899 = {dataGroup_lo_hi_899, dataGroup_lo_lo_899};
  wire [1023:0] dataGroup_hi_899 = {dataGroup_hi_hi_899, dataGroup_hi_lo_899};
  wire [7:0]    dataGroup_3_28 = dataGroup_lo_899[199:192];
  wire [1023:0] dataGroup_lo_900 = {dataGroup_lo_hi_900, dataGroup_lo_lo_900};
  wire [1023:0] dataGroup_hi_900 = {dataGroup_hi_hi_900, dataGroup_hi_lo_900};
  wire [7:0]    dataGroup_4_28 = dataGroup_lo_900[263:256];
  wire [1023:0] dataGroup_lo_901 = {dataGroup_lo_hi_901, dataGroup_lo_lo_901};
  wire [1023:0] dataGroup_hi_901 = {dataGroup_hi_hi_901, dataGroup_hi_lo_901};
  wire [7:0]    dataGroup_5_28 = dataGroup_lo_901[327:320];
  wire [1023:0] dataGroup_lo_902 = {dataGroup_lo_hi_902, dataGroup_lo_lo_902};
  wire [1023:0] dataGroup_hi_902 = {dataGroup_hi_hi_902, dataGroup_hi_lo_902};
  wire [7:0]    dataGroup_6_28 = dataGroup_lo_902[391:384];
  wire [1023:0] dataGroup_lo_903 = {dataGroup_lo_hi_903, dataGroup_lo_lo_903};
  wire [1023:0] dataGroup_hi_903 = {dataGroup_hi_hi_903, dataGroup_hi_lo_903};
  wire [7:0]    dataGroup_7_28 = dataGroup_lo_903[455:448];
  wire [1023:0] dataGroup_lo_904 = {dataGroup_lo_hi_904, dataGroup_lo_lo_904};
  wire [1023:0] dataGroup_hi_904 = {dataGroup_hi_hi_904, dataGroup_hi_lo_904};
  wire [7:0]    dataGroup_8_28 = dataGroup_lo_904[519:512];
  wire [1023:0] dataGroup_lo_905 = {dataGroup_lo_hi_905, dataGroup_lo_lo_905};
  wire [1023:0] dataGroup_hi_905 = {dataGroup_hi_hi_905, dataGroup_hi_lo_905};
  wire [7:0]    dataGroup_9_28 = dataGroup_lo_905[583:576];
  wire [1023:0] dataGroup_lo_906 = {dataGroup_lo_hi_906, dataGroup_lo_lo_906};
  wire [1023:0] dataGroup_hi_906 = {dataGroup_hi_hi_906, dataGroup_hi_lo_906};
  wire [7:0]    dataGroup_10_28 = dataGroup_lo_906[647:640];
  wire [1023:0] dataGroup_lo_907 = {dataGroup_lo_hi_907, dataGroup_lo_lo_907};
  wire [1023:0] dataGroup_hi_907 = {dataGroup_hi_hi_907, dataGroup_hi_lo_907};
  wire [7:0]    dataGroup_11_28 = dataGroup_lo_907[711:704];
  wire [1023:0] dataGroup_lo_908 = {dataGroup_lo_hi_908, dataGroup_lo_lo_908};
  wire [1023:0] dataGroup_hi_908 = {dataGroup_hi_hi_908, dataGroup_hi_lo_908};
  wire [7:0]    dataGroup_12_28 = dataGroup_lo_908[775:768];
  wire [1023:0] dataGroup_lo_909 = {dataGroup_lo_hi_909, dataGroup_lo_lo_909};
  wire [1023:0] dataGroup_hi_909 = {dataGroup_hi_hi_909, dataGroup_hi_lo_909};
  wire [7:0]    dataGroup_13_28 = dataGroup_lo_909[839:832];
  wire [1023:0] dataGroup_lo_910 = {dataGroup_lo_hi_910, dataGroup_lo_lo_910};
  wire [1023:0] dataGroup_hi_910 = {dataGroup_hi_hi_910, dataGroup_hi_lo_910};
  wire [7:0]    dataGroup_14_28 = dataGroup_lo_910[903:896];
  wire [1023:0] dataGroup_lo_911 = {dataGroup_lo_hi_911, dataGroup_lo_lo_911};
  wire [1023:0] dataGroup_hi_911 = {dataGroup_hi_hi_911, dataGroup_hi_lo_911};
  wire [7:0]    dataGroup_15_28 = dataGroup_lo_911[967:960];
  wire [1023:0] dataGroup_lo_912 = {dataGroup_lo_hi_912, dataGroup_lo_lo_912};
  wire [1023:0] dataGroup_hi_912 = {dataGroup_hi_hi_912, dataGroup_hi_lo_912};
  wire [7:0]    dataGroup_16_28 = dataGroup_hi_912[7:0];
  wire [1023:0] dataGroup_lo_913 = {dataGroup_lo_hi_913, dataGroup_lo_lo_913};
  wire [1023:0] dataGroup_hi_913 = {dataGroup_hi_hi_913, dataGroup_hi_lo_913};
  wire [7:0]    dataGroup_17_28 = dataGroup_hi_913[71:64];
  wire [1023:0] dataGroup_lo_914 = {dataGroup_lo_hi_914, dataGroup_lo_lo_914};
  wire [1023:0] dataGroup_hi_914 = {dataGroup_hi_hi_914, dataGroup_hi_lo_914};
  wire [7:0]    dataGroup_18_28 = dataGroup_hi_914[135:128];
  wire [1023:0] dataGroup_lo_915 = {dataGroup_lo_hi_915, dataGroup_lo_lo_915};
  wire [1023:0] dataGroup_hi_915 = {dataGroup_hi_hi_915, dataGroup_hi_lo_915};
  wire [7:0]    dataGroup_19_28 = dataGroup_hi_915[199:192];
  wire [1023:0] dataGroup_lo_916 = {dataGroup_lo_hi_916, dataGroup_lo_lo_916};
  wire [1023:0] dataGroup_hi_916 = {dataGroup_hi_hi_916, dataGroup_hi_lo_916};
  wire [7:0]    dataGroup_20_28 = dataGroup_hi_916[263:256];
  wire [1023:0] dataGroup_lo_917 = {dataGroup_lo_hi_917, dataGroup_lo_lo_917};
  wire [1023:0] dataGroup_hi_917 = {dataGroup_hi_hi_917, dataGroup_hi_lo_917};
  wire [7:0]    dataGroup_21_28 = dataGroup_hi_917[327:320];
  wire [1023:0] dataGroup_lo_918 = {dataGroup_lo_hi_918, dataGroup_lo_lo_918};
  wire [1023:0] dataGroup_hi_918 = {dataGroup_hi_hi_918, dataGroup_hi_lo_918};
  wire [7:0]    dataGroup_22_28 = dataGroup_hi_918[391:384];
  wire [1023:0] dataGroup_lo_919 = {dataGroup_lo_hi_919, dataGroup_lo_lo_919};
  wire [1023:0] dataGroup_hi_919 = {dataGroup_hi_hi_919, dataGroup_hi_lo_919};
  wire [7:0]    dataGroup_23_28 = dataGroup_hi_919[455:448];
  wire [1023:0] dataGroup_lo_920 = {dataGroup_lo_hi_920, dataGroup_lo_lo_920};
  wire [1023:0] dataGroup_hi_920 = {dataGroup_hi_hi_920, dataGroup_hi_lo_920};
  wire [7:0]    dataGroup_24_28 = dataGroup_hi_920[519:512];
  wire [1023:0] dataGroup_lo_921 = {dataGroup_lo_hi_921, dataGroup_lo_lo_921};
  wire [1023:0] dataGroup_hi_921 = {dataGroup_hi_hi_921, dataGroup_hi_lo_921};
  wire [7:0]    dataGroup_25_28 = dataGroup_hi_921[583:576];
  wire [1023:0] dataGroup_lo_922 = {dataGroup_lo_hi_922, dataGroup_lo_lo_922};
  wire [1023:0] dataGroup_hi_922 = {dataGroup_hi_hi_922, dataGroup_hi_lo_922};
  wire [7:0]    dataGroup_26_28 = dataGroup_hi_922[647:640];
  wire [1023:0] dataGroup_lo_923 = {dataGroup_lo_hi_923, dataGroup_lo_lo_923};
  wire [1023:0] dataGroup_hi_923 = {dataGroup_hi_hi_923, dataGroup_hi_lo_923};
  wire [7:0]    dataGroup_27_28 = dataGroup_hi_923[711:704];
  wire [1023:0] dataGroup_lo_924 = {dataGroup_lo_hi_924, dataGroup_lo_lo_924};
  wire [1023:0] dataGroup_hi_924 = {dataGroup_hi_hi_924, dataGroup_hi_lo_924};
  wire [7:0]    dataGroup_28_28 = dataGroup_hi_924[775:768];
  wire [1023:0] dataGroup_lo_925 = {dataGroup_lo_hi_925, dataGroup_lo_lo_925};
  wire [1023:0] dataGroup_hi_925 = {dataGroup_hi_hi_925, dataGroup_hi_lo_925};
  wire [7:0]    dataGroup_29_28 = dataGroup_hi_925[839:832];
  wire [1023:0] dataGroup_lo_926 = {dataGroup_lo_hi_926, dataGroup_lo_lo_926};
  wire [1023:0] dataGroup_hi_926 = {dataGroup_hi_hi_926, dataGroup_hi_lo_926};
  wire [7:0]    dataGroup_30_28 = dataGroup_hi_926[903:896];
  wire [1023:0] dataGroup_lo_927 = {dataGroup_lo_hi_927, dataGroup_lo_lo_927};
  wire [1023:0] dataGroup_hi_927 = {dataGroup_hi_hi_927, dataGroup_hi_lo_927};
  wire [7:0]    dataGroup_31_28 = dataGroup_hi_927[967:960];
  wire [15:0]   res_lo_lo_lo_lo_28 = {dataGroup_1_28, dataGroup_0_28};
  wire [15:0]   res_lo_lo_lo_hi_28 = {dataGroup_3_28, dataGroup_2_28};
  wire [31:0]   res_lo_lo_lo_28 = {res_lo_lo_lo_hi_28, res_lo_lo_lo_lo_28};
  wire [15:0]   res_lo_lo_hi_lo_28 = {dataGroup_5_28, dataGroup_4_28};
  wire [15:0]   res_lo_lo_hi_hi_28 = {dataGroup_7_28, dataGroup_6_28};
  wire [31:0]   res_lo_lo_hi_28 = {res_lo_lo_hi_hi_28, res_lo_lo_hi_lo_28};
  wire [63:0]   res_lo_lo_28 = {res_lo_lo_hi_28, res_lo_lo_lo_28};
  wire [15:0]   res_lo_hi_lo_lo_28 = {dataGroup_9_28, dataGroup_8_28};
  wire [15:0]   res_lo_hi_lo_hi_28 = {dataGroup_11_28, dataGroup_10_28};
  wire [31:0]   res_lo_hi_lo_28 = {res_lo_hi_lo_hi_28, res_lo_hi_lo_lo_28};
  wire [15:0]   res_lo_hi_hi_lo_28 = {dataGroup_13_28, dataGroup_12_28};
  wire [15:0]   res_lo_hi_hi_hi_28 = {dataGroup_15_28, dataGroup_14_28};
  wire [31:0]   res_lo_hi_hi_28 = {res_lo_hi_hi_hi_28, res_lo_hi_hi_lo_28};
  wire [63:0]   res_lo_hi_28 = {res_lo_hi_hi_28, res_lo_hi_lo_28};
  wire [127:0]  res_lo_28 = {res_lo_hi_28, res_lo_lo_28};
  wire [15:0]   res_hi_lo_lo_lo_28 = {dataGroup_17_28, dataGroup_16_28};
  wire [15:0]   res_hi_lo_lo_hi_28 = {dataGroup_19_28, dataGroup_18_28};
  wire [31:0]   res_hi_lo_lo_28 = {res_hi_lo_lo_hi_28, res_hi_lo_lo_lo_28};
  wire [15:0]   res_hi_lo_hi_lo_28 = {dataGroup_21_28, dataGroup_20_28};
  wire [15:0]   res_hi_lo_hi_hi_28 = {dataGroup_23_28, dataGroup_22_28};
  wire [31:0]   res_hi_lo_hi_28 = {res_hi_lo_hi_hi_28, res_hi_lo_hi_lo_28};
  wire [63:0]   res_hi_lo_28 = {res_hi_lo_hi_28, res_hi_lo_lo_28};
  wire [15:0]   res_hi_hi_lo_lo_28 = {dataGroup_25_28, dataGroup_24_28};
  wire [15:0]   res_hi_hi_lo_hi_28 = {dataGroup_27_28, dataGroup_26_28};
  wire [31:0]   res_hi_hi_lo_28 = {res_hi_hi_lo_hi_28, res_hi_hi_lo_lo_28};
  wire [15:0]   res_hi_hi_hi_lo_28 = {dataGroup_29_28, dataGroup_28_28};
  wire [15:0]   res_hi_hi_hi_hi_28 = {dataGroup_31_28, dataGroup_30_28};
  wire [31:0]   res_hi_hi_hi_28 = {res_hi_hi_hi_hi_28, res_hi_hi_hi_lo_28};
  wire [63:0]   res_hi_hi_28 = {res_hi_hi_hi_28, res_hi_hi_lo_28};
  wire [127:0]  res_hi_28 = {res_hi_hi_28, res_hi_lo_28};
  wire [255:0]  res_56 = {res_hi_28, res_lo_28};
  wire [1023:0] dataGroup_lo_928 = {dataGroup_lo_hi_928, dataGroup_lo_lo_928};
  wire [1023:0] dataGroup_hi_928 = {dataGroup_hi_hi_928, dataGroup_hi_lo_928};
  wire [7:0]    dataGroup_0_29 = dataGroup_lo_928[15:8];
  wire [1023:0] dataGroup_lo_929 = {dataGroup_lo_hi_929, dataGroup_lo_lo_929};
  wire [1023:0] dataGroup_hi_929 = {dataGroup_hi_hi_929, dataGroup_hi_lo_929};
  wire [7:0]    dataGroup_1_29 = dataGroup_lo_929[79:72];
  wire [1023:0] dataGroup_lo_930 = {dataGroup_lo_hi_930, dataGroup_lo_lo_930};
  wire [1023:0] dataGroup_hi_930 = {dataGroup_hi_hi_930, dataGroup_hi_lo_930};
  wire [7:0]    dataGroup_2_29 = dataGroup_lo_930[143:136];
  wire [1023:0] dataGroup_lo_931 = {dataGroup_lo_hi_931, dataGroup_lo_lo_931};
  wire [1023:0] dataGroup_hi_931 = {dataGroup_hi_hi_931, dataGroup_hi_lo_931};
  wire [7:0]    dataGroup_3_29 = dataGroup_lo_931[207:200];
  wire [1023:0] dataGroup_lo_932 = {dataGroup_lo_hi_932, dataGroup_lo_lo_932};
  wire [1023:0] dataGroup_hi_932 = {dataGroup_hi_hi_932, dataGroup_hi_lo_932};
  wire [7:0]    dataGroup_4_29 = dataGroup_lo_932[271:264];
  wire [1023:0] dataGroup_lo_933 = {dataGroup_lo_hi_933, dataGroup_lo_lo_933};
  wire [1023:0] dataGroup_hi_933 = {dataGroup_hi_hi_933, dataGroup_hi_lo_933};
  wire [7:0]    dataGroup_5_29 = dataGroup_lo_933[335:328];
  wire [1023:0] dataGroup_lo_934 = {dataGroup_lo_hi_934, dataGroup_lo_lo_934};
  wire [1023:0] dataGroup_hi_934 = {dataGroup_hi_hi_934, dataGroup_hi_lo_934};
  wire [7:0]    dataGroup_6_29 = dataGroup_lo_934[399:392];
  wire [1023:0] dataGroup_lo_935 = {dataGroup_lo_hi_935, dataGroup_lo_lo_935};
  wire [1023:0] dataGroup_hi_935 = {dataGroup_hi_hi_935, dataGroup_hi_lo_935};
  wire [7:0]    dataGroup_7_29 = dataGroup_lo_935[463:456];
  wire [1023:0] dataGroup_lo_936 = {dataGroup_lo_hi_936, dataGroup_lo_lo_936};
  wire [1023:0] dataGroup_hi_936 = {dataGroup_hi_hi_936, dataGroup_hi_lo_936};
  wire [7:0]    dataGroup_8_29 = dataGroup_lo_936[527:520];
  wire [1023:0] dataGroup_lo_937 = {dataGroup_lo_hi_937, dataGroup_lo_lo_937};
  wire [1023:0] dataGroup_hi_937 = {dataGroup_hi_hi_937, dataGroup_hi_lo_937};
  wire [7:0]    dataGroup_9_29 = dataGroup_lo_937[591:584];
  wire [1023:0] dataGroup_lo_938 = {dataGroup_lo_hi_938, dataGroup_lo_lo_938};
  wire [1023:0] dataGroup_hi_938 = {dataGroup_hi_hi_938, dataGroup_hi_lo_938};
  wire [7:0]    dataGroup_10_29 = dataGroup_lo_938[655:648];
  wire [1023:0] dataGroup_lo_939 = {dataGroup_lo_hi_939, dataGroup_lo_lo_939};
  wire [1023:0] dataGroup_hi_939 = {dataGroup_hi_hi_939, dataGroup_hi_lo_939};
  wire [7:0]    dataGroup_11_29 = dataGroup_lo_939[719:712];
  wire [1023:0] dataGroup_lo_940 = {dataGroup_lo_hi_940, dataGroup_lo_lo_940};
  wire [1023:0] dataGroup_hi_940 = {dataGroup_hi_hi_940, dataGroup_hi_lo_940};
  wire [7:0]    dataGroup_12_29 = dataGroup_lo_940[783:776];
  wire [1023:0] dataGroup_lo_941 = {dataGroup_lo_hi_941, dataGroup_lo_lo_941};
  wire [1023:0] dataGroup_hi_941 = {dataGroup_hi_hi_941, dataGroup_hi_lo_941};
  wire [7:0]    dataGroup_13_29 = dataGroup_lo_941[847:840];
  wire [1023:0] dataGroup_lo_942 = {dataGroup_lo_hi_942, dataGroup_lo_lo_942};
  wire [1023:0] dataGroup_hi_942 = {dataGroup_hi_hi_942, dataGroup_hi_lo_942};
  wire [7:0]    dataGroup_14_29 = dataGroup_lo_942[911:904];
  wire [1023:0] dataGroup_lo_943 = {dataGroup_lo_hi_943, dataGroup_lo_lo_943};
  wire [1023:0] dataGroup_hi_943 = {dataGroup_hi_hi_943, dataGroup_hi_lo_943};
  wire [7:0]    dataGroup_15_29 = dataGroup_lo_943[975:968];
  wire [1023:0] dataGroup_lo_944 = {dataGroup_lo_hi_944, dataGroup_lo_lo_944};
  wire [1023:0] dataGroup_hi_944 = {dataGroup_hi_hi_944, dataGroup_hi_lo_944};
  wire [7:0]    dataGroup_16_29 = dataGroup_hi_944[15:8];
  wire [1023:0] dataGroup_lo_945 = {dataGroup_lo_hi_945, dataGroup_lo_lo_945};
  wire [1023:0] dataGroup_hi_945 = {dataGroup_hi_hi_945, dataGroup_hi_lo_945};
  wire [7:0]    dataGroup_17_29 = dataGroup_hi_945[79:72];
  wire [1023:0] dataGroup_lo_946 = {dataGroup_lo_hi_946, dataGroup_lo_lo_946};
  wire [1023:0] dataGroup_hi_946 = {dataGroup_hi_hi_946, dataGroup_hi_lo_946};
  wire [7:0]    dataGroup_18_29 = dataGroup_hi_946[143:136];
  wire [1023:0] dataGroup_lo_947 = {dataGroup_lo_hi_947, dataGroup_lo_lo_947};
  wire [1023:0] dataGroup_hi_947 = {dataGroup_hi_hi_947, dataGroup_hi_lo_947};
  wire [7:0]    dataGroup_19_29 = dataGroup_hi_947[207:200];
  wire [1023:0] dataGroup_lo_948 = {dataGroup_lo_hi_948, dataGroup_lo_lo_948};
  wire [1023:0] dataGroup_hi_948 = {dataGroup_hi_hi_948, dataGroup_hi_lo_948};
  wire [7:0]    dataGroup_20_29 = dataGroup_hi_948[271:264];
  wire [1023:0] dataGroup_lo_949 = {dataGroup_lo_hi_949, dataGroup_lo_lo_949};
  wire [1023:0] dataGroup_hi_949 = {dataGroup_hi_hi_949, dataGroup_hi_lo_949};
  wire [7:0]    dataGroup_21_29 = dataGroup_hi_949[335:328];
  wire [1023:0] dataGroup_lo_950 = {dataGroup_lo_hi_950, dataGroup_lo_lo_950};
  wire [1023:0] dataGroup_hi_950 = {dataGroup_hi_hi_950, dataGroup_hi_lo_950};
  wire [7:0]    dataGroup_22_29 = dataGroup_hi_950[399:392];
  wire [1023:0] dataGroup_lo_951 = {dataGroup_lo_hi_951, dataGroup_lo_lo_951};
  wire [1023:0] dataGroup_hi_951 = {dataGroup_hi_hi_951, dataGroup_hi_lo_951};
  wire [7:0]    dataGroup_23_29 = dataGroup_hi_951[463:456];
  wire [1023:0] dataGroup_lo_952 = {dataGroup_lo_hi_952, dataGroup_lo_lo_952};
  wire [1023:0] dataGroup_hi_952 = {dataGroup_hi_hi_952, dataGroup_hi_lo_952};
  wire [7:0]    dataGroup_24_29 = dataGroup_hi_952[527:520];
  wire [1023:0] dataGroup_lo_953 = {dataGroup_lo_hi_953, dataGroup_lo_lo_953};
  wire [1023:0] dataGroup_hi_953 = {dataGroup_hi_hi_953, dataGroup_hi_lo_953};
  wire [7:0]    dataGroup_25_29 = dataGroup_hi_953[591:584];
  wire [1023:0] dataGroup_lo_954 = {dataGroup_lo_hi_954, dataGroup_lo_lo_954};
  wire [1023:0] dataGroup_hi_954 = {dataGroup_hi_hi_954, dataGroup_hi_lo_954};
  wire [7:0]    dataGroup_26_29 = dataGroup_hi_954[655:648];
  wire [1023:0] dataGroup_lo_955 = {dataGroup_lo_hi_955, dataGroup_lo_lo_955};
  wire [1023:0] dataGroup_hi_955 = {dataGroup_hi_hi_955, dataGroup_hi_lo_955};
  wire [7:0]    dataGroup_27_29 = dataGroup_hi_955[719:712];
  wire [1023:0] dataGroup_lo_956 = {dataGroup_lo_hi_956, dataGroup_lo_lo_956};
  wire [1023:0] dataGroup_hi_956 = {dataGroup_hi_hi_956, dataGroup_hi_lo_956};
  wire [7:0]    dataGroup_28_29 = dataGroup_hi_956[783:776];
  wire [1023:0] dataGroup_lo_957 = {dataGroup_lo_hi_957, dataGroup_lo_lo_957};
  wire [1023:0] dataGroup_hi_957 = {dataGroup_hi_hi_957, dataGroup_hi_lo_957};
  wire [7:0]    dataGroup_29_29 = dataGroup_hi_957[847:840];
  wire [1023:0] dataGroup_lo_958 = {dataGroup_lo_hi_958, dataGroup_lo_lo_958};
  wire [1023:0] dataGroup_hi_958 = {dataGroup_hi_hi_958, dataGroup_hi_lo_958};
  wire [7:0]    dataGroup_30_29 = dataGroup_hi_958[911:904];
  wire [1023:0] dataGroup_lo_959 = {dataGroup_lo_hi_959, dataGroup_lo_lo_959};
  wire [1023:0] dataGroup_hi_959 = {dataGroup_hi_hi_959, dataGroup_hi_lo_959};
  wire [7:0]    dataGroup_31_29 = dataGroup_hi_959[975:968];
  wire [15:0]   res_lo_lo_lo_lo_29 = {dataGroup_1_29, dataGroup_0_29};
  wire [15:0]   res_lo_lo_lo_hi_29 = {dataGroup_3_29, dataGroup_2_29};
  wire [31:0]   res_lo_lo_lo_29 = {res_lo_lo_lo_hi_29, res_lo_lo_lo_lo_29};
  wire [15:0]   res_lo_lo_hi_lo_29 = {dataGroup_5_29, dataGroup_4_29};
  wire [15:0]   res_lo_lo_hi_hi_29 = {dataGroup_7_29, dataGroup_6_29};
  wire [31:0]   res_lo_lo_hi_29 = {res_lo_lo_hi_hi_29, res_lo_lo_hi_lo_29};
  wire [63:0]   res_lo_lo_29 = {res_lo_lo_hi_29, res_lo_lo_lo_29};
  wire [15:0]   res_lo_hi_lo_lo_29 = {dataGroup_9_29, dataGroup_8_29};
  wire [15:0]   res_lo_hi_lo_hi_29 = {dataGroup_11_29, dataGroup_10_29};
  wire [31:0]   res_lo_hi_lo_29 = {res_lo_hi_lo_hi_29, res_lo_hi_lo_lo_29};
  wire [15:0]   res_lo_hi_hi_lo_29 = {dataGroup_13_29, dataGroup_12_29};
  wire [15:0]   res_lo_hi_hi_hi_29 = {dataGroup_15_29, dataGroup_14_29};
  wire [31:0]   res_lo_hi_hi_29 = {res_lo_hi_hi_hi_29, res_lo_hi_hi_lo_29};
  wire [63:0]   res_lo_hi_29 = {res_lo_hi_hi_29, res_lo_hi_lo_29};
  wire [127:0]  res_lo_29 = {res_lo_hi_29, res_lo_lo_29};
  wire [15:0]   res_hi_lo_lo_lo_29 = {dataGroup_17_29, dataGroup_16_29};
  wire [15:0]   res_hi_lo_lo_hi_29 = {dataGroup_19_29, dataGroup_18_29};
  wire [31:0]   res_hi_lo_lo_29 = {res_hi_lo_lo_hi_29, res_hi_lo_lo_lo_29};
  wire [15:0]   res_hi_lo_hi_lo_29 = {dataGroup_21_29, dataGroup_20_29};
  wire [15:0]   res_hi_lo_hi_hi_29 = {dataGroup_23_29, dataGroup_22_29};
  wire [31:0]   res_hi_lo_hi_29 = {res_hi_lo_hi_hi_29, res_hi_lo_hi_lo_29};
  wire [63:0]   res_hi_lo_29 = {res_hi_lo_hi_29, res_hi_lo_lo_29};
  wire [15:0]   res_hi_hi_lo_lo_29 = {dataGroup_25_29, dataGroup_24_29};
  wire [15:0]   res_hi_hi_lo_hi_29 = {dataGroup_27_29, dataGroup_26_29};
  wire [31:0]   res_hi_hi_lo_29 = {res_hi_hi_lo_hi_29, res_hi_hi_lo_lo_29};
  wire [15:0]   res_hi_hi_hi_lo_29 = {dataGroup_29_29, dataGroup_28_29};
  wire [15:0]   res_hi_hi_hi_hi_29 = {dataGroup_31_29, dataGroup_30_29};
  wire [31:0]   res_hi_hi_hi_29 = {res_hi_hi_hi_hi_29, res_hi_hi_hi_lo_29};
  wire [63:0]   res_hi_hi_29 = {res_hi_hi_hi_29, res_hi_hi_lo_29};
  wire [127:0]  res_hi_29 = {res_hi_hi_29, res_hi_lo_29};
  wire [255:0]  res_57 = {res_hi_29, res_lo_29};
  wire [1023:0] dataGroup_lo_960 = {dataGroup_lo_hi_960, dataGroup_lo_lo_960};
  wire [1023:0] dataGroup_hi_960 = {dataGroup_hi_hi_960, dataGroup_hi_lo_960};
  wire [7:0]    dataGroup_0_30 = dataGroup_lo_960[23:16];
  wire [1023:0] dataGroup_lo_961 = {dataGroup_lo_hi_961, dataGroup_lo_lo_961};
  wire [1023:0] dataGroup_hi_961 = {dataGroup_hi_hi_961, dataGroup_hi_lo_961};
  wire [7:0]    dataGroup_1_30 = dataGroup_lo_961[87:80];
  wire [1023:0] dataGroup_lo_962 = {dataGroup_lo_hi_962, dataGroup_lo_lo_962};
  wire [1023:0] dataGroup_hi_962 = {dataGroup_hi_hi_962, dataGroup_hi_lo_962};
  wire [7:0]    dataGroup_2_30 = dataGroup_lo_962[151:144];
  wire [1023:0] dataGroup_lo_963 = {dataGroup_lo_hi_963, dataGroup_lo_lo_963};
  wire [1023:0] dataGroup_hi_963 = {dataGroup_hi_hi_963, dataGroup_hi_lo_963};
  wire [7:0]    dataGroup_3_30 = dataGroup_lo_963[215:208];
  wire [1023:0] dataGroup_lo_964 = {dataGroup_lo_hi_964, dataGroup_lo_lo_964};
  wire [1023:0] dataGroup_hi_964 = {dataGroup_hi_hi_964, dataGroup_hi_lo_964};
  wire [7:0]    dataGroup_4_30 = dataGroup_lo_964[279:272];
  wire [1023:0] dataGroup_lo_965 = {dataGroup_lo_hi_965, dataGroup_lo_lo_965};
  wire [1023:0] dataGroup_hi_965 = {dataGroup_hi_hi_965, dataGroup_hi_lo_965};
  wire [7:0]    dataGroup_5_30 = dataGroup_lo_965[343:336];
  wire [1023:0] dataGroup_lo_966 = {dataGroup_lo_hi_966, dataGroup_lo_lo_966};
  wire [1023:0] dataGroup_hi_966 = {dataGroup_hi_hi_966, dataGroup_hi_lo_966};
  wire [7:0]    dataGroup_6_30 = dataGroup_lo_966[407:400];
  wire [1023:0] dataGroup_lo_967 = {dataGroup_lo_hi_967, dataGroup_lo_lo_967};
  wire [1023:0] dataGroup_hi_967 = {dataGroup_hi_hi_967, dataGroup_hi_lo_967};
  wire [7:0]    dataGroup_7_30 = dataGroup_lo_967[471:464];
  wire [1023:0] dataGroup_lo_968 = {dataGroup_lo_hi_968, dataGroup_lo_lo_968};
  wire [1023:0] dataGroup_hi_968 = {dataGroup_hi_hi_968, dataGroup_hi_lo_968};
  wire [7:0]    dataGroup_8_30 = dataGroup_lo_968[535:528];
  wire [1023:0] dataGroup_lo_969 = {dataGroup_lo_hi_969, dataGroup_lo_lo_969};
  wire [1023:0] dataGroup_hi_969 = {dataGroup_hi_hi_969, dataGroup_hi_lo_969};
  wire [7:0]    dataGroup_9_30 = dataGroup_lo_969[599:592];
  wire [1023:0] dataGroup_lo_970 = {dataGroup_lo_hi_970, dataGroup_lo_lo_970};
  wire [1023:0] dataGroup_hi_970 = {dataGroup_hi_hi_970, dataGroup_hi_lo_970};
  wire [7:0]    dataGroup_10_30 = dataGroup_lo_970[663:656];
  wire [1023:0] dataGroup_lo_971 = {dataGroup_lo_hi_971, dataGroup_lo_lo_971};
  wire [1023:0] dataGroup_hi_971 = {dataGroup_hi_hi_971, dataGroup_hi_lo_971};
  wire [7:0]    dataGroup_11_30 = dataGroup_lo_971[727:720];
  wire [1023:0] dataGroup_lo_972 = {dataGroup_lo_hi_972, dataGroup_lo_lo_972};
  wire [1023:0] dataGroup_hi_972 = {dataGroup_hi_hi_972, dataGroup_hi_lo_972};
  wire [7:0]    dataGroup_12_30 = dataGroup_lo_972[791:784];
  wire [1023:0] dataGroup_lo_973 = {dataGroup_lo_hi_973, dataGroup_lo_lo_973};
  wire [1023:0] dataGroup_hi_973 = {dataGroup_hi_hi_973, dataGroup_hi_lo_973};
  wire [7:0]    dataGroup_13_30 = dataGroup_lo_973[855:848];
  wire [1023:0] dataGroup_lo_974 = {dataGroup_lo_hi_974, dataGroup_lo_lo_974};
  wire [1023:0] dataGroup_hi_974 = {dataGroup_hi_hi_974, dataGroup_hi_lo_974};
  wire [7:0]    dataGroup_14_30 = dataGroup_lo_974[919:912];
  wire [1023:0] dataGroup_lo_975 = {dataGroup_lo_hi_975, dataGroup_lo_lo_975};
  wire [1023:0] dataGroup_hi_975 = {dataGroup_hi_hi_975, dataGroup_hi_lo_975};
  wire [7:0]    dataGroup_15_30 = dataGroup_lo_975[983:976];
  wire [1023:0] dataGroup_lo_976 = {dataGroup_lo_hi_976, dataGroup_lo_lo_976};
  wire [1023:0] dataGroup_hi_976 = {dataGroup_hi_hi_976, dataGroup_hi_lo_976};
  wire [7:0]    dataGroup_16_30 = dataGroup_hi_976[23:16];
  wire [1023:0] dataGroup_lo_977 = {dataGroup_lo_hi_977, dataGroup_lo_lo_977};
  wire [1023:0] dataGroup_hi_977 = {dataGroup_hi_hi_977, dataGroup_hi_lo_977};
  wire [7:0]    dataGroup_17_30 = dataGroup_hi_977[87:80];
  wire [1023:0] dataGroup_lo_978 = {dataGroup_lo_hi_978, dataGroup_lo_lo_978};
  wire [1023:0] dataGroup_hi_978 = {dataGroup_hi_hi_978, dataGroup_hi_lo_978};
  wire [7:0]    dataGroup_18_30 = dataGroup_hi_978[151:144];
  wire [1023:0] dataGroup_lo_979 = {dataGroup_lo_hi_979, dataGroup_lo_lo_979};
  wire [1023:0] dataGroup_hi_979 = {dataGroup_hi_hi_979, dataGroup_hi_lo_979};
  wire [7:0]    dataGroup_19_30 = dataGroup_hi_979[215:208];
  wire [1023:0] dataGroup_lo_980 = {dataGroup_lo_hi_980, dataGroup_lo_lo_980};
  wire [1023:0] dataGroup_hi_980 = {dataGroup_hi_hi_980, dataGroup_hi_lo_980};
  wire [7:0]    dataGroup_20_30 = dataGroup_hi_980[279:272];
  wire [1023:0] dataGroup_lo_981 = {dataGroup_lo_hi_981, dataGroup_lo_lo_981};
  wire [1023:0] dataGroup_hi_981 = {dataGroup_hi_hi_981, dataGroup_hi_lo_981};
  wire [7:0]    dataGroup_21_30 = dataGroup_hi_981[343:336];
  wire [1023:0] dataGroup_lo_982 = {dataGroup_lo_hi_982, dataGroup_lo_lo_982};
  wire [1023:0] dataGroup_hi_982 = {dataGroup_hi_hi_982, dataGroup_hi_lo_982};
  wire [7:0]    dataGroup_22_30 = dataGroup_hi_982[407:400];
  wire [1023:0] dataGroup_lo_983 = {dataGroup_lo_hi_983, dataGroup_lo_lo_983};
  wire [1023:0] dataGroup_hi_983 = {dataGroup_hi_hi_983, dataGroup_hi_lo_983};
  wire [7:0]    dataGroup_23_30 = dataGroup_hi_983[471:464];
  wire [1023:0] dataGroup_lo_984 = {dataGroup_lo_hi_984, dataGroup_lo_lo_984};
  wire [1023:0] dataGroup_hi_984 = {dataGroup_hi_hi_984, dataGroup_hi_lo_984};
  wire [7:0]    dataGroup_24_30 = dataGroup_hi_984[535:528];
  wire [1023:0] dataGroup_lo_985 = {dataGroup_lo_hi_985, dataGroup_lo_lo_985};
  wire [1023:0] dataGroup_hi_985 = {dataGroup_hi_hi_985, dataGroup_hi_lo_985};
  wire [7:0]    dataGroup_25_30 = dataGroup_hi_985[599:592];
  wire [1023:0] dataGroup_lo_986 = {dataGroup_lo_hi_986, dataGroup_lo_lo_986};
  wire [1023:0] dataGroup_hi_986 = {dataGroup_hi_hi_986, dataGroup_hi_lo_986};
  wire [7:0]    dataGroup_26_30 = dataGroup_hi_986[663:656];
  wire [1023:0] dataGroup_lo_987 = {dataGroup_lo_hi_987, dataGroup_lo_lo_987};
  wire [1023:0] dataGroup_hi_987 = {dataGroup_hi_hi_987, dataGroup_hi_lo_987};
  wire [7:0]    dataGroup_27_30 = dataGroup_hi_987[727:720];
  wire [1023:0] dataGroup_lo_988 = {dataGroup_lo_hi_988, dataGroup_lo_lo_988};
  wire [1023:0] dataGroup_hi_988 = {dataGroup_hi_hi_988, dataGroup_hi_lo_988};
  wire [7:0]    dataGroup_28_30 = dataGroup_hi_988[791:784];
  wire [1023:0] dataGroup_lo_989 = {dataGroup_lo_hi_989, dataGroup_lo_lo_989};
  wire [1023:0] dataGroup_hi_989 = {dataGroup_hi_hi_989, dataGroup_hi_lo_989};
  wire [7:0]    dataGroup_29_30 = dataGroup_hi_989[855:848];
  wire [1023:0] dataGroup_lo_990 = {dataGroup_lo_hi_990, dataGroup_lo_lo_990};
  wire [1023:0] dataGroup_hi_990 = {dataGroup_hi_hi_990, dataGroup_hi_lo_990};
  wire [7:0]    dataGroup_30_30 = dataGroup_hi_990[919:912];
  wire [1023:0] dataGroup_lo_991 = {dataGroup_lo_hi_991, dataGroup_lo_lo_991};
  wire [1023:0] dataGroup_hi_991 = {dataGroup_hi_hi_991, dataGroup_hi_lo_991};
  wire [7:0]    dataGroup_31_30 = dataGroup_hi_991[983:976];
  wire [15:0]   res_lo_lo_lo_lo_30 = {dataGroup_1_30, dataGroup_0_30};
  wire [15:0]   res_lo_lo_lo_hi_30 = {dataGroup_3_30, dataGroup_2_30};
  wire [31:0]   res_lo_lo_lo_30 = {res_lo_lo_lo_hi_30, res_lo_lo_lo_lo_30};
  wire [15:0]   res_lo_lo_hi_lo_30 = {dataGroup_5_30, dataGroup_4_30};
  wire [15:0]   res_lo_lo_hi_hi_30 = {dataGroup_7_30, dataGroup_6_30};
  wire [31:0]   res_lo_lo_hi_30 = {res_lo_lo_hi_hi_30, res_lo_lo_hi_lo_30};
  wire [63:0]   res_lo_lo_30 = {res_lo_lo_hi_30, res_lo_lo_lo_30};
  wire [15:0]   res_lo_hi_lo_lo_30 = {dataGroup_9_30, dataGroup_8_30};
  wire [15:0]   res_lo_hi_lo_hi_30 = {dataGroup_11_30, dataGroup_10_30};
  wire [31:0]   res_lo_hi_lo_30 = {res_lo_hi_lo_hi_30, res_lo_hi_lo_lo_30};
  wire [15:0]   res_lo_hi_hi_lo_30 = {dataGroup_13_30, dataGroup_12_30};
  wire [15:0]   res_lo_hi_hi_hi_30 = {dataGroup_15_30, dataGroup_14_30};
  wire [31:0]   res_lo_hi_hi_30 = {res_lo_hi_hi_hi_30, res_lo_hi_hi_lo_30};
  wire [63:0]   res_lo_hi_30 = {res_lo_hi_hi_30, res_lo_hi_lo_30};
  wire [127:0]  res_lo_30 = {res_lo_hi_30, res_lo_lo_30};
  wire [15:0]   res_hi_lo_lo_lo_30 = {dataGroup_17_30, dataGroup_16_30};
  wire [15:0]   res_hi_lo_lo_hi_30 = {dataGroup_19_30, dataGroup_18_30};
  wire [31:0]   res_hi_lo_lo_30 = {res_hi_lo_lo_hi_30, res_hi_lo_lo_lo_30};
  wire [15:0]   res_hi_lo_hi_lo_30 = {dataGroup_21_30, dataGroup_20_30};
  wire [15:0]   res_hi_lo_hi_hi_30 = {dataGroup_23_30, dataGroup_22_30};
  wire [31:0]   res_hi_lo_hi_30 = {res_hi_lo_hi_hi_30, res_hi_lo_hi_lo_30};
  wire [63:0]   res_hi_lo_30 = {res_hi_lo_hi_30, res_hi_lo_lo_30};
  wire [15:0]   res_hi_hi_lo_lo_30 = {dataGroup_25_30, dataGroup_24_30};
  wire [15:0]   res_hi_hi_lo_hi_30 = {dataGroup_27_30, dataGroup_26_30};
  wire [31:0]   res_hi_hi_lo_30 = {res_hi_hi_lo_hi_30, res_hi_hi_lo_lo_30};
  wire [15:0]   res_hi_hi_hi_lo_30 = {dataGroup_29_30, dataGroup_28_30};
  wire [15:0]   res_hi_hi_hi_hi_30 = {dataGroup_31_30, dataGroup_30_30};
  wire [31:0]   res_hi_hi_hi_30 = {res_hi_hi_hi_hi_30, res_hi_hi_hi_lo_30};
  wire [63:0]   res_hi_hi_30 = {res_hi_hi_hi_30, res_hi_hi_lo_30};
  wire [127:0]  res_hi_30 = {res_hi_hi_30, res_hi_lo_30};
  wire [255:0]  res_58 = {res_hi_30, res_lo_30};
  wire [1023:0] dataGroup_lo_992 = {dataGroup_lo_hi_992, dataGroup_lo_lo_992};
  wire [1023:0] dataGroup_hi_992 = {dataGroup_hi_hi_992, dataGroup_hi_lo_992};
  wire [7:0]    dataGroup_0_31 = dataGroup_lo_992[31:24];
  wire [1023:0] dataGroup_lo_993 = {dataGroup_lo_hi_993, dataGroup_lo_lo_993};
  wire [1023:0] dataGroup_hi_993 = {dataGroup_hi_hi_993, dataGroup_hi_lo_993};
  wire [7:0]    dataGroup_1_31 = dataGroup_lo_993[95:88];
  wire [1023:0] dataGroup_lo_994 = {dataGroup_lo_hi_994, dataGroup_lo_lo_994};
  wire [1023:0] dataGroup_hi_994 = {dataGroup_hi_hi_994, dataGroup_hi_lo_994};
  wire [7:0]    dataGroup_2_31 = dataGroup_lo_994[159:152];
  wire [1023:0] dataGroup_lo_995 = {dataGroup_lo_hi_995, dataGroup_lo_lo_995};
  wire [1023:0] dataGroup_hi_995 = {dataGroup_hi_hi_995, dataGroup_hi_lo_995};
  wire [7:0]    dataGroup_3_31 = dataGroup_lo_995[223:216];
  wire [1023:0] dataGroup_lo_996 = {dataGroup_lo_hi_996, dataGroup_lo_lo_996};
  wire [1023:0] dataGroup_hi_996 = {dataGroup_hi_hi_996, dataGroup_hi_lo_996};
  wire [7:0]    dataGroup_4_31 = dataGroup_lo_996[287:280];
  wire [1023:0] dataGroup_lo_997 = {dataGroup_lo_hi_997, dataGroup_lo_lo_997};
  wire [1023:0] dataGroup_hi_997 = {dataGroup_hi_hi_997, dataGroup_hi_lo_997};
  wire [7:0]    dataGroup_5_31 = dataGroup_lo_997[351:344];
  wire [1023:0] dataGroup_lo_998 = {dataGroup_lo_hi_998, dataGroup_lo_lo_998};
  wire [1023:0] dataGroup_hi_998 = {dataGroup_hi_hi_998, dataGroup_hi_lo_998};
  wire [7:0]    dataGroup_6_31 = dataGroup_lo_998[415:408];
  wire [1023:0] dataGroup_lo_999 = {dataGroup_lo_hi_999, dataGroup_lo_lo_999};
  wire [1023:0] dataGroup_hi_999 = {dataGroup_hi_hi_999, dataGroup_hi_lo_999};
  wire [7:0]    dataGroup_7_31 = dataGroup_lo_999[479:472];
  wire [1023:0] dataGroup_lo_1000 = {dataGroup_lo_hi_1000, dataGroup_lo_lo_1000};
  wire [1023:0] dataGroup_hi_1000 = {dataGroup_hi_hi_1000, dataGroup_hi_lo_1000};
  wire [7:0]    dataGroup_8_31 = dataGroup_lo_1000[543:536];
  wire [1023:0] dataGroup_lo_1001 = {dataGroup_lo_hi_1001, dataGroup_lo_lo_1001};
  wire [1023:0] dataGroup_hi_1001 = {dataGroup_hi_hi_1001, dataGroup_hi_lo_1001};
  wire [7:0]    dataGroup_9_31 = dataGroup_lo_1001[607:600];
  wire [1023:0] dataGroup_lo_1002 = {dataGroup_lo_hi_1002, dataGroup_lo_lo_1002};
  wire [1023:0] dataGroup_hi_1002 = {dataGroup_hi_hi_1002, dataGroup_hi_lo_1002};
  wire [7:0]    dataGroup_10_31 = dataGroup_lo_1002[671:664];
  wire [1023:0] dataGroup_lo_1003 = {dataGroup_lo_hi_1003, dataGroup_lo_lo_1003};
  wire [1023:0] dataGroup_hi_1003 = {dataGroup_hi_hi_1003, dataGroup_hi_lo_1003};
  wire [7:0]    dataGroup_11_31 = dataGroup_lo_1003[735:728];
  wire [1023:0] dataGroup_lo_1004 = {dataGroup_lo_hi_1004, dataGroup_lo_lo_1004};
  wire [1023:0] dataGroup_hi_1004 = {dataGroup_hi_hi_1004, dataGroup_hi_lo_1004};
  wire [7:0]    dataGroup_12_31 = dataGroup_lo_1004[799:792];
  wire [1023:0] dataGroup_lo_1005 = {dataGroup_lo_hi_1005, dataGroup_lo_lo_1005};
  wire [1023:0] dataGroup_hi_1005 = {dataGroup_hi_hi_1005, dataGroup_hi_lo_1005};
  wire [7:0]    dataGroup_13_31 = dataGroup_lo_1005[863:856];
  wire [1023:0] dataGroup_lo_1006 = {dataGroup_lo_hi_1006, dataGroup_lo_lo_1006};
  wire [1023:0] dataGroup_hi_1006 = {dataGroup_hi_hi_1006, dataGroup_hi_lo_1006};
  wire [7:0]    dataGroup_14_31 = dataGroup_lo_1006[927:920];
  wire [1023:0] dataGroup_lo_1007 = {dataGroup_lo_hi_1007, dataGroup_lo_lo_1007};
  wire [1023:0] dataGroup_hi_1007 = {dataGroup_hi_hi_1007, dataGroup_hi_lo_1007};
  wire [7:0]    dataGroup_15_31 = dataGroup_lo_1007[991:984];
  wire [1023:0] dataGroup_lo_1008 = {dataGroup_lo_hi_1008, dataGroup_lo_lo_1008};
  wire [1023:0] dataGroup_hi_1008 = {dataGroup_hi_hi_1008, dataGroup_hi_lo_1008};
  wire [7:0]    dataGroup_16_31 = dataGroup_hi_1008[31:24];
  wire [1023:0] dataGroup_lo_1009 = {dataGroup_lo_hi_1009, dataGroup_lo_lo_1009};
  wire [1023:0] dataGroup_hi_1009 = {dataGroup_hi_hi_1009, dataGroup_hi_lo_1009};
  wire [7:0]    dataGroup_17_31 = dataGroup_hi_1009[95:88];
  wire [1023:0] dataGroup_lo_1010 = {dataGroup_lo_hi_1010, dataGroup_lo_lo_1010};
  wire [1023:0] dataGroup_hi_1010 = {dataGroup_hi_hi_1010, dataGroup_hi_lo_1010};
  wire [7:0]    dataGroup_18_31 = dataGroup_hi_1010[159:152];
  wire [1023:0] dataGroup_lo_1011 = {dataGroup_lo_hi_1011, dataGroup_lo_lo_1011};
  wire [1023:0] dataGroup_hi_1011 = {dataGroup_hi_hi_1011, dataGroup_hi_lo_1011};
  wire [7:0]    dataGroup_19_31 = dataGroup_hi_1011[223:216];
  wire [1023:0] dataGroup_lo_1012 = {dataGroup_lo_hi_1012, dataGroup_lo_lo_1012};
  wire [1023:0] dataGroup_hi_1012 = {dataGroup_hi_hi_1012, dataGroup_hi_lo_1012};
  wire [7:0]    dataGroup_20_31 = dataGroup_hi_1012[287:280];
  wire [1023:0] dataGroup_lo_1013 = {dataGroup_lo_hi_1013, dataGroup_lo_lo_1013};
  wire [1023:0] dataGroup_hi_1013 = {dataGroup_hi_hi_1013, dataGroup_hi_lo_1013};
  wire [7:0]    dataGroup_21_31 = dataGroup_hi_1013[351:344];
  wire [1023:0] dataGroup_lo_1014 = {dataGroup_lo_hi_1014, dataGroup_lo_lo_1014};
  wire [1023:0] dataGroup_hi_1014 = {dataGroup_hi_hi_1014, dataGroup_hi_lo_1014};
  wire [7:0]    dataGroup_22_31 = dataGroup_hi_1014[415:408];
  wire [1023:0] dataGroup_lo_1015 = {dataGroup_lo_hi_1015, dataGroup_lo_lo_1015};
  wire [1023:0] dataGroup_hi_1015 = {dataGroup_hi_hi_1015, dataGroup_hi_lo_1015};
  wire [7:0]    dataGroup_23_31 = dataGroup_hi_1015[479:472];
  wire [1023:0] dataGroup_lo_1016 = {dataGroup_lo_hi_1016, dataGroup_lo_lo_1016};
  wire [1023:0] dataGroup_hi_1016 = {dataGroup_hi_hi_1016, dataGroup_hi_lo_1016};
  wire [7:0]    dataGroup_24_31 = dataGroup_hi_1016[543:536];
  wire [1023:0] dataGroup_lo_1017 = {dataGroup_lo_hi_1017, dataGroup_lo_lo_1017};
  wire [1023:0] dataGroup_hi_1017 = {dataGroup_hi_hi_1017, dataGroup_hi_lo_1017};
  wire [7:0]    dataGroup_25_31 = dataGroup_hi_1017[607:600];
  wire [1023:0] dataGroup_lo_1018 = {dataGroup_lo_hi_1018, dataGroup_lo_lo_1018};
  wire [1023:0] dataGroup_hi_1018 = {dataGroup_hi_hi_1018, dataGroup_hi_lo_1018};
  wire [7:0]    dataGroup_26_31 = dataGroup_hi_1018[671:664];
  wire [1023:0] dataGroup_lo_1019 = {dataGroup_lo_hi_1019, dataGroup_lo_lo_1019};
  wire [1023:0] dataGroup_hi_1019 = {dataGroup_hi_hi_1019, dataGroup_hi_lo_1019};
  wire [7:0]    dataGroup_27_31 = dataGroup_hi_1019[735:728];
  wire [1023:0] dataGroup_lo_1020 = {dataGroup_lo_hi_1020, dataGroup_lo_lo_1020};
  wire [1023:0] dataGroup_hi_1020 = {dataGroup_hi_hi_1020, dataGroup_hi_lo_1020};
  wire [7:0]    dataGroup_28_31 = dataGroup_hi_1020[799:792];
  wire [1023:0] dataGroup_lo_1021 = {dataGroup_lo_hi_1021, dataGroup_lo_lo_1021};
  wire [1023:0] dataGroup_hi_1021 = {dataGroup_hi_hi_1021, dataGroup_hi_lo_1021};
  wire [7:0]    dataGroup_29_31 = dataGroup_hi_1021[863:856];
  wire [1023:0] dataGroup_lo_1022 = {dataGroup_lo_hi_1022, dataGroup_lo_lo_1022};
  wire [1023:0] dataGroup_hi_1022 = {dataGroup_hi_hi_1022, dataGroup_hi_lo_1022};
  wire [7:0]    dataGroup_30_31 = dataGroup_hi_1022[927:920];
  wire [1023:0] dataGroup_lo_1023 = {dataGroup_lo_hi_1023, dataGroup_lo_lo_1023};
  wire [1023:0] dataGroup_hi_1023 = {dataGroup_hi_hi_1023, dataGroup_hi_lo_1023};
  wire [7:0]    dataGroup_31_31 = dataGroup_hi_1023[991:984];
  wire [15:0]   res_lo_lo_lo_lo_31 = {dataGroup_1_31, dataGroup_0_31};
  wire [15:0]   res_lo_lo_lo_hi_31 = {dataGroup_3_31, dataGroup_2_31};
  wire [31:0]   res_lo_lo_lo_31 = {res_lo_lo_lo_hi_31, res_lo_lo_lo_lo_31};
  wire [15:0]   res_lo_lo_hi_lo_31 = {dataGroup_5_31, dataGroup_4_31};
  wire [15:0]   res_lo_lo_hi_hi_31 = {dataGroup_7_31, dataGroup_6_31};
  wire [31:0]   res_lo_lo_hi_31 = {res_lo_lo_hi_hi_31, res_lo_lo_hi_lo_31};
  wire [63:0]   res_lo_lo_31 = {res_lo_lo_hi_31, res_lo_lo_lo_31};
  wire [15:0]   res_lo_hi_lo_lo_31 = {dataGroup_9_31, dataGroup_8_31};
  wire [15:0]   res_lo_hi_lo_hi_31 = {dataGroup_11_31, dataGroup_10_31};
  wire [31:0]   res_lo_hi_lo_31 = {res_lo_hi_lo_hi_31, res_lo_hi_lo_lo_31};
  wire [15:0]   res_lo_hi_hi_lo_31 = {dataGroup_13_31, dataGroup_12_31};
  wire [15:0]   res_lo_hi_hi_hi_31 = {dataGroup_15_31, dataGroup_14_31};
  wire [31:0]   res_lo_hi_hi_31 = {res_lo_hi_hi_hi_31, res_lo_hi_hi_lo_31};
  wire [63:0]   res_lo_hi_31 = {res_lo_hi_hi_31, res_lo_hi_lo_31};
  wire [127:0]  res_lo_31 = {res_lo_hi_31, res_lo_lo_31};
  wire [15:0]   res_hi_lo_lo_lo_31 = {dataGroup_17_31, dataGroup_16_31};
  wire [15:0]   res_hi_lo_lo_hi_31 = {dataGroup_19_31, dataGroup_18_31};
  wire [31:0]   res_hi_lo_lo_31 = {res_hi_lo_lo_hi_31, res_hi_lo_lo_lo_31};
  wire [15:0]   res_hi_lo_hi_lo_31 = {dataGroup_21_31, dataGroup_20_31};
  wire [15:0]   res_hi_lo_hi_hi_31 = {dataGroup_23_31, dataGroup_22_31};
  wire [31:0]   res_hi_lo_hi_31 = {res_hi_lo_hi_hi_31, res_hi_lo_hi_lo_31};
  wire [63:0]   res_hi_lo_31 = {res_hi_lo_hi_31, res_hi_lo_lo_31};
  wire [15:0]   res_hi_hi_lo_lo_31 = {dataGroup_25_31, dataGroup_24_31};
  wire [15:0]   res_hi_hi_lo_hi_31 = {dataGroup_27_31, dataGroup_26_31};
  wire [31:0]   res_hi_hi_lo_31 = {res_hi_hi_lo_hi_31, res_hi_hi_lo_lo_31};
  wire [15:0]   res_hi_hi_hi_lo_31 = {dataGroup_29_31, dataGroup_28_31};
  wire [15:0]   res_hi_hi_hi_hi_31 = {dataGroup_31_31, dataGroup_30_31};
  wire [31:0]   res_hi_hi_hi_31 = {res_hi_hi_hi_hi_31, res_hi_hi_hi_lo_31};
  wire [63:0]   res_hi_hi_31 = {res_hi_hi_hi_31, res_hi_hi_lo_31};
  wire [127:0]  res_hi_31 = {res_hi_hi_31, res_hi_lo_31};
  wire [255:0]  res_59 = {res_hi_31, res_lo_31};
  wire [1023:0] dataGroup_lo_1024 = {dataGroup_lo_hi_1024, dataGroup_lo_lo_1024};
  wire [1023:0] dataGroup_hi_1024 = {dataGroup_hi_hi_1024, dataGroup_hi_lo_1024};
  wire [7:0]    dataGroup_0_32 = dataGroup_lo_1024[39:32];
  wire [1023:0] dataGroup_lo_1025 = {dataGroup_lo_hi_1025, dataGroup_lo_lo_1025};
  wire [1023:0] dataGroup_hi_1025 = {dataGroup_hi_hi_1025, dataGroup_hi_lo_1025};
  wire [7:0]    dataGroup_1_32 = dataGroup_lo_1025[103:96];
  wire [1023:0] dataGroup_lo_1026 = {dataGroup_lo_hi_1026, dataGroup_lo_lo_1026};
  wire [1023:0] dataGroup_hi_1026 = {dataGroup_hi_hi_1026, dataGroup_hi_lo_1026};
  wire [7:0]    dataGroup_2_32 = dataGroup_lo_1026[167:160];
  wire [1023:0] dataGroup_lo_1027 = {dataGroup_lo_hi_1027, dataGroup_lo_lo_1027};
  wire [1023:0] dataGroup_hi_1027 = {dataGroup_hi_hi_1027, dataGroup_hi_lo_1027};
  wire [7:0]    dataGroup_3_32 = dataGroup_lo_1027[231:224];
  wire [1023:0] dataGroup_lo_1028 = {dataGroup_lo_hi_1028, dataGroup_lo_lo_1028};
  wire [1023:0] dataGroup_hi_1028 = {dataGroup_hi_hi_1028, dataGroup_hi_lo_1028};
  wire [7:0]    dataGroup_4_32 = dataGroup_lo_1028[295:288];
  wire [1023:0] dataGroup_lo_1029 = {dataGroup_lo_hi_1029, dataGroup_lo_lo_1029};
  wire [1023:0] dataGroup_hi_1029 = {dataGroup_hi_hi_1029, dataGroup_hi_lo_1029};
  wire [7:0]    dataGroup_5_32 = dataGroup_lo_1029[359:352];
  wire [1023:0] dataGroup_lo_1030 = {dataGroup_lo_hi_1030, dataGroup_lo_lo_1030};
  wire [1023:0] dataGroup_hi_1030 = {dataGroup_hi_hi_1030, dataGroup_hi_lo_1030};
  wire [7:0]    dataGroup_6_32 = dataGroup_lo_1030[423:416];
  wire [1023:0] dataGroup_lo_1031 = {dataGroup_lo_hi_1031, dataGroup_lo_lo_1031};
  wire [1023:0] dataGroup_hi_1031 = {dataGroup_hi_hi_1031, dataGroup_hi_lo_1031};
  wire [7:0]    dataGroup_7_32 = dataGroup_lo_1031[487:480];
  wire [1023:0] dataGroup_lo_1032 = {dataGroup_lo_hi_1032, dataGroup_lo_lo_1032};
  wire [1023:0] dataGroup_hi_1032 = {dataGroup_hi_hi_1032, dataGroup_hi_lo_1032};
  wire [7:0]    dataGroup_8_32 = dataGroup_lo_1032[551:544];
  wire [1023:0] dataGroup_lo_1033 = {dataGroup_lo_hi_1033, dataGroup_lo_lo_1033};
  wire [1023:0] dataGroup_hi_1033 = {dataGroup_hi_hi_1033, dataGroup_hi_lo_1033};
  wire [7:0]    dataGroup_9_32 = dataGroup_lo_1033[615:608];
  wire [1023:0] dataGroup_lo_1034 = {dataGroup_lo_hi_1034, dataGroup_lo_lo_1034};
  wire [1023:0] dataGroup_hi_1034 = {dataGroup_hi_hi_1034, dataGroup_hi_lo_1034};
  wire [7:0]    dataGroup_10_32 = dataGroup_lo_1034[679:672];
  wire [1023:0] dataGroup_lo_1035 = {dataGroup_lo_hi_1035, dataGroup_lo_lo_1035};
  wire [1023:0] dataGroup_hi_1035 = {dataGroup_hi_hi_1035, dataGroup_hi_lo_1035};
  wire [7:0]    dataGroup_11_32 = dataGroup_lo_1035[743:736];
  wire [1023:0] dataGroup_lo_1036 = {dataGroup_lo_hi_1036, dataGroup_lo_lo_1036};
  wire [1023:0] dataGroup_hi_1036 = {dataGroup_hi_hi_1036, dataGroup_hi_lo_1036};
  wire [7:0]    dataGroup_12_32 = dataGroup_lo_1036[807:800];
  wire [1023:0] dataGroup_lo_1037 = {dataGroup_lo_hi_1037, dataGroup_lo_lo_1037};
  wire [1023:0] dataGroup_hi_1037 = {dataGroup_hi_hi_1037, dataGroup_hi_lo_1037};
  wire [7:0]    dataGroup_13_32 = dataGroup_lo_1037[871:864];
  wire [1023:0] dataGroup_lo_1038 = {dataGroup_lo_hi_1038, dataGroup_lo_lo_1038};
  wire [1023:0] dataGroup_hi_1038 = {dataGroup_hi_hi_1038, dataGroup_hi_lo_1038};
  wire [7:0]    dataGroup_14_32 = dataGroup_lo_1038[935:928];
  wire [1023:0] dataGroup_lo_1039 = {dataGroup_lo_hi_1039, dataGroup_lo_lo_1039};
  wire [1023:0] dataGroup_hi_1039 = {dataGroup_hi_hi_1039, dataGroup_hi_lo_1039};
  wire [7:0]    dataGroup_15_32 = dataGroup_lo_1039[999:992];
  wire [1023:0] dataGroup_lo_1040 = {dataGroup_lo_hi_1040, dataGroup_lo_lo_1040};
  wire [1023:0] dataGroup_hi_1040 = {dataGroup_hi_hi_1040, dataGroup_hi_lo_1040};
  wire [7:0]    dataGroup_16_32 = dataGroup_hi_1040[39:32];
  wire [1023:0] dataGroup_lo_1041 = {dataGroup_lo_hi_1041, dataGroup_lo_lo_1041};
  wire [1023:0] dataGroup_hi_1041 = {dataGroup_hi_hi_1041, dataGroup_hi_lo_1041};
  wire [7:0]    dataGroup_17_32 = dataGroup_hi_1041[103:96];
  wire [1023:0] dataGroup_lo_1042 = {dataGroup_lo_hi_1042, dataGroup_lo_lo_1042};
  wire [1023:0] dataGroup_hi_1042 = {dataGroup_hi_hi_1042, dataGroup_hi_lo_1042};
  wire [7:0]    dataGroup_18_32 = dataGroup_hi_1042[167:160];
  wire [1023:0] dataGroup_lo_1043 = {dataGroup_lo_hi_1043, dataGroup_lo_lo_1043};
  wire [1023:0] dataGroup_hi_1043 = {dataGroup_hi_hi_1043, dataGroup_hi_lo_1043};
  wire [7:0]    dataGroup_19_32 = dataGroup_hi_1043[231:224];
  wire [1023:0] dataGroup_lo_1044 = {dataGroup_lo_hi_1044, dataGroup_lo_lo_1044};
  wire [1023:0] dataGroup_hi_1044 = {dataGroup_hi_hi_1044, dataGroup_hi_lo_1044};
  wire [7:0]    dataGroup_20_32 = dataGroup_hi_1044[295:288];
  wire [1023:0] dataGroup_lo_1045 = {dataGroup_lo_hi_1045, dataGroup_lo_lo_1045};
  wire [1023:0] dataGroup_hi_1045 = {dataGroup_hi_hi_1045, dataGroup_hi_lo_1045};
  wire [7:0]    dataGroup_21_32 = dataGroup_hi_1045[359:352];
  wire [1023:0] dataGroup_lo_1046 = {dataGroup_lo_hi_1046, dataGroup_lo_lo_1046};
  wire [1023:0] dataGroup_hi_1046 = {dataGroup_hi_hi_1046, dataGroup_hi_lo_1046};
  wire [7:0]    dataGroup_22_32 = dataGroup_hi_1046[423:416];
  wire [1023:0] dataGroup_lo_1047 = {dataGroup_lo_hi_1047, dataGroup_lo_lo_1047};
  wire [1023:0] dataGroup_hi_1047 = {dataGroup_hi_hi_1047, dataGroup_hi_lo_1047};
  wire [7:0]    dataGroup_23_32 = dataGroup_hi_1047[487:480];
  wire [1023:0] dataGroup_lo_1048 = {dataGroup_lo_hi_1048, dataGroup_lo_lo_1048};
  wire [1023:0] dataGroup_hi_1048 = {dataGroup_hi_hi_1048, dataGroup_hi_lo_1048};
  wire [7:0]    dataGroup_24_32 = dataGroup_hi_1048[551:544];
  wire [1023:0] dataGroup_lo_1049 = {dataGroup_lo_hi_1049, dataGroup_lo_lo_1049};
  wire [1023:0] dataGroup_hi_1049 = {dataGroup_hi_hi_1049, dataGroup_hi_lo_1049};
  wire [7:0]    dataGroup_25_32 = dataGroup_hi_1049[615:608];
  wire [1023:0] dataGroup_lo_1050 = {dataGroup_lo_hi_1050, dataGroup_lo_lo_1050};
  wire [1023:0] dataGroup_hi_1050 = {dataGroup_hi_hi_1050, dataGroup_hi_lo_1050};
  wire [7:0]    dataGroup_26_32 = dataGroup_hi_1050[679:672];
  wire [1023:0] dataGroup_lo_1051 = {dataGroup_lo_hi_1051, dataGroup_lo_lo_1051};
  wire [1023:0] dataGroup_hi_1051 = {dataGroup_hi_hi_1051, dataGroup_hi_lo_1051};
  wire [7:0]    dataGroup_27_32 = dataGroup_hi_1051[743:736];
  wire [1023:0] dataGroup_lo_1052 = {dataGroup_lo_hi_1052, dataGroup_lo_lo_1052};
  wire [1023:0] dataGroup_hi_1052 = {dataGroup_hi_hi_1052, dataGroup_hi_lo_1052};
  wire [7:0]    dataGroup_28_32 = dataGroup_hi_1052[807:800];
  wire [1023:0] dataGroup_lo_1053 = {dataGroup_lo_hi_1053, dataGroup_lo_lo_1053};
  wire [1023:0] dataGroup_hi_1053 = {dataGroup_hi_hi_1053, dataGroup_hi_lo_1053};
  wire [7:0]    dataGroup_29_32 = dataGroup_hi_1053[871:864];
  wire [1023:0] dataGroup_lo_1054 = {dataGroup_lo_hi_1054, dataGroup_lo_lo_1054};
  wire [1023:0] dataGroup_hi_1054 = {dataGroup_hi_hi_1054, dataGroup_hi_lo_1054};
  wire [7:0]    dataGroup_30_32 = dataGroup_hi_1054[935:928];
  wire [1023:0] dataGroup_lo_1055 = {dataGroup_lo_hi_1055, dataGroup_lo_lo_1055};
  wire [1023:0] dataGroup_hi_1055 = {dataGroup_hi_hi_1055, dataGroup_hi_lo_1055};
  wire [7:0]    dataGroup_31_32 = dataGroup_hi_1055[999:992];
  wire [15:0]   res_lo_lo_lo_lo_32 = {dataGroup_1_32, dataGroup_0_32};
  wire [15:0]   res_lo_lo_lo_hi_32 = {dataGroup_3_32, dataGroup_2_32};
  wire [31:0]   res_lo_lo_lo_32 = {res_lo_lo_lo_hi_32, res_lo_lo_lo_lo_32};
  wire [15:0]   res_lo_lo_hi_lo_32 = {dataGroup_5_32, dataGroup_4_32};
  wire [15:0]   res_lo_lo_hi_hi_32 = {dataGroup_7_32, dataGroup_6_32};
  wire [31:0]   res_lo_lo_hi_32 = {res_lo_lo_hi_hi_32, res_lo_lo_hi_lo_32};
  wire [63:0]   res_lo_lo_32 = {res_lo_lo_hi_32, res_lo_lo_lo_32};
  wire [15:0]   res_lo_hi_lo_lo_32 = {dataGroup_9_32, dataGroup_8_32};
  wire [15:0]   res_lo_hi_lo_hi_32 = {dataGroup_11_32, dataGroup_10_32};
  wire [31:0]   res_lo_hi_lo_32 = {res_lo_hi_lo_hi_32, res_lo_hi_lo_lo_32};
  wire [15:0]   res_lo_hi_hi_lo_32 = {dataGroup_13_32, dataGroup_12_32};
  wire [15:0]   res_lo_hi_hi_hi_32 = {dataGroup_15_32, dataGroup_14_32};
  wire [31:0]   res_lo_hi_hi_32 = {res_lo_hi_hi_hi_32, res_lo_hi_hi_lo_32};
  wire [63:0]   res_lo_hi_32 = {res_lo_hi_hi_32, res_lo_hi_lo_32};
  wire [127:0]  res_lo_32 = {res_lo_hi_32, res_lo_lo_32};
  wire [15:0]   res_hi_lo_lo_lo_32 = {dataGroup_17_32, dataGroup_16_32};
  wire [15:0]   res_hi_lo_lo_hi_32 = {dataGroup_19_32, dataGroup_18_32};
  wire [31:0]   res_hi_lo_lo_32 = {res_hi_lo_lo_hi_32, res_hi_lo_lo_lo_32};
  wire [15:0]   res_hi_lo_hi_lo_32 = {dataGroup_21_32, dataGroup_20_32};
  wire [15:0]   res_hi_lo_hi_hi_32 = {dataGroup_23_32, dataGroup_22_32};
  wire [31:0]   res_hi_lo_hi_32 = {res_hi_lo_hi_hi_32, res_hi_lo_hi_lo_32};
  wire [63:0]   res_hi_lo_32 = {res_hi_lo_hi_32, res_hi_lo_lo_32};
  wire [15:0]   res_hi_hi_lo_lo_32 = {dataGroup_25_32, dataGroup_24_32};
  wire [15:0]   res_hi_hi_lo_hi_32 = {dataGroup_27_32, dataGroup_26_32};
  wire [31:0]   res_hi_hi_lo_32 = {res_hi_hi_lo_hi_32, res_hi_hi_lo_lo_32};
  wire [15:0]   res_hi_hi_hi_lo_32 = {dataGroup_29_32, dataGroup_28_32};
  wire [15:0]   res_hi_hi_hi_hi_32 = {dataGroup_31_32, dataGroup_30_32};
  wire [31:0]   res_hi_hi_hi_32 = {res_hi_hi_hi_hi_32, res_hi_hi_hi_lo_32};
  wire [63:0]   res_hi_hi_32 = {res_hi_hi_hi_32, res_hi_hi_lo_32};
  wire [127:0]  res_hi_32 = {res_hi_hi_32, res_hi_lo_32};
  wire [255:0]  res_60 = {res_hi_32, res_lo_32};
  wire [1023:0] dataGroup_lo_1056 = {dataGroup_lo_hi_1056, dataGroup_lo_lo_1056};
  wire [1023:0] dataGroup_hi_1056 = {dataGroup_hi_hi_1056, dataGroup_hi_lo_1056};
  wire [7:0]    dataGroup_0_33 = dataGroup_lo_1056[47:40];
  wire [1023:0] dataGroup_lo_1057 = {dataGroup_lo_hi_1057, dataGroup_lo_lo_1057};
  wire [1023:0] dataGroup_hi_1057 = {dataGroup_hi_hi_1057, dataGroup_hi_lo_1057};
  wire [7:0]    dataGroup_1_33 = dataGroup_lo_1057[111:104];
  wire [1023:0] dataGroup_lo_1058 = {dataGroup_lo_hi_1058, dataGroup_lo_lo_1058};
  wire [1023:0] dataGroup_hi_1058 = {dataGroup_hi_hi_1058, dataGroup_hi_lo_1058};
  wire [7:0]    dataGroup_2_33 = dataGroup_lo_1058[175:168];
  wire [1023:0] dataGroup_lo_1059 = {dataGroup_lo_hi_1059, dataGroup_lo_lo_1059};
  wire [1023:0] dataGroup_hi_1059 = {dataGroup_hi_hi_1059, dataGroup_hi_lo_1059};
  wire [7:0]    dataGroup_3_33 = dataGroup_lo_1059[239:232];
  wire [1023:0] dataGroup_lo_1060 = {dataGroup_lo_hi_1060, dataGroup_lo_lo_1060};
  wire [1023:0] dataGroup_hi_1060 = {dataGroup_hi_hi_1060, dataGroup_hi_lo_1060};
  wire [7:0]    dataGroup_4_33 = dataGroup_lo_1060[303:296];
  wire [1023:0] dataGroup_lo_1061 = {dataGroup_lo_hi_1061, dataGroup_lo_lo_1061};
  wire [1023:0] dataGroup_hi_1061 = {dataGroup_hi_hi_1061, dataGroup_hi_lo_1061};
  wire [7:0]    dataGroup_5_33 = dataGroup_lo_1061[367:360];
  wire [1023:0] dataGroup_lo_1062 = {dataGroup_lo_hi_1062, dataGroup_lo_lo_1062};
  wire [1023:0] dataGroup_hi_1062 = {dataGroup_hi_hi_1062, dataGroup_hi_lo_1062};
  wire [7:0]    dataGroup_6_33 = dataGroup_lo_1062[431:424];
  wire [1023:0] dataGroup_lo_1063 = {dataGroup_lo_hi_1063, dataGroup_lo_lo_1063};
  wire [1023:0] dataGroup_hi_1063 = {dataGroup_hi_hi_1063, dataGroup_hi_lo_1063};
  wire [7:0]    dataGroup_7_33 = dataGroup_lo_1063[495:488];
  wire [1023:0] dataGroup_lo_1064 = {dataGroup_lo_hi_1064, dataGroup_lo_lo_1064};
  wire [1023:0] dataGroup_hi_1064 = {dataGroup_hi_hi_1064, dataGroup_hi_lo_1064};
  wire [7:0]    dataGroup_8_33 = dataGroup_lo_1064[559:552];
  wire [1023:0] dataGroup_lo_1065 = {dataGroup_lo_hi_1065, dataGroup_lo_lo_1065};
  wire [1023:0] dataGroup_hi_1065 = {dataGroup_hi_hi_1065, dataGroup_hi_lo_1065};
  wire [7:0]    dataGroup_9_33 = dataGroup_lo_1065[623:616];
  wire [1023:0] dataGroup_lo_1066 = {dataGroup_lo_hi_1066, dataGroup_lo_lo_1066};
  wire [1023:0] dataGroup_hi_1066 = {dataGroup_hi_hi_1066, dataGroup_hi_lo_1066};
  wire [7:0]    dataGroup_10_33 = dataGroup_lo_1066[687:680];
  wire [1023:0] dataGroup_lo_1067 = {dataGroup_lo_hi_1067, dataGroup_lo_lo_1067};
  wire [1023:0] dataGroup_hi_1067 = {dataGroup_hi_hi_1067, dataGroup_hi_lo_1067};
  wire [7:0]    dataGroup_11_33 = dataGroup_lo_1067[751:744];
  wire [1023:0] dataGroup_lo_1068 = {dataGroup_lo_hi_1068, dataGroup_lo_lo_1068};
  wire [1023:0] dataGroup_hi_1068 = {dataGroup_hi_hi_1068, dataGroup_hi_lo_1068};
  wire [7:0]    dataGroup_12_33 = dataGroup_lo_1068[815:808];
  wire [1023:0] dataGroup_lo_1069 = {dataGroup_lo_hi_1069, dataGroup_lo_lo_1069};
  wire [1023:0] dataGroup_hi_1069 = {dataGroup_hi_hi_1069, dataGroup_hi_lo_1069};
  wire [7:0]    dataGroup_13_33 = dataGroup_lo_1069[879:872];
  wire [1023:0] dataGroup_lo_1070 = {dataGroup_lo_hi_1070, dataGroup_lo_lo_1070};
  wire [1023:0] dataGroup_hi_1070 = {dataGroup_hi_hi_1070, dataGroup_hi_lo_1070};
  wire [7:0]    dataGroup_14_33 = dataGroup_lo_1070[943:936];
  wire [1023:0] dataGroup_lo_1071 = {dataGroup_lo_hi_1071, dataGroup_lo_lo_1071};
  wire [1023:0] dataGroup_hi_1071 = {dataGroup_hi_hi_1071, dataGroup_hi_lo_1071};
  wire [7:0]    dataGroup_15_33 = dataGroup_lo_1071[1007:1000];
  wire [1023:0] dataGroup_lo_1072 = {dataGroup_lo_hi_1072, dataGroup_lo_lo_1072};
  wire [1023:0] dataGroup_hi_1072 = {dataGroup_hi_hi_1072, dataGroup_hi_lo_1072};
  wire [7:0]    dataGroup_16_33 = dataGroup_hi_1072[47:40];
  wire [1023:0] dataGroup_lo_1073 = {dataGroup_lo_hi_1073, dataGroup_lo_lo_1073};
  wire [1023:0] dataGroup_hi_1073 = {dataGroup_hi_hi_1073, dataGroup_hi_lo_1073};
  wire [7:0]    dataGroup_17_33 = dataGroup_hi_1073[111:104];
  wire [1023:0] dataGroup_lo_1074 = {dataGroup_lo_hi_1074, dataGroup_lo_lo_1074};
  wire [1023:0] dataGroup_hi_1074 = {dataGroup_hi_hi_1074, dataGroup_hi_lo_1074};
  wire [7:0]    dataGroup_18_33 = dataGroup_hi_1074[175:168];
  wire [1023:0] dataGroup_lo_1075 = {dataGroup_lo_hi_1075, dataGroup_lo_lo_1075};
  wire [1023:0] dataGroup_hi_1075 = {dataGroup_hi_hi_1075, dataGroup_hi_lo_1075};
  wire [7:0]    dataGroup_19_33 = dataGroup_hi_1075[239:232];
  wire [1023:0] dataGroup_lo_1076 = {dataGroup_lo_hi_1076, dataGroup_lo_lo_1076};
  wire [1023:0] dataGroup_hi_1076 = {dataGroup_hi_hi_1076, dataGroup_hi_lo_1076};
  wire [7:0]    dataGroup_20_33 = dataGroup_hi_1076[303:296];
  wire [1023:0] dataGroup_lo_1077 = {dataGroup_lo_hi_1077, dataGroup_lo_lo_1077};
  wire [1023:0] dataGroup_hi_1077 = {dataGroup_hi_hi_1077, dataGroup_hi_lo_1077};
  wire [7:0]    dataGroup_21_33 = dataGroup_hi_1077[367:360];
  wire [1023:0] dataGroup_lo_1078 = {dataGroup_lo_hi_1078, dataGroup_lo_lo_1078};
  wire [1023:0] dataGroup_hi_1078 = {dataGroup_hi_hi_1078, dataGroup_hi_lo_1078};
  wire [7:0]    dataGroup_22_33 = dataGroup_hi_1078[431:424];
  wire [1023:0] dataGroup_lo_1079 = {dataGroup_lo_hi_1079, dataGroup_lo_lo_1079};
  wire [1023:0] dataGroup_hi_1079 = {dataGroup_hi_hi_1079, dataGroup_hi_lo_1079};
  wire [7:0]    dataGroup_23_33 = dataGroup_hi_1079[495:488];
  wire [1023:0] dataGroup_lo_1080 = {dataGroup_lo_hi_1080, dataGroup_lo_lo_1080};
  wire [1023:0] dataGroup_hi_1080 = {dataGroup_hi_hi_1080, dataGroup_hi_lo_1080};
  wire [7:0]    dataGroup_24_33 = dataGroup_hi_1080[559:552];
  wire [1023:0] dataGroup_lo_1081 = {dataGroup_lo_hi_1081, dataGroup_lo_lo_1081};
  wire [1023:0] dataGroup_hi_1081 = {dataGroup_hi_hi_1081, dataGroup_hi_lo_1081};
  wire [7:0]    dataGroup_25_33 = dataGroup_hi_1081[623:616];
  wire [1023:0] dataGroup_lo_1082 = {dataGroup_lo_hi_1082, dataGroup_lo_lo_1082};
  wire [1023:0] dataGroup_hi_1082 = {dataGroup_hi_hi_1082, dataGroup_hi_lo_1082};
  wire [7:0]    dataGroup_26_33 = dataGroup_hi_1082[687:680];
  wire [1023:0] dataGroup_lo_1083 = {dataGroup_lo_hi_1083, dataGroup_lo_lo_1083};
  wire [1023:0] dataGroup_hi_1083 = {dataGroup_hi_hi_1083, dataGroup_hi_lo_1083};
  wire [7:0]    dataGroup_27_33 = dataGroup_hi_1083[751:744];
  wire [1023:0] dataGroup_lo_1084 = {dataGroup_lo_hi_1084, dataGroup_lo_lo_1084};
  wire [1023:0] dataGroup_hi_1084 = {dataGroup_hi_hi_1084, dataGroup_hi_lo_1084};
  wire [7:0]    dataGroup_28_33 = dataGroup_hi_1084[815:808];
  wire [1023:0] dataGroup_lo_1085 = {dataGroup_lo_hi_1085, dataGroup_lo_lo_1085};
  wire [1023:0] dataGroup_hi_1085 = {dataGroup_hi_hi_1085, dataGroup_hi_lo_1085};
  wire [7:0]    dataGroup_29_33 = dataGroup_hi_1085[879:872];
  wire [1023:0] dataGroup_lo_1086 = {dataGroup_lo_hi_1086, dataGroup_lo_lo_1086};
  wire [1023:0] dataGroup_hi_1086 = {dataGroup_hi_hi_1086, dataGroup_hi_lo_1086};
  wire [7:0]    dataGroup_30_33 = dataGroup_hi_1086[943:936];
  wire [1023:0] dataGroup_lo_1087 = {dataGroup_lo_hi_1087, dataGroup_lo_lo_1087};
  wire [1023:0] dataGroup_hi_1087 = {dataGroup_hi_hi_1087, dataGroup_hi_lo_1087};
  wire [7:0]    dataGroup_31_33 = dataGroup_hi_1087[1007:1000];
  wire [15:0]   res_lo_lo_lo_lo_33 = {dataGroup_1_33, dataGroup_0_33};
  wire [15:0]   res_lo_lo_lo_hi_33 = {dataGroup_3_33, dataGroup_2_33};
  wire [31:0]   res_lo_lo_lo_33 = {res_lo_lo_lo_hi_33, res_lo_lo_lo_lo_33};
  wire [15:0]   res_lo_lo_hi_lo_33 = {dataGroup_5_33, dataGroup_4_33};
  wire [15:0]   res_lo_lo_hi_hi_33 = {dataGroup_7_33, dataGroup_6_33};
  wire [31:0]   res_lo_lo_hi_33 = {res_lo_lo_hi_hi_33, res_lo_lo_hi_lo_33};
  wire [63:0]   res_lo_lo_33 = {res_lo_lo_hi_33, res_lo_lo_lo_33};
  wire [15:0]   res_lo_hi_lo_lo_33 = {dataGroup_9_33, dataGroup_8_33};
  wire [15:0]   res_lo_hi_lo_hi_33 = {dataGroup_11_33, dataGroup_10_33};
  wire [31:0]   res_lo_hi_lo_33 = {res_lo_hi_lo_hi_33, res_lo_hi_lo_lo_33};
  wire [15:0]   res_lo_hi_hi_lo_33 = {dataGroup_13_33, dataGroup_12_33};
  wire [15:0]   res_lo_hi_hi_hi_33 = {dataGroup_15_33, dataGroup_14_33};
  wire [31:0]   res_lo_hi_hi_33 = {res_lo_hi_hi_hi_33, res_lo_hi_hi_lo_33};
  wire [63:0]   res_lo_hi_33 = {res_lo_hi_hi_33, res_lo_hi_lo_33};
  wire [127:0]  res_lo_33 = {res_lo_hi_33, res_lo_lo_33};
  wire [15:0]   res_hi_lo_lo_lo_33 = {dataGroup_17_33, dataGroup_16_33};
  wire [15:0]   res_hi_lo_lo_hi_33 = {dataGroup_19_33, dataGroup_18_33};
  wire [31:0]   res_hi_lo_lo_33 = {res_hi_lo_lo_hi_33, res_hi_lo_lo_lo_33};
  wire [15:0]   res_hi_lo_hi_lo_33 = {dataGroup_21_33, dataGroup_20_33};
  wire [15:0]   res_hi_lo_hi_hi_33 = {dataGroup_23_33, dataGroup_22_33};
  wire [31:0]   res_hi_lo_hi_33 = {res_hi_lo_hi_hi_33, res_hi_lo_hi_lo_33};
  wire [63:0]   res_hi_lo_33 = {res_hi_lo_hi_33, res_hi_lo_lo_33};
  wire [15:0]   res_hi_hi_lo_lo_33 = {dataGroup_25_33, dataGroup_24_33};
  wire [15:0]   res_hi_hi_lo_hi_33 = {dataGroup_27_33, dataGroup_26_33};
  wire [31:0]   res_hi_hi_lo_33 = {res_hi_hi_lo_hi_33, res_hi_hi_lo_lo_33};
  wire [15:0]   res_hi_hi_hi_lo_33 = {dataGroup_29_33, dataGroup_28_33};
  wire [15:0]   res_hi_hi_hi_hi_33 = {dataGroup_31_33, dataGroup_30_33};
  wire [31:0]   res_hi_hi_hi_33 = {res_hi_hi_hi_hi_33, res_hi_hi_hi_lo_33};
  wire [63:0]   res_hi_hi_33 = {res_hi_hi_hi_33, res_hi_hi_lo_33};
  wire [127:0]  res_hi_33 = {res_hi_hi_33, res_hi_lo_33};
  wire [255:0]  res_61 = {res_hi_33, res_lo_33};
  wire [1023:0] dataGroup_lo_1088 = {dataGroup_lo_hi_1088, dataGroup_lo_lo_1088};
  wire [1023:0] dataGroup_hi_1088 = {dataGroup_hi_hi_1088, dataGroup_hi_lo_1088};
  wire [7:0]    dataGroup_0_34 = dataGroup_lo_1088[55:48];
  wire [1023:0] dataGroup_lo_1089 = {dataGroup_lo_hi_1089, dataGroup_lo_lo_1089};
  wire [1023:0] dataGroup_hi_1089 = {dataGroup_hi_hi_1089, dataGroup_hi_lo_1089};
  wire [7:0]    dataGroup_1_34 = dataGroup_lo_1089[119:112];
  wire [1023:0] dataGroup_lo_1090 = {dataGroup_lo_hi_1090, dataGroup_lo_lo_1090};
  wire [1023:0] dataGroup_hi_1090 = {dataGroup_hi_hi_1090, dataGroup_hi_lo_1090};
  wire [7:0]    dataGroup_2_34 = dataGroup_lo_1090[183:176];
  wire [1023:0] dataGroup_lo_1091 = {dataGroup_lo_hi_1091, dataGroup_lo_lo_1091};
  wire [1023:0] dataGroup_hi_1091 = {dataGroup_hi_hi_1091, dataGroup_hi_lo_1091};
  wire [7:0]    dataGroup_3_34 = dataGroup_lo_1091[247:240];
  wire [1023:0] dataGroup_lo_1092 = {dataGroup_lo_hi_1092, dataGroup_lo_lo_1092};
  wire [1023:0] dataGroup_hi_1092 = {dataGroup_hi_hi_1092, dataGroup_hi_lo_1092};
  wire [7:0]    dataGroup_4_34 = dataGroup_lo_1092[311:304];
  wire [1023:0] dataGroup_lo_1093 = {dataGroup_lo_hi_1093, dataGroup_lo_lo_1093};
  wire [1023:0] dataGroup_hi_1093 = {dataGroup_hi_hi_1093, dataGroup_hi_lo_1093};
  wire [7:0]    dataGroup_5_34 = dataGroup_lo_1093[375:368];
  wire [1023:0] dataGroup_lo_1094 = {dataGroup_lo_hi_1094, dataGroup_lo_lo_1094};
  wire [1023:0] dataGroup_hi_1094 = {dataGroup_hi_hi_1094, dataGroup_hi_lo_1094};
  wire [7:0]    dataGroup_6_34 = dataGroup_lo_1094[439:432];
  wire [1023:0] dataGroup_lo_1095 = {dataGroup_lo_hi_1095, dataGroup_lo_lo_1095};
  wire [1023:0] dataGroup_hi_1095 = {dataGroup_hi_hi_1095, dataGroup_hi_lo_1095};
  wire [7:0]    dataGroup_7_34 = dataGroup_lo_1095[503:496];
  wire [1023:0] dataGroup_lo_1096 = {dataGroup_lo_hi_1096, dataGroup_lo_lo_1096};
  wire [1023:0] dataGroup_hi_1096 = {dataGroup_hi_hi_1096, dataGroup_hi_lo_1096};
  wire [7:0]    dataGroup_8_34 = dataGroup_lo_1096[567:560];
  wire [1023:0] dataGroup_lo_1097 = {dataGroup_lo_hi_1097, dataGroup_lo_lo_1097};
  wire [1023:0] dataGroup_hi_1097 = {dataGroup_hi_hi_1097, dataGroup_hi_lo_1097};
  wire [7:0]    dataGroup_9_34 = dataGroup_lo_1097[631:624];
  wire [1023:0] dataGroup_lo_1098 = {dataGroup_lo_hi_1098, dataGroup_lo_lo_1098};
  wire [1023:0] dataGroup_hi_1098 = {dataGroup_hi_hi_1098, dataGroup_hi_lo_1098};
  wire [7:0]    dataGroup_10_34 = dataGroup_lo_1098[695:688];
  wire [1023:0] dataGroup_lo_1099 = {dataGroup_lo_hi_1099, dataGroup_lo_lo_1099};
  wire [1023:0] dataGroup_hi_1099 = {dataGroup_hi_hi_1099, dataGroup_hi_lo_1099};
  wire [7:0]    dataGroup_11_34 = dataGroup_lo_1099[759:752];
  wire [1023:0] dataGroup_lo_1100 = {dataGroup_lo_hi_1100, dataGroup_lo_lo_1100};
  wire [1023:0] dataGroup_hi_1100 = {dataGroup_hi_hi_1100, dataGroup_hi_lo_1100};
  wire [7:0]    dataGroup_12_34 = dataGroup_lo_1100[823:816];
  wire [1023:0] dataGroup_lo_1101 = {dataGroup_lo_hi_1101, dataGroup_lo_lo_1101};
  wire [1023:0] dataGroup_hi_1101 = {dataGroup_hi_hi_1101, dataGroup_hi_lo_1101};
  wire [7:0]    dataGroup_13_34 = dataGroup_lo_1101[887:880];
  wire [1023:0] dataGroup_lo_1102 = {dataGroup_lo_hi_1102, dataGroup_lo_lo_1102};
  wire [1023:0] dataGroup_hi_1102 = {dataGroup_hi_hi_1102, dataGroup_hi_lo_1102};
  wire [7:0]    dataGroup_14_34 = dataGroup_lo_1102[951:944];
  wire [1023:0] dataGroup_lo_1103 = {dataGroup_lo_hi_1103, dataGroup_lo_lo_1103};
  wire [1023:0] dataGroup_hi_1103 = {dataGroup_hi_hi_1103, dataGroup_hi_lo_1103};
  wire [7:0]    dataGroup_15_34 = dataGroup_lo_1103[1015:1008];
  wire [1023:0] dataGroup_lo_1104 = {dataGroup_lo_hi_1104, dataGroup_lo_lo_1104};
  wire [1023:0] dataGroup_hi_1104 = {dataGroup_hi_hi_1104, dataGroup_hi_lo_1104};
  wire [7:0]    dataGroup_16_34 = dataGroup_hi_1104[55:48];
  wire [1023:0] dataGroup_lo_1105 = {dataGroup_lo_hi_1105, dataGroup_lo_lo_1105};
  wire [1023:0] dataGroup_hi_1105 = {dataGroup_hi_hi_1105, dataGroup_hi_lo_1105};
  wire [7:0]    dataGroup_17_34 = dataGroup_hi_1105[119:112];
  wire [1023:0] dataGroup_lo_1106 = {dataGroup_lo_hi_1106, dataGroup_lo_lo_1106};
  wire [1023:0] dataGroup_hi_1106 = {dataGroup_hi_hi_1106, dataGroup_hi_lo_1106};
  wire [7:0]    dataGroup_18_34 = dataGroup_hi_1106[183:176];
  wire [1023:0] dataGroup_lo_1107 = {dataGroup_lo_hi_1107, dataGroup_lo_lo_1107};
  wire [1023:0] dataGroup_hi_1107 = {dataGroup_hi_hi_1107, dataGroup_hi_lo_1107};
  wire [7:0]    dataGroup_19_34 = dataGroup_hi_1107[247:240];
  wire [1023:0] dataGroup_lo_1108 = {dataGroup_lo_hi_1108, dataGroup_lo_lo_1108};
  wire [1023:0] dataGroup_hi_1108 = {dataGroup_hi_hi_1108, dataGroup_hi_lo_1108};
  wire [7:0]    dataGroup_20_34 = dataGroup_hi_1108[311:304];
  wire [1023:0] dataGroup_lo_1109 = {dataGroup_lo_hi_1109, dataGroup_lo_lo_1109};
  wire [1023:0] dataGroup_hi_1109 = {dataGroup_hi_hi_1109, dataGroup_hi_lo_1109};
  wire [7:0]    dataGroup_21_34 = dataGroup_hi_1109[375:368];
  wire [1023:0] dataGroup_lo_1110 = {dataGroup_lo_hi_1110, dataGroup_lo_lo_1110};
  wire [1023:0] dataGroup_hi_1110 = {dataGroup_hi_hi_1110, dataGroup_hi_lo_1110};
  wire [7:0]    dataGroup_22_34 = dataGroup_hi_1110[439:432];
  wire [1023:0] dataGroup_lo_1111 = {dataGroup_lo_hi_1111, dataGroup_lo_lo_1111};
  wire [1023:0] dataGroup_hi_1111 = {dataGroup_hi_hi_1111, dataGroup_hi_lo_1111};
  wire [7:0]    dataGroup_23_34 = dataGroup_hi_1111[503:496];
  wire [1023:0] dataGroup_lo_1112 = {dataGroup_lo_hi_1112, dataGroup_lo_lo_1112};
  wire [1023:0] dataGroup_hi_1112 = {dataGroup_hi_hi_1112, dataGroup_hi_lo_1112};
  wire [7:0]    dataGroup_24_34 = dataGroup_hi_1112[567:560];
  wire [1023:0] dataGroup_lo_1113 = {dataGroup_lo_hi_1113, dataGroup_lo_lo_1113};
  wire [1023:0] dataGroup_hi_1113 = {dataGroup_hi_hi_1113, dataGroup_hi_lo_1113};
  wire [7:0]    dataGroup_25_34 = dataGroup_hi_1113[631:624];
  wire [1023:0] dataGroup_lo_1114 = {dataGroup_lo_hi_1114, dataGroup_lo_lo_1114};
  wire [1023:0] dataGroup_hi_1114 = {dataGroup_hi_hi_1114, dataGroup_hi_lo_1114};
  wire [7:0]    dataGroup_26_34 = dataGroup_hi_1114[695:688];
  wire [1023:0] dataGroup_lo_1115 = {dataGroup_lo_hi_1115, dataGroup_lo_lo_1115};
  wire [1023:0] dataGroup_hi_1115 = {dataGroup_hi_hi_1115, dataGroup_hi_lo_1115};
  wire [7:0]    dataGroup_27_34 = dataGroup_hi_1115[759:752];
  wire [1023:0] dataGroup_lo_1116 = {dataGroup_lo_hi_1116, dataGroup_lo_lo_1116};
  wire [1023:0] dataGroup_hi_1116 = {dataGroup_hi_hi_1116, dataGroup_hi_lo_1116};
  wire [7:0]    dataGroup_28_34 = dataGroup_hi_1116[823:816];
  wire [1023:0] dataGroup_lo_1117 = {dataGroup_lo_hi_1117, dataGroup_lo_lo_1117};
  wire [1023:0] dataGroup_hi_1117 = {dataGroup_hi_hi_1117, dataGroup_hi_lo_1117};
  wire [7:0]    dataGroup_29_34 = dataGroup_hi_1117[887:880];
  wire [1023:0] dataGroup_lo_1118 = {dataGroup_lo_hi_1118, dataGroup_lo_lo_1118};
  wire [1023:0] dataGroup_hi_1118 = {dataGroup_hi_hi_1118, dataGroup_hi_lo_1118};
  wire [7:0]    dataGroup_30_34 = dataGroup_hi_1118[951:944];
  wire [1023:0] dataGroup_lo_1119 = {dataGroup_lo_hi_1119, dataGroup_lo_lo_1119};
  wire [1023:0] dataGroup_hi_1119 = {dataGroup_hi_hi_1119, dataGroup_hi_lo_1119};
  wire [7:0]    dataGroup_31_34 = dataGroup_hi_1119[1015:1008];
  wire [15:0]   res_lo_lo_lo_lo_34 = {dataGroup_1_34, dataGroup_0_34};
  wire [15:0]   res_lo_lo_lo_hi_34 = {dataGroup_3_34, dataGroup_2_34};
  wire [31:0]   res_lo_lo_lo_34 = {res_lo_lo_lo_hi_34, res_lo_lo_lo_lo_34};
  wire [15:0]   res_lo_lo_hi_lo_34 = {dataGroup_5_34, dataGroup_4_34};
  wire [15:0]   res_lo_lo_hi_hi_34 = {dataGroup_7_34, dataGroup_6_34};
  wire [31:0]   res_lo_lo_hi_34 = {res_lo_lo_hi_hi_34, res_lo_lo_hi_lo_34};
  wire [63:0]   res_lo_lo_34 = {res_lo_lo_hi_34, res_lo_lo_lo_34};
  wire [15:0]   res_lo_hi_lo_lo_34 = {dataGroup_9_34, dataGroup_8_34};
  wire [15:0]   res_lo_hi_lo_hi_34 = {dataGroup_11_34, dataGroup_10_34};
  wire [31:0]   res_lo_hi_lo_34 = {res_lo_hi_lo_hi_34, res_lo_hi_lo_lo_34};
  wire [15:0]   res_lo_hi_hi_lo_34 = {dataGroup_13_34, dataGroup_12_34};
  wire [15:0]   res_lo_hi_hi_hi_34 = {dataGroup_15_34, dataGroup_14_34};
  wire [31:0]   res_lo_hi_hi_34 = {res_lo_hi_hi_hi_34, res_lo_hi_hi_lo_34};
  wire [63:0]   res_lo_hi_34 = {res_lo_hi_hi_34, res_lo_hi_lo_34};
  wire [127:0]  res_lo_34 = {res_lo_hi_34, res_lo_lo_34};
  wire [15:0]   res_hi_lo_lo_lo_34 = {dataGroup_17_34, dataGroup_16_34};
  wire [15:0]   res_hi_lo_lo_hi_34 = {dataGroup_19_34, dataGroup_18_34};
  wire [31:0]   res_hi_lo_lo_34 = {res_hi_lo_lo_hi_34, res_hi_lo_lo_lo_34};
  wire [15:0]   res_hi_lo_hi_lo_34 = {dataGroup_21_34, dataGroup_20_34};
  wire [15:0]   res_hi_lo_hi_hi_34 = {dataGroup_23_34, dataGroup_22_34};
  wire [31:0]   res_hi_lo_hi_34 = {res_hi_lo_hi_hi_34, res_hi_lo_hi_lo_34};
  wire [63:0]   res_hi_lo_34 = {res_hi_lo_hi_34, res_hi_lo_lo_34};
  wire [15:0]   res_hi_hi_lo_lo_34 = {dataGroup_25_34, dataGroup_24_34};
  wire [15:0]   res_hi_hi_lo_hi_34 = {dataGroup_27_34, dataGroup_26_34};
  wire [31:0]   res_hi_hi_lo_34 = {res_hi_hi_lo_hi_34, res_hi_hi_lo_lo_34};
  wire [15:0]   res_hi_hi_hi_lo_34 = {dataGroup_29_34, dataGroup_28_34};
  wire [15:0]   res_hi_hi_hi_hi_34 = {dataGroup_31_34, dataGroup_30_34};
  wire [31:0]   res_hi_hi_hi_34 = {res_hi_hi_hi_hi_34, res_hi_hi_hi_lo_34};
  wire [63:0]   res_hi_hi_34 = {res_hi_hi_hi_34, res_hi_hi_lo_34};
  wire [127:0]  res_hi_34 = {res_hi_hi_34, res_hi_lo_34};
  wire [255:0]  res_62 = {res_hi_34, res_lo_34};
  wire [1023:0] dataGroup_lo_1120 = {dataGroup_lo_hi_1120, dataGroup_lo_lo_1120};
  wire [1023:0] dataGroup_hi_1120 = {dataGroup_hi_hi_1120, dataGroup_hi_lo_1120};
  wire [7:0]    dataGroup_0_35 = dataGroup_lo_1120[63:56];
  wire [1023:0] dataGroup_lo_1121 = {dataGroup_lo_hi_1121, dataGroup_lo_lo_1121};
  wire [1023:0] dataGroup_hi_1121 = {dataGroup_hi_hi_1121, dataGroup_hi_lo_1121};
  wire [7:0]    dataGroup_1_35 = dataGroup_lo_1121[127:120];
  wire [1023:0] dataGroup_lo_1122 = {dataGroup_lo_hi_1122, dataGroup_lo_lo_1122};
  wire [1023:0] dataGroup_hi_1122 = {dataGroup_hi_hi_1122, dataGroup_hi_lo_1122};
  wire [7:0]    dataGroup_2_35 = dataGroup_lo_1122[191:184];
  wire [1023:0] dataGroup_lo_1123 = {dataGroup_lo_hi_1123, dataGroup_lo_lo_1123};
  wire [1023:0] dataGroup_hi_1123 = {dataGroup_hi_hi_1123, dataGroup_hi_lo_1123};
  wire [7:0]    dataGroup_3_35 = dataGroup_lo_1123[255:248];
  wire [1023:0] dataGroup_lo_1124 = {dataGroup_lo_hi_1124, dataGroup_lo_lo_1124};
  wire [1023:0] dataGroup_hi_1124 = {dataGroup_hi_hi_1124, dataGroup_hi_lo_1124};
  wire [7:0]    dataGroup_4_35 = dataGroup_lo_1124[319:312];
  wire [1023:0] dataGroup_lo_1125 = {dataGroup_lo_hi_1125, dataGroup_lo_lo_1125};
  wire [1023:0] dataGroup_hi_1125 = {dataGroup_hi_hi_1125, dataGroup_hi_lo_1125};
  wire [7:0]    dataGroup_5_35 = dataGroup_lo_1125[383:376];
  wire [1023:0] dataGroup_lo_1126 = {dataGroup_lo_hi_1126, dataGroup_lo_lo_1126};
  wire [1023:0] dataGroup_hi_1126 = {dataGroup_hi_hi_1126, dataGroup_hi_lo_1126};
  wire [7:0]    dataGroup_6_35 = dataGroup_lo_1126[447:440];
  wire [1023:0] dataGroup_lo_1127 = {dataGroup_lo_hi_1127, dataGroup_lo_lo_1127};
  wire [1023:0] dataGroup_hi_1127 = {dataGroup_hi_hi_1127, dataGroup_hi_lo_1127};
  wire [7:0]    dataGroup_7_35 = dataGroup_lo_1127[511:504];
  wire [1023:0] dataGroup_lo_1128 = {dataGroup_lo_hi_1128, dataGroup_lo_lo_1128};
  wire [1023:0] dataGroup_hi_1128 = {dataGroup_hi_hi_1128, dataGroup_hi_lo_1128};
  wire [7:0]    dataGroup_8_35 = dataGroup_lo_1128[575:568];
  wire [1023:0] dataGroup_lo_1129 = {dataGroup_lo_hi_1129, dataGroup_lo_lo_1129};
  wire [1023:0] dataGroup_hi_1129 = {dataGroup_hi_hi_1129, dataGroup_hi_lo_1129};
  wire [7:0]    dataGroup_9_35 = dataGroup_lo_1129[639:632];
  wire [1023:0] dataGroup_lo_1130 = {dataGroup_lo_hi_1130, dataGroup_lo_lo_1130};
  wire [1023:0] dataGroup_hi_1130 = {dataGroup_hi_hi_1130, dataGroup_hi_lo_1130};
  wire [7:0]    dataGroup_10_35 = dataGroup_lo_1130[703:696];
  wire [1023:0] dataGroup_lo_1131 = {dataGroup_lo_hi_1131, dataGroup_lo_lo_1131};
  wire [1023:0] dataGroup_hi_1131 = {dataGroup_hi_hi_1131, dataGroup_hi_lo_1131};
  wire [7:0]    dataGroup_11_35 = dataGroup_lo_1131[767:760];
  wire [1023:0] dataGroup_lo_1132 = {dataGroup_lo_hi_1132, dataGroup_lo_lo_1132};
  wire [1023:0] dataGroup_hi_1132 = {dataGroup_hi_hi_1132, dataGroup_hi_lo_1132};
  wire [7:0]    dataGroup_12_35 = dataGroup_lo_1132[831:824];
  wire [1023:0] dataGroup_lo_1133 = {dataGroup_lo_hi_1133, dataGroup_lo_lo_1133};
  wire [1023:0] dataGroup_hi_1133 = {dataGroup_hi_hi_1133, dataGroup_hi_lo_1133};
  wire [7:0]    dataGroup_13_35 = dataGroup_lo_1133[895:888];
  wire [1023:0] dataGroup_lo_1134 = {dataGroup_lo_hi_1134, dataGroup_lo_lo_1134};
  wire [1023:0] dataGroup_hi_1134 = {dataGroup_hi_hi_1134, dataGroup_hi_lo_1134};
  wire [7:0]    dataGroup_14_35 = dataGroup_lo_1134[959:952];
  wire [1023:0] dataGroup_lo_1135 = {dataGroup_lo_hi_1135, dataGroup_lo_lo_1135};
  wire [1023:0] dataGroup_hi_1135 = {dataGroup_hi_hi_1135, dataGroup_hi_lo_1135};
  wire [7:0]    dataGroup_15_35 = dataGroup_lo_1135[1023:1016];
  wire [1023:0] dataGroup_lo_1136 = {dataGroup_lo_hi_1136, dataGroup_lo_lo_1136};
  wire [1023:0] dataGroup_hi_1136 = {dataGroup_hi_hi_1136, dataGroup_hi_lo_1136};
  wire [7:0]    dataGroup_16_35 = dataGroup_hi_1136[63:56];
  wire [1023:0] dataGroup_lo_1137 = {dataGroup_lo_hi_1137, dataGroup_lo_lo_1137};
  wire [1023:0] dataGroup_hi_1137 = {dataGroup_hi_hi_1137, dataGroup_hi_lo_1137};
  wire [7:0]    dataGroup_17_35 = dataGroup_hi_1137[127:120];
  wire [1023:0] dataGroup_lo_1138 = {dataGroup_lo_hi_1138, dataGroup_lo_lo_1138};
  wire [1023:0] dataGroup_hi_1138 = {dataGroup_hi_hi_1138, dataGroup_hi_lo_1138};
  wire [7:0]    dataGroup_18_35 = dataGroup_hi_1138[191:184];
  wire [1023:0] dataGroup_lo_1139 = {dataGroup_lo_hi_1139, dataGroup_lo_lo_1139};
  wire [1023:0] dataGroup_hi_1139 = {dataGroup_hi_hi_1139, dataGroup_hi_lo_1139};
  wire [7:0]    dataGroup_19_35 = dataGroup_hi_1139[255:248];
  wire [1023:0] dataGroup_lo_1140 = {dataGroup_lo_hi_1140, dataGroup_lo_lo_1140};
  wire [1023:0] dataGroup_hi_1140 = {dataGroup_hi_hi_1140, dataGroup_hi_lo_1140};
  wire [7:0]    dataGroup_20_35 = dataGroup_hi_1140[319:312];
  wire [1023:0] dataGroup_lo_1141 = {dataGroup_lo_hi_1141, dataGroup_lo_lo_1141};
  wire [1023:0] dataGroup_hi_1141 = {dataGroup_hi_hi_1141, dataGroup_hi_lo_1141};
  wire [7:0]    dataGroup_21_35 = dataGroup_hi_1141[383:376];
  wire [1023:0] dataGroup_lo_1142 = {dataGroup_lo_hi_1142, dataGroup_lo_lo_1142};
  wire [1023:0] dataGroup_hi_1142 = {dataGroup_hi_hi_1142, dataGroup_hi_lo_1142};
  wire [7:0]    dataGroup_22_35 = dataGroup_hi_1142[447:440];
  wire [1023:0] dataGroup_lo_1143 = {dataGroup_lo_hi_1143, dataGroup_lo_lo_1143};
  wire [1023:0] dataGroup_hi_1143 = {dataGroup_hi_hi_1143, dataGroup_hi_lo_1143};
  wire [7:0]    dataGroup_23_35 = dataGroup_hi_1143[511:504];
  wire [1023:0] dataGroup_lo_1144 = {dataGroup_lo_hi_1144, dataGroup_lo_lo_1144};
  wire [1023:0] dataGroup_hi_1144 = {dataGroup_hi_hi_1144, dataGroup_hi_lo_1144};
  wire [7:0]    dataGroup_24_35 = dataGroup_hi_1144[575:568];
  wire [1023:0] dataGroup_lo_1145 = {dataGroup_lo_hi_1145, dataGroup_lo_lo_1145};
  wire [1023:0] dataGroup_hi_1145 = {dataGroup_hi_hi_1145, dataGroup_hi_lo_1145};
  wire [7:0]    dataGroup_25_35 = dataGroup_hi_1145[639:632];
  wire [1023:0] dataGroup_lo_1146 = {dataGroup_lo_hi_1146, dataGroup_lo_lo_1146};
  wire [1023:0] dataGroup_hi_1146 = {dataGroup_hi_hi_1146, dataGroup_hi_lo_1146};
  wire [7:0]    dataGroup_26_35 = dataGroup_hi_1146[703:696];
  wire [1023:0] dataGroup_lo_1147 = {dataGroup_lo_hi_1147, dataGroup_lo_lo_1147};
  wire [1023:0] dataGroup_hi_1147 = {dataGroup_hi_hi_1147, dataGroup_hi_lo_1147};
  wire [7:0]    dataGroup_27_35 = dataGroup_hi_1147[767:760];
  wire [1023:0] dataGroup_lo_1148 = {dataGroup_lo_hi_1148, dataGroup_lo_lo_1148};
  wire [1023:0] dataGroup_hi_1148 = {dataGroup_hi_hi_1148, dataGroup_hi_lo_1148};
  wire [7:0]    dataGroup_28_35 = dataGroup_hi_1148[831:824];
  wire [1023:0] dataGroup_lo_1149 = {dataGroup_lo_hi_1149, dataGroup_lo_lo_1149};
  wire [1023:0] dataGroup_hi_1149 = {dataGroup_hi_hi_1149, dataGroup_hi_lo_1149};
  wire [7:0]    dataGroup_29_35 = dataGroup_hi_1149[895:888];
  wire [1023:0] dataGroup_lo_1150 = {dataGroup_lo_hi_1150, dataGroup_lo_lo_1150};
  wire [1023:0] dataGroup_hi_1150 = {dataGroup_hi_hi_1150, dataGroup_hi_lo_1150};
  wire [7:0]    dataGroup_30_35 = dataGroup_hi_1150[959:952];
  wire [1023:0] dataGroup_lo_1151 = {dataGroup_lo_hi_1151, dataGroup_lo_lo_1151};
  wire [1023:0] dataGroup_hi_1151 = {dataGroup_hi_hi_1151, dataGroup_hi_lo_1151};
  wire [7:0]    dataGroup_31_35 = dataGroup_hi_1151[1023:1016];
  wire [15:0]   res_lo_lo_lo_lo_35 = {dataGroup_1_35, dataGroup_0_35};
  wire [15:0]   res_lo_lo_lo_hi_35 = {dataGroup_3_35, dataGroup_2_35};
  wire [31:0]   res_lo_lo_lo_35 = {res_lo_lo_lo_hi_35, res_lo_lo_lo_lo_35};
  wire [15:0]   res_lo_lo_hi_lo_35 = {dataGroup_5_35, dataGroup_4_35};
  wire [15:0]   res_lo_lo_hi_hi_35 = {dataGroup_7_35, dataGroup_6_35};
  wire [31:0]   res_lo_lo_hi_35 = {res_lo_lo_hi_hi_35, res_lo_lo_hi_lo_35};
  wire [63:0]   res_lo_lo_35 = {res_lo_lo_hi_35, res_lo_lo_lo_35};
  wire [15:0]   res_lo_hi_lo_lo_35 = {dataGroup_9_35, dataGroup_8_35};
  wire [15:0]   res_lo_hi_lo_hi_35 = {dataGroup_11_35, dataGroup_10_35};
  wire [31:0]   res_lo_hi_lo_35 = {res_lo_hi_lo_hi_35, res_lo_hi_lo_lo_35};
  wire [15:0]   res_lo_hi_hi_lo_35 = {dataGroup_13_35, dataGroup_12_35};
  wire [15:0]   res_lo_hi_hi_hi_35 = {dataGroup_15_35, dataGroup_14_35};
  wire [31:0]   res_lo_hi_hi_35 = {res_lo_hi_hi_hi_35, res_lo_hi_hi_lo_35};
  wire [63:0]   res_lo_hi_35 = {res_lo_hi_hi_35, res_lo_hi_lo_35};
  wire [127:0]  res_lo_35 = {res_lo_hi_35, res_lo_lo_35};
  wire [15:0]   res_hi_lo_lo_lo_35 = {dataGroup_17_35, dataGroup_16_35};
  wire [15:0]   res_hi_lo_lo_hi_35 = {dataGroup_19_35, dataGroup_18_35};
  wire [31:0]   res_hi_lo_lo_35 = {res_hi_lo_lo_hi_35, res_hi_lo_lo_lo_35};
  wire [15:0]   res_hi_lo_hi_lo_35 = {dataGroup_21_35, dataGroup_20_35};
  wire [15:0]   res_hi_lo_hi_hi_35 = {dataGroup_23_35, dataGroup_22_35};
  wire [31:0]   res_hi_lo_hi_35 = {res_hi_lo_hi_hi_35, res_hi_lo_hi_lo_35};
  wire [63:0]   res_hi_lo_35 = {res_hi_lo_hi_35, res_hi_lo_lo_35};
  wire [15:0]   res_hi_hi_lo_lo_35 = {dataGroup_25_35, dataGroup_24_35};
  wire [15:0]   res_hi_hi_lo_hi_35 = {dataGroup_27_35, dataGroup_26_35};
  wire [31:0]   res_hi_hi_lo_35 = {res_hi_hi_lo_hi_35, res_hi_hi_lo_lo_35};
  wire [15:0]   res_hi_hi_hi_lo_35 = {dataGroup_29_35, dataGroup_28_35};
  wire [15:0]   res_hi_hi_hi_hi_35 = {dataGroup_31_35, dataGroup_30_35};
  wire [31:0]   res_hi_hi_hi_35 = {res_hi_hi_hi_hi_35, res_hi_hi_hi_lo_35};
  wire [63:0]   res_hi_hi_35 = {res_hi_hi_hi_35, res_hi_hi_lo_35};
  wire [127:0]  res_hi_35 = {res_hi_hi_35, res_hi_lo_35};
  wire [255:0]  res_63 = {res_hi_35, res_lo_35};
  wire [511:0]  lo_lo_7 = {res_57, res_56};
  wire [511:0]  lo_hi_7 = {res_59, res_58};
  wire [1023:0] lo_7 = {lo_hi_7, lo_lo_7};
  wire [511:0]  hi_lo_7 = {res_61, res_60};
  wire [511:0]  hi_hi_7 = {res_63, res_62};
  wire [1023:0] hi_7 = {hi_hi_7, hi_lo_7};
  wire [2047:0] regroupLoadData_0_7 = {hi_7, lo_7};
  wire [1023:0] dataGroup_lo_1152 = {dataGroup_lo_hi_1152, dataGroup_lo_lo_1152};
  wire [1023:0] dataGroup_hi_1152 = {dataGroup_hi_hi_1152, dataGroup_hi_lo_1152};
  wire [15:0]   dataGroup_0_36 = dataGroup_lo_1152[15:0];
  wire [1023:0] dataGroup_lo_1153 = {dataGroup_lo_hi_1153, dataGroup_lo_lo_1153};
  wire [1023:0] dataGroup_hi_1153 = {dataGroup_hi_hi_1153, dataGroup_hi_lo_1153};
  wire [15:0]   dataGroup_1_36 = dataGroup_lo_1153[31:16];
  wire [1023:0] dataGroup_lo_1154 = {dataGroup_lo_hi_1154, dataGroup_lo_lo_1154};
  wire [1023:0] dataGroup_hi_1154 = {dataGroup_hi_hi_1154, dataGroup_hi_lo_1154};
  wire [15:0]   dataGroup_2_36 = dataGroup_lo_1154[47:32];
  wire [1023:0] dataGroup_lo_1155 = {dataGroup_lo_hi_1155, dataGroup_lo_lo_1155};
  wire [1023:0] dataGroup_hi_1155 = {dataGroup_hi_hi_1155, dataGroup_hi_lo_1155};
  wire [15:0]   dataGroup_3_36 = dataGroup_lo_1155[63:48];
  wire [1023:0] dataGroup_lo_1156 = {dataGroup_lo_hi_1156, dataGroup_lo_lo_1156};
  wire [1023:0] dataGroup_hi_1156 = {dataGroup_hi_hi_1156, dataGroup_hi_lo_1156};
  wire [15:0]   dataGroup_4_36 = dataGroup_lo_1156[79:64];
  wire [1023:0] dataGroup_lo_1157 = {dataGroup_lo_hi_1157, dataGroup_lo_lo_1157};
  wire [1023:0] dataGroup_hi_1157 = {dataGroup_hi_hi_1157, dataGroup_hi_lo_1157};
  wire [15:0]   dataGroup_5_36 = dataGroup_lo_1157[95:80];
  wire [1023:0] dataGroup_lo_1158 = {dataGroup_lo_hi_1158, dataGroup_lo_lo_1158};
  wire [1023:0] dataGroup_hi_1158 = {dataGroup_hi_hi_1158, dataGroup_hi_lo_1158};
  wire [15:0]   dataGroup_6_36 = dataGroup_lo_1158[111:96];
  wire [1023:0] dataGroup_lo_1159 = {dataGroup_lo_hi_1159, dataGroup_lo_lo_1159};
  wire [1023:0] dataGroup_hi_1159 = {dataGroup_hi_hi_1159, dataGroup_hi_lo_1159};
  wire [15:0]   dataGroup_7_36 = dataGroup_lo_1159[127:112];
  wire [1023:0] dataGroup_lo_1160 = {dataGroup_lo_hi_1160, dataGroup_lo_lo_1160};
  wire [1023:0] dataGroup_hi_1160 = {dataGroup_hi_hi_1160, dataGroup_hi_lo_1160};
  wire [15:0]   dataGroup_8_36 = dataGroup_lo_1160[143:128];
  wire [1023:0] dataGroup_lo_1161 = {dataGroup_lo_hi_1161, dataGroup_lo_lo_1161};
  wire [1023:0] dataGroup_hi_1161 = {dataGroup_hi_hi_1161, dataGroup_hi_lo_1161};
  wire [15:0]   dataGroup_9_36 = dataGroup_lo_1161[159:144];
  wire [1023:0] dataGroup_lo_1162 = {dataGroup_lo_hi_1162, dataGroup_lo_lo_1162};
  wire [1023:0] dataGroup_hi_1162 = {dataGroup_hi_hi_1162, dataGroup_hi_lo_1162};
  wire [15:0]   dataGroup_10_36 = dataGroup_lo_1162[175:160];
  wire [1023:0] dataGroup_lo_1163 = {dataGroup_lo_hi_1163, dataGroup_lo_lo_1163};
  wire [1023:0] dataGroup_hi_1163 = {dataGroup_hi_hi_1163, dataGroup_hi_lo_1163};
  wire [15:0]   dataGroup_11_36 = dataGroup_lo_1163[191:176];
  wire [1023:0] dataGroup_lo_1164 = {dataGroup_lo_hi_1164, dataGroup_lo_lo_1164};
  wire [1023:0] dataGroup_hi_1164 = {dataGroup_hi_hi_1164, dataGroup_hi_lo_1164};
  wire [15:0]   dataGroup_12_36 = dataGroup_lo_1164[207:192];
  wire [1023:0] dataGroup_lo_1165 = {dataGroup_lo_hi_1165, dataGroup_lo_lo_1165};
  wire [1023:0] dataGroup_hi_1165 = {dataGroup_hi_hi_1165, dataGroup_hi_lo_1165};
  wire [15:0]   dataGroup_13_36 = dataGroup_lo_1165[223:208];
  wire [1023:0] dataGroup_lo_1166 = {dataGroup_lo_hi_1166, dataGroup_lo_lo_1166};
  wire [1023:0] dataGroup_hi_1166 = {dataGroup_hi_hi_1166, dataGroup_hi_lo_1166};
  wire [15:0]   dataGroup_14_36 = dataGroup_lo_1166[239:224];
  wire [1023:0] dataGroup_lo_1167 = {dataGroup_lo_hi_1167, dataGroup_lo_lo_1167};
  wire [1023:0] dataGroup_hi_1167 = {dataGroup_hi_hi_1167, dataGroup_hi_lo_1167};
  wire [15:0]   dataGroup_15_36 = dataGroup_lo_1167[255:240];
  wire [31:0]   res_lo_lo_lo_36 = {dataGroup_1_36, dataGroup_0_36};
  wire [31:0]   res_lo_lo_hi_36 = {dataGroup_3_36, dataGroup_2_36};
  wire [63:0]   res_lo_lo_36 = {res_lo_lo_hi_36, res_lo_lo_lo_36};
  wire [31:0]   res_lo_hi_lo_36 = {dataGroup_5_36, dataGroup_4_36};
  wire [31:0]   res_lo_hi_hi_36 = {dataGroup_7_36, dataGroup_6_36};
  wire [63:0]   res_lo_hi_36 = {res_lo_hi_hi_36, res_lo_hi_lo_36};
  wire [127:0]  res_lo_36 = {res_lo_hi_36, res_lo_lo_36};
  wire [31:0]   res_hi_lo_lo_36 = {dataGroup_9_36, dataGroup_8_36};
  wire [31:0]   res_hi_lo_hi_36 = {dataGroup_11_36, dataGroup_10_36};
  wire [63:0]   res_hi_lo_36 = {res_hi_lo_hi_36, res_hi_lo_lo_36};
  wire [31:0]   res_hi_hi_lo_36 = {dataGroup_13_36, dataGroup_12_36};
  wire [31:0]   res_hi_hi_hi_36 = {dataGroup_15_36, dataGroup_14_36};
  wire [63:0]   res_hi_hi_36 = {res_hi_hi_hi_36, res_hi_hi_lo_36};
  wire [127:0]  res_hi_36 = {res_hi_hi_36, res_hi_lo_36};
  wire [255:0]  res_64 = {res_hi_36, res_lo_36};
  wire [511:0]  lo_lo_8 = {256'h0, res_64};
  wire [1023:0] lo_8 = {512'h0, lo_lo_8};
  wire [2047:0] regroupLoadData_1_0 = {1024'h0, lo_8};
  wire [1023:0] dataGroup_lo_1168 = {dataGroup_lo_hi_1168, dataGroup_lo_lo_1168};
  wire [1023:0] dataGroup_hi_1168 = {dataGroup_hi_hi_1168, dataGroup_hi_lo_1168};
  wire [15:0]   dataGroup_0_37 = dataGroup_lo_1168[15:0];
  wire [1023:0] dataGroup_lo_1169 = {dataGroup_lo_hi_1169, dataGroup_lo_lo_1169};
  wire [1023:0] dataGroup_hi_1169 = {dataGroup_hi_hi_1169, dataGroup_hi_lo_1169};
  wire [15:0]   dataGroup_1_37 = dataGroup_lo_1169[47:32];
  wire [1023:0] dataGroup_lo_1170 = {dataGroup_lo_hi_1170, dataGroup_lo_lo_1170};
  wire [1023:0] dataGroup_hi_1170 = {dataGroup_hi_hi_1170, dataGroup_hi_lo_1170};
  wire [15:0]   dataGroup_2_37 = dataGroup_lo_1170[79:64];
  wire [1023:0] dataGroup_lo_1171 = {dataGroup_lo_hi_1171, dataGroup_lo_lo_1171};
  wire [1023:0] dataGroup_hi_1171 = {dataGroup_hi_hi_1171, dataGroup_hi_lo_1171};
  wire [15:0]   dataGroup_3_37 = dataGroup_lo_1171[111:96];
  wire [1023:0] dataGroup_lo_1172 = {dataGroup_lo_hi_1172, dataGroup_lo_lo_1172};
  wire [1023:0] dataGroup_hi_1172 = {dataGroup_hi_hi_1172, dataGroup_hi_lo_1172};
  wire [15:0]   dataGroup_4_37 = dataGroup_lo_1172[143:128];
  wire [1023:0] dataGroup_lo_1173 = {dataGroup_lo_hi_1173, dataGroup_lo_lo_1173};
  wire [1023:0] dataGroup_hi_1173 = {dataGroup_hi_hi_1173, dataGroup_hi_lo_1173};
  wire [15:0]   dataGroup_5_37 = dataGroup_lo_1173[175:160];
  wire [1023:0] dataGroup_lo_1174 = {dataGroup_lo_hi_1174, dataGroup_lo_lo_1174};
  wire [1023:0] dataGroup_hi_1174 = {dataGroup_hi_hi_1174, dataGroup_hi_lo_1174};
  wire [15:0]   dataGroup_6_37 = dataGroup_lo_1174[207:192];
  wire [1023:0] dataGroup_lo_1175 = {dataGroup_lo_hi_1175, dataGroup_lo_lo_1175};
  wire [1023:0] dataGroup_hi_1175 = {dataGroup_hi_hi_1175, dataGroup_hi_lo_1175};
  wire [15:0]   dataGroup_7_37 = dataGroup_lo_1175[239:224];
  wire [1023:0] dataGroup_lo_1176 = {dataGroup_lo_hi_1176, dataGroup_lo_lo_1176};
  wire [1023:0] dataGroup_hi_1176 = {dataGroup_hi_hi_1176, dataGroup_hi_lo_1176};
  wire [15:0]   dataGroup_8_37 = dataGroup_lo_1176[271:256];
  wire [1023:0] dataGroup_lo_1177 = {dataGroup_lo_hi_1177, dataGroup_lo_lo_1177};
  wire [1023:0] dataGroup_hi_1177 = {dataGroup_hi_hi_1177, dataGroup_hi_lo_1177};
  wire [15:0]   dataGroup_9_37 = dataGroup_lo_1177[303:288];
  wire [1023:0] dataGroup_lo_1178 = {dataGroup_lo_hi_1178, dataGroup_lo_lo_1178};
  wire [1023:0] dataGroup_hi_1178 = {dataGroup_hi_hi_1178, dataGroup_hi_lo_1178};
  wire [15:0]   dataGroup_10_37 = dataGroup_lo_1178[335:320];
  wire [1023:0] dataGroup_lo_1179 = {dataGroup_lo_hi_1179, dataGroup_lo_lo_1179};
  wire [1023:0] dataGroup_hi_1179 = {dataGroup_hi_hi_1179, dataGroup_hi_lo_1179};
  wire [15:0]   dataGroup_11_37 = dataGroup_lo_1179[367:352];
  wire [1023:0] dataGroup_lo_1180 = {dataGroup_lo_hi_1180, dataGroup_lo_lo_1180};
  wire [1023:0] dataGroup_hi_1180 = {dataGroup_hi_hi_1180, dataGroup_hi_lo_1180};
  wire [15:0]   dataGroup_12_37 = dataGroup_lo_1180[399:384];
  wire [1023:0] dataGroup_lo_1181 = {dataGroup_lo_hi_1181, dataGroup_lo_lo_1181};
  wire [1023:0] dataGroup_hi_1181 = {dataGroup_hi_hi_1181, dataGroup_hi_lo_1181};
  wire [15:0]   dataGroup_13_37 = dataGroup_lo_1181[431:416];
  wire [1023:0] dataGroup_lo_1182 = {dataGroup_lo_hi_1182, dataGroup_lo_lo_1182};
  wire [1023:0] dataGroup_hi_1182 = {dataGroup_hi_hi_1182, dataGroup_hi_lo_1182};
  wire [15:0]   dataGroup_14_37 = dataGroup_lo_1182[463:448];
  wire [1023:0] dataGroup_lo_1183 = {dataGroup_lo_hi_1183, dataGroup_lo_lo_1183};
  wire [1023:0] dataGroup_hi_1183 = {dataGroup_hi_hi_1183, dataGroup_hi_lo_1183};
  wire [15:0]   dataGroup_15_37 = dataGroup_lo_1183[495:480];
  wire [31:0]   res_lo_lo_lo_37 = {dataGroup_1_37, dataGroup_0_37};
  wire [31:0]   res_lo_lo_hi_37 = {dataGroup_3_37, dataGroup_2_37};
  wire [63:0]   res_lo_lo_37 = {res_lo_lo_hi_37, res_lo_lo_lo_37};
  wire [31:0]   res_lo_hi_lo_37 = {dataGroup_5_37, dataGroup_4_37};
  wire [31:0]   res_lo_hi_hi_37 = {dataGroup_7_37, dataGroup_6_37};
  wire [63:0]   res_lo_hi_37 = {res_lo_hi_hi_37, res_lo_hi_lo_37};
  wire [127:0]  res_lo_37 = {res_lo_hi_37, res_lo_lo_37};
  wire [31:0]   res_hi_lo_lo_37 = {dataGroup_9_37, dataGroup_8_37};
  wire [31:0]   res_hi_lo_hi_37 = {dataGroup_11_37, dataGroup_10_37};
  wire [63:0]   res_hi_lo_37 = {res_hi_lo_hi_37, res_hi_lo_lo_37};
  wire [31:0]   res_hi_hi_lo_37 = {dataGroup_13_37, dataGroup_12_37};
  wire [31:0]   res_hi_hi_hi_37 = {dataGroup_15_37, dataGroup_14_37};
  wire [63:0]   res_hi_hi_37 = {res_hi_hi_hi_37, res_hi_hi_lo_37};
  wire [127:0]  res_hi_37 = {res_hi_hi_37, res_hi_lo_37};
  wire [255:0]  res_72 = {res_hi_37, res_lo_37};
  wire [1023:0] dataGroup_lo_1184 = {dataGroup_lo_hi_1184, dataGroup_lo_lo_1184};
  wire [1023:0] dataGroup_hi_1184 = {dataGroup_hi_hi_1184, dataGroup_hi_lo_1184};
  wire [15:0]   dataGroup_0_38 = dataGroup_lo_1184[31:16];
  wire [1023:0] dataGroup_lo_1185 = {dataGroup_lo_hi_1185, dataGroup_lo_lo_1185};
  wire [1023:0] dataGroup_hi_1185 = {dataGroup_hi_hi_1185, dataGroup_hi_lo_1185};
  wire [15:0]   dataGroup_1_38 = dataGroup_lo_1185[63:48];
  wire [1023:0] dataGroup_lo_1186 = {dataGroup_lo_hi_1186, dataGroup_lo_lo_1186};
  wire [1023:0] dataGroup_hi_1186 = {dataGroup_hi_hi_1186, dataGroup_hi_lo_1186};
  wire [15:0]   dataGroup_2_38 = dataGroup_lo_1186[95:80];
  wire [1023:0] dataGroup_lo_1187 = {dataGroup_lo_hi_1187, dataGroup_lo_lo_1187};
  wire [1023:0] dataGroup_hi_1187 = {dataGroup_hi_hi_1187, dataGroup_hi_lo_1187};
  wire [15:0]   dataGroup_3_38 = dataGroup_lo_1187[127:112];
  wire [1023:0] dataGroup_lo_1188 = {dataGroup_lo_hi_1188, dataGroup_lo_lo_1188};
  wire [1023:0] dataGroup_hi_1188 = {dataGroup_hi_hi_1188, dataGroup_hi_lo_1188};
  wire [15:0]   dataGroup_4_38 = dataGroup_lo_1188[159:144];
  wire [1023:0] dataGroup_lo_1189 = {dataGroup_lo_hi_1189, dataGroup_lo_lo_1189};
  wire [1023:0] dataGroup_hi_1189 = {dataGroup_hi_hi_1189, dataGroup_hi_lo_1189};
  wire [15:0]   dataGroup_5_38 = dataGroup_lo_1189[191:176];
  wire [1023:0] dataGroup_lo_1190 = {dataGroup_lo_hi_1190, dataGroup_lo_lo_1190};
  wire [1023:0] dataGroup_hi_1190 = {dataGroup_hi_hi_1190, dataGroup_hi_lo_1190};
  wire [15:0]   dataGroup_6_38 = dataGroup_lo_1190[223:208];
  wire [1023:0] dataGroup_lo_1191 = {dataGroup_lo_hi_1191, dataGroup_lo_lo_1191};
  wire [1023:0] dataGroup_hi_1191 = {dataGroup_hi_hi_1191, dataGroup_hi_lo_1191};
  wire [15:0]   dataGroup_7_38 = dataGroup_lo_1191[255:240];
  wire [1023:0] dataGroup_lo_1192 = {dataGroup_lo_hi_1192, dataGroup_lo_lo_1192};
  wire [1023:0] dataGroup_hi_1192 = {dataGroup_hi_hi_1192, dataGroup_hi_lo_1192};
  wire [15:0]   dataGroup_8_38 = dataGroup_lo_1192[287:272];
  wire [1023:0] dataGroup_lo_1193 = {dataGroup_lo_hi_1193, dataGroup_lo_lo_1193};
  wire [1023:0] dataGroup_hi_1193 = {dataGroup_hi_hi_1193, dataGroup_hi_lo_1193};
  wire [15:0]   dataGroup_9_38 = dataGroup_lo_1193[319:304];
  wire [1023:0] dataGroup_lo_1194 = {dataGroup_lo_hi_1194, dataGroup_lo_lo_1194};
  wire [1023:0] dataGroup_hi_1194 = {dataGroup_hi_hi_1194, dataGroup_hi_lo_1194};
  wire [15:0]   dataGroup_10_38 = dataGroup_lo_1194[351:336];
  wire [1023:0] dataGroup_lo_1195 = {dataGroup_lo_hi_1195, dataGroup_lo_lo_1195};
  wire [1023:0] dataGroup_hi_1195 = {dataGroup_hi_hi_1195, dataGroup_hi_lo_1195};
  wire [15:0]   dataGroup_11_38 = dataGroup_lo_1195[383:368];
  wire [1023:0] dataGroup_lo_1196 = {dataGroup_lo_hi_1196, dataGroup_lo_lo_1196};
  wire [1023:0] dataGroup_hi_1196 = {dataGroup_hi_hi_1196, dataGroup_hi_lo_1196};
  wire [15:0]   dataGroup_12_38 = dataGroup_lo_1196[415:400];
  wire [1023:0] dataGroup_lo_1197 = {dataGroup_lo_hi_1197, dataGroup_lo_lo_1197};
  wire [1023:0] dataGroup_hi_1197 = {dataGroup_hi_hi_1197, dataGroup_hi_lo_1197};
  wire [15:0]   dataGroup_13_38 = dataGroup_lo_1197[447:432];
  wire [1023:0] dataGroup_lo_1198 = {dataGroup_lo_hi_1198, dataGroup_lo_lo_1198};
  wire [1023:0] dataGroup_hi_1198 = {dataGroup_hi_hi_1198, dataGroup_hi_lo_1198};
  wire [15:0]   dataGroup_14_38 = dataGroup_lo_1198[479:464];
  wire [1023:0] dataGroup_lo_1199 = {dataGroup_lo_hi_1199, dataGroup_lo_lo_1199};
  wire [1023:0] dataGroup_hi_1199 = {dataGroup_hi_hi_1199, dataGroup_hi_lo_1199};
  wire [15:0]   dataGroup_15_38 = dataGroup_lo_1199[511:496];
  wire [31:0]   res_lo_lo_lo_38 = {dataGroup_1_38, dataGroup_0_38};
  wire [31:0]   res_lo_lo_hi_38 = {dataGroup_3_38, dataGroup_2_38};
  wire [63:0]   res_lo_lo_38 = {res_lo_lo_hi_38, res_lo_lo_lo_38};
  wire [31:0]   res_lo_hi_lo_38 = {dataGroup_5_38, dataGroup_4_38};
  wire [31:0]   res_lo_hi_hi_38 = {dataGroup_7_38, dataGroup_6_38};
  wire [63:0]   res_lo_hi_38 = {res_lo_hi_hi_38, res_lo_hi_lo_38};
  wire [127:0]  res_lo_38 = {res_lo_hi_38, res_lo_lo_38};
  wire [31:0]   res_hi_lo_lo_38 = {dataGroup_9_38, dataGroup_8_38};
  wire [31:0]   res_hi_lo_hi_38 = {dataGroup_11_38, dataGroup_10_38};
  wire [63:0]   res_hi_lo_38 = {res_hi_lo_hi_38, res_hi_lo_lo_38};
  wire [31:0]   res_hi_hi_lo_38 = {dataGroup_13_38, dataGroup_12_38};
  wire [31:0]   res_hi_hi_hi_38 = {dataGroup_15_38, dataGroup_14_38};
  wire [63:0]   res_hi_hi_38 = {res_hi_hi_hi_38, res_hi_hi_lo_38};
  wire [127:0]  res_hi_38 = {res_hi_hi_38, res_hi_lo_38};
  wire [255:0]  res_73 = {res_hi_38, res_lo_38};
  wire [511:0]  lo_lo_9 = {res_73, res_72};
  wire [1023:0] lo_9 = {512'h0, lo_lo_9};
  wire [2047:0] regroupLoadData_1_1 = {1024'h0, lo_9};
  wire [1023:0] dataGroup_lo_1200 = {dataGroup_lo_hi_1200, dataGroup_lo_lo_1200};
  wire [1023:0] dataGroup_hi_1200 = {dataGroup_hi_hi_1200, dataGroup_hi_lo_1200};
  wire [15:0]   dataGroup_0_39 = dataGroup_lo_1200[15:0];
  wire [1023:0] dataGroup_lo_1201 = {dataGroup_lo_hi_1201, dataGroup_lo_lo_1201};
  wire [1023:0] dataGroup_hi_1201 = {dataGroup_hi_hi_1201, dataGroup_hi_lo_1201};
  wire [15:0]   dataGroup_1_39 = dataGroup_lo_1201[63:48];
  wire [1023:0] dataGroup_lo_1202 = {dataGroup_lo_hi_1202, dataGroup_lo_lo_1202};
  wire [1023:0] dataGroup_hi_1202 = {dataGroup_hi_hi_1202, dataGroup_hi_lo_1202};
  wire [15:0]   dataGroup_2_39 = dataGroup_lo_1202[111:96];
  wire [1023:0] dataGroup_lo_1203 = {dataGroup_lo_hi_1203, dataGroup_lo_lo_1203};
  wire [1023:0] dataGroup_hi_1203 = {dataGroup_hi_hi_1203, dataGroup_hi_lo_1203};
  wire [15:0]   dataGroup_3_39 = dataGroup_lo_1203[159:144];
  wire [1023:0] dataGroup_lo_1204 = {dataGroup_lo_hi_1204, dataGroup_lo_lo_1204};
  wire [1023:0] dataGroup_hi_1204 = {dataGroup_hi_hi_1204, dataGroup_hi_lo_1204};
  wire [15:0]   dataGroup_4_39 = dataGroup_lo_1204[207:192];
  wire [1023:0] dataGroup_lo_1205 = {dataGroup_lo_hi_1205, dataGroup_lo_lo_1205};
  wire [1023:0] dataGroup_hi_1205 = {dataGroup_hi_hi_1205, dataGroup_hi_lo_1205};
  wire [15:0]   dataGroup_5_39 = dataGroup_lo_1205[255:240];
  wire [1023:0] dataGroup_lo_1206 = {dataGroup_lo_hi_1206, dataGroup_lo_lo_1206};
  wire [1023:0] dataGroup_hi_1206 = {dataGroup_hi_hi_1206, dataGroup_hi_lo_1206};
  wire [15:0]   dataGroup_6_39 = dataGroup_lo_1206[303:288];
  wire [1023:0] dataGroup_lo_1207 = {dataGroup_lo_hi_1207, dataGroup_lo_lo_1207};
  wire [1023:0] dataGroup_hi_1207 = {dataGroup_hi_hi_1207, dataGroup_hi_lo_1207};
  wire [15:0]   dataGroup_7_39 = dataGroup_lo_1207[351:336];
  wire [1023:0] dataGroup_lo_1208 = {dataGroup_lo_hi_1208, dataGroup_lo_lo_1208};
  wire [1023:0] dataGroup_hi_1208 = {dataGroup_hi_hi_1208, dataGroup_hi_lo_1208};
  wire [15:0]   dataGroup_8_39 = dataGroup_lo_1208[399:384];
  wire [1023:0] dataGroup_lo_1209 = {dataGroup_lo_hi_1209, dataGroup_lo_lo_1209};
  wire [1023:0] dataGroup_hi_1209 = {dataGroup_hi_hi_1209, dataGroup_hi_lo_1209};
  wire [15:0]   dataGroup_9_39 = dataGroup_lo_1209[447:432];
  wire [1023:0] dataGroup_lo_1210 = {dataGroup_lo_hi_1210, dataGroup_lo_lo_1210};
  wire [1023:0] dataGroup_hi_1210 = {dataGroup_hi_hi_1210, dataGroup_hi_lo_1210};
  wire [15:0]   dataGroup_10_39 = dataGroup_lo_1210[495:480];
  wire [1023:0] dataGroup_lo_1211 = {dataGroup_lo_hi_1211, dataGroup_lo_lo_1211};
  wire [1023:0] dataGroup_hi_1211 = {dataGroup_hi_hi_1211, dataGroup_hi_lo_1211};
  wire [15:0]   dataGroup_11_39 = dataGroup_lo_1211[543:528];
  wire [1023:0] dataGroup_lo_1212 = {dataGroup_lo_hi_1212, dataGroup_lo_lo_1212};
  wire [1023:0] dataGroup_hi_1212 = {dataGroup_hi_hi_1212, dataGroup_hi_lo_1212};
  wire [15:0]   dataGroup_12_39 = dataGroup_lo_1212[591:576];
  wire [1023:0] dataGroup_lo_1213 = {dataGroup_lo_hi_1213, dataGroup_lo_lo_1213};
  wire [1023:0] dataGroup_hi_1213 = {dataGroup_hi_hi_1213, dataGroup_hi_lo_1213};
  wire [15:0]   dataGroup_13_39 = dataGroup_lo_1213[639:624];
  wire [1023:0] dataGroup_lo_1214 = {dataGroup_lo_hi_1214, dataGroup_lo_lo_1214};
  wire [1023:0] dataGroup_hi_1214 = {dataGroup_hi_hi_1214, dataGroup_hi_lo_1214};
  wire [15:0]   dataGroup_14_39 = dataGroup_lo_1214[687:672];
  wire [1023:0] dataGroup_lo_1215 = {dataGroup_lo_hi_1215, dataGroup_lo_lo_1215};
  wire [1023:0] dataGroup_hi_1215 = {dataGroup_hi_hi_1215, dataGroup_hi_lo_1215};
  wire [15:0]   dataGroup_15_39 = dataGroup_lo_1215[735:720];
  wire [31:0]   res_lo_lo_lo_39 = {dataGroup_1_39, dataGroup_0_39};
  wire [31:0]   res_lo_lo_hi_39 = {dataGroup_3_39, dataGroup_2_39};
  wire [63:0]   res_lo_lo_39 = {res_lo_lo_hi_39, res_lo_lo_lo_39};
  wire [31:0]   res_lo_hi_lo_39 = {dataGroup_5_39, dataGroup_4_39};
  wire [31:0]   res_lo_hi_hi_39 = {dataGroup_7_39, dataGroup_6_39};
  wire [63:0]   res_lo_hi_39 = {res_lo_hi_hi_39, res_lo_hi_lo_39};
  wire [127:0]  res_lo_39 = {res_lo_hi_39, res_lo_lo_39};
  wire [31:0]   res_hi_lo_lo_39 = {dataGroup_9_39, dataGroup_8_39};
  wire [31:0]   res_hi_lo_hi_39 = {dataGroup_11_39, dataGroup_10_39};
  wire [63:0]   res_hi_lo_39 = {res_hi_lo_hi_39, res_hi_lo_lo_39};
  wire [31:0]   res_hi_hi_lo_39 = {dataGroup_13_39, dataGroup_12_39};
  wire [31:0]   res_hi_hi_hi_39 = {dataGroup_15_39, dataGroup_14_39};
  wire [63:0]   res_hi_hi_39 = {res_hi_hi_hi_39, res_hi_hi_lo_39};
  wire [127:0]  res_hi_39 = {res_hi_hi_39, res_hi_lo_39};
  wire [255:0]  res_80 = {res_hi_39, res_lo_39};
  wire [1023:0] dataGroup_lo_1216 = {dataGroup_lo_hi_1216, dataGroup_lo_lo_1216};
  wire [1023:0] dataGroup_hi_1216 = {dataGroup_hi_hi_1216, dataGroup_hi_lo_1216};
  wire [15:0]   dataGroup_0_40 = dataGroup_lo_1216[31:16];
  wire [1023:0] dataGroup_lo_1217 = {dataGroup_lo_hi_1217, dataGroup_lo_lo_1217};
  wire [1023:0] dataGroup_hi_1217 = {dataGroup_hi_hi_1217, dataGroup_hi_lo_1217};
  wire [15:0]   dataGroup_1_40 = dataGroup_lo_1217[79:64];
  wire [1023:0] dataGroup_lo_1218 = {dataGroup_lo_hi_1218, dataGroup_lo_lo_1218};
  wire [1023:0] dataGroup_hi_1218 = {dataGroup_hi_hi_1218, dataGroup_hi_lo_1218};
  wire [15:0]   dataGroup_2_40 = dataGroup_lo_1218[127:112];
  wire [1023:0] dataGroup_lo_1219 = {dataGroup_lo_hi_1219, dataGroup_lo_lo_1219};
  wire [1023:0] dataGroup_hi_1219 = {dataGroup_hi_hi_1219, dataGroup_hi_lo_1219};
  wire [15:0]   dataGroup_3_40 = dataGroup_lo_1219[175:160];
  wire [1023:0] dataGroup_lo_1220 = {dataGroup_lo_hi_1220, dataGroup_lo_lo_1220};
  wire [1023:0] dataGroup_hi_1220 = {dataGroup_hi_hi_1220, dataGroup_hi_lo_1220};
  wire [15:0]   dataGroup_4_40 = dataGroup_lo_1220[223:208];
  wire [1023:0] dataGroup_lo_1221 = {dataGroup_lo_hi_1221, dataGroup_lo_lo_1221};
  wire [1023:0] dataGroup_hi_1221 = {dataGroup_hi_hi_1221, dataGroup_hi_lo_1221};
  wire [15:0]   dataGroup_5_40 = dataGroup_lo_1221[271:256];
  wire [1023:0] dataGroup_lo_1222 = {dataGroup_lo_hi_1222, dataGroup_lo_lo_1222};
  wire [1023:0] dataGroup_hi_1222 = {dataGroup_hi_hi_1222, dataGroup_hi_lo_1222};
  wire [15:0]   dataGroup_6_40 = dataGroup_lo_1222[319:304];
  wire [1023:0] dataGroup_lo_1223 = {dataGroup_lo_hi_1223, dataGroup_lo_lo_1223};
  wire [1023:0] dataGroup_hi_1223 = {dataGroup_hi_hi_1223, dataGroup_hi_lo_1223};
  wire [15:0]   dataGroup_7_40 = dataGroup_lo_1223[367:352];
  wire [1023:0] dataGroup_lo_1224 = {dataGroup_lo_hi_1224, dataGroup_lo_lo_1224};
  wire [1023:0] dataGroup_hi_1224 = {dataGroup_hi_hi_1224, dataGroup_hi_lo_1224};
  wire [15:0]   dataGroup_8_40 = dataGroup_lo_1224[415:400];
  wire [1023:0] dataGroup_lo_1225 = {dataGroup_lo_hi_1225, dataGroup_lo_lo_1225};
  wire [1023:0] dataGroup_hi_1225 = {dataGroup_hi_hi_1225, dataGroup_hi_lo_1225};
  wire [15:0]   dataGroup_9_40 = dataGroup_lo_1225[463:448];
  wire [1023:0] dataGroup_lo_1226 = {dataGroup_lo_hi_1226, dataGroup_lo_lo_1226};
  wire [1023:0] dataGroup_hi_1226 = {dataGroup_hi_hi_1226, dataGroup_hi_lo_1226};
  wire [15:0]   dataGroup_10_40 = dataGroup_lo_1226[511:496];
  wire [1023:0] dataGroup_lo_1227 = {dataGroup_lo_hi_1227, dataGroup_lo_lo_1227};
  wire [1023:0] dataGroup_hi_1227 = {dataGroup_hi_hi_1227, dataGroup_hi_lo_1227};
  wire [15:0]   dataGroup_11_40 = dataGroup_lo_1227[559:544];
  wire [1023:0] dataGroup_lo_1228 = {dataGroup_lo_hi_1228, dataGroup_lo_lo_1228};
  wire [1023:0] dataGroup_hi_1228 = {dataGroup_hi_hi_1228, dataGroup_hi_lo_1228};
  wire [15:0]   dataGroup_12_40 = dataGroup_lo_1228[607:592];
  wire [1023:0] dataGroup_lo_1229 = {dataGroup_lo_hi_1229, dataGroup_lo_lo_1229};
  wire [1023:0] dataGroup_hi_1229 = {dataGroup_hi_hi_1229, dataGroup_hi_lo_1229};
  wire [15:0]   dataGroup_13_40 = dataGroup_lo_1229[655:640];
  wire [1023:0] dataGroup_lo_1230 = {dataGroup_lo_hi_1230, dataGroup_lo_lo_1230};
  wire [1023:0] dataGroup_hi_1230 = {dataGroup_hi_hi_1230, dataGroup_hi_lo_1230};
  wire [15:0]   dataGroup_14_40 = dataGroup_lo_1230[703:688];
  wire [1023:0] dataGroup_lo_1231 = {dataGroup_lo_hi_1231, dataGroup_lo_lo_1231};
  wire [1023:0] dataGroup_hi_1231 = {dataGroup_hi_hi_1231, dataGroup_hi_lo_1231};
  wire [15:0]   dataGroup_15_40 = dataGroup_lo_1231[751:736];
  wire [31:0]   res_lo_lo_lo_40 = {dataGroup_1_40, dataGroup_0_40};
  wire [31:0]   res_lo_lo_hi_40 = {dataGroup_3_40, dataGroup_2_40};
  wire [63:0]   res_lo_lo_40 = {res_lo_lo_hi_40, res_lo_lo_lo_40};
  wire [31:0]   res_lo_hi_lo_40 = {dataGroup_5_40, dataGroup_4_40};
  wire [31:0]   res_lo_hi_hi_40 = {dataGroup_7_40, dataGroup_6_40};
  wire [63:0]   res_lo_hi_40 = {res_lo_hi_hi_40, res_lo_hi_lo_40};
  wire [127:0]  res_lo_40 = {res_lo_hi_40, res_lo_lo_40};
  wire [31:0]   res_hi_lo_lo_40 = {dataGroup_9_40, dataGroup_8_40};
  wire [31:0]   res_hi_lo_hi_40 = {dataGroup_11_40, dataGroup_10_40};
  wire [63:0]   res_hi_lo_40 = {res_hi_lo_hi_40, res_hi_lo_lo_40};
  wire [31:0]   res_hi_hi_lo_40 = {dataGroup_13_40, dataGroup_12_40};
  wire [31:0]   res_hi_hi_hi_40 = {dataGroup_15_40, dataGroup_14_40};
  wire [63:0]   res_hi_hi_40 = {res_hi_hi_hi_40, res_hi_hi_lo_40};
  wire [127:0]  res_hi_40 = {res_hi_hi_40, res_hi_lo_40};
  wire [255:0]  res_81 = {res_hi_40, res_lo_40};
  wire [1023:0] dataGroup_lo_1232 = {dataGroup_lo_hi_1232, dataGroup_lo_lo_1232};
  wire [1023:0] dataGroup_hi_1232 = {dataGroup_hi_hi_1232, dataGroup_hi_lo_1232};
  wire [15:0]   dataGroup_0_41 = dataGroup_lo_1232[47:32];
  wire [1023:0] dataGroup_lo_1233 = {dataGroup_lo_hi_1233, dataGroup_lo_lo_1233};
  wire [1023:0] dataGroup_hi_1233 = {dataGroup_hi_hi_1233, dataGroup_hi_lo_1233};
  wire [15:0]   dataGroup_1_41 = dataGroup_lo_1233[95:80];
  wire [1023:0] dataGroup_lo_1234 = {dataGroup_lo_hi_1234, dataGroup_lo_lo_1234};
  wire [1023:0] dataGroup_hi_1234 = {dataGroup_hi_hi_1234, dataGroup_hi_lo_1234};
  wire [15:0]   dataGroup_2_41 = dataGroup_lo_1234[143:128];
  wire [1023:0] dataGroup_lo_1235 = {dataGroup_lo_hi_1235, dataGroup_lo_lo_1235};
  wire [1023:0] dataGroup_hi_1235 = {dataGroup_hi_hi_1235, dataGroup_hi_lo_1235};
  wire [15:0]   dataGroup_3_41 = dataGroup_lo_1235[191:176];
  wire [1023:0] dataGroup_lo_1236 = {dataGroup_lo_hi_1236, dataGroup_lo_lo_1236};
  wire [1023:0] dataGroup_hi_1236 = {dataGroup_hi_hi_1236, dataGroup_hi_lo_1236};
  wire [15:0]   dataGroup_4_41 = dataGroup_lo_1236[239:224];
  wire [1023:0] dataGroup_lo_1237 = {dataGroup_lo_hi_1237, dataGroup_lo_lo_1237};
  wire [1023:0] dataGroup_hi_1237 = {dataGroup_hi_hi_1237, dataGroup_hi_lo_1237};
  wire [15:0]   dataGroup_5_41 = dataGroup_lo_1237[287:272];
  wire [1023:0] dataGroup_lo_1238 = {dataGroup_lo_hi_1238, dataGroup_lo_lo_1238};
  wire [1023:0] dataGroup_hi_1238 = {dataGroup_hi_hi_1238, dataGroup_hi_lo_1238};
  wire [15:0]   dataGroup_6_41 = dataGroup_lo_1238[335:320];
  wire [1023:0] dataGroup_lo_1239 = {dataGroup_lo_hi_1239, dataGroup_lo_lo_1239};
  wire [1023:0] dataGroup_hi_1239 = {dataGroup_hi_hi_1239, dataGroup_hi_lo_1239};
  wire [15:0]   dataGroup_7_41 = dataGroup_lo_1239[383:368];
  wire [1023:0] dataGroup_lo_1240 = {dataGroup_lo_hi_1240, dataGroup_lo_lo_1240};
  wire [1023:0] dataGroup_hi_1240 = {dataGroup_hi_hi_1240, dataGroup_hi_lo_1240};
  wire [15:0]   dataGroup_8_41 = dataGroup_lo_1240[431:416];
  wire [1023:0] dataGroup_lo_1241 = {dataGroup_lo_hi_1241, dataGroup_lo_lo_1241};
  wire [1023:0] dataGroup_hi_1241 = {dataGroup_hi_hi_1241, dataGroup_hi_lo_1241};
  wire [15:0]   dataGroup_9_41 = dataGroup_lo_1241[479:464];
  wire [1023:0] dataGroup_lo_1242 = {dataGroup_lo_hi_1242, dataGroup_lo_lo_1242};
  wire [1023:0] dataGroup_hi_1242 = {dataGroup_hi_hi_1242, dataGroup_hi_lo_1242};
  wire [15:0]   dataGroup_10_41 = dataGroup_lo_1242[527:512];
  wire [1023:0] dataGroup_lo_1243 = {dataGroup_lo_hi_1243, dataGroup_lo_lo_1243};
  wire [1023:0] dataGroup_hi_1243 = {dataGroup_hi_hi_1243, dataGroup_hi_lo_1243};
  wire [15:0]   dataGroup_11_41 = dataGroup_lo_1243[575:560];
  wire [1023:0] dataGroup_lo_1244 = {dataGroup_lo_hi_1244, dataGroup_lo_lo_1244};
  wire [1023:0] dataGroup_hi_1244 = {dataGroup_hi_hi_1244, dataGroup_hi_lo_1244};
  wire [15:0]   dataGroup_12_41 = dataGroup_lo_1244[623:608];
  wire [1023:0] dataGroup_lo_1245 = {dataGroup_lo_hi_1245, dataGroup_lo_lo_1245};
  wire [1023:0] dataGroup_hi_1245 = {dataGroup_hi_hi_1245, dataGroup_hi_lo_1245};
  wire [15:0]   dataGroup_13_41 = dataGroup_lo_1245[671:656];
  wire [1023:0] dataGroup_lo_1246 = {dataGroup_lo_hi_1246, dataGroup_lo_lo_1246};
  wire [1023:0] dataGroup_hi_1246 = {dataGroup_hi_hi_1246, dataGroup_hi_lo_1246};
  wire [15:0]   dataGroup_14_41 = dataGroup_lo_1246[719:704];
  wire [1023:0] dataGroup_lo_1247 = {dataGroup_lo_hi_1247, dataGroup_lo_lo_1247};
  wire [1023:0] dataGroup_hi_1247 = {dataGroup_hi_hi_1247, dataGroup_hi_lo_1247};
  wire [15:0]   dataGroup_15_41 = dataGroup_lo_1247[767:752];
  wire [31:0]   res_lo_lo_lo_41 = {dataGroup_1_41, dataGroup_0_41};
  wire [31:0]   res_lo_lo_hi_41 = {dataGroup_3_41, dataGroup_2_41};
  wire [63:0]   res_lo_lo_41 = {res_lo_lo_hi_41, res_lo_lo_lo_41};
  wire [31:0]   res_lo_hi_lo_41 = {dataGroup_5_41, dataGroup_4_41};
  wire [31:0]   res_lo_hi_hi_41 = {dataGroup_7_41, dataGroup_6_41};
  wire [63:0]   res_lo_hi_41 = {res_lo_hi_hi_41, res_lo_hi_lo_41};
  wire [127:0]  res_lo_41 = {res_lo_hi_41, res_lo_lo_41};
  wire [31:0]   res_hi_lo_lo_41 = {dataGroup_9_41, dataGroup_8_41};
  wire [31:0]   res_hi_lo_hi_41 = {dataGroup_11_41, dataGroup_10_41};
  wire [63:0]   res_hi_lo_41 = {res_hi_lo_hi_41, res_hi_lo_lo_41};
  wire [31:0]   res_hi_hi_lo_41 = {dataGroup_13_41, dataGroup_12_41};
  wire [31:0]   res_hi_hi_hi_41 = {dataGroup_15_41, dataGroup_14_41};
  wire [63:0]   res_hi_hi_41 = {res_hi_hi_hi_41, res_hi_hi_lo_41};
  wire [127:0]  res_hi_41 = {res_hi_hi_41, res_hi_lo_41};
  wire [255:0]  res_82 = {res_hi_41, res_lo_41};
  wire [511:0]  lo_lo_10 = {res_81, res_80};
  wire [511:0]  lo_hi_10 = {256'h0, res_82};
  wire [1023:0] lo_10 = {lo_hi_10, lo_lo_10};
  wire [2047:0] regroupLoadData_1_2 = {1024'h0, lo_10};
  wire [1023:0] dataGroup_lo_1248 = {dataGroup_lo_hi_1248, dataGroup_lo_lo_1248};
  wire [1023:0] dataGroup_hi_1248 = {dataGroup_hi_hi_1248, dataGroup_hi_lo_1248};
  wire [15:0]   dataGroup_0_42 = dataGroup_lo_1248[15:0];
  wire [1023:0] dataGroup_lo_1249 = {dataGroup_lo_hi_1249, dataGroup_lo_lo_1249};
  wire [1023:0] dataGroup_hi_1249 = {dataGroup_hi_hi_1249, dataGroup_hi_lo_1249};
  wire [15:0]   dataGroup_1_42 = dataGroup_lo_1249[79:64];
  wire [1023:0] dataGroup_lo_1250 = {dataGroup_lo_hi_1250, dataGroup_lo_lo_1250};
  wire [1023:0] dataGroup_hi_1250 = {dataGroup_hi_hi_1250, dataGroup_hi_lo_1250};
  wire [15:0]   dataGroup_2_42 = dataGroup_lo_1250[143:128];
  wire [1023:0] dataGroup_lo_1251 = {dataGroup_lo_hi_1251, dataGroup_lo_lo_1251};
  wire [1023:0] dataGroup_hi_1251 = {dataGroup_hi_hi_1251, dataGroup_hi_lo_1251};
  wire [15:0]   dataGroup_3_42 = dataGroup_lo_1251[207:192];
  wire [1023:0] dataGroup_lo_1252 = {dataGroup_lo_hi_1252, dataGroup_lo_lo_1252};
  wire [1023:0] dataGroup_hi_1252 = {dataGroup_hi_hi_1252, dataGroup_hi_lo_1252};
  wire [15:0]   dataGroup_4_42 = dataGroup_lo_1252[271:256];
  wire [1023:0] dataGroup_lo_1253 = {dataGroup_lo_hi_1253, dataGroup_lo_lo_1253};
  wire [1023:0] dataGroup_hi_1253 = {dataGroup_hi_hi_1253, dataGroup_hi_lo_1253};
  wire [15:0]   dataGroup_5_42 = dataGroup_lo_1253[335:320];
  wire [1023:0] dataGroup_lo_1254 = {dataGroup_lo_hi_1254, dataGroup_lo_lo_1254};
  wire [1023:0] dataGroup_hi_1254 = {dataGroup_hi_hi_1254, dataGroup_hi_lo_1254};
  wire [15:0]   dataGroup_6_42 = dataGroup_lo_1254[399:384];
  wire [1023:0] dataGroup_lo_1255 = {dataGroup_lo_hi_1255, dataGroup_lo_lo_1255};
  wire [1023:0] dataGroup_hi_1255 = {dataGroup_hi_hi_1255, dataGroup_hi_lo_1255};
  wire [15:0]   dataGroup_7_42 = dataGroup_lo_1255[463:448];
  wire [1023:0] dataGroup_lo_1256 = {dataGroup_lo_hi_1256, dataGroup_lo_lo_1256};
  wire [1023:0] dataGroup_hi_1256 = {dataGroup_hi_hi_1256, dataGroup_hi_lo_1256};
  wire [15:0]   dataGroup_8_42 = dataGroup_lo_1256[527:512];
  wire [1023:0] dataGroup_lo_1257 = {dataGroup_lo_hi_1257, dataGroup_lo_lo_1257};
  wire [1023:0] dataGroup_hi_1257 = {dataGroup_hi_hi_1257, dataGroup_hi_lo_1257};
  wire [15:0]   dataGroup_9_42 = dataGroup_lo_1257[591:576];
  wire [1023:0] dataGroup_lo_1258 = {dataGroup_lo_hi_1258, dataGroup_lo_lo_1258};
  wire [1023:0] dataGroup_hi_1258 = {dataGroup_hi_hi_1258, dataGroup_hi_lo_1258};
  wire [15:0]   dataGroup_10_42 = dataGroup_lo_1258[655:640];
  wire [1023:0] dataGroup_lo_1259 = {dataGroup_lo_hi_1259, dataGroup_lo_lo_1259};
  wire [1023:0] dataGroup_hi_1259 = {dataGroup_hi_hi_1259, dataGroup_hi_lo_1259};
  wire [15:0]   dataGroup_11_42 = dataGroup_lo_1259[719:704];
  wire [1023:0] dataGroup_lo_1260 = {dataGroup_lo_hi_1260, dataGroup_lo_lo_1260};
  wire [1023:0] dataGroup_hi_1260 = {dataGroup_hi_hi_1260, dataGroup_hi_lo_1260};
  wire [15:0]   dataGroup_12_42 = dataGroup_lo_1260[783:768];
  wire [1023:0] dataGroup_lo_1261 = {dataGroup_lo_hi_1261, dataGroup_lo_lo_1261};
  wire [1023:0] dataGroup_hi_1261 = {dataGroup_hi_hi_1261, dataGroup_hi_lo_1261};
  wire [15:0]   dataGroup_13_42 = dataGroup_lo_1261[847:832];
  wire [1023:0] dataGroup_lo_1262 = {dataGroup_lo_hi_1262, dataGroup_lo_lo_1262};
  wire [1023:0] dataGroup_hi_1262 = {dataGroup_hi_hi_1262, dataGroup_hi_lo_1262};
  wire [15:0]   dataGroup_14_42 = dataGroup_lo_1262[911:896];
  wire [1023:0] dataGroup_lo_1263 = {dataGroup_lo_hi_1263, dataGroup_lo_lo_1263};
  wire [1023:0] dataGroup_hi_1263 = {dataGroup_hi_hi_1263, dataGroup_hi_lo_1263};
  wire [15:0]   dataGroup_15_42 = dataGroup_lo_1263[975:960];
  wire [31:0]   res_lo_lo_lo_42 = {dataGroup_1_42, dataGroup_0_42};
  wire [31:0]   res_lo_lo_hi_42 = {dataGroup_3_42, dataGroup_2_42};
  wire [63:0]   res_lo_lo_42 = {res_lo_lo_hi_42, res_lo_lo_lo_42};
  wire [31:0]   res_lo_hi_lo_42 = {dataGroup_5_42, dataGroup_4_42};
  wire [31:0]   res_lo_hi_hi_42 = {dataGroup_7_42, dataGroup_6_42};
  wire [63:0]   res_lo_hi_42 = {res_lo_hi_hi_42, res_lo_hi_lo_42};
  wire [127:0]  res_lo_42 = {res_lo_hi_42, res_lo_lo_42};
  wire [31:0]   res_hi_lo_lo_42 = {dataGroup_9_42, dataGroup_8_42};
  wire [31:0]   res_hi_lo_hi_42 = {dataGroup_11_42, dataGroup_10_42};
  wire [63:0]   res_hi_lo_42 = {res_hi_lo_hi_42, res_hi_lo_lo_42};
  wire [31:0]   res_hi_hi_lo_42 = {dataGroup_13_42, dataGroup_12_42};
  wire [31:0]   res_hi_hi_hi_42 = {dataGroup_15_42, dataGroup_14_42};
  wire [63:0]   res_hi_hi_42 = {res_hi_hi_hi_42, res_hi_hi_lo_42};
  wire [127:0]  res_hi_42 = {res_hi_hi_42, res_hi_lo_42};
  wire [255:0]  res_88 = {res_hi_42, res_lo_42};
  wire [1023:0] dataGroup_lo_1264 = {dataGroup_lo_hi_1264, dataGroup_lo_lo_1264};
  wire [1023:0] dataGroup_hi_1264 = {dataGroup_hi_hi_1264, dataGroup_hi_lo_1264};
  wire [15:0]   dataGroup_0_43 = dataGroup_lo_1264[31:16];
  wire [1023:0] dataGroup_lo_1265 = {dataGroup_lo_hi_1265, dataGroup_lo_lo_1265};
  wire [1023:0] dataGroup_hi_1265 = {dataGroup_hi_hi_1265, dataGroup_hi_lo_1265};
  wire [15:0]   dataGroup_1_43 = dataGroup_lo_1265[95:80];
  wire [1023:0] dataGroup_lo_1266 = {dataGroup_lo_hi_1266, dataGroup_lo_lo_1266};
  wire [1023:0] dataGroup_hi_1266 = {dataGroup_hi_hi_1266, dataGroup_hi_lo_1266};
  wire [15:0]   dataGroup_2_43 = dataGroup_lo_1266[159:144];
  wire [1023:0] dataGroup_lo_1267 = {dataGroup_lo_hi_1267, dataGroup_lo_lo_1267};
  wire [1023:0] dataGroup_hi_1267 = {dataGroup_hi_hi_1267, dataGroup_hi_lo_1267};
  wire [15:0]   dataGroup_3_43 = dataGroup_lo_1267[223:208];
  wire [1023:0] dataGroup_lo_1268 = {dataGroup_lo_hi_1268, dataGroup_lo_lo_1268};
  wire [1023:0] dataGroup_hi_1268 = {dataGroup_hi_hi_1268, dataGroup_hi_lo_1268};
  wire [15:0]   dataGroup_4_43 = dataGroup_lo_1268[287:272];
  wire [1023:0] dataGroup_lo_1269 = {dataGroup_lo_hi_1269, dataGroup_lo_lo_1269};
  wire [1023:0] dataGroup_hi_1269 = {dataGroup_hi_hi_1269, dataGroup_hi_lo_1269};
  wire [15:0]   dataGroup_5_43 = dataGroup_lo_1269[351:336];
  wire [1023:0] dataGroup_lo_1270 = {dataGroup_lo_hi_1270, dataGroup_lo_lo_1270};
  wire [1023:0] dataGroup_hi_1270 = {dataGroup_hi_hi_1270, dataGroup_hi_lo_1270};
  wire [15:0]   dataGroup_6_43 = dataGroup_lo_1270[415:400];
  wire [1023:0] dataGroup_lo_1271 = {dataGroup_lo_hi_1271, dataGroup_lo_lo_1271};
  wire [1023:0] dataGroup_hi_1271 = {dataGroup_hi_hi_1271, dataGroup_hi_lo_1271};
  wire [15:0]   dataGroup_7_43 = dataGroup_lo_1271[479:464];
  wire [1023:0] dataGroup_lo_1272 = {dataGroup_lo_hi_1272, dataGroup_lo_lo_1272};
  wire [1023:0] dataGroup_hi_1272 = {dataGroup_hi_hi_1272, dataGroup_hi_lo_1272};
  wire [15:0]   dataGroup_8_43 = dataGroup_lo_1272[543:528];
  wire [1023:0] dataGroup_lo_1273 = {dataGroup_lo_hi_1273, dataGroup_lo_lo_1273};
  wire [1023:0] dataGroup_hi_1273 = {dataGroup_hi_hi_1273, dataGroup_hi_lo_1273};
  wire [15:0]   dataGroup_9_43 = dataGroup_lo_1273[607:592];
  wire [1023:0] dataGroup_lo_1274 = {dataGroup_lo_hi_1274, dataGroup_lo_lo_1274};
  wire [1023:0] dataGroup_hi_1274 = {dataGroup_hi_hi_1274, dataGroup_hi_lo_1274};
  wire [15:0]   dataGroup_10_43 = dataGroup_lo_1274[671:656];
  wire [1023:0] dataGroup_lo_1275 = {dataGroup_lo_hi_1275, dataGroup_lo_lo_1275};
  wire [1023:0] dataGroup_hi_1275 = {dataGroup_hi_hi_1275, dataGroup_hi_lo_1275};
  wire [15:0]   dataGroup_11_43 = dataGroup_lo_1275[735:720];
  wire [1023:0] dataGroup_lo_1276 = {dataGroup_lo_hi_1276, dataGroup_lo_lo_1276};
  wire [1023:0] dataGroup_hi_1276 = {dataGroup_hi_hi_1276, dataGroup_hi_lo_1276};
  wire [15:0]   dataGroup_12_43 = dataGroup_lo_1276[799:784];
  wire [1023:0] dataGroup_lo_1277 = {dataGroup_lo_hi_1277, dataGroup_lo_lo_1277};
  wire [1023:0] dataGroup_hi_1277 = {dataGroup_hi_hi_1277, dataGroup_hi_lo_1277};
  wire [15:0]   dataGroup_13_43 = dataGroup_lo_1277[863:848];
  wire [1023:0] dataGroup_lo_1278 = {dataGroup_lo_hi_1278, dataGroup_lo_lo_1278};
  wire [1023:0] dataGroup_hi_1278 = {dataGroup_hi_hi_1278, dataGroup_hi_lo_1278};
  wire [15:0]   dataGroup_14_43 = dataGroup_lo_1278[927:912];
  wire [1023:0] dataGroup_lo_1279 = {dataGroup_lo_hi_1279, dataGroup_lo_lo_1279};
  wire [1023:0] dataGroup_hi_1279 = {dataGroup_hi_hi_1279, dataGroup_hi_lo_1279};
  wire [15:0]   dataGroup_15_43 = dataGroup_lo_1279[991:976];
  wire [31:0]   res_lo_lo_lo_43 = {dataGroup_1_43, dataGroup_0_43};
  wire [31:0]   res_lo_lo_hi_43 = {dataGroup_3_43, dataGroup_2_43};
  wire [63:0]   res_lo_lo_43 = {res_lo_lo_hi_43, res_lo_lo_lo_43};
  wire [31:0]   res_lo_hi_lo_43 = {dataGroup_5_43, dataGroup_4_43};
  wire [31:0]   res_lo_hi_hi_43 = {dataGroup_7_43, dataGroup_6_43};
  wire [63:0]   res_lo_hi_43 = {res_lo_hi_hi_43, res_lo_hi_lo_43};
  wire [127:0]  res_lo_43 = {res_lo_hi_43, res_lo_lo_43};
  wire [31:0]   res_hi_lo_lo_43 = {dataGroup_9_43, dataGroup_8_43};
  wire [31:0]   res_hi_lo_hi_43 = {dataGroup_11_43, dataGroup_10_43};
  wire [63:0]   res_hi_lo_43 = {res_hi_lo_hi_43, res_hi_lo_lo_43};
  wire [31:0]   res_hi_hi_lo_43 = {dataGroup_13_43, dataGroup_12_43};
  wire [31:0]   res_hi_hi_hi_43 = {dataGroup_15_43, dataGroup_14_43};
  wire [63:0]   res_hi_hi_43 = {res_hi_hi_hi_43, res_hi_hi_lo_43};
  wire [127:0]  res_hi_43 = {res_hi_hi_43, res_hi_lo_43};
  wire [255:0]  res_89 = {res_hi_43, res_lo_43};
  wire [1023:0] dataGroup_lo_1280 = {dataGroup_lo_hi_1280, dataGroup_lo_lo_1280};
  wire [1023:0] dataGroup_hi_1280 = {dataGroup_hi_hi_1280, dataGroup_hi_lo_1280};
  wire [15:0]   dataGroup_0_44 = dataGroup_lo_1280[47:32];
  wire [1023:0] dataGroup_lo_1281 = {dataGroup_lo_hi_1281, dataGroup_lo_lo_1281};
  wire [1023:0] dataGroup_hi_1281 = {dataGroup_hi_hi_1281, dataGroup_hi_lo_1281};
  wire [15:0]   dataGroup_1_44 = dataGroup_lo_1281[111:96];
  wire [1023:0] dataGroup_lo_1282 = {dataGroup_lo_hi_1282, dataGroup_lo_lo_1282};
  wire [1023:0] dataGroup_hi_1282 = {dataGroup_hi_hi_1282, dataGroup_hi_lo_1282};
  wire [15:0]   dataGroup_2_44 = dataGroup_lo_1282[175:160];
  wire [1023:0] dataGroup_lo_1283 = {dataGroup_lo_hi_1283, dataGroup_lo_lo_1283};
  wire [1023:0] dataGroup_hi_1283 = {dataGroup_hi_hi_1283, dataGroup_hi_lo_1283};
  wire [15:0]   dataGroup_3_44 = dataGroup_lo_1283[239:224];
  wire [1023:0] dataGroup_lo_1284 = {dataGroup_lo_hi_1284, dataGroup_lo_lo_1284};
  wire [1023:0] dataGroup_hi_1284 = {dataGroup_hi_hi_1284, dataGroup_hi_lo_1284};
  wire [15:0]   dataGroup_4_44 = dataGroup_lo_1284[303:288];
  wire [1023:0] dataGroup_lo_1285 = {dataGroup_lo_hi_1285, dataGroup_lo_lo_1285};
  wire [1023:0] dataGroup_hi_1285 = {dataGroup_hi_hi_1285, dataGroup_hi_lo_1285};
  wire [15:0]   dataGroup_5_44 = dataGroup_lo_1285[367:352];
  wire [1023:0] dataGroup_lo_1286 = {dataGroup_lo_hi_1286, dataGroup_lo_lo_1286};
  wire [1023:0] dataGroup_hi_1286 = {dataGroup_hi_hi_1286, dataGroup_hi_lo_1286};
  wire [15:0]   dataGroup_6_44 = dataGroup_lo_1286[431:416];
  wire [1023:0] dataGroup_lo_1287 = {dataGroup_lo_hi_1287, dataGroup_lo_lo_1287};
  wire [1023:0] dataGroup_hi_1287 = {dataGroup_hi_hi_1287, dataGroup_hi_lo_1287};
  wire [15:0]   dataGroup_7_44 = dataGroup_lo_1287[495:480];
  wire [1023:0] dataGroup_lo_1288 = {dataGroup_lo_hi_1288, dataGroup_lo_lo_1288};
  wire [1023:0] dataGroup_hi_1288 = {dataGroup_hi_hi_1288, dataGroup_hi_lo_1288};
  wire [15:0]   dataGroup_8_44 = dataGroup_lo_1288[559:544];
  wire [1023:0] dataGroup_lo_1289 = {dataGroup_lo_hi_1289, dataGroup_lo_lo_1289};
  wire [1023:0] dataGroup_hi_1289 = {dataGroup_hi_hi_1289, dataGroup_hi_lo_1289};
  wire [15:0]   dataGroup_9_44 = dataGroup_lo_1289[623:608];
  wire [1023:0] dataGroup_lo_1290 = {dataGroup_lo_hi_1290, dataGroup_lo_lo_1290};
  wire [1023:0] dataGroup_hi_1290 = {dataGroup_hi_hi_1290, dataGroup_hi_lo_1290};
  wire [15:0]   dataGroup_10_44 = dataGroup_lo_1290[687:672];
  wire [1023:0] dataGroup_lo_1291 = {dataGroup_lo_hi_1291, dataGroup_lo_lo_1291};
  wire [1023:0] dataGroup_hi_1291 = {dataGroup_hi_hi_1291, dataGroup_hi_lo_1291};
  wire [15:0]   dataGroup_11_44 = dataGroup_lo_1291[751:736];
  wire [1023:0] dataGroup_lo_1292 = {dataGroup_lo_hi_1292, dataGroup_lo_lo_1292};
  wire [1023:0] dataGroup_hi_1292 = {dataGroup_hi_hi_1292, dataGroup_hi_lo_1292};
  wire [15:0]   dataGroup_12_44 = dataGroup_lo_1292[815:800];
  wire [1023:0] dataGroup_lo_1293 = {dataGroup_lo_hi_1293, dataGroup_lo_lo_1293};
  wire [1023:0] dataGroup_hi_1293 = {dataGroup_hi_hi_1293, dataGroup_hi_lo_1293};
  wire [15:0]   dataGroup_13_44 = dataGroup_lo_1293[879:864];
  wire [1023:0] dataGroup_lo_1294 = {dataGroup_lo_hi_1294, dataGroup_lo_lo_1294};
  wire [1023:0] dataGroup_hi_1294 = {dataGroup_hi_hi_1294, dataGroup_hi_lo_1294};
  wire [15:0]   dataGroup_14_44 = dataGroup_lo_1294[943:928];
  wire [1023:0] dataGroup_lo_1295 = {dataGroup_lo_hi_1295, dataGroup_lo_lo_1295};
  wire [1023:0] dataGroup_hi_1295 = {dataGroup_hi_hi_1295, dataGroup_hi_lo_1295};
  wire [15:0]   dataGroup_15_44 = dataGroup_lo_1295[1007:992];
  wire [31:0]   res_lo_lo_lo_44 = {dataGroup_1_44, dataGroup_0_44};
  wire [31:0]   res_lo_lo_hi_44 = {dataGroup_3_44, dataGroup_2_44};
  wire [63:0]   res_lo_lo_44 = {res_lo_lo_hi_44, res_lo_lo_lo_44};
  wire [31:0]   res_lo_hi_lo_44 = {dataGroup_5_44, dataGroup_4_44};
  wire [31:0]   res_lo_hi_hi_44 = {dataGroup_7_44, dataGroup_6_44};
  wire [63:0]   res_lo_hi_44 = {res_lo_hi_hi_44, res_lo_hi_lo_44};
  wire [127:0]  res_lo_44 = {res_lo_hi_44, res_lo_lo_44};
  wire [31:0]   res_hi_lo_lo_44 = {dataGroup_9_44, dataGroup_8_44};
  wire [31:0]   res_hi_lo_hi_44 = {dataGroup_11_44, dataGroup_10_44};
  wire [63:0]   res_hi_lo_44 = {res_hi_lo_hi_44, res_hi_lo_lo_44};
  wire [31:0]   res_hi_hi_lo_44 = {dataGroup_13_44, dataGroup_12_44};
  wire [31:0]   res_hi_hi_hi_44 = {dataGroup_15_44, dataGroup_14_44};
  wire [63:0]   res_hi_hi_44 = {res_hi_hi_hi_44, res_hi_hi_lo_44};
  wire [127:0]  res_hi_44 = {res_hi_hi_44, res_hi_lo_44};
  wire [255:0]  res_90 = {res_hi_44, res_lo_44};
  wire [1023:0] dataGroup_lo_1296 = {dataGroup_lo_hi_1296, dataGroup_lo_lo_1296};
  wire [1023:0] dataGroup_hi_1296 = {dataGroup_hi_hi_1296, dataGroup_hi_lo_1296};
  wire [15:0]   dataGroup_0_45 = dataGroup_lo_1296[63:48];
  wire [1023:0] dataGroup_lo_1297 = {dataGroup_lo_hi_1297, dataGroup_lo_lo_1297};
  wire [1023:0] dataGroup_hi_1297 = {dataGroup_hi_hi_1297, dataGroup_hi_lo_1297};
  wire [15:0]   dataGroup_1_45 = dataGroup_lo_1297[127:112];
  wire [1023:0] dataGroup_lo_1298 = {dataGroup_lo_hi_1298, dataGroup_lo_lo_1298};
  wire [1023:0] dataGroup_hi_1298 = {dataGroup_hi_hi_1298, dataGroup_hi_lo_1298};
  wire [15:0]   dataGroup_2_45 = dataGroup_lo_1298[191:176];
  wire [1023:0] dataGroup_lo_1299 = {dataGroup_lo_hi_1299, dataGroup_lo_lo_1299};
  wire [1023:0] dataGroup_hi_1299 = {dataGroup_hi_hi_1299, dataGroup_hi_lo_1299};
  wire [15:0]   dataGroup_3_45 = dataGroup_lo_1299[255:240];
  wire [1023:0] dataGroup_lo_1300 = {dataGroup_lo_hi_1300, dataGroup_lo_lo_1300};
  wire [1023:0] dataGroup_hi_1300 = {dataGroup_hi_hi_1300, dataGroup_hi_lo_1300};
  wire [15:0]   dataGroup_4_45 = dataGroup_lo_1300[319:304];
  wire [1023:0] dataGroup_lo_1301 = {dataGroup_lo_hi_1301, dataGroup_lo_lo_1301};
  wire [1023:0] dataGroup_hi_1301 = {dataGroup_hi_hi_1301, dataGroup_hi_lo_1301};
  wire [15:0]   dataGroup_5_45 = dataGroup_lo_1301[383:368];
  wire [1023:0] dataGroup_lo_1302 = {dataGroup_lo_hi_1302, dataGroup_lo_lo_1302};
  wire [1023:0] dataGroup_hi_1302 = {dataGroup_hi_hi_1302, dataGroup_hi_lo_1302};
  wire [15:0]   dataGroup_6_45 = dataGroup_lo_1302[447:432];
  wire [1023:0] dataGroup_lo_1303 = {dataGroup_lo_hi_1303, dataGroup_lo_lo_1303};
  wire [1023:0] dataGroup_hi_1303 = {dataGroup_hi_hi_1303, dataGroup_hi_lo_1303};
  wire [15:0]   dataGroup_7_45 = dataGroup_lo_1303[511:496];
  wire [1023:0] dataGroup_lo_1304 = {dataGroup_lo_hi_1304, dataGroup_lo_lo_1304};
  wire [1023:0] dataGroup_hi_1304 = {dataGroup_hi_hi_1304, dataGroup_hi_lo_1304};
  wire [15:0]   dataGroup_8_45 = dataGroup_lo_1304[575:560];
  wire [1023:0] dataGroup_lo_1305 = {dataGroup_lo_hi_1305, dataGroup_lo_lo_1305};
  wire [1023:0] dataGroup_hi_1305 = {dataGroup_hi_hi_1305, dataGroup_hi_lo_1305};
  wire [15:0]   dataGroup_9_45 = dataGroup_lo_1305[639:624];
  wire [1023:0] dataGroup_lo_1306 = {dataGroup_lo_hi_1306, dataGroup_lo_lo_1306};
  wire [1023:0] dataGroup_hi_1306 = {dataGroup_hi_hi_1306, dataGroup_hi_lo_1306};
  wire [15:0]   dataGroup_10_45 = dataGroup_lo_1306[703:688];
  wire [1023:0] dataGroup_lo_1307 = {dataGroup_lo_hi_1307, dataGroup_lo_lo_1307};
  wire [1023:0] dataGroup_hi_1307 = {dataGroup_hi_hi_1307, dataGroup_hi_lo_1307};
  wire [15:0]   dataGroup_11_45 = dataGroup_lo_1307[767:752];
  wire [1023:0] dataGroup_lo_1308 = {dataGroup_lo_hi_1308, dataGroup_lo_lo_1308};
  wire [1023:0] dataGroup_hi_1308 = {dataGroup_hi_hi_1308, dataGroup_hi_lo_1308};
  wire [15:0]   dataGroup_12_45 = dataGroup_lo_1308[831:816];
  wire [1023:0] dataGroup_lo_1309 = {dataGroup_lo_hi_1309, dataGroup_lo_lo_1309};
  wire [1023:0] dataGroup_hi_1309 = {dataGroup_hi_hi_1309, dataGroup_hi_lo_1309};
  wire [15:0]   dataGroup_13_45 = dataGroup_lo_1309[895:880];
  wire [1023:0] dataGroup_lo_1310 = {dataGroup_lo_hi_1310, dataGroup_lo_lo_1310};
  wire [1023:0] dataGroup_hi_1310 = {dataGroup_hi_hi_1310, dataGroup_hi_lo_1310};
  wire [15:0]   dataGroup_14_45 = dataGroup_lo_1310[959:944];
  wire [1023:0] dataGroup_lo_1311 = {dataGroup_lo_hi_1311, dataGroup_lo_lo_1311};
  wire [1023:0] dataGroup_hi_1311 = {dataGroup_hi_hi_1311, dataGroup_hi_lo_1311};
  wire [15:0]   dataGroup_15_45 = dataGroup_lo_1311[1023:1008];
  wire [31:0]   res_lo_lo_lo_45 = {dataGroup_1_45, dataGroup_0_45};
  wire [31:0]   res_lo_lo_hi_45 = {dataGroup_3_45, dataGroup_2_45};
  wire [63:0]   res_lo_lo_45 = {res_lo_lo_hi_45, res_lo_lo_lo_45};
  wire [31:0]   res_lo_hi_lo_45 = {dataGroup_5_45, dataGroup_4_45};
  wire [31:0]   res_lo_hi_hi_45 = {dataGroup_7_45, dataGroup_6_45};
  wire [63:0]   res_lo_hi_45 = {res_lo_hi_hi_45, res_lo_hi_lo_45};
  wire [127:0]  res_lo_45 = {res_lo_hi_45, res_lo_lo_45};
  wire [31:0]   res_hi_lo_lo_45 = {dataGroup_9_45, dataGroup_8_45};
  wire [31:0]   res_hi_lo_hi_45 = {dataGroup_11_45, dataGroup_10_45};
  wire [63:0]   res_hi_lo_45 = {res_hi_lo_hi_45, res_hi_lo_lo_45};
  wire [31:0]   res_hi_hi_lo_45 = {dataGroup_13_45, dataGroup_12_45};
  wire [31:0]   res_hi_hi_hi_45 = {dataGroup_15_45, dataGroup_14_45};
  wire [63:0]   res_hi_hi_45 = {res_hi_hi_hi_45, res_hi_hi_lo_45};
  wire [127:0]  res_hi_45 = {res_hi_hi_45, res_hi_lo_45};
  wire [255:0]  res_91 = {res_hi_45, res_lo_45};
  wire [511:0]  lo_lo_11 = {res_89, res_88};
  wire [511:0]  lo_hi_11 = {res_91, res_90};
  wire [1023:0] lo_11 = {lo_hi_11, lo_lo_11};
  wire [2047:0] regroupLoadData_1_3 = {1024'h0, lo_11};
  wire [1023:0] dataGroup_lo_1312 = {dataGroup_lo_hi_1312, dataGroup_lo_lo_1312};
  wire [1023:0] dataGroup_hi_1312 = {dataGroup_hi_hi_1312, dataGroup_hi_lo_1312};
  wire [15:0]   dataGroup_0_46 = dataGroup_lo_1312[15:0];
  wire [1023:0] dataGroup_lo_1313 = {dataGroup_lo_hi_1313, dataGroup_lo_lo_1313};
  wire [1023:0] dataGroup_hi_1313 = {dataGroup_hi_hi_1313, dataGroup_hi_lo_1313};
  wire [15:0]   dataGroup_1_46 = dataGroup_lo_1313[95:80];
  wire [1023:0] dataGroup_lo_1314 = {dataGroup_lo_hi_1314, dataGroup_lo_lo_1314};
  wire [1023:0] dataGroup_hi_1314 = {dataGroup_hi_hi_1314, dataGroup_hi_lo_1314};
  wire [15:0]   dataGroup_2_46 = dataGroup_lo_1314[175:160];
  wire [1023:0] dataGroup_lo_1315 = {dataGroup_lo_hi_1315, dataGroup_lo_lo_1315};
  wire [1023:0] dataGroup_hi_1315 = {dataGroup_hi_hi_1315, dataGroup_hi_lo_1315};
  wire [15:0]   dataGroup_3_46 = dataGroup_lo_1315[255:240];
  wire [1023:0] dataGroup_lo_1316 = {dataGroup_lo_hi_1316, dataGroup_lo_lo_1316};
  wire [1023:0] dataGroup_hi_1316 = {dataGroup_hi_hi_1316, dataGroup_hi_lo_1316};
  wire [15:0]   dataGroup_4_46 = dataGroup_lo_1316[335:320];
  wire [1023:0] dataGroup_lo_1317 = {dataGroup_lo_hi_1317, dataGroup_lo_lo_1317};
  wire [1023:0] dataGroup_hi_1317 = {dataGroup_hi_hi_1317, dataGroup_hi_lo_1317};
  wire [15:0]   dataGroup_5_46 = dataGroup_lo_1317[415:400];
  wire [1023:0] dataGroup_lo_1318 = {dataGroup_lo_hi_1318, dataGroup_lo_lo_1318};
  wire [1023:0] dataGroup_hi_1318 = {dataGroup_hi_hi_1318, dataGroup_hi_lo_1318};
  wire [15:0]   dataGroup_6_46 = dataGroup_lo_1318[495:480];
  wire [1023:0] dataGroup_lo_1319 = {dataGroup_lo_hi_1319, dataGroup_lo_lo_1319};
  wire [1023:0] dataGroup_hi_1319 = {dataGroup_hi_hi_1319, dataGroup_hi_lo_1319};
  wire [15:0]   dataGroup_7_46 = dataGroup_lo_1319[575:560];
  wire [1023:0] dataGroup_lo_1320 = {dataGroup_lo_hi_1320, dataGroup_lo_lo_1320};
  wire [1023:0] dataGroup_hi_1320 = {dataGroup_hi_hi_1320, dataGroup_hi_lo_1320};
  wire [15:0]   dataGroup_8_46 = dataGroup_lo_1320[655:640];
  wire [1023:0] dataGroup_lo_1321 = {dataGroup_lo_hi_1321, dataGroup_lo_lo_1321};
  wire [1023:0] dataGroup_hi_1321 = {dataGroup_hi_hi_1321, dataGroup_hi_lo_1321};
  wire [15:0]   dataGroup_9_46 = dataGroup_lo_1321[735:720];
  wire [1023:0] dataGroup_lo_1322 = {dataGroup_lo_hi_1322, dataGroup_lo_lo_1322};
  wire [1023:0] dataGroup_hi_1322 = {dataGroup_hi_hi_1322, dataGroup_hi_lo_1322};
  wire [15:0]   dataGroup_10_46 = dataGroup_lo_1322[815:800];
  wire [1023:0] dataGroup_lo_1323 = {dataGroup_lo_hi_1323, dataGroup_lo_lo_1323};
  wire [1023:0] dataGroup_hi_1323 = {dataGroup_hi_hi_1323, dataGroup_hi_lo_1323};
  wire [15:0]   dataGroup_11_46 = dataGroup_lo_1323[895:880];
  wire [1023:0] dataGroup_lo_1324 = {dataGroup_lo_hi_1324, dataGroup_lo_lo_1324};
  wire [1023:0] dataGroup_hi_1324 = {dataGroup_hi_hi_1324, dataGroup_hi_lo_1324};
  wire [15:0]   dataGroup_12_46 = dataGroup_lo_1324[975:960];
  wire [1023:0] dataGroup_lo_1325 = {dataGroup_lo_hi_1325, dataGroup_lo_lo_1325};
  wire [1023:0] dataGroup_hi_1325 = {dataGroup_hi_hi_1325, dataGroup_hi_lo_1325};
  wire [15:0]   dataGroup_13_46 = dataGroup_hi_1325[31:16];
  wire [1023:0] dataGroup_lo_1326 = {dataGroup_lo_hi_1326, dataGroup_lo_lo_1326};
  wire [1023:0] dataGroup_hi_1326 = {dataGroup_hi_hi_1326, dataGroup_hi_lo_1326};
  wire [15:0]   dataGroup_14_46 = dataGroup_hi_1326[111:96];
  wire [1023:0] dataGroup_lo_1327 = {dataGroup_lo_hi_1327, dataGroup_lo_lo_1327};
  wire [1023:0] dataGroup_hi_1327 = {dataGroup_hi_hi_1327, dataGroup_hi_lo_1327};
  wire [15:0]   dataGroup_15_46 = dataGroup_hi_1327[191:176];
  wire [31:0]   res_lo_lo_lo_46 = {dataGroup_1_46, dataGroup_0_46};
  wire [31:0]   res_lo_lo_hi_46 = {dataGroup_3_46, dataGroup_2_46};
  wire [63:0]   res_lo_lo_46 = {res_lo_lo_hi_46, res_lo_lo_lo_46};
  wire [31:0]   res_lo_hi_lo_46 = {dataGroup_5_46, dataGroup_4_46};
  wire [31:0]   res_lo_hi_hi_46 = {dataGroup_7_46, dataGroup_6_46};
  wire [63:0]   res_lo_hi_46 = {res_lo_hi_hi_46, res_lo_hi_lo_46};
  wire [127:0]  res_lo_46 = {res_lo_hi_46, res_lo_lo_46};
  wire [31:0]   res_hi_lo_lo_46 = {dataGroup_9_46, dataGroup_8_46};
  wire [31:0]   res_hi_lo_hi_46 = {dataGroup_11_46, dataGroup_10_46};
  wire [63:0]   res_hi_lo_46 = {res_hi_lo_hi_46, res_hi_lo_lo_46};
  wire [31:0]   res_hi_hi_lo_46 = {dataGroup_13_46, dataGroup_12_46};
  wire [31:0]   res_hi_hi_hi_46 = {dataGroup_15_46, dataGroup_14_46};
  wire [63:0]   res_hi_hi_46 = {res_hi_hi_hi_46, res_hi_hi_lo_46};
  wire [127:0]  res_hi_46 = {res_hi_hi_46, res_hi_lo_46};
  wire [255:0]  res_96 = {res_hi_46, res_lo_46};
  wire [1023:0] dataGroup_lo_1328 = {dataGroup_lo_hi_1328, dataGroup_lo_lo_1328};
  wire [1023:0] dataGroup_hi_1328 = {dataGroup_hi_hi_1328, dataGroup_hi_lo_1328};
  wire [15:0]   dataGroup_0_47 = dataGroup_lo_1328[31:16];
  wire [1023:0] dataGroup_lo_1329 = {dataGroup_lo_hi_1329, dataGroup_lo_lo_1329};
  wire [1023:0] dataGroup_hi_1329 = {dataGroup_hi_hi_1329, dataGroup_hi_lo_1329};
  wire [15:0]   dataGroup_1_47 = dataGroup_lo_1329[111:96];
  wire [1023:0] dataGroup_lo_1330 = {dataGroup_lo_hi_1330, dataGroup_lo_lo_1330};
  wire [1023:0] dataGroup_hi_1330 = {dataGroup_hi_hi_1330, dataGroup_hi_lo_1330};
  wire [15:0]   dataGroup_2_47 = dataGroup_lo_1330[191:176];
  wire [1023:0] dataGroup_lo_1331 = {dataGroup_lo_hi_1331, dataGroup_lo_lo_1331};
  wire [1023:0] dataGroup_hi_1331 = {dataGroup_hi_hi_1331, dataGroup_hi_lo_1331};
  wire [15:0]   dataGroup_3_47 = dataGroup_lo_1331[271:256];
  wire [1023:0] dataGroup_lo_1332 = {dataGroup_lo_hi_1332, dataGroup_lo_lo_1332};
  wire [1023:0] dataGroup_hi_1332 = {dataGroup_hi_hi_1332, dataGroup_hi_lo_1332};
  wire [15:0]   dataGroup_4_47 = dataGroup_lo_1332[351:336];
  wire [1023:0] dataGroup_lo_1333 = {dataGroup_lo_hi_1333, dataGroup_lo_lo_1333};
  wire [1023:0] dataGroup_hi_1333 = {dataGroup_hi_hi_1333, dataGroup_hi_lo_1333};
  wire [15:0]   dataGroup_5_47 = dataGroup_lo_1333[431:416];
  wire [1023:0] dataGroup_lo_1334 = {dataGroup_lo_hi_1334, dataGroup_lo_lo_1334};
  wire [1023:0] dataGroup_hi_1334 = {dataGroup_hi_hi_1334, dataGroup_hi_lo_1334};
  wire [15:0]   dataGroup_6_47 = dataGroup_lo_1334[511:496];
  wire [1023:0] dataGroup_lo_1335 = {dataGroup_lo_hi_1335, dataGroup_lo_lo_1335};
  wire [1023:0] dataGroup_hi_1335 = {dataGroup_hi_hi_1335, dataGroup_hi_lo_1335};
  wire [15:0]   dataGroup_7_47 = dataGroup_lo_1335[591:576];
  wire [1023:0] dataGroup_lo_1336 = {dataGroup_lo_hi_1336, dataGroup_lo_lo_1336};
  wire [1023:0] dataGroup_hi_1336 = {dataGroup_hi_hi_1336, dataGroup_hi_lo_1336};
  wire [15:0]   dataGroup_8_47 = dataGroup_lo_1336[671:656];
  wire [1023:0] dataGroup_lo_1337 = {dataGroup_lo_hi_1337, dataGroup_lo_lo_1337};
  wire [1023:0] dataGroup_hi_1337 = {dataGroup_hi_hi_1337, dataGroup_hi_lo_1337};
  wire [15:0]   dataGroup_9_47 = dataGroup_lo_1337[751:736];
  wire [1023:0] dataGroup_lo_1338 = {dataGroup_lo_hi_1338, dataGroup_lo_lo_1338};
  wire [1023:0] dataGroup_hi_1338 = {dataGroup_hi_hi_1338, dataGroup_hi_lo_1338};
  wire [15:0]   dataGroup_10_47 = dataGroup_lo_1338[831:816];
  wire [1023:0] dataGroup_lo_1339 = {dataGroup_lo_hi_1339, dataGroup_lo_lo_1339};
  wire [1023:0] dataGroup_hi_1339 = {dataGroup_hi_hi_1339, dataGroup_hi_lo_1339};
  wire [15:0]   dataGroup_11_47 = dataGroup_lo_1339[911:896];
  wire [1023:0] dataGroup_lo_1340 = {dataGroup_lo_hi_1340, dataGroup_lo_lo_1340};
  wire [1023:0] dataGroup_hi_1340 = {dataGroup_hi_hi_1340, dataGroup_hi_lo_1340};
  wire [15:0]   dataGroup_12_47 = dataGroup_lo_1340[991:976];
  wire [1023:0] dataGroup_lo_1341 = {dataGroup_lo_hi_1341, dataGroup_lo_lo_1341};
  wire [1023:0] dataGroup_hi_1341 = {dataGroup_hi_hi_1341, dataGroup_hi_lo_1341};
  wire [15:0]   dataGroup_13_47 = dataGroup_hi_1341[47:32];
  wire [1023:0] dataGroup_lo_1342 = {dataGroup_lo_hi_1342, dataGroup_lo_lo_1342};
  wire [1023:0] dataGroup_hi_1342 = {dataGroup_hi_hi_1342, dataGroup_hi_lo_1342};
  wire [15:0]   dataGroup_14_47 = dataGroup_hi_1342[127:112];
  wire [1023:0] dataGroup_lo_1343 = {dataGroup_lo_hi_1343, dataGroup_lo_lo_1343};
  wire [1023:0] dataGroup_hi_1343 = {dataGroup_hi_hi_1343, dataGroup_hi_lo_1343};
  wire [15:0]   dataGroup_15_47 = dataGroup_hi_1343[207:192];
  wire [31:0]   res_lo_lo_lo_47 = {dataGroup_1_47, dataGroup_0_47};
  wire [31:0]   res_lo_lo_hi_47 = {dataGroup_3_47, dataGroup_2_47};
  wire [63:0]   res_lo_lo_47 = {res_lo_lo_hi_47, res_lo_lo_lo_47};
  wire [31:0]   res_lo_hi_lo_47 = {dataGroup_5_47, dataGroup_4_47};
  wire [31:0]   res_lo_hi_hi_47 = {dataGroup_7_47, dataGroup_6_47};
  wire [63:0]   res_lo_hi_47 = {res_lo_hi_hi_47, res_lo_hi_lo_47};
  wire [127:0]  res_lo_47 = {res_lo_hi_47, res_lo_lo_47};
  wire [31:0]   res_hi_lo_lo_47 = {dataGroup_9_47, dataGroup_8_47};
  wire [31:0]   res_hi_lo_hi_47 = {dataGroup_11_47, dataGroup_10_47};
  wire [63:0]   res_hi_lo_47 = {res_hi_lo_hi_47, res_hi_lo_lo_47};
  wire [31:0]   res_hi_hi_lo_47 = {dataGroup_13_47, dataGroup_12_47};
  wire [31:0]   res_hi_hi_hi_47 = {dataGroup_15_47, dataGroup_14_47};
  wire [63:0]   res_hi_hi_47 = {res_hi_hi_hi_47, res_hi_hi_lo_47};
  wire [127:0]  res_hi_47 = {res_hi_hi_47, res_hi_lo_47};
  wire [255:0]  res_97 = {res_hi_47, res_lo_47};
  wire [1023:0] dataGroup_lo_1344 = {dataGroup_lo_hi_1344, dataGroup_lo_lo_1344};
  wire [1023:0] dataGroup_hi_1344 = {dataGroup_hi_hi_1344, dataGroup_hi_lo_1344};
  wire [15:0]   dataGroup_0_48 = dataGroup_lo_1344[47:32];
  wire [1023:0] dataGroup_lo_1345 = {dataGroup_lo_hi_1345, dataGroup_lo_lo_1345};
  wire [1023:0] dataGroup_hi_1345 = {dataGroup_hi_hi_1345, dataGroup_hi_lo_1345};
  wire [15:0]   dataGroup_1_48 = dataGroup_lo_1345[127:112];
  wire [1023:0] dataGroup_lo_1346 = {dataGroup_lo_hi_1346, dataGroup_lo_lo_1346};
  wire [1023:0] dataGroup_hi_1346 = {dataGroup_hi_hi_1346, dataGroup_hi_lo_1346};
  wire [15:0]   dataGroup_2_48 = dataGroup_lo_1346[207:192];
  wire [1023:0] dataGroup_lo_1347 = {dataGroup_lo_hi_1347, dataGroup_lo_lo_1347};
  wire [1023:0] dataGroup_hi_1347 = {dataGroup_hi_hi_1347, dataGroup_hi_lo_1347};
  wire [15:0]   dataGroup_3_48 = dataGroup_lo_1347[287:272];
  wire [1023:0] dataGroup_lo_1348 = {dataGroup_lo_hi_1348, dataGroup_lo_lo_1348};
  wire [1023:0] dataGroup_hi_1348 = {dataGroup_hi_hi_1348, dataGroup_hi_lo_1348};
  wire [15:0]   dataGroup_4_48 = dataGroup_lo_1348[367:352];
  wire [1023:0] dataGroup_lo_1349 = {dataGroup_lo_hi_1349, dataGroup_lo_lo_1349};
  wire [1023:0] dataGroup_hi_1349 = {dataGroup_hi_hi_1349, dataGroup_hi_lo_1349};
  wire [15:0]   dataGroup_5_48 = dataGroup_lo_1349[447:432];
  wire [1023:0] dataGroup_lo_1350 = {dataGroup_lo_hi_1350, dataGroup_lo_lo_1350};
  wire [1023:0] dataGroup_hi_1350 = {dataGroup_hi_hi_1350, dataGroup_hi_lo_1350};
  wire [15:0]   dataGroup_6_48 = dataGroup_lo_1350[527:512];
  wire [1023:0] dataGroup_lo_1351 = {dataGroup_lo_hi_1351, dataGroup_lo_lo_1351};
  wire [1023:0] dataGroup_hi_1351 = {dataGroup_hi_hi_1351, dataGroup_hi_lo_1351};
  wire [15:0]   dataGroup_7_48 = dataGroup_lo_1351[607:592];
  wire [1023:0] dataGroup_lo_1352 = {dataGroup_lo_hi_1352, dataGroup_lo_lo_1352};
  wire [1023:0] dataGroup_hi_1352 = {dataGroup_hi_hi_1352, dataGroup_hi_lo_1352};
  wire [15:0]   dataGroup_8_48 = dataGroup_lo_1352[687:672];
  wire [1023:0] dataGroup_lo_1353 = {dataGroup_lo_hi_1353, dataGroup_lo_lo_1353};
  wire [1023:0] dataGroup_hi_1353 = {dataGroup_hi_hi_1353, dataGroup_hi_lo_1353};
  wire [15:0]   dataGroup_9_48 = dataGroup_lo_1353[767:752];
  wire [1023:0] dataGroup_lo_1354 = {dataGroup_lo_hi_1354, dataGroup_lo_lo_1354};
  wire [1023:0] dataGroup_hi_1354 = {dataGroup_hi_hi_1354, dataGroup_hi_lo_1354};
  wire [15:0]   dataGroup_10_48 = dataGroup_lo_1354[847:832];
  wire [1023:0] dataGroup_lo_1355 = {dataGroup_lo_hi_1355, dataGroup_lo_lo_1355};
  wire [1023:0] dataGroup_hi_1355 = {dataGroup_hi_hi_1355, dataGroup_hi_lo_1355};
  wire [15:0]   dataGroup_11_48 = dataGroup_lo_1355[927:912];
  wire [1023:0] dataGroup_lo_1356 = {dataGroup_lo_hi_1356, dataGroup_lo_lo_1356};
  wire [1023:0] dataGroup_hi_1356 = {dataGroup_hi_hi_1356, dataGroup_hi_lo_1356};
  wire [15:0]   dataGroup_12_48 = dataGroup_lo_1356[1007:992];
  wire [1023:0] dataGroup_lo_1357 = {dataGroup_lo_hi_1357, dataGroup_lo_lo_1357};
  wire [1023:0] dataGroup_hi_1357 = {dataGroup_hi_hi_1357, dataGroup_hi_lo_1357};
  wire [15:0]   dataGroup_13_48 = dataGroup_hi_1357[63:48];
  wire [1023:0] dataGroup_lo_1358 = {dataGroup_lo_hi_1358, dataGroup_lo_lo_1358};
  wire [1023:0] dataGroup_hi_1358 = {dataGroup_hi_hi_1358, dataGroup_hi_lo_1358};
  wire [15:0]   dataGroup_14_48 = dataGroup_hi_1358[143:128];
  wire [1023:0] dataGroup_lo_1359 = {dataGroup_lo_hi_1359, dataGroup_lo_lo_1359};
  wire [1023:0] dataGroup_hi_1359 = {dataGroup_hi_hi_1359, dataGroup_hi_lo_1359};
  wire [15:0]   dataGroup_15_48 = dataGroup_hi_1359[223:208];
  wire [31:0]   res_lo_lo_lo_48 = {dataGroup_1_48, dataGroup_0_48};
  wire [31:0]   res_lo_lo_hi_48 = {dataGroup_3_48, dataGroup_2_48};
  wire [63:0]   res_lo_lo_48 = {res_lo_lo_hi_48, res_lo_lo_lo_48};
  wire [31:0]   res_lo_hi_lo_48 = {dataGroup_5_48, dataGroup_4_48};
  wire [31:0]   res_lo_hi_hi_48 = {dataGroup_7_48, dataGroup_6_48};
  wire [63:0]   res_lo_hi_48 = {res_lo_hi_hi_48, res_lo_hi_lo_48};
  wire [127:0]  res_lo_48 = {res_lo_hi_48, res_lo_lo_48};
  wire [31:0]   res_hi_lo_lo_48 = {dataGroup_9_48, dataGroup_8_48};
  wire [31:0]   res_hi_lo_hi_48 = {dataGroup_11_48, dataGroup_10_48};
  wire [63:0]   res_hi_lo_48 = {res_hi_lo_hi_48, res_hi_lo_lo_48};
  wire [31:0]   res_hi_hi_lo_48 = {dataGroup_13_48, dataGroup_12_48};
  wire [31:0]   res_hi_hi_hi_48 = {dataGroup_15_48, dataGroup_14_48};
  wire [63:0]   res_hi_hi_48 = {res_hi_hi_hi_48, res_hi_hi_lo_48};
  wire [127:0]  res_hi_48 = {res_hi_hi_48, res_hi_lo_48};
  wire [255:0]  res_98 = {res_hi_48, res_lo_48};
  wire [1023:0] dataGroup_lo_1360 = {dataGroup_lo_hi_1360, dataGroup_lo_lo_1360};
  wire [1023:0] dataGroup_hi_1360 = {dataGroup_hi_hi_1360, dataGroup_hi_lo_1360};
  wire [15:0]   dataGroup_0_49 = dataGroup_lo_1360[63:48];
  wire [1023:0] dataGroup_lo_1361 = {dataGroup_lo_hi_1361, dataGroup_lo_lo_1361};
  wire [1023:0] dataGroup_hi_1361 = {dataGroup_hi_hi_1361, dataGroup_hi_lo_1361};
  wire [15:0]   dataGroup_1_49 = dataGroup_lo_1361[143:128];
  wire [1023:0] dataGroup_lo_1362 = {dataGroup_lo_hi_1362, dataGroup_lo_lo_1362};
  wire [1023:0] dataGroup_hi_1362 = {dataGroup_hi_hi_1362, dataGroup_hi_lo_1362};
  wire [15:0]   dataGroup_2_49 = dataGroup_lo_1362[223:208];
  wire [1023:0] dataGroup_lo_1363 = {dataGroup_lo_hi_1363, dataGroup_lo_lo_1363};
  wire [1023:0] dataGroup_hi_1363 = {dataGroup_hi_hi_1363, dataGroup_hi_lo_1363};
  wire [15:0]   dataGroup_3_49 = dataGroup_lo_1363[303:288];
  wire [1023:0] dataGroup_lo_1364 = {dataGroup_lo_hi_1364, dataGroup_lo_lo_1364};
  wire [1023:0] dataGroup_hi_1364 = {dataGroup_hi_hi_1364, dataGroup_hi_lo_1364};
  wire [15:0]   dataGroup_4_49 = dataGroup_lo_1364[383:368];
  wire [1023:0] dataGroup_lo_1365 = {dataGroup_lo_hi_1365, dataGroup_lo_lo_1365};
  wire [1023:0] dataGroup_hi_1365 = {dataGroup_hi_hi_1365, dataGroup_hi_lo_1365};
  wire [15:0]   dataGroup_5_49 = dataGroup_lo_1365[463:448];
  wire [1023:0] dataGroup_lo_1366 = {dataGroup_lo_hi_1366, dataGroup_lo_lo_1366};
  wire [1023:0] dataGroup_hi_1366 = {dataGroup_hi_hi_1366, dataGroup_hi_lo_1366};
  wire [15:0]   dataGroup_6_49 = dataGroup_lo_1366[543:528];
  wire [1023:0] dataGroup_lo_1367 = {dataGroup_lo_hi_1367, dataGroup_lo_lo_1367};
  wire [1023:0] dataGroup_hi_1367 = {dataGroup_hi_hi_1367, dataGroup_hi_lo_1367};
  wire [15:0]   dataGroup_7_49 = dataGroup_lo_1367[623:608];
  wire [1023:0] dataGroup_lo_1368 = {dataGroup_lo_hi_1368, dataGroup_lo_lo_1368};
  wire [1023:0] dataGroup_hi_1368 = {dataGroup_hi_hi_1368, dataGroup_hi_lo_1368};
  wire [15:0]   dataGroup_8_49 = dataGroup_lo_1368[703:688];
  wire [1023:0] dataGroup_lo_1369 = {dataGroup_lo_hi_1369, dataGroup_lo_lo_1369};
  wire [1023:0] dataGroup_hi_1369 = {dataGroup_hi_hi_1369, dataGroup_hi_lo_1369};
  wire [15:0]   dataGroup_9_49 = dataGroup_lo_1369[783:768];
  wire [1023:0] dataGroup_lo_1370 = {dataGroup_lo_hi_1370, dataGroup_lo_lo_1370};
  wire [1023:0] dataGroup_hi_1370 = {dataGroup_hi_hi_1370, dataGroup_hi_lo_1370};
  wire [15:0]   dataGroup_10_49 = dataGroup_lo_1370[863:848];
  wire [1023:0] dataGroup_lo_1371 = {dataGroup_lo_hi_1371, dataGroup_lo_lo_1371};
  wire [1023:0] dataGroup_hi_1371 = {dataGroup_hi_hi_1371, dataGroup_hi_lo_1371};
  wire [15:0]   dataGroup_11_49 = dataGroup_lo_1371[943:928];
  wire [1023:0] dataGroup_lo_1372 = {dataGroup_lo_hi_1372, dataGroup_lo_lo_1372};
  wire [1023:0] dataGroup_hi_1372 = {dataGroup_hi_hi_1372, dataGroup_hi_lo_1372};
  wire [15:0]   dataGroup_12_49 = dataGroup_lo_1372[1023:1008];
  wire [1023:0] dataGroup_lo_1373 = {dataGroup_lo_hi_1373, dataGroup_lo_lo_1373};
  wire [1023:0] dataGroup_hi_1373 = {dataGroup_hi_hi_1373, dataGroup_hi_lo_1373};
  wire [15:0]   dataGroup_13_49 = dataGroup_hi_1373[79:64];
  wire [1023:0] dataGroup_lo_1374 = {dataGroup_lo_hi_1374, dataGroup_lo_lo_1374};
  wire [1023:0] dataGroup_hi_1374 = {dataGroup_hi_hi_1374, dataGroup_hi_lo_1374};
  wire [15:0]   dataGroup_14_49 = dataGroup_hi_1374[159:144];
  wire [1023:0] dataGroup_lo_1375 = {dataGroup_lo_hi_1375, dataGroup_lo_lo_1375};
  wire [1023:0] dataGroup_hi_1375 = {dataGroup_hi_hi_1375, dataGroup_hi_lo_1375};
  wire [15:0]   dataGroup_15_49 = dataGroup_hi_1375[239:224];
  wire [31:0]   res_lo_lo_lo_49 = {dataGroup_1_49, dataGroup_0_49};
  wire [31:0]   res_lo_lo_hi_49 = {dataGroup_3_49, dataGroup_2_49};
  wire [63:0]   res_lo_lo_49 = {res_lo_lo_hi_49, res_lo_lo_lo_49};
  wire [31:0]   res_lo_hi_lo_49 = {dataGroup_5_49, dataGroup_4_49};
  wire [31:0]   res_lo_hi_hi_49 = {dataGroup_7_49, dataGroup_6_49};
  wire [63:0]   res_lo_hi_49 = {res_lo_hi_hi_49, res_lo_hi_lo_49};
  wire [127:0]  res_lo_49 = {res_lo_hi_49, res_lo_lo_49};
  wire [31:0]   res_hi_lo_lo_49 = {dataGroup_9_49, dataGroup_8_49};
  wire [31:0]   res_hi_lo_hi_49 = {dataGroup_11_49, dataGroup_10_49};
  wire [63:0]   res_hi_lo_49 = {res_hi_lo_hi_49, res_hi_lo_lo_49};
  wire [31:0]   res_hi_hi_lo_49 = {dataGroup_13_49, dataGroup_12_49};
  wire [31:0]   res_hi_hi_hi_49 = {dataGroup_15_49, dataGroup_14_49};
  wire [63:0]   res_hi_hi_49 = {res_hi_hi_hi_49, res_hi_hi_lo_49};
  wire [127:0]  res_hi_49 = {res_hi_hi_49, res_hi_lo_49};
  wire [255:0]  res_99 = {res_hi_49, res_lo_49};
  wire [1023:0] dataGroup_lo_1376 = {dataGroup_lo_hi_1376, dataGroup_lo_lo_1376};
  wire [1023:0] dataGroup_hi_1376 = {dataGroup_hi_hi_1376, dataGroup_hi_lo_1376};
  wire [15:0]   dataGroup_0_50 = dataGroup_lo_1376[79:64];
  wire [1023:0] dataGroup_lo_1377 = {dataGroup_lo_hi_1377, dataGroup_lo_lo_1377};
  wire [1023:0] dataGroup_hi_1377 = {dataGroup_hi_hi_1377, dataGroup_hi_lo_1377};
  wire [15:0]   dataGroup_1_50 = dataGroup_lo_1377[159:144];
  wire [1023:0] dataGroup_lo_1378 = {dataGroup_lo_hi_1378, dataGroup_lo_lo_1378};
  wire [1023:0] dataGroup_hi_1378 = {dataGroup_hi_hi_1378, dataGroup_hi_lo_1378};
  wire [15:0]   dataGroup_2_50 = dataGroup_lo_1378[239:224];
  wire [1023:0] dataGroup_lo_1379 = {dataGroup_lo_hi_1379, dataGroup_lo_lo_1379};
  wire [1023:0] dataGroup_hi_1379 = {dataGroup_hi_hi_1379, dataGroup_hi_lo_1379};
  wire [15:0]   dataGroup_3_50 = dataGroup_lo_1379[319:304];
  wire [1023:0] dataGroup_lo_1380 = {dataGroup_lo_hi_1380, dataGroup_lo_lo_1380};
  wire [1023:0] dataGroup_hi_1380 = {dataGroup_hi_hi_1380, dataGroup_hi_lo_1380};
  wire [15:0]   dataGroup_4_50 = dataGroup_lo_1380[399:384];
  wire [1023:0] dataGroup_lo_1381 = {dataGroup_lo_hi_1381, dataGroup_lo_lo_1381};
  wire [1023:0] dataGroup_hi_1381 = {dataGroup_hi_hi_1381, dataGroup_hi_lo_1381};
  wire [15:0]   dataGroup_5_50 = dataGroup_lo_1381[479:464];
  wire [1023:0] dataGroup_lo_1382 = {dataGroup_lo_hi_1382, dataGroup_lo_lo_1382};
  wire [1023:0] dataGroup_hi_1382 = {dataGroup_hi_hi_1382, dataGroup_hi_lo_1382};
  wire [15:0]   dataGroup_6_50 = dataGroup_lo_1382[559:544];
  wire [1023:0] dataGroup_lo_1383 = {dataGroup_lo_hi_1383, dataGroup_lo_lo_1383};
  wire [1023:0] dataGroup_hi_1383 = {dataGroup_hi_hi_1383, dataGroup_hi_lo_1383};
  wire [15:0]   dataGroup_7_50 = dataGroup_lo_1383[639:624];
  wire [1023:0] dataGroup_lo_1384 = {dataGroup_lo_hi_1384, dataGroup_lo_lo_1384};
  wire [1023:0] dataGroup_hi_1384 = {dataGroup_hi_hi_1384, dataGroup_hi_lo_1384};
  wire [15:0]   dataGroup_8_50 = dataGroup_lo_1384[719:704];
  wire [1023:0] dataGroup_lo_1385 = {dataGroup_lo_hi_1385, dataGroup_lo_lo_1385};
  wire [1023:0] dataGroup_hi_1385 = {dataGroup_hi_hi_1385, dataGroup_hi_lo_1385};
  wire [15:0]   dataGroup_9_50 = dataGroup_lo_1385[799:784];
  wire [1023:0] dataGroup_lo_1386 = {dataGroup_lo_hi_1386, dataGroup_lo_lo_1386};
  wire [1023:0] dataGroup_hi_1386 = {dataGroup_hi_hi_1386, dataGroup_hi_lo_1386};
  wire [15:0]   dataGroup_10_50 = dataGroup_lo_1386[879:864];
  wire [1023:0] dataGroup_lo_1387 = {dataGroup_lo_hi_1387, dataGroup_lo_lo_1387};
  wire [1023:0] dataGroup_hi_1387 = {dataGroup_hi_hi_1387, dataGroup_hi_lo_1387};
  wire [15:0]   dataGroup_11_50 = dataGroup_lo_1387[959:944];
  wire [1023:0] dataGroup_lo_1388 = {dataGroup_lo_hi_1388, dataGroup_lo_lo_1388};
  wire [1023:0] dataGroup_hi_1388 = {dataGroup_hi_hi_1388, dataGroup_hi_lo_1388};
  wire [15:0]   dataGroup_12_50 = dataGroup_hi_1388[15:0];
  wire [1023:0] dataGroup_lo_1389 = {dataGroup_lo_hi_1389, dataGroup_lo_lo_1389};
  wire [1023:0] dataGroup_hi_1389 = {dataGroup_hi_hi_1389, dataGroup_hi_lo_1389};
  wire [15:0]   dataGroup_13_50 = dataGroup_hi_1389[95:80];
  wire [1023:0] dataGroup_lo_1390 = {dataGroup_lo_hi_1390, dataGroup_lo_lo_1390};
  wire [1023:0] dataGroup_hi_1390 = {dataGroup_hi_hi_1390, dataGroup_hi_lo_1390};
  wire [15:0]   dataGroup_14_50 = dataGroup_hi_1390[175:160];
  wire [1023:0] dataGroup_lo_1391 = {dataGroup_lo_hi_1391, dataGroup_lo_lo_1391};
  wire [1023:0] dataGroup_hi_1391 = {dataGroup_hi_hi_1391, dataGroup_hi_lo_1391};
  wire [15:0]   dataGroup_15_50 = dataGroup_hi_1391[255:240];
  wire [31:0]   res_lo_lo_lo_50 = {dataGroup_1_50, dataGroup_0_50};
  wire [31:0]   res_lo_lo_hi_50 = {dataGroup_3_50, dataGroup_2_50};
  wire [63:0]   res_lo_lo_50 = {res_lo_lo_hi_50, res_lo_lo_lo_50};
  wire [31:0]   res_lo_hi_lo_50 = {dataGroup_5_50, dataGroup_4_50};
  wire [31:0]   res_lo_hi_hi_50 = {dataGroup_7_50, dataGroup_6_50};
  wire [63:0]   res_lo_hi_50 = {res_lo_hi_hi_50, res_lo_hi_lo_50};
  wire [127:0]  res_lo_50 = {res_lo_hi_50, res_lo_lo_50};
  wire [31:0]   res_hi_lo_lo_50 = {dataGroup_9_50, dataGroup_8_50};
  wire [31:0]   res_hi_lo_hi_50 = {dataGroup_11_50, dataGroup_10_50};
  wire [63:0]   res_hi_lo_50 = {res_hi_lo_hi_50, res_hi_lo_lo_50};
  wire [31:0]   res_hi_hi_lo_50 = {dataGroup_13_50, dataGroup_12_50};
  wire [31:0]   res_hi_hi_hi_50 = {dataGroup_15_50, dataGroup_14_50};
  wire [63:0]   res_hi_hi_50 = {res_hi_hi_hi_50, res_hi_hi_lo_50};
  wire [127:0]  res_hi_50 = {res_hi_hi_50, res_hi_lo_50};
  wire [255:0]  res_100 = {res_hi_50, res_lo_50};
  wire [511:0]  lo_lo_12 = {res_97, res_96};
  wire [511:0]  lo_hi_12 = {res_99, res_98};
  wire [1023:0] lo_12 = {lo_hi_12, lo_lo_12};
  wire [511:0]  hi_lo_12 = {256'h0, res_100};
  wire [1023:0] hi_12 = {512'h0, hi_lo_12};
  wire [2047:0] regroupLoadData_1_4 = {hi_12, lo_12};
  wire [1023:0] dataGroup_lo_1392 = {dataGroup_lo_hi_1392, dataGroup_lo_lo_1392};
  wire [1023:0] dataGroup_hi_1392 = {dataGroup_hi_hi_1392, dataGroup_hi_lo_1392};
  wire [15:0]   dataGroup_0_51 = dataGroup_lo_1392[15:0];
  wire [1023:0] dataGroup_lo_1393 = {dataGroup_lo_hi_1393, dataGroup_lo_lo_1393};
  wire [1023:0] dataGroup_hi_1393 = {dataGroup_hi_hi_1393, dataGroup_hi_lo_1393};
  wire [15:0]   dataGroup_1_51 = dataGroup_lo_1393[111:96];
  wire [1023:0] dataGroup_lo_1394 = {dataGroup_lo_hi_1394, dataGroup_lo_lo_1394};
  wire [1023:0] dataGroup_hi_1394 = {dataGroup_hi_hi_1394, dataGroup_hi_lo_1394};
  wire [15:0]   dataGroup_2_51 = dataGroup_lo_1394[207:192];
  wire [1023:0] dataGroup_lo_1395 = {dataGroup_lo_hi_1395, dataGroup_lo_lo_1395};
  wire [1023:0] dataGroup_hi_1395 = {dataGroup_hi_hi_1395, dataGroup_hi_lo_1395};
  wire [15:0]   dataGroup_3_51 = dataGroup_lo_1395[303:288];
  wire [1023:0] dataGroup_lo_1396 = {dataGroup_lo_hi_1396, dataGroup_lo_lo_1396};
  wire [1023:0] dataGroup_hi_1396 = {dataGroup_hi_hi_1396, dataGroup_hi_lo_1396};
  wire [15:0]   dataGroup_4_51 = dataGroup_lo_1396[399:384];
  wire [1023:0] dataGroup_lo_1397 = {dataGroup_lo_hi_1397, dataGroup_lo_lo_1397};
  wire [1023:0] dataGroup_hi_1397 = {dataGroup_hi_hi_1397, dataGroup_hi_lo_1397};
  wire [15:0]   dataGroup_5_51 = dataGroup_lo_1397[495:480];
  wire [1023:0] dataGroup_lo_1398 = {dataGroup_lo_hi_1398, dataGroup_lo_lo_1398};
  wire [1023:0] dataGroup_hi_1398 = {dataGroup_hi_hi_1398, dataGroup_hi_lo_1398};
  wire [15:0]   dataGroup_6_51 = dataGroup_lo_1398[591:576];
  wire [1023:0] dataGroup_lo_1399 = {dataGroup_lo_hi_1399, dataGroup_lo_lo_1399};
  wire [1023:0] dataGroup_hi_1399 = {dataGroup_hi_hi_1399, dataGroup_hi_lo_1399};
  wire [15:0]   dataGroup_7_51 = dataGroup_lo_1399[687:672];
  wire [1023:0] dataGroup_lo_1400 = {dataGroup_lo_hi_1400, dataGroup_lo_lo_1400};
  wire [1023:0] dataGroup_hi_1400 = {dataGroup_hi_hi_1400, dataGroup_hi_lo_1400};
  wire [15:0]   dataGroup_8_51 = dataGroup_lo_1400[783:768];
  wire [1023:0] dataGroup_lo_1401 = {dataGroup_lo_hi_1401, dataGroup_lo_lo_1401};
  wire [1023:0] dataGroup_hi_1401 = {dataGroup_hi_hi_1401, dataGroup_hi_lo_1401};
  wire [15:0]   dataGroup_9_51 = dataGroup_lo_1401[879:864];
  wire [1023:0] dataGroup_lo_1402 = {dataGroup_lo_hi_1402, dataGroup_lo_lo_1402};
  wire [1023:0] dataGroup_hi_1402 = {dataGroup_hi_hi_1402, dataGroup_hi_lo_1402};
  wire [15:0]   dataGroup_10_51 = dataGroup_lo_1402[975:960];
  wire [1023:0] dataGroup_lo_1403 = {dataGroup_lo_hi_1403, dataGroup_lo_lo_1403};
  wire [1023:0] dataGroup_hi_1403 = {dataGroup_hi_hi_1403, dataGroup_hi_lo_1403};
  wire [15:0]   dataGroup_11_51 = dataGroup_hi_1403[47:32];
  wire [1023:0] dataGroup_lo_1404 = {dataGroup_lo_hi_1404, dataGroup_lo_lo_1404};
  wire [1023:0] dataGroup_hi_1404 = {dataGroup_hi_hi_1404, dataGroup_hi_lo_1404};
  wire [15:0]   dataGroup_12_51 = dataGroup_hi_1404[143:128];
  wire [1023:0] dataGroup_lo_1405 = {dataGroup_lo_hi_1405, dataGroup_lo_lo_1405};
  wire [1023:0] dataGroup_hi_1405 = {dataGroup_hi_hi_1405, dataGroup_hi_lo_1405};
  wire [15:0]   dataGroup_13_51 = dataGroup_hi_1405[239:224];
  wire [1023:0] dataGroup_lo_1406 = {dataGroup_lo_hi_1406, dataGroup_lo_lo_1406};
  wire [1023:0] dataGroup_hi_1406 = {dataGroup_hi_hi_1406, dataGroup_hi_lo_1406};
  wire [15:0]   dataGroup_14_51 = dataGroup_hi_1406[335:320];
  wire [1023:0] dataGroup_lo_1407 = {dataGroup_lo_hi_1407, dataGroup_lo_lo_1407};
  wire [1023:0] dataGroup_hi_1407 = {dataGroup_hi_hi_1407, dataGroup_hi_lo_1407};
  wire [15:0]   dataGroup_15_51 = dataGroup_hi_1407[431:416];
  wire [31:0]   res_lo_lo_lo_51 = {dataGroup_1_51, dataGroup_0_51};
  wire [31:0]   res_lo_lo_hi_51 = {dataGroup_3_51, dataGroup_2_51};
  wire [63:0]   res_lo_lo_51 = {res_lo_lo_hi_51, res_lo_lo_lo_51};
  wire [31:0]   res_lo_hi_lo_51 = {dataGroup_5_51, dataGroup_4_51};
  wire [31:0]   res_lo_hi_hi_51 = {dataGroup_7_51, dataGroup_6_51};
  wire [63:0]   res_lo_hi_51 = {res_lo_hi_hi_51, res_lo_hi_lo_51};
  wire [127:0]  res_lo_51 = {res_lo_hi_51, res_lo_lo_51};
  wire [31:0]   res_hi_lo_lo_51 = {dataGroup_9_51, dataGroup_8_51};
  wire [31:0]   res_hi_lo_hi_51 = {dataGroup_11_51, dataGroup_10_51};
  wire [63:0]   res_hi_lo_51 = {res_hi_lo_hi_51, res_hi_lo_lo_51};
  wire [31:0]   res_hi_hi_lo_51 = {dataGroup_13_51, dataGroup_12_51};
  wire [31:0]   res_hi_hi_hi_51 = {dataGroup_15_51, dataGroup_14_51};
  wire [63:0]   res_hi_hi_51 = {res_hi_hi_hi_51, res_hi_hi_lo_51};
  wire [127:0]  res_hi_51 = {res_hi_hi_51, res_hi_lo_51};
  wire [255:0]  res_104 = {res_hi_51, res_lo_51};
  wire [1023:0] dataGroup_lo_1408 = {dataGroup_lo_hi_1408, dataGroup_lo_lo_1408};
  wire [1023:0] dataGroup_hi_1408 = {dataGroup_hi_hi_1408, dataGroup_hi_lo_1408};
  wire [15:0]   dataGroup_0_52 = dataGroup_lo_1408[31:16];
  wire [1023:0] dataGroup_lo_1409 = {dataGroup_lo_hi_1409, dataGroup_lo_lo_1409};
  wire [1023:0] dataGroup_hi_1409 = {dataGroup_hi_hi_1409, dataGroup_hi_lo_1409};
  wire [15:0]   dataGroup_1_52 = dataGroup_lo_1409[127:112];
  wire [1023:0] dataGroup_lo_1410 = {dataGroup_lo_hi_1410, dataGroup_lo_lo_1410};
  wire [1023:0] dataGroup_hi_1410 = {dataGroup_hi_hi_1410, dataGroup_hi_lo_1410};
  wire [15:0]   dataGroup_2_52 = dataGroup_lo_1410[223:208];
  wire [1023:0] dataGroup_lo_1411 = {dataGroup_lo_hi_1411, dataGroup_lo_lo_1411};
  wire [1023:0] dataGroup_hi_1411 = {dataGroup_hi_hi_1411, dataGroup_hi_lo_1411};
  wire [15:0]   dataGroup_3_52 = dataGroup_lo_1411[319:304];
  wire [1023:0] dataGroup_lo_1412 = {dataGroup_lo_hi_1412, dataGroup_lo_lo_1412};
  wire [1023:0] dataGroup_hi_1412 = {dataGroup_hi_hi_1412, dataGroup_hi_lo_1412};
  wire [15:0]   dataGroup_4_52 = dataGroup_lo_1412[415:400];
  wire [1023:0] dataGroup_lo_1413 = {dataGroup_lo_hi_1413, dataGroup_lo_lo_1413};
  wire [1023:0] dataGroup_hi_1413 = {dataGroup_hi_hi_1413, dataGroup_hi_lo_1413};
  wire [15:0]   dataGroup_5_52 = dataGroup_lo_1413[511:496];
  wire [1023:0] dataGroup_lo_1414 = {dataGroup_lo_hi_1414, dataGroup_lo_lo_1414};
  wire [1023:0] dataGroup_hi_1414 = {dataGroup_hi_hi_1414, dataGroup_hi_lo_1414};
  wire [15:0]   dataGroup_6_52 = dataGroup_lo_1414[607:592];
  wire [1023:0] dataGroup_lo_1415 = {dataGroup_lo_hi_1415, dataGroup_lo_lo_1415};
  wire [1023:0] dataGroup_hi_1415 = {dataGroup_hi_hi_1415, dataGroup_hi_lo_1415};
  wire [15:0]   dataGroup_7_52 = dataGroup_lo_1415[703:688];
  wire [1023:0] dataGroup_lo_1416 = {dataGroup_lo_hi_1416, dataGroup_lo_lo_1416};
  wire [1023:0] dataGroup_hi_1416 = {dataGroup_hi_hi_1416, dataGroup_hi_lo_1416};
  wire [15:0]   dataGroup_8_52 = dataGroup_lo_1416[799:784];
  wire [1023:0] dataGroup_lo_1417 = {dataGroup_lo_hi_1417, dataGroup_lo_lo_1417};
  wire [1023:0] dataGroup_hi_1417 = {dataGroup_hi_hi_1417, dataGroup_hi_lo_1417};
  wire [15:0]   dataGroup_9_52 = dataGroup_lo_1417[895:880];
  wire [1023:0] dataGroup_lo_1418 = {dataGroup_lo_hi_1418, dataGroup_lo_lo_1418};
  wire [1023:0] dataGroup_hi_1418 = {dataGroup_hi_hi_1418, dataGroup_hi_lo_1418};
  wire [15:0]   dataGroup_10_52 = dataGroup_lo_1418[991:976];
  wire [1023:0] dataGroup_lo_1419 = {dataGroup_lo_hi_1419, dataGroup_lo_lo_1419};
  wire [1023:0] dataGroup_hi_1419 = {dataGroup_hi_hi_1419, dataGroup_hi_lo_1419};
  wire [15:0]   dataGroup_11_52 = dataGroup_hi_1419[63:48];
  wire [1023:0] dataGroup_lo_1420 = {dataGroup_lo_hi_1420, dataGroup_lo_lo_1420};
  wire [1023:0] dataGroup_hi_1420 = {dataGroup_hi_hi_1420, dataGroup_hi_lo_1420};
  wire [15:0]   dataGroup_12_52 = dataGroup_hi_1420[159:144];
  wire [1023:0] dataGroup_lo_1421 = {dataGroup_lo_hi_1421, dataGroup_lo_lo_1421};
  wire [1023:0] dataGroup_hi_1421 = {dataGroup_hi_hi_1421, dataGroup_hi_lo_1421};
  wire [15:0]   dataGroup_13_52 = dataGroup_hi_1421[255:240];
  wire [1023:0] dataGroup_lo_1422 = {dataGroup_lo_hi_1422, dataGroup_lo_lo_1422};
  wire [1023:0] dataGroup_hi_1422 = {dataGroup_hi_hi_1422, dataGroup_hi_lo_1422};
  wire [15:0]   dataGroup_14_52 = dataGroup_hi_1422[351:336];
  wire [1023:0] dataGroup_lo_1423 = {dataGroup_lo_hi_1423, dataGroup_lo_lo_1423};
  wire [1023:0] dataGroup_hi_1423 = {dataGroup_hi_hi_1423, dataGroup_hi_lo_1423};
  wire [15:0]   dataGroup_15_52 = dataGroup_hi_1423[447:432];
  wire [31:0]   res_lo_lo_lo_52 = {dataGroup_1_52, dataGroup_0_52};
  wire [31:0]   res_lo_lo_hi_52 = {dataGroup_3_52, dataGroup_2_52};
  wire [63:0]   res_lo_lo_52 = {res_lo_lo_hi_52, res_lo_lo_lo_52};
  wire [31:0]   res_lo_hi_lo_52 = {dataGroup_5_52, dataGroup_4_52};
  wire [31:0]   res_lo_hi_hi_52 = {dataGroup_7_52, dataGroup_6_52};
  wire [63:0]   res_lo_hi_52 = {res_lo_hi_hi_52, res_lo_hi_lo_52};
  wire [127:0]  res_lo_52 = {res_lo_hi_52, res_lo_lo_52};
  wire [31:0]   res_hi_lo_lo_52 = {dataGroup_9_52, dataGroup_8_52};
  wire [31:0]   res_hi_lo_hi_52 = {dataGroup_11_52, dataGroup_10_52};
  wire [63:0]   res_hi_lo_52 = {res_hi_lo_hi_52, res_hi_lo_lo_52};
  wire [31:0]   res_hi_hi_lo_52 = {dataGroup_13_52, dataGroup_12_52};
  wire [31:0]   res_hi_hi_hi_52 = {dataGroup_15_52, dataGroup_14_52};
  wire [63:0]   res_hi_hi_52 = {res_hi_hi_hi_52, res_hi_hi_lo_52};
  wire [127:0]  res_hi_52 = {res_hi_hi_52, res_hi_lo_52};
  wire [255:0]  res_105 = {res_hi_52, res_lo_52};
  wire [1023:0] dataGroup_lo_1424 = {dataGroup_lo_hi_1424, dataGroup_lo_lo_1424};
  wire [1023:0] dataGroup_hi_1424 = {dataGroup_hi_hi_1424, dataGroup_hi_lo_1424};
  wire [15:0]   dataGroup_0_53 = dataGroup_lo_1424[47:32];
  wire [1023:0] dataGroup_lo_1425 = {dataGroup_lo_hi_1425, dataGroup_lo_lo_1425};
  wire [1023:0] dataGroup_hi_1425 = {dataGroup_hi_hi_1425, dataGroup_hi_lo_1425};
  wire [15:0]   dataGroup_1_53 = dataGroup_lo_1425[143:128];
  wire [1023:0] dataGroup_lo_1426 = {dataGroup_lo_hi_1426, dataGroup_lo_lo_1426};
  wire [1023:0] dataGroup_hi_1426 = {dataGroup_hi_hi_1426, dataGroup_hi_lo_1426};
  wire [15:0]   dataGroup_2_53 = dataGroup_lo_1426[239:224];
  wire [1023:0] dataGroup_lo_1427 = {dataGroup_lo_hi_1427, dataGroup_lo_lo_1427};
  wire [1023:0] dataGroup_hi_1427 = {dataGroup_hi_hi_1427, dataGroup_hi_lo_1427};
  wire [15:0]   dataGroup_3_53 = dataGroup_lo_1427[335:320];
  wire [1023:0] dataGroup_lo_1428 = {dataGroup_lo_hi_1428, dataGroup_lo_lo_1428};
  wire [1023:0] dataGroup_hi_1428 = {dataGroup_hi_hi_1428, dataGroup_hi_lo_1428};
  wire [15:0]   dataGroup_4_53 = dataGroup_lo_1428[431:416];
  wire [1023:0] dataGroup_lo_1429 = {dataGroup_lo_hi_1429, dataGroup_lo_lo_1429};
  wire [1023:0] dataGroup_hi_1429 = {dataGroup_hi_hi_1429, dataGroup_hi_lo_1429};
  wire [15:0]   dataGroup_5_53 = dataGroup_lo_1429[527:512];
  wire [1023:0] dataGroup_lo_1430 = {dataGroup_lo_hi_1430, dataGroup_lo_lo_1430};
  wire [1023:0] dataGroup_hi_1430 = {dataGroup_hi_hi_1430, dataGroup_hi_lo_1430};
  wire [15:0]   dataGroup_6_53 = dataGroup_lo_1430[623:608];
  wire [1023:0] dataGroup_lo_1431 = {dataGroup_lo_hi_1431, dataGroup_lo_lo_1431};
  wire [1023:0] dataGroup_hi_1431 = {dataGroup_hi_hi_1431, dataGroup_hi_lo_1431};
  wire [15:0]   dataGroup_7_53 = dataGroup_lo_1431[719:704];
  wire [1023:0] dataGroup_lo_1432 = {dataGroup_lo_hi_1432, dataGroup_lo_lo_1432};
  wire [1023:0] dataGroup_hi_1432 = {dataGroup_hi_hi_1432, dataGroup_hi_lo_1432};
  wire [15:0]   dataGroup_8_53 = dataGroup_lo_1432[815:800];
  wire [1023:0] dataGroup_lo_1433 = {dataGroup_lo_hi_1433, dataGroup_lo_lo_1433};
  wire [1023:0] dataGroup_hi_1433 = {dataGroup_hi_hi_1433, dataGroup_hi_lo_1433};
  wire [15:0]   dataGroup_9_53 = dataGroup_lo_1433[911:896];
  wire [1023:0] dataGroup_lo_1434 = {dataGroup_lo_hi_1434, dataGroup_lo_lo_1434};
  wire [1023:0] dataGroup_hi_1434 = {dataGroup_hi_hi_1434, dataGroup_hi_lo_1434};
  wire [15:0]   dataGroup_10_53 = dataGroup_lo_1434[1007:992];
  wire [1023:0] dataGroup_lo_1435 = {dataGroup_lo_hi_1435, dataGroup_lo_lo_1435};
  wire [1023:0] dataGroup_hi_1435 = {dataGroup_hi_hi_1435, dataGroup_hi_lo_1435};
  wire [15:0]   dataGroup_11_53 = dataGroup_hi_1435[79:64];
  wire [1023:0] dataGroup_lo_1436 = {dataGroup_lo_hi_1436, dataGroup_lo_lo_1436};
  wire [1023:0] dataGroup_hi_1436 = {dataGroup_hi_hi_1436, dataGroup_hi_lo_1436};
  wire [15:0]   dataGroup_12_53 = dataGroup_hi_1436[175:160];
  wire [1023:0] dataGroup_lo_1437 = {dataGroup_lo_hi_1437, dataGroup_lo_lo_1437};
  wire [1023:0] dataGroup_hi_1437 = {dataGroup_hi_hi_1437, dataGroup_hi_lo_1437};
  wire [15:0]   dataGroup_13_53 = dataGroup_hi_1437[271:256];
  wire [1023:0] dataGroup_lo_1438 = {dataGroup_lo_hi_1438, dataGroup_lo_lo_1438};
  wire [1023:0] dataGroup_hi_1438 = {dataGroup_hi_hi_1438, dataGroup_hi_lo_1438};
  wire [15:0]   dataGroup_14_53 = dataGroup_hi_1438[367:352];
  wire [1023:0] dataGroup_lo_1439 = {dataGroup_lo_hi_1439, dataGroup_lo_lo_1439};
  wire [1023:0] dataGroup_hi_1439 = {dataGroup_hi_hi_1439, dataGroup_hi_lo_1439};
  wire [15:0]   dataGroup_15_53 = dataGroup_hi_1439[463:448];
  wire [31:0]   res_lo_lo_lo_53 = {dataGroup_1_53, dataGroup_0_53};
  wire [31:0]   res_lo_lo_hi_53 = {dataGroup_3_53, dataGroup_2_53};
  wire [63:0]   res_lo_lo_53 = {res_lo_lo_hi_53, res_lo_lo_lo_53};
  wire [31:0]   res_lo_hi_lo_53 = {dataGroup_5_53, dataGroup_4_53};
  wire [31:0]   res_lo_hi_hi_53 = {dataGroup_7_53, dataGroup_6_53};
  wire [63:0]   res_lo_hi_53 = {res_lo_hi_hi_53, res_lo_hi_lo_53};
  wire [127:0]  res_lo_53 = {res_lo_hi_53, res_lo_lo_53};
  wire [31:0]   res_hi_lo_lo_53 = {dataGroup_9_53, dataGroup_8_53};
  wire [31:0]   res_hi_lo_hi_53 = {dataGroup_11_53, dataGroup_10_53};
  wire [63:0]   res_hi_lo_53 = {res_hi_lo_hi_53, res_hi_lo_lo_53};
  wire [31:0]   res_hi_hi_lo_53 = {dataGroup_13_53, dataGroup_12_53};
  wire [31:0]   res_hi_hi_hi_53 = {dataGroup_15_53, dataGroup_14_53};
  wire [63:0]   res_hi_hi_53 = {res_hi_hi_hi_53, res_hi_hi_lo_53};
  wire [127:0]  res_hi_53 = {res_hi_hi_53, res_hi_lo_53};
  wire [255:0]  res_106 = {res_hi_53, res_lo_53};
  wire [1023:0] dataGroup_lo_1440 = {dataGroup_lo_hi_1440, dataGroup_lo_lo_1440};
  wire [1023:0] dataGroup_hi_1440 = {dataGroup_hi_hi_1440, dataGroup_hi_lo_1440};
  wire [15:0]   dataGroup_0_54 = dataGroup_lo_1440[63:48];
  wire [1023:0] dataGroup_lo_1441 = {dataGroup_lo_hi_1441, dataGroup_lo_lo_1441};
  wire [1023:0] dataGroup_hi_1441 = {dataGroup_hi_hi_1441, dataGroup_hi_lo_1441};
  wire [15:0]   dataGroup_1_54 = dataGroup_lo_1441[159:144];
  wire [1023:0] dataGroup_lo_1442 = {dataGroup_lo_hi_1442, dataGroup_lo_lo_1442};
  wire [1023:0] dataGroup_hi_1442 = {dataGroup_hi_hi_1442, dataGroup_hi_lo_1442};
  wire [15:0]   dataGroup_2_54 = dataGroup_lo_1442[255:240];
  wire [1023:0] dataGroup_lo_1443 = {dataGroup_lo_hi_1443, dataGroup_lo_lo_1443};
  wire [1023:0] dataGroup_hi_1443 = {dataGroup_hi_hi_1443, dataGroup_hi_lo_1443};
  wire [15:0]   dataGroup_3_54 = dataGroup_lo_1443[351:336];
  wire [1023:0] dataGroup_lo_1444 = {dataGroup_lo_hi_1444, dataGroup_lo_lo_1444};
  wire [1023:0] dataGroup_hi_1444 = {dataGroup_hi_hi_1444, dataGroup_hi_lo_1444};
  wire [15:0]   dataGroup_4_54 = dataGroup_lo_1444[447:432];
  wire [1023:0] dataGroup_lo_1445 = {dataGroup_lo_hi_1445, dataGroup_lo_lo_1445};
  wire [1023:0] dataGroup_hi_1445 = {dataGroup_hi_hi_1445, dataGroup_hi_lo_1445};
  wire [15:0]   dataGroup_5_54 = dataGroup_lo_1445[543:528];
  wire [1023:0] dataGroup_lo_1446 = {dataGroup_lo_hi_1446, dataGroup_lo_lo_1446};
  wire [1023:0] dataGroup_hi_1446 = {dataGroup_hi_hi_1446, dataGroup_hi_lo_1446};
  wire [15:0]   dataGroup_6_54 = dataGroup_lo_1446[639:624];
  wire [1023:0] dataGroup_lo_1447 = {dataGroup_lo_hi_1447, dataGroup_lo_lo_1447};
  wire [1023:0] dataGroup_hi_1447 = {dataGroup_hi_hi_1447, dataGroup_hi_lo_1447};
  wire [15:0]   dataGroup_7_54 = dataGroup_lo_1447[735:720];
  wire [1023:0] dataGroup_lo_1448 = {dataGroup_lo_hi_1448, dataGroup_lo_lo_1448};
  wire [1023:0] dataGroup_hi_1448 = {dataGroup_hi_hi_1448, dataGroup_hi_lo_1448};
  wire [15:0]   dataGroup_8_54 = dataGroup_lo_1448[831:816];
  wire [1023:0] dataGroup_lo_1449 = {dataGroup_lo_hi_1449, dataGroup_lo_lo_1449};
  wire [1023:0] dataGroup_hi_1449 = {dataGroup_hi_hi_1449, dataGroup_hi_lo_1449};
  wire [15:0]   dataGroup_9_54 = dataGroup_lo_1449[927:912];
  wire [1023:0] dataGroup_lo_1450 = {dataGroup_lo_hi_1450, dataGroup_lo_lo_1450};
  wire [1023:0] dataGroup_hi_1450 = {dataGroup_hi_hi_1450, dataGroup_hi_lo_1450};
  wire [15:0]   dataGroup_10_54 = dataGroup_lo_1450[1023:1008];
  wire [1023:0] dataGroup_lo_1451 = {dataGroup_lo_hi_1451, dataGroup_lo_lo_1451};
  wire [1023:0] dataGroup_hi_1451 = {dataGroup_hi_hi_1451, dataGroup_hi_lo_1451};
  wire [15:0]   dataGroup_11_54 = dataGroup_hi_1451[95:80];
  wire [1023:0] dataGroup_lo_1452 = {dataGroup_lo_hi_1452, dataGroup_lo_lo_1452};
  wire [1023:0] dataGroup_hi_1452 = {dataGroup_hi_hi_1452, dataGroup_hi_lo_1452};
  wire [15:0]   dataGroup_12_54 = dataGroup_hi_1452[191:176];
  wire [1023:0] dataGroup_lo_1453 = {dataGroup_lo_hi_1453, dataGroup_lo_lo_1453};
  wire [1023:0] dataGroup_hi_1453 = {dataGroup_hi_hi_1453, dataGroup_hi_lo_1453};
  wire [15:0]   dataGroup_13_54 = dataGroup_hi_1453[287:272];
  wire [1023:0] dataGroup_lo_1454 = {dataGroup_lo_hi_1454, dataGroup_lo_lo_1454};
  wire [1023:0] dataGroup_hi_1454 = {dataGroup_hi_hi_1454, dataGroup_hi_lo_1454};
  wire [15:0]   dataGroup_14_54 = dataGroup_hi_1454[383:368];
  wire [1023:0] dataGroup_lo_1455 = {dataGroup_lo_hi_1455, dataGroup_lo_lo_1455};
  wire [1023:0] dataGroup_hi_1455 = {dataGroup_hi_hi_1455, dataGroup_hi_lo_1455};
  wire [15:0]   dataGroup_15_54 = dataGroup_hi_1455[479:464];
  wire [31:0]   res_lo_lo_lo_54 = {dataGroup_1_54, dataGroup_0_54};
  wire [31:0]   res_lo_lo_hi_54 = {dataGroup_3_54, dataGroup_2_54};
  wire [63:0]   res_lo_lo_54 = {res_lo_lo_hi_54, res_lo_lo_lo_54};
  wire [31:0]   res_lo_hi_lo_54 = {dataGroup_5_54, dataGroup_4_54};
  wire [31:0]   res_lo_hi_hi_54 = {dataGroup_7_54, dataGroup_6_54};
  wire [63:0]   res_lo_hi_54 = {res_lo_hi_hi_54, res_lo_hi_lo_54};
  wire [127:0]  res_lo_54 = {res_lo_hi_54, res_lo_lo_54};
  wire [31:0]   res_hi_lo_lo_54 = {dataGroup_9_54, dataGroup_8_54};
  wire [31:0]   res_hi_lo_hi_54 = {dataGroup_11_54, dataGroup_10_54};
  wire [63:0]   res_hi_lo_54 = {res_hi_lo_hi_54, res_hi_lo_lo_54};
  wire [31:0]   res_hi_hi_lo_54 = {dataGroup_13_54, dataGroup_12_54};
  wire [31:0]   res_hi_hi_hi_54 = {dataGroup_15_54, dataGroup_14_54};
  wire [63:0]   res_hi_hi_54 = {res_hi_hi_hi_54, res_hi_hi_lo_54};
  wire [127:0]  res_hi_54 = {res_hi_hi_54, res_hi_lo_54};
  wire [255:0]  res_107 = {res_hi_54, res_lo_54};
  wire [1023:0] dataGroup_lo_1456 = {dataGroup_lo_hi_1456, dataGroup_lo_lo_1456};
  wire [1023:0] dataGroup_hi_1456 = {dataGroup_hi_hi_1456, dataGroup_hi_lo_1456};
  wire [15:0]   dataGroup_0_55 = dataGroup_lo_1456[79:64];
  wire [1023:0] dataGroup_lo_1457 = {dataGroup_lo_hi_1457, dataGroup_lo_lo_1457};
  wire [1023:0] dataGroup_hi_1457 = {dataGroup_hi_hi_1457, dataGroup_hi_lo_1457};
  wire [15:0]   dataGroup_1_55 = dataGroup_lo_1457[175:160];
  wire [1023:0] dataGroup_lo_1458 = {dataGroup_lo_hi_1458, dataGroup_lo_lo_1458};
  wire [1023:0] dataGroup_hi_1458 = {dataGroup_hi_hi_1458, dataGroup_hi_lo_1458};
  wire [15:0]   dataGroup_2_55 = dataGroup_lo_1458[271:256];
  wire [1023:0] dataGroup_lo_1459 = {dataGroup_lo_hi_1459, dataGroup_lo_lo_1459};
  wire [1023:0] dataGroup_hi_1459 = {dataGroup_hi_hi_1459, dataGroup_hi_lo_1459};
  wire [15:0]   dataGroup_3_55 = dataGroup_lo_1459[367:352];
  wire [1023:0] dataGroup_lo_1460 = {dataGroup_lo_hi_1460, dataGroup_lo_lo_1460};
  wire [1023:0] dataGroup_hi_1460 = {dataGroup_hi_hi_1460, dataGroup_hi_lo_1460};
  wire [15:0]   dataGroup_4_55 = dataGroup_lo_1460[463:448];
  wire [1023:0] dataGroup_lo_1461 = {dataGroup_lo_hi_1461, dataGroup_lo_lo_1461};
  wire [1023:0] dataGroup_hi_1461 = {dataGroup_hi_hi_1461, dataGroup_hi_lo_1461};
  wire [15:0]   dataGroup_5_55 = dataGroup_lo_1461[559:544];
  wire [1023:0] dataGroup_lo_1462 = {dataGroup_lo_hi_1462, dataGroup_lo_lo_1462};
  wire [1023:0] dataGroup_hi_1462 = {dataGroup_hi_hi_1462, dataGroup_hi_lo_1462};
  wire [15:0]   dataGroup_6_55 = dataGroup_lo_1462[655:640];
  wire [1023:0] dataGroup_lo_1463 = {dataGroup_lo_hi_1463, dataGroup_lo_lo_1463};
  wire [1023:0] dataGroup_hi_1463 = {dataGroup_hi_hi_1463, dataGroup_hi_lo_1463};
  wire [15:0]   dataGroup_7_55 = dataGroup_lo_1463[751:736];
  wire [1023:0] dataGroup_lo_1464 = {dataGroup_lo_hi_1464, dataGroup_lo_lo_1464};
  wire [1023:0] dataGroup_hi_1464 = {dataGroup_hi_hi_1464, dataGroup_hi_lo_1464};
  wire [15:0]   dataGroup_8_55 = dataGroup_lo_1464[847:832];
  wire [1023:0] dataGroup_lo_1465 = {dataGroup_lo_hi_1465, dataGroup_lo_lo_1465};
  wire [1023:0] dataGroup_hi_1465 = {dataGroup_hi_hi_1465, dataGroup_hi_lo_1465};
  wire [15:0]   dataGroup_9_55 = dataGroup_lo_1465[943:928];
  wire [1023:0] dataGroup_lo_1466 = {dataGroup_lo_hi_1466, dataGroup_lo_lo_1466};
  wire [1023:0] dataGroup_hi_1466 = {dataGroup_hi_hi_1466, dataGroup_hi_lo_1466};
  wire [15:0]   dataGroup_10_55 = dataGroup_hi_1466[15:0];
  wire [1023:0] dataGroup_lo_1467 = {dataGroup_lo_hi_1467, dataGroup_lo_lo_1467};
  wire [1023:0] dataGroup_hi_1467 = {dataGroup_hi_hi_1467, dataGroup_hi_lo_1467};
  wire [15:0]   dataGroup_11_55 = dataGroup_hi_1467[111:96];
  wire [1023:0] dataGroup_lo_1468 = {dataGroup_lo_hi_1468, dataGroup_lo_lo_1468};
  wire [1023:0] dataGroup_hi_1468 = {dataGroup_hi_hi_1468, dataGroup_hi_lo_1468};
  wire [15:0]   dataGroup_12_55 = dataGroup_hi_1468[207:192];
  wire [1023:0] dataGroup_lo_1469 = {dataGroup_lo_hi_1469, dataGroup_lo_lo_1469};
  wire [1023:0] dataGroup_hi_1469 = {dataGroup_hi_hi_1469, dataGroup_hi_lo_1469};
  wire [15:0]   dataGroup_13_55 = dataGroup_hi_1469[303:288];
  wire [1023:0] dataGroup_lo_1470 = {dataGroup_lo_hi_1470, dataGroup_lo_lo_1470};
  wire [1023:0] dataGroup_hi_1470 = {dataGroup_hi_hi_1470, dataGroup_hi_lo_1470};
  wire [15:0]   dataGroup_14_55 = dataGroup_hi_1470[399:384];
  wire [1023:0] dataGroup_lo_1471 = {dataGroup_lo_hi_1471, dataGroup_lo_lo_1471};
  wire [1023:0] dataGroup_hi_1471 = {dataGroup_hi_hi_1471, dataGroup_hi_lo_1471};
  wire [15:0]   dataGroup_15_55 = dataGroup_hi_1471[495:480];
  wire [31:0]   res_lo_lo_lo_55 = {dataGroup_1_55, dataGroup_0_55};
  wire [31:0]   res_lo_lo_hi_55 = {dataGroup_3_55, dataGroup_2_55};
  wire [63:0]   res_lo_lo_55 = {res_lo_lo_hi_55, res_lo_lo_lo_55};
  wire [31:0]   res_lo_hi_lo_55 = {dataGroup_5_55, dataGroup_4_55};
  wire [31:0]   res_lo_hi_hi_55 = {dataGroup_7_55, dataGroup_6_55};
  wire [63:0]   res_lo_hi_55 = {res_lo_hi_hi_55, res_lo_hi_lo_55};
  wire [127:0]  res_lo_55 = {res_lo_hi_55, res_lo_lo_55};
  wire [31:0]   res_hi_lo_lo_55 = {dataGroup_9_55, dataGroup_8_55};
  wire [31:0]   res_hi_lo_hi_55 = {dataGroup_11_55, dataGroup_10_55};
  wire [63:0]   res_hi_lo_55 = {res_hi_lo_hi_55, res_hi_lo_lo_55};
  wire [31:0]   res_hi_hi_lo_55 = {dataGroup_13_55, dataGroup_12_55};
  wire [31:0]   res_hi_hi_hi_55 = {dataGroup_15_55, dataGroup_14_55};
  wire [63:0]   res_hi_hi_55 = {res_hi_hi_hi_55, res_hi_hi_lo_55};
  wire [127:0]  res_hi_55 = {res_hi_hi_55, res_hi_lo_55};
  wire [255:0]  res_108 = {res_hi_55, res_lo_55};
  wire [1023:0] dataGroup_lo_1472 = {dataGroup_lo_hi_1472, dataGroup_lo_lo_1472};
  wire [1023:0] dataGroup_hi_1472 = {dataGroup_hi_hi_1472, dataGroup_hi_lo_1472};
  wire [15:0]   dataGroup_0_56 = dataGroup_lo_1472[95:80];
  wire [1023:0] dataGroup_lo_1473 = {dataGroup_lo_hi_1473, dataGroup_lo_lo_1473};
  wire [1023:0] dataGroup_hi_1473 = {dataGroup_hi_hi_1473, dataGroup_hi_lo_1473};
  wire [15:0]   dataGroup_1_56 = dataGroup_lo_1473[191:176];
  wire [1023:0] dataGroup_lo_1474 = {dataGroup_lo_hi_1474, dataGroup_lo_lo_1474};
  wire [1023:0] dataGroup_hi_1474 = {dataGroup_hi_hi_1474, dataGroup_hi_lo_1474};
  wire [15:0]   dataGroup_2_56 = dataGroup_lo_1474[287:272];
  wire [1023:0] dataGroup_lo_1475 = {dataGroup_lo_hi_1475, dataGroup_lo_lo_1475};
  wire [1023:0] dataGroup_hi_1475 = {dataGroup_hi_hi_1475, dataGroup_hi_lo_1475};
  wire [15:0]   dataGroup_3_56 = dataGroup_lo_1475[383:368];
  wire [1023:0] dataGroup_lo_1476 = {dataGroup_lo_hi_1476, dataGroup_lo_lo_1476};
  wire [1023:0] dataGroup_hi_1476 = {dataGroup_hi_hi_1476, dataGroup_hi_lo_1476};
  wire [15:0]   dataGroup_4_56 = dataGroup_lo_1476[479:464];
  wire [1023:0] dataGroup_lo_1477 = {dataGroup_lo_hi_1477, dataGroup_lo_lo_1477};
  wire [1023:0] dataGroup_hi_1477 = {dataGroup_hi_hi_1477, dataGroup_hi_lo_1477};
  wire [15:0]   dataGroup_5_56 = dataGroup_lo_1477[575:560];
  wire [1023:0] dataGroup_lo_1478 = {dataGroup_lo_hi_1478, dataGroup_lo_lo_1478};
  wire [1023:0] dataGroup_hi_1478 = {dataGroup_hi_hi_1478, dataGroup_hi_lo_1478};
  wire [15:0]   dataGroup_6_56 = dataGroup_lo_1478[671:656];
  wire [1023:0] dataGroup_lo_1479 = {dataGroup_lo_hi_1479, dataGroup_lo_lo_1479};
  wire [1023:0] dataGroup_hi_1479 = {dataGroup_hi_hi_1479, dataGroup_hi_lo_1479};
  wire [15:0]   dataGroup_7_56 = dataGroup_lo_1479[767:752];
  wire [1023:0] dataGroup_lo_1480 = {dataGroup_lo_hi_1480, dataGroup_lo_lo_1480};
  wire [1023:0] dataGroup_hi_1480 = {dataGroup_hi_hi_1480, dataGroup_hi_lo_1480};
  wire [15:0]   dataGroup_8_56 = dataGroup_lo_1480[863:848];
  wire [1023:0] dataGroup_lo_1481 = {dataGroup_lo_hi_1481, dataGroup_lo_lo_1481};
  wire [1023:0] dataGroup_hi_1481 = {dataGroup_hi_hi_1481, dataGroup_hi_lo_1481};
  wire [15:0]   dataGroup_9_56 = dataGroup_lo_1481[959:944];
  wire [1023:0] dataGroup_lo_1482 = {dataGroup_lo_hi_1482, dataGroup_lo_lo_1482};
  wire [1023:0] dataGroup_hi_1482 = {dataGroup_hi_hi_1482, dataGroup_hi_lo_1482};
  wire [15:0]   dataGroup_10_56 = dataGroup_hi_1482[31:16];
  wire [1023:0] dataGroup_lo_1483 = {dataGroup_lo_hi_1483, dataGroup_lo_lo_1483};
  wire [1023:0] dataGroup_hi_1483 = {dataGroup_hi_hi_1483, dataGroup_hi_lo_1483};
  wire [15:0]   dataGroup_11_56 = dataGroup_hi_1483[127:112];
  wire [1023:0] dataGroup_lo_1484 = {dataGroup_lo_hi_1484, dataGroup_lo_lo_1484};
  wire [1023:0] dataGroup_hi_1484 = {dataGroup_hi_hi_1484, dataGroup_hi_lo_1484};
  wire [15:0]   dataGroup_12_56 = dataGroup_hi_1484[223:208];
  wire [1023:0] dataGroup_lo_1485 = {dataGroup_lo_hi_1485, dataGroup_lo_lo_1485};
  wire [1023:0] dataGroup_hi_1485 = {dataGroup_hi_hi_1485, dataGroup_hi_lo_1485};
  wire [15:0]   dataGroup_13_56 = dataGroup_hi_1485[319:304];
  wire [1023:0] dataGroup_lo_1486 = {dataGroup_lo_hi_1486, dataGroup_lo_lo_1486};
  wire [1023:0] dataGroup_hi_1486 = {dataGroup_hi_hi_1486, dataGroup_hi_lo_1486};
  wire [15:0]   dataGroup_14_56 = dataGroup_hi_1486[415:400];
  wire [1023:0] dataGroup_lo_1487 = {dataGroup_lo_hi_1487, dataGroup_lo_lo_1487};
  wire [1023:0] dataGroup_hi_1487 = {dataGroup_hi_hi_1487, dataGroup_hi_lo_1487};
  wire [15:0]   dataGroup_15_56 = dataGroup_hi_1487[511:496];
  wire [31:0]   res_lo_lo_lo_56 = {dataGroup_1_56, dataGroup_0_56};
  wire [31:0]   res_lo_lo_hi_56 = {dataGroup_3_56, dataGroup_2_56};
  wire [63:0]   res_lo_lo_56 = {res_lo_lo_hi_56, res_lo_lo_lo_56};
  wire [31:0]   res_lo_hi_lo_56 = {dataGroup_5_56, dataGroup_4_56};
  wire [31:0]   res_lo_hi_hi_56 = {dataGroup_7_56, dataGroup_6_56};
  wire [63:0]   res_lo_hi_56 = {res_lo_hi_hi_56, res_lo_hi_lo_56};
  wire [127:0]  res_lo_56 = {res_lo_hi_56, res_lo_lo_56};
  wire [31:0]   res_hi_lo_lo_56 = {dataGroup_9_56, dataGroup_8_56};
  wire [31:0]   res_hi_lo_hi_56 = {dataGroup_11_56, dataGroup_10_56};
  wire [63:0]   res_hi_lo_56 = {res_hi_lo_hi_56, res_hi_lo_lo_56};
  wire [31:0]   res_hi_hi_lo_56 = {dataGroup_13_56, dataGroup_12_56};
  wire [31:0]   res_hi_hi_hi_56 = {dataGroup_15_56, dataGroup_14_56};
  wire [63:0]   res_hi_hi_56 = {res_hi_hi_hi_56, res_hi_hi_lo_56};
  wire [127:0]  res_hi_56 = {res_hi_hi_56, res_hi_lo_56};
  wire [255:0]  res_109 = {res_hi_56, res_lo_56};
  wire [511:0]  lo_lo_13 = {res_105, res_104};
  wire [511:0]  lo_hi_13 = {res_107, res_106};
  wire [1023:0] lo_13 = {lo_hi_13, lo_lo_13};
  wire [511:0]  hi_lo_13 = {res_109, res_108};
  wire [1023:0] hi_13 = {512'h0, hi_lo_13};
  wire [2047:0] regroupLoadData_1_5 = {hi_13, lo_13};
  wire [1023:0] dataGroup_lo_1488 = {dataGroup_lo_hi_1488, dataGroup_lo_lo_1488};
  wire [1023:0] dataGroup_hi_1488 = {dataGroup_hi_hi_1488, dataGroup_hi_lo_1488};
  wire [15:0]   dataGroup_0_57 = dataGroup_lo_1488[15:0];
  wire [1023:0] dataGroup_lo_1489 = {dataGroup_lo_hi_1489, dataGroup_lo_lo_1489};
  wire [1023:0] dataGroup_hi_1489 = {dataGroup_hi_hi_1489, dataGroup_hi_lo_1489};
  wire [15:0]   dataGroup_1_57 = dataGroup_lo_1489[127:112];
  wire [1023:0] dataGroup_lo_1490 = {dataGroup_lo_hi_1490, dataGroup_lo_lo_1490};
  wire [1023:0] dataGroup_hi_1490 = {dataGroup_hi_hi_1490, dataGroup_hi_lo_1490};
  wire [15:0]   dataGroup_2_57 = dataGroup_lo_1490[239:224];
  wire [1023:0] dataGroup_lo_1491 = {dataGroup_lo_hi_1491, dataGroup_lo_lo_1491};
  wire [1023:0] dataGroup_hi_1491 = {dataGroup_hi_hi_1491, dataGroup_hi_lo_1491};
  wire [15:0]   dataGroup_3_57 = dataGroup_lo_1491[351:336];
  wire [1023:0] dataGroup_lo_1492 = {dataGroup_lo_hi_1492, dataGroup_lo_lo_1492};
  wire [1023:0] dataGroup_hi_1492 = {dataGroup_hi_hi_1492, dataGroup_hi_lo_1492};
  wire [15:0]   dataGroup_4_57 = dataGroup_lo_1492[463:448];
  wire [1023:0] dataGroup_lo_1493 = {dataGroup_lo_hi_1493, dataGroup_lo_lo_1493};
  wire [1023:0] dataGroup_hi_1493 = {dataGroup_hi_hi_1493, dataGroup_hi_lo_1493};
  wire [15:0]   dataGroup_5_57 = dataGroup_lo_1493[575:560];
  wire [1023:0] dataGroup_lo_1494 = {dataGroup_lo_hi_1494, dataGroup_lo_lo_1494};
  wire [1023:0] dataGroup_hi_1494 = {dataGroup_hi_hi_1494, dataGroup_hi_lo_1494};
  wire [15:0]   dataGroup_6_57 = dataGroup_lo_1494[687:672];
  wire [1023:0] dataGroup_lo_1495 = {dataGroup_lo_hi_1495, dataGroup_lo_lo_1495};
  wire [1023:0] dataGroup_hi_1495 = {dataGroup_hi_hi_1495, dataGroup_hi_lo_1495};
  wire [15:0]   dataGroup_7_57 = dataGroup_lo_1495[799:784];
  wire [1023:0] dataGroup_lo_1496 = {dataGroup_lo_hi_1496, dataGroup_lo_lo_1496};
  wire [1023:0] dataGroup_hi_1496 = {dataGroup_hi_hi_1496, dataGroup_hi_lo_1496};
  wire [15:0]   dataGroup_8_57 = dataGroup_lo_1496[911:896];
  wire [1023:0] dataGroup_lo_1497 = {dataGroup_lo_hi_1497, dataGroup_lo_lo_1497};
  wire [1023:0] dataGroup_hi_1497 = {dataGroup_hi_hi_1497, dataGroup_hi_lo_1497};
  wire [15:0]   dataGroup_9_57 = dataGroup_lo_1497[1023:1008];
  wire [1023:0] dataGroup_lo_1498 = {dataGroup_lo_hi_1498, dataGroup_lo_lo_1498};
  wire [1023:0] dataGroup_hi_1498 = {dataGroup_hi_hi_1498, dataGroup_hi_lo_1498};
  wire [15:0]   dataGroup_10_57 = dataGroup_hi_1498[111:96];
  wire [1023:0] dataGroup_lo_1499 = {dataGroup_lo_hi_1499, dataGroup_lo_lo_1499};
  wire [1023:0] dataGroup_hi_1499 = {dataGroup_hi_hi_1499, dataGroup_hi_lo_1499};
  wire [15:0]   dataGroup_11_57 = dataGroup_hi_1499[223:208];
  wire [1023:0] dataGroup_lo_1500 = {dataGroup_lo_hi_1500, dataGroup_lo_lo_1500};
  wire [1023:0] dataGroup_hi_1500 = {dataGroup_hi_hi_1500, dataGroup_hi_lo_1500};
  wire [15:0]   dataGroup_12_57 = dataGroup_hi_1500[335:320];
  wire [1023:0] dataGroup_lo_1501 = {dataGroup_lo_hi_1501, dataGroup_lo_lo_1501};
  wire [1023:0] dataGroup_hi_1501 = {dataGroup_hi_hi_1501, dataGroup_hi_lo_1501};
  wire [15:0]   dataGroup_13_57 = dataGroup_hi_1501[447:432];
  wire [1023:0] dataGroup_lo_1502 = {dataGroup_lo_hi_1502, dataGroup_lo_lo_1502};
  wire [1023:0] dataGroup_hi_1502 = {dataGroup_hi_hi_1502, dataGroup_hi_lo_1502};
  wire [15:0]   dataGroup_14_57 = dataGroup_hi_1502[559:544];
  wire [1023:0] dataGroup_lo_1503 = {dataGroup_lo_hi_1503, dataGroup_lo_lo_1503};
  wire [1023:0] dataGroup_hi_1503 = {dataGroup_hi_hi_1503, dataGroup_hi_lo_1503};
  wire [15:0]   dataGroup_15_57 = dataGroup_hi_1503[671:656];
  wire [31:0]   res_lo_lo_lo_57 = {dataGroup_1_57, dataGroup_0_57};
  wire [31:0]   res_lo_lo_hi_57 = {dataGroup_3_57, dataGroup_2_57};
  wire [63:0]   res_lo_lo_57 = {res_lo_lo_hi_57, res_lo_lo_lo_57};
  wire [31:0]   res_lo_hi_lo_57 = {dataGroup_5_57, dataGroup_4_57};
  wire [31:0]   res_lo_hi_hi_57 = {dataGroup_7_57, dataGroup_6_57};
  wire [63:0]   res_lo_hi_57 = {res_lo_hi_hi_57, res_lo_hi_lo_57};
  wire [127:0]  res_lo_57 = {res_lo_hi_57, res_lo_lo_57};
  wire [31:0]   res_hi_lo_lo_57 = {dataGroup_9_57, dataGroup_8_57};
  wire [31:0]   res_hi_lo_hi_57 = {dataGroup_11_57, dataGroup_10_57};
  wire [63:0]   res_hi_lo_57 = {res_hi_lo_hi_57, res_hi_lo_lo_57};
  wire [31:0]   res_hi_hi_lo_57 = {dataGroup_13_57, dataGroup_12_57};
  wire [31:0]   res_hi_hi_hi_57 = {dataGroup_15_57, dataGroup_14_57};
  wire [63:0]   res_hi_hi_57 = {res_hi_hi_hi_57, res_hi_hi_lo_57};
  wire [127:0]  res_hi_57 = {res_hi_hi_57, res_hi_lo_57};
  wire [255:0]  res_112 = {res_hi_57, res_lo_57};
  wire [1023:0] dataGroup_lo_1504 = {dataGroup_lo_hi_1504, dataGroup_lo_lo_1504};
  wire [1023:0] dataGroup_hi_1504 = {dataGroup_hi_hi_1504, dataGroup_hi_lo_1504};
  wire [15:0]   dataGroup_0_58 = dataGroup_lo_1504[31:16];
  wire [1023:0] dataGroup_lo_1505 = {dataGroup_lo_hi_1505, dataGroup_lo_lo_1505};
  wire [1023:0] dataGroup_hi_1505 = {dataGroup_hi_hi_1505, dataGroup_hi_lo_1505};
  wire [15:0]   dataGroup_1_58 = dataGroup_lo_1505[143:128];
  wire [1023:0] dataGroup_lo_1506 = {dataGroup_lo_hi_1506, dataGroup_lo_lo_1506};
  wire [1023:0] dataGroup_hi_1506 = {dataGroup_hi_hi_1506, dataGroup_hi_lo_1506};
  wire [15:0]   dataGroup_2_58 = dataGroup_lo_1506[255:240];
  wire [1023:0] dataGroup_lo_1507 = {dataGroup_lo_hi_1507, dataGroup_lo_lo_1507};
  wire [1023:0] dataGroup_hi_1507 = {dataGroup_hi_hi_1507, dataGroup_hi_lo_1507};
  wire [15:0]   dataGroup_3_58 = dataGroup_lo_1507[367:352];
  wire [1023:0] dataGroup_lo_1508 = {dataGroup_lo_hi_1508, dataGroup_lo_lo_1508};
  wire [1023:0] dataGroup_hi_1508 = {dataGroup_hi_hi_1508, dataGroup_hi_lo_1508};
  wire [15:0]   dataGroup_4_58 = dataGroup_lo_1508[479:464];
  wire [1023:0] dataGroup_lo_1509 = {dataGroup_lo_hi_1509, dataGroup_lo_lo_1509};
  wire [1023:0] dataGroup_hi_1509 = {dataGroup_hi_hi_1509, dataGroup_hi_lo_1509};
  wire [15:0]   dataGroup_5_58 = dataGroup_lo_1509[591:576];
  wire [1023:0] dataGroup_lo_1510 = {dataGroup_lo_hi_1510, dataGroup_lo_lo_1510};
  wire [1023:0] dataGroup_hi_1510 = {dataGroup_hi_hi_1510, dataGroup_hi_lo_1510};
  wire [15:0]   dataGroup_6_58 = dataGroup_lo_1510[703:688];
  wire [1023:0] dataGroup_lo_1511 = {dataGroup_lo_hi_1511, dataGroup_lo_lo_1511};
  wire [1023:0] dataGroup_hi_1511 = {dataGroup_hi_hi_1511, dataGroup_hi_lo_1511};
  wire [15:0]   dataGroup_7_58 = dataGroup_lo_1511[815:800];
  wire [1023:0] dataGroup_lo_1512 = {dataGroup_lo_hi_1512, dataGroup_lo_lo_1512};
  wire [1023:0] dataGroup_hi_1512 = {dataGroup_hi_hi_1512, dataGroup_hi_lo_1512};
  wire [15:0]   dataGroup_8_58 = dataGroup_lo_1512[927:912];
  wire [1023:0] dataGroup_lo_1513 = {dataGroup_lo_hi_1513, dataGroup_lo_lo_1513};
  wire [1023:0] dataGroup_hi_1513 = {dataGroup_hi_hi_1513, dataGroup_hi_lo_1513};
  wire [15:0]   dataGroup_9_58 = dataGroup_hi_1513[15:0];
  wire [1023:0] dataGroup_lo_1514 = {dataGroup_lo_hi_1514, dataGroup_lo_lo_1514};
  wire [1023:0] dataGroup_hi_1514 = {dataGroup_hi_hi_1514, dataGroup_hi_lo_1514};
  wire [15:0]   dataGroup_10_58 = dataGroup_hi_1514[127:112];
  wire [1023:0] dataGroup_lo_1515 = {dataGroup_lo_hi_1515, dataGroup_lo_lo_1515};
  wire [1023:0] dataGroup_hi_1515 = {dataGroup_hi_hi_1515, dataGroup_hi_lo_1515};
  wire [15:0]   dataGroup_11_58 = dataGroup_hi_1515[239:224];
  wire [1023:0] dataGroup_lo_1516 = {dataGroup_lo_hi_1516, dataGroup_lo_lo_1516};
  wire [1023:0] dataGroup_hi_1516 = {dataGroup_hi_hi_1516, dataGroup_hi_lo_1516};
  wire [15:0]   dataGroup_12_58 = dataGroup_hi_1516[351:336];
  wire [1023:0] dataGroup_lo_1517 = {dataGroup_lo_hi_1517, dataGroup_lo_lo_1517};
  wire [1023:0] dataGroup_hi_1517 = {dataGroup_hi_hi_1517, dataGroup_hi_lo_1517};
  wire [15:0]   dataGroup_13_58 = dataGroup_hi_1517[463:448];
  wire [1023:0] dataGroup_lo_1518 = {dataGroup_lo_hi_1518, dataGroup_lo_lo_1518};
  wire [1023:0] dataGroup_hi_1518 = {dataGroup_hi_hi_1518, dataGroup_hi_lo_1518};
  wire [15:0]   dataGroup_14_58 = dataGroup_hi_1518[575:560];
  wire [1023:0] dataGroup_lo_1519 = {dataGroup_lo_hi_1519, dataGroup_lo_lo_1519};
  wire [1023:0] dataGroup_hi_1519 = {dataGroup_hi_hi_1519, dataGroup_hi_lo_1519};
  wire [15:0]   dataGroup_15_58 = dataGroup_hi_1519[687:672];
  wire [31:0]   res_lo_lo_lo_58 = {dataGroup_1_58, dataGroup_0_58};
  wire [31:0]   res_lo_lo_hi_58 = {dataGroup_3_58, dataGroup_2_58};
  wire [63:0]   res_lo_lo_58 = {res_lo_lo_hi_58, res_lo_lo_lo_58};
  wire [31:0]   res_lo_hi_lo_58 = {dataGroup_5_58, dataGroup_4_58};
  wire [31:0]   res_lo_hi_hi_58 = {dataGroup_7_58, dataGroup_6_58};
  wire [63:0]   res_lo_hi_58 = {res_lo_hi_hi_58, res_lo_hi_lo_58};
  wire [127:0]  res_lo_58 = {res_lo_hi_58, res_lo_lo_58};
  wire [31:0]   res_hi_lo_lo_58 = {dataGroup_9_58, dataGroup_8_58};
  wire [31:0]   res_hi_lo_hi_58 = {dataGroup_11_58, dataGroup_10_58};
  wire [63:0]   res_hi_lo_58 = {res_hi_lo_hi_58, res_hi_lo_lo_58};
  wire [31:0]   res_hi_hi_lo_58 = {dataGroup_13_58, dataGroup_12_58};
  wire [31:0]   res_hi_hi_hi_58 = {dataGroup_15_58, dataGroup_14_58};
  wire [63:0]   res_hi_hi_58 = {res_hi_hi_hi_58, res_hi_hi_lo_58};
  wire [127:0]  res_hi_58 = {res_hi_hi_58, res_hi_lo_58};
  wire [255:0]  res_113 = {res_hi_58, res_lo_58};
  wire [1023:0] dataGroup_lo_1520 = {dataGroup_lo_hi_1520, dataGroup_lo_lo_1520};
  wire [1023:0] dataGroup_hi_1520 = {dataGroup_hi_hi_1520, dataGroup_hi_lo_1520};
  wire [15:0]   dataGroup_0_59 = dataGroup_lo_1520[47:32];
  wire [1023:0] dataGroup_lo_1521 = {dataGroup_lo_hi_1521, dataGroup_lo_lo_1521};
  wire [1023:0] dataGroup_hi_1521 = {dataGroup_hi_hi_1521, dataGroup_hi_lo_1521};
  wire [15:0]   dataGroup_1_59 = dataGroup_lo_1521[159:144];
  wire [1023:0] dataGroup_lo_1522 = {dataGroup_lo_hi_1522, dataGroup_lo_lo_1522};
  wire [1023:0] dataGroup_hi_1522 = {dataGroup_hi_hi_1522, dataGroup_hi_lo_1522};
  wire [15:0]   dataGroup_2_59 = dataGroup_lo_1522[271:256];
  wire [1023:0] dataGroup_lo_1523 = {dataGroup_lo_hi_1523, dataGroup_lo_lo_1523};
  wire [1023:0] dataGroup_hi_1523 = {dataGroup_hi_hi_1523, dataGroup_hi_lo_1523};
  wire [15:0]   dataGroup_3_59 = dataGroup_lo_1523[383:368];
  wire [1023:0] dataGroup_lo_1524 = {dataGroup_lo_hi_1524, dataGroup_lo_lo_1524};
  wire [1023:0] dataGroup_hi_1524 = {dataGroup_hi_hi_1524, dataGroup_hi_lo_1524};
  wire [15:0]   dataGroup_4_59 = dataGroup_lo_1524[495:480];
  wire [1023:0] dataGroup_lo_1525 = {dataGroup_lo_hi_1525, dataGroup_lo_lo_1525};
  wire [1023:0] dataGroup_hi_1525 = {dataGroup_hi_hi_1525, dataGroup_hi_lo_1525};
  wire [15:0]   dataGroup_5_59 = dataGroup_lo_1525[607:592];
  wire [1023:0] dataGroup_lo_1526 = {dataGroup_lo_hi_1526, dataGroup_lo_lo_1526};
  wire [1023:0] dataGroup_hi_1526 = {dataGroup_hi_hi_1526, dataGroup_hi_lo_1526};
  wire [15:0]   dataGroup_6_59 = dataGroup_lo_1526[719:704];
  wire [1023:0] dataGroup_lo_1527 = {dataGroup_lo_hi_1527, dataGroup_lo_lo_1527};
  wire [1023:0] dataGroup_hi_1527 = {dataGroup_hi_hi_1527, dataGroup_hi_lo_1527};
  wire [15:0]   dataGroup_7_59 = dataGroup_lo_1527[831:816];
  wire [1023:0] dataGroup_lo_1528 = {dataGroup_lo_hi_1528, dataGroup_lo_lo_1528};
  wire [1023:0] dataGroup_hi_1528 = {dataGroup_hi_hi_1528, dataGroup_hi_lo_1528};
  wire [15:0]   dataGroup_8_59 = dataGroup_lo_1528[943:928];
  wire [1023:0] dataGroup_lo_1529 = {dataGroup_lo_hi_1529, dataGroup_lo_lo_1529};
  wire [1023:0] dataGroup_hi_1529 = {dataGroup_hi_hi_1529, dataGroup_hi_lo_1529};
  wire [15:0]   dataGroup_9_59 = dataGroup_hi_1529[31:16];
  wire [1023:0] dataGroup_lo_1530 = {dataGroup_lo_hi_1530, dataGroup_lo_lo_1530};
  wire [1023:0] dataGroup_hi_1530 = {dataGroup_hi_hi_1530, dataGroup_hi_lo_1530};
  wire [15:0]   dataGroup_10_59 = dataGroup_hi_1530[143:128];
  wire [1023:0] dataGroup_lo_1531 = {dataGroup_lo_hi_1531, dataGroup_lo_lo_1531};
  wire [1023:0] dataGroup_hi_1531 = {dataGroup_hi_hi_1531, dataGroup_hi_lo_1531};
  wire [15:0]   dataGroup_11_59 = dataGroup_hi_1531[255:240];
  wire [1023:0] dataGroup_lo_1532 = {dataGroup_lo_hi_1532, dataGroup_lo_lo_1532};
  wire [1023:0] dataGroup_hi_1532 = {dataGroup_hi_hi_1532, dataGroup_hi_lo_1532};
  wire [15:0]   dataGroup_12_59 = dataGroup_hi_1532[367:352];
  wire [1023:0] dataGroup_lo_1533 = {dataGroup_lo_hi_1533, dataGroup_lo_lo_1533};
  wire [1023:0] dataGroup_hi_1533 = {dataGroup_hi_hi_1533, dataGroup_hi_lo_1533};
  wire [15:0]   dataGroup_13_59 = dataGroup_hi_1533[479:464];
  wire [1023:0] dataGroup_lo_1534 = {dataGroup_lo_hi_1534, dataGroup_lo_lo_1534};
  wire [1023:0] dataGroup_hi_1534 = {dataGroup_hi_hi_1534, dataGroup_hi_lo_1534};
  wire [15:0]   dataGroup_14_59 = dataGroup_hi_1534[591:576];
  wire [1023:0] dataGroup_lo_1535 = {dataGroup_lo_hi_1535, dataGroup_lo_lo_1535};
  wire [1023:0] dataGroup_hi_1535 = {dataGroup_hi_hi_1535, dataGroup_hi_lo_1535};
  wire [15:0]   dataGroup_15_59 = dataGroup_hi_1535[703:688];
  wire [31:0]   res_lo_lo_lo_59 = {dataGroup_1_59, dataGroup_0_59};
  wire [31:0]   res_lo_lo_hi_59 = {dataGroup_3_59, dataGroup_2_59};
  wire [63:0]   res_lo_lo_59 = {res_lo_lo_hi_59, res_lo_lo_lo_59};
  wire [31:0]   res_lo_hi_lo_59 = {dataGroup_5_59, dataGroup_4_59};
  wire [31:0]   res_lo_hi_hi_59 = {dataGroup_7_59, dataGroup_6_59};
  wire [63:0]   res_lo_hi_59 = {res_lo_hi_hi_59, res_lo_hi_lo_59};
  wire [127:0]  res_lo_59 = {res_lo_hi_59, res_lo_lo_59};
  wire [31:0]   res_hi_lo_lo_59 = {dataGroup_9_59, dataGroup_8_59};
  wire [31:0]   res_hi_lo_hi_59 = {dataGroup_11_59, dataGroup_10_59};
  wire [63:0]   res_hi_lo_59 = {res_hi_lo_hi_59, res_hi_lo_lo_59};
  wire [31:0]   res_hi_hi_lo_59 = {dataGroup_13_59, dataGroup_12_59};
  wire [31:0]   res_hi_hi_hi_59 = {dataGroup_15_59, dataGroup_14_59};
  wire [63:0]   res_hi_hi_59 = {res_hi_hi_hi_59, res_hi_hi_lo_59};
  wire [127:0]  res_hi_59 = {res_hi_hi_59, res_hi_lo_59};
  wire [255:0]  res_114 = {res_hi_59, res_lo_59};
  wire [1023:0] dataGroup_lo_1536 = {dataGroup_lo_hi_1536, dataGroup_lo_lo_1536};
  wire [1023:0] dataGroup_hi_1536 = {dataGroup_hi_hi_1536, dataGroup_hi_lo_1536};
  wire [15:0]   dataGroup_0_60 = dataGroup_lo_1536[63:48];
  wire [1023:0] dataGroup_lo_1537 = {dataGroup_lo_hi_1537, dataGroup_lo_lo_1537};
  wire [1023:0] dataGroup_hi_1537 = {dataGroup_hi_hi_1537, dataGroup_hi_lo_1537};
  wire [15:0]   dataGroup_1_60 = dataGroup_lo_1537[175:160];
  wire [1023:0] dataGroup_lo_1538 = {dataGroup_lo_hi_1538, dataGroup_lo_lo_1538};
  wire [1023:0] dataGroup_hi_1538 = {dataGroup_hi_hi_1538, dataGroup_hi_lo_1538};
  wire [15:0]   dataGroup_2_60 = dataGroup_lo_1538[287:272];
  wire [1023:0] dataGroup_lo_1539 = {dataGroup_lo_hi_1539, dataGroup_lo_lo_1539};
  wire [1023:0] dataGroup_hi_1539 = {dataGroup_hi_hi_1539, dataGroup_hi_lo_1539};
  wire [15:0]   dataGroup_3_60 = dataGroup_lo_1539[399:384];
  wire [1023:0] dataGroup_lo_1540 = {dataGroup_lo_hi_1540, dataGroup_lo_lo_1540};
  wire [1023:0] dataGroup_hi_1540 = {dataGroup_hi_hi_1540, dataGroup_hi_lo_1540};
  wire [15:0]   dataGroup_4_60 = dataGroup_lo_1540[511:496];
  wire [1023:0] dataGroup_lo_1541 = {dataGroup_lo_hi_1541, dataGroup_lo_lo_1541};
  wire [1023:0] dataGroup_hi_1541 = {dataGroup_hi_hi_1541, dataGroup_hi_lo_1541};
  wire [15:0]   dataGroup_5_60 = dataGroup_lo_1541[623:608];
  wire [1023:0] dataGroup_lo_1542 = {dataGroup_lo_hi_1542, dataGroup_lo_lo_1542};
  wire [1023:0] dataGroup_hi_1542 = {dataGroup_hi_hi_1542, dataGroup_hi_lo_1542};
  wire [15:0]   dataGroup_6_60 = dataGroup_lo_1542[735:720];
  wire [1023:0] dataGroup_lo_1543 = {dataGroup_lo_hi_1543, dataGroup_lo_lo_1543};
  wire [1023:0] dataGroup_hi_1543 = {dataGroup_hi_hi_1543, dataGroup_hi_lo_1543};
  wire [15:0]   dataGroup_7_60 = dataGroup_lo_1543[847:832];
  wire [1023:0] dataGroup_lo_1544 = {dataGroup_lo_hi_1544, dataGroup_lo_lo_1544};
  wire [1023:0] dataGroup_hi_1544 = {dataGroup_hi_hi_1544, dataGroup_hi_lo_1544};
  wire [15:0]   dataGroup_8_60 = dataGroup_lo_1544[959:944];
  wire [1023:0] dataGroup_lo_1545 = {dataGroup_lo_hi_1545, dataGroup_lo_lo_1545};
  wire [1023:0] dataGroup_hi_1545 = {dataGroup_hi_hi_1545, dataGroup_hi_lo_1545};
  wire [15:0]   dataGroup_9_60 = dataGroup_hi_1545[47:32];
  wire [1023:0] dataGroup_lo_1546 = {dataGroup_lo_hi_1546, dataGroup_lo_lo_1546};
  wire [1023:0] dataGroup_hi_1546 = {dataGroup_hi_hi_1546, dataGroup_hi_lo_1546};
  wire [15:0]   dataGroup_10_60 = dataGroup_hi_1546[159:144];
  wire [1023:0] dataGroup_lo_1547 = {dataGroup_lo_hi_1547, dataGroup_lo_lo_1547};
  wire [1023:0] dataGroup_hi_1547 = {dataGroup_hi_hi_1547, dataGroup_hi_lo_1547};
  wire [15:0]   dataGroup_11_60 = dataGroup_hi_1547[271:256];
  wire [1023:0] dataGroup_lo_1548 = {dataGroup_lo_hi_1548, dataGroup_lo_lo_1548};
  wire [1023:0] dataGroup_hi_1548 = {dataGroup_hi_hi_1548, dataGroup_hi_lo_1548};
  wire [15:0]   dataGroup_12_60 = dataGroup_hi_1548[383:368];
  wire [1023:0] dataGroup_lo_1549 = {dataGroup_lo_hi_1549, dataGroup_lo_lo_1549};
  wire [1023:0] dataGroup_hi_1549 = {dataGroup_hi_hi_1549, dataGroup_hi_lo_1549};
  wire [15:0]   dataGroup_13_60 = dataGroup_hi_1549[495:480];
  wire [1023:0] dataGroup_lo_1550 = {dataGroup_lo_hi_1550, dataGroup_lo_lo_1550};
  wire [1023:0] dataGroup_hi_1550 = {dataGroup_hi_hi_1550, dataGroup_hi_lo_1550};
  wire [15:0]   dataGroup_14_60 = dataGroup_hi_1550[607:592];
  wire [1023:0] dataGroup_lo_1551 = {dataGroup_lo_hi_1551, dataGroup_lo_lo_1551};
  wire [1023:0] dataGroup_hi_1551 = {dataGroup_hi_hi_1551, dataGroup_hi_lo_1551};
  wire [15:0]   dataGroup_15_60 = dataGroup_hi_1551[719:704];
  wire [31:0]   res_lo_lo_lo_60 = {dataGroup_1_60, dataGroup_0_60};
  wire [31:0]   res_lo_lo_hi_60 = {dataGroup_3_60, dataGroup_2_60};
  wire [63:0]   res_lo_lo_60 = {res_lo_lo_hi_60, res_lo_lo_lo_60};
  wire [31:0]   res_lo_hi_lo_60 = {dataGroup_5_60, dataGroup_4_60};
  wire [31:0]   res_lo_hi_hi_60 = {dataGroup_7_60, dataGroup_6_60};
  wire [63:0]   res_lo_hi_60 = {res_lo_hi_hi_60, res_lo_hi_lo_60};
  wire [127:0]  res_lo_60 = {res_lo_hi_60, res_lo_lo_60};
  wire [31:0]   res_hi_lo_lo_60 = {dataGroup_9_60, dataGroup_8_60};
  wire [31:0]   res_hi_lo_hi_60 = {dataGroup_11_60, dataGroup_10_60};
  wire [63:0]   res_hi_lo_60 = {res_hi_lo_hi_60, res_hi_lo_lo_60};
  wire [31:0]   res_hi_hi_lo_60 = {dataGroup_13_60, dataGroup_12_60};
  wire [31:0]   res_hi_hi_hi_60 = {dataGroup_15_60, dataGroup_14_60};
  wire [63:0]   res_hi_hi_60 = {res_hi_hi_hi_60, res_hi_hi_lo_60};
  wire [127:0]  res_hi_60 = {res_hi_hi_60, res_hi_lo_60};
  wire [255:0]  res_115 = {res_hi_60, res_lo_60};
  wire [1023:0] dataGroup_lo_1552 = {dataGroup_lo_hi_1552, dataGroup_lo_lo_1552};
  wire [1023:0] dataGroup_hi_1552 = {dataGroup_hi_hi_1552, dataGroup_hi_lo_1552};
  wire [15:0]   dataGroup_0_61 = dataGroup_lo_1552[79:64];
  wire [1023:0] dataGroup_lo_1553 = {dataGroup_lo_hi_1553, dataGroup_lo_lo_1553};
  wire [1023:0] dataGroup_hi_1553 = {dataGroup_hi_hi_1553, dataGroup_hi_lo_1553};
  wire [15:0]   dataGroup_1_61 = dataGroup_lo_1553[191:176];
  wire [1023:0] dataGroup_lo_1554 = {dataGroup_lo_hi_1554, dataGroup_lo_lo_1554};
  wire [1023:0] dataGroup_hi_1554 = {dataGroup_hi_hi_1554, dataGroup_hi_lo_1554};
  wire [15:0]   dataGroup_2_61 = dataGroup_lo_1554[303:288];
  wire [1023:0] dataGroup_lo_1555 = {dataGroup_lo_hi_1555, dataGroup_lo_lo_1555};
  wire [1023:0] dataGroup_hi_1555 = {dataGroup_hi_hi_1555, dataGroup_hi_lo_1555};
  wire [15:0]   dataGroup_3_61 = dataGroup_lo_1555[415:400];
  wire [1023:0] dataGroup_lo_1556 = {dataGroup_lo_hi_1556, dataGroup_lo_lo_1556};
  wire [1023:0] dataGroup_hi_1556 = {dataGroup_hi_hi_1556, dataGroup_hi_lo_1556};
  wire [15:0]   dataGroup_4_61 = dataGroup_lo_1556[527:512];
  wire [1023:0] dataGroup_lo_1557 = {dataGroup_lo_hi_1557, dataGroup_lo_lo_1557};
  wire [1023:0] dataGroup_hi_1557 = {dataGroup_hi_hi_1557, dataGroup_hi_lo_1557};
  wire [15:0]   dataGroup_5_61 = dataGroup_lo_1557[639:624];
  wire [1023:0] dataGroup_lo_1558 = {dataGroup_lo_hi_1558, dataGroup_lo_lo_1558};
  wire [1023:0] dataGroup_hi_1558 = {dataGroup_hi_hi_1558, dataGroup_hi_lo_1558};
  wire [15:0]   dataGroup_6_61 = dataGroup_lo_1558[751:736];
  wire [1023:0] dataGroup_lo_1559 = {dataGroup_lo_hi_1559, dataGroup_lo_lo_1559};
  wire [1023:0] dataGroup_hi_1559 = {dataGroup_hi_hi_1559, dataGroup_hi_lo_1559};
  wire [15:0]   dataGroup_7_61 = dataGroup_lo_1559[863:848];
  wire [1023:0] dataGroup_lo_1560 = {dataGroup_lo_hi_1560, dataGroup_lo_lo_1560};
  wire [1023:0] dataGroup_hi_1560 = {dataGroup_hi_hi_1560, dataGroup_hi_lo_1560};
  wire [15:0]   dataGroup_8_61 = dataGroup_lo_1560[975:960];
  wire [1023:0] dataGroup_lo_1561 = {dataGroup_lo_hi_1561, dataGroup_lo_lo_1561};
  wire [1023:0] dataGroup_hi_1561 = {dataGroup_hi_hi_1561, dataGroup_hi_lo_1561};
  wire [15:0]   dataGroup_9_61 = dataGroup_hi_1561[63:48];
  wire [1023:0] dataGroup_lo_1562 = {dataGroup_lo_hi_1562, dataGroup_lo_lo_1562};
  wire [1023:0] dataGroup_hi_1562 = {dataGroup_hi_hi_1562, dataGroup_hi_lo_1562};
  wire [15:0]   dataGroup_10_61 = dataGroup_hi_1562[175:160];
  wire [1023:0] dataGroup_lo_1563 = {dataGroup_lo_hi_1563, dataGroup_lo_lo_1563};
  wire [1023:0] dataGroup_hi_1563 = {dataGroup_hi_hi_1563, dataGroup_hi_lo_1563};
  wire [15:0]   dataGroup_11_61 = dataGroup_hi_1563[287:272];
  wire [1023:0] dataGroup_lo_1564 = {dataGroup_lo_hi_1564, dataGroup_lo_lo_1564};
  wire [1023:0] dataGroup_hi_1564 = {dataGroup_hi_hi_1564, dataGroup_hi_lo_1564};
  wire [15:0]   dataGroup_12_61 = dataGroup_hi_1564[399:384];
  wire [1023:0] dataGroup_lo_1565 = {dataGroup_lo_hi_1565, dataGroup_lo_lo_1565};
  wire [1023:0] dataGroup_hi_1565 = {dataGroup_hi_hi_1565, dataGroup_hi_lo_1565};
  wire [15:0]   dataGroup_13_61 = dataGroup_hi_1565[511:496];
  wire [1023:0] dataGroup_lo_1566 = {dataGroup_lo_hi_1566, dataGroup_lo_lo_1566};
  wire [1023:0] dataGroup_hi_1566 = {dataGroup_hi_hi_1566, dataGroup_hi_lo_1566};
  wire [15:0]   dataGroup_14_61 = dataGroup_hi_1566[623:608];
  wire [1023:0] dataGroup_lo_1567 = {dataGroup_lo_hi_1567, dataGroup_lo_lo_1567};
  wire [1023:0] dataGroup_hi_1567 = {dataGroup_hi_hi_1567, dataGroup_hi_lo_1567};
  wire [15:0]   dataGroup_15_61 = dataGroup_hi_1567[735:720];
  wire [31:0]   res_lo_lo_lo_61 = {dataGroup_1_61, dataGroup_0_61};
  wire [31:0]   res_lo_lo_hi_61 = {dataGroup_3_61, dataGroup_2_61};
  wire [63:0]   res_lo_lo_61 = {res_lo_lo_hi_61, res_lo_lo_lo_61};
  wire [31:0]   res_lo_hi_lo_61 = {dataGroup_5_61, dataGroup_4_61};
  wire [31:0]   res_lo_hi_hi_61 = {dataGroup_7_61, dataGroup_6_61};
  wire [63:0]   res_lo_hi_61 = {res_lo_hi_hi_61, res_lo_hi_lo_61};
  wire [127:0]  res_lo_61 = {res_lo_hi_61, res_lo_lo_61};
  wire [31:0]   res_hi_lo_lo_61 = {dataGroup_9_61, dataGroup_8_61};
  wire [31:0]   res_hi_lo_hi_61 = {dataGroup_11_61, dataGroup_10_61};
  wire [63:0]   res_hi_lo_61 = {res_hi_lo_hi_61, res_hi_lo_lo_61};
  wire [31:0]   res_hi_hi_lo_61 = {dataGroup_13_61, dataGroup_12_61};
  wire [31:0]   res_hi_hi_hi_61 = {dataGroup_15_61, dataGroup_14_61};
  wire [63:0]   res_hi_hi_61 = {res_hi_hi_hi_61, res_hi_hi_lo_61};
  wire [127:0]  res_hi_61 = {res_hi_hi_61, res_hi_lo_61};
  wire [255:0]  res_116 = {res_hi_61, res_lo_61};
  wire [1023:0] dataGroup_lo_1568 = {dataGroup_lo_hi_1568, dataGroup_lo_lo_1568};
  wire [1023:0] dataGroup_hi_1568 = {dataGroup_hi_hi_1568, dataGroup_hi_lo_1568};
  wire [15:0]   dataGroup_0_62 = dataGroup_lo_1568[95:80];
  wire [1023:0] dataGroup_lo_1569 = {dataGroup_lo_hi_1569, dataGroup_lo_lo_1569};
  wire [1023:0] dataGroup_hi_1569 = {dataGroup_hi_hi_1569, dataGroup_hi_lo_1569};
  wire [15:0]   dataGroup_1_62 = dataGroup_lo_1569[207:192];
  wire [1023:0] dataGroup_lo_1570 = {dataGroup_lo_hi_1570, dataGroup_lo_lo_1570};
  wire [1023:0] dataGroup_hi_1570 = {dataGroup_hi_hi_1570, dataGroup_hi_lo_1570};
  wire [15:0]   dataGroup_2_62 = dataGroup_lo_1570[319:304];
  wire [1023:0] dataGroup_lo_1571 = {dataGroup_lo_hi_1571, dataGroup_lo_lo_1571};
  wire [1023:0] dataGroup_hi_1571 = {dataGroup_hi_hi_1571, dataGroup_hi_lo_1571};
  wire [15:0]   dataGroup_3_62 = dataGroup_lo_1571[431:416];
  wire [1023:0] dataGroup_lo_1572 = {dataGroup_lo_hi_1572, dataGroup_lo_lo_1572};
  wire [1023:0] dataGroup_hi_1572 = {dataGroup_hi_hi_1572, dataGroup_hi_lo_1572};
  wire [15:0]   dataGroup_4_62 = dataGroup_lo_1572[543:528];
  wire [1023:0] dataGroup_lo_1573 = {dataGroup_lo_hi_1573, dataGroup_lo_lo_1573};
  wire [1023:0] dataGroup_hi_1573 = {dataGroup_hi_hi_1573, dataGroup_hi_lo_1573};
  wire [15:0]   dataGroup_5_62 = dataGroup_lo_1573[655:640];
  wire [1023:0] dataGroup_lo_1574 = {dataGroup_lo_hi_1574, dataGroup_lo_lo_1574};
  wire [1023:0] dataGroup_hi_1574 = {dataGroup_hi_hi_1574, dataGroup_hi_lo_1574};
  wire [15:0]   dataGroup_6_62 = dataGroup_lo_1574[767:752];
  wire [1023:0] dataGroup_lo_1575 = {dataGroup_lo_hi_1575, dataGroup_lo_lo_1575};
  wire [1023:0] dataGroup_hi_1575 = {dataGroup_hi_hi_1575, dataGroup_hi_lo_1575};
  wire [15:0]   dataGroup_7_62 = dataGroup_lo_1575[879:864];
  wire [1023:0] dataGroup_lo_1576 = {dataGroup_lo_hi_1576, dataGroup_lo_lo_1576};
  wire [1023:0] dataGroup_hi_1576 = {dataGroup_hi_hi_1576, dataGroup_hi_lo_1576};
  wire [15:0]   dataGroup_8_62 = dataGroup_lo_1576[991:976];
  wire [1023:0] dataGroup_lo_1577 = {dataGroup_lo_hi_1577, dataGroup_lo_lo_1577};
  wire [1023:0] dataGroup_hi_1577 = {dataGroup_hi_hi_1577, dataGroup_hi_lo_1577};
  wire [15:0]   dataGroup_9_62 = dataGroup_hi_1577[79:64];
  wire [1023:0] dataGroup_lo_1578 = {dataGroup_lo_hi_1578, dataGroup_lo_lo_1578};
  wire [1023:0] dataGroup_hi_1578 = {dataGroup_hi_hi_1578, dataGroup_hi_lo_1578};
  wire [15:0]   dataGroup_10_62 = dataGroup_hi_1578[191:176];
  wire [1023:0] dataGroup_lo_1579 = {dataGroup_lo_hi_1579, dataGroup_lo_lo_1579};
  wire [1023:0] dataGroup_hi_1579 = {dataGroup_hi_hi_1579, dataGroup_hi_lo_1579};
  wire [15:0]   dataGroup_11_62 = dataGroup_hi_1579[303:288];
  wire [1023:0] dataGroup_lo_1580 = {dataGroup_lo_hi_1580, dataGroup_lo_lo_1580};
  wire [1023:0] dataGroup_hi_1580 = {dataGroup_hi_hi_1580, dataGroup_hi_lo_1580};
  wire [15:0]   dataGroup_12_62 = dataGroup_hi_1580[415:400];
  wire [1023:0] dataGroup_lo_1581 = {dataGroup_lo_hi_1581, dataGroup_lo_lo_1581};
  wire [1023:0] dataGroup_hi_1581 = {dataGroup_hi_hi_1581, dataGroup_hi_lo_1581};
  wire [15:0]   dataGroup_13_62 = dataGroup_hi_1581[527:512];
  wire [1023:0] dataGroup_lo_1582 = {dataGroup_lo_hi_1582, dataGroup_lo_lo_1582};
  wire [1023:0] dataGroup_hi_1582 = {dataGroup_hi_hi_1582, dataGroup_hi_lo_1582};
  wire [15:0]   dataGroup_14_62 = dataGroup_hi_1582[639:624];
  wire [1023:0] dataGroup_lo_1583 = {dataGroup_lo_hi_1583, dataGroup_lo_lo_1583};
  wire [1023:0] dataGroup_hi_1583 = {dataGroup_hi_hi_1583, dataGroup_hi_lo_1583};
  wire [15:0]   dataGroup_15_62 = dataGroup_hi_1583[751:736];
  wire [31:0]   res_lo_lo_lo_62 = {dataGroup_1_62, dataGroup_0_62};
  wire [31:0]   res_lo_lo_hi_62 = {dataGroup_3_62, dataGroup_2_62};
  wire [63:0]   res_lo_lo_62 = {res_lo_lo_hi_62, res_lo_lo_lo_62};
  wire [31:0]   res_lo_hi_lo_62 = {dataGroup_5_62, dataGroup_4_62};
  wire [31:0]   res_lo_hi_hi_62 = {dataGroup_7_62, dataGroup_6_62};
  wire [63:0]   res_lo_hi_62 = {res_lo_hi_hi_62, res_lo_hi_lo_62};
  wire [127:0]  res_lo_62 = {res_lo_hi_62, res_lo_lo_62};
  wire [31:0]   res_hi_lo_lo_62 = {dataGroup_9_62, dataGroup_8_62};
  wire [31:0]   res_hi_lo_hi_62 = {dataGroup_11_62, dataGroup_10_62};
  wire [63:0]   res_hi_lo_62 = {res_hi_lo_hi_62, res_hi_lo_lo_62};
  wire [31:0]   res_hi_hi_lo_62 = {dataGroup_13_62, dataGroup_12_62};
  wire [31:0]   res_hi_hi_hi_62 = {dataGroup_15_62, dataGroup_14_62};
  wire [63:0]   res_hi_hi_62 = {res_hi_hi_hi_62, res_hi_hi_lo_62};
  wire [127:0]  res_hi_62 = {res_hi_hi_62, res_hi_lo_62};
  wire [255:0]  res_117 = {res_hi_62, res_lo_62};
  wire [1023:0] dataGroup_lo_1584 = {dataGroup_lo_hi_1584, dataGroup_lo_lo_1584};
  wire [1023:0] dataGroup_hi_1584 = {dataGroup_hi_hi_1584, dataGroup_hi_lo_1584};
  wire [15:0]   dataGroup_0_63 = dataGroup_lo_1584[111:96];
  wire [1023:0] dataGroup_lo_1585 = {dataGroup_lo_hi_1585, dataGroup_lo_lo_1585};
  wire [1023:0] dataGroup_hi_1585 = {dataGroup_hi_hi_1585, dataGroup_hi_lo_1585};
  wire [15:0]   dataGroup_1_63 = dataGroup_lo_1585[223:208];
  wire [1023:0] dataGroup_lo_1586 = {dataGroup_lo_hi_1586, dataGroup_lo_lo_1586};
  wire [1023:0] dataGroup_hi_1586 = {dataGroup_hi_hi_1586, dataGroup_hi_lo_1586};
  wire [15:0]   dataGroup_2_63 = dataGroup_lo_1586[335:320];
  wire [1023:0] dataGroup_lo_1587 = {dataGroup_lo_hi_1587, dataGroup_lo_lo_1587};
  wire [1023:0] dataGroup_hi_1587 = {dataGroup_hi_hi_1587, dataGroup_hi_lo_1587};
  wire [15:0]   dataGroup_3_63 = dataGroup_lo_1587[447:432];
  wire [1023:0] dataGroup_lo_1588 = {dataGroup_lo_hi_1588, dataGroup_lo_lo_1588};
  wire [1023:0] dataGroup_hi_1588 = {dataGroup_hi_hi_1588, dataGroup_hi_lo_1588};
  wire [15:0]   dataGroup_4_63 = dataGroup_lo_1588[559:544];
  wire [1023:0] dataGroup_lo_1589 = {dataGroup_lo_hi_1589, dataGroup_lo_lo_1589};
  wire [1023:0] dataGroup_hi_1589 = {dataGroup_hi_hi_1589, dataGroup_hi_lo_1589};
  wire [15:0]   dataGroup_5_63 = dataGroup_lo_1589[671:656];
  wire [1023:0] dataGroup_lo_1590 = {dataGroup_lo_hi_1590, dataGroup_lo_lo_1590};
  wire [1023:0] dataGroup_hi_1590 = {dataGroup_hi_hi_1590, dataGroup_hi_lo_1590};
  wire [15:0]   dataGroup_6_63 = dataGroup_lo_1590[783:768];
  wire [1023:0] dataGroup_lo_1591 = {dataGroup_lo_hi_1591, dataGroup_lo_lo_1591};
  wire [1023:0] dataGroup_hi_1591 = {dataGroup_hi_hi_1591, dataGroup_hi_lo_1591};
  wire [15:0]   dataGroup_7_63 = dataGroup_lo_1591[895:880];
  wire [1023:0] dataGroup_lo_1592 = {dataGroup_lo_hi_1592, dataGroup_lo_lo_1592};
  wire [1023:0] dataGroup_hi_1592 = {dataGroup_hi_hi_1592, dataGroup_hi_lo_1592};
  wire [15:0]   dataGroup_8_63 = dataGroup_lo_1592[1007:992];
  wire [1023:0] dataGroup_lo_1593 = {dataGroup_lo_hi_1593, dataGroup_lo_lo_1593};
  wire [1023:0] dataGroup_hi_1593 = {dataGroup_hi_hi_1593, dataGroup_hi_lo_1593};
  wire [15:0]   dataGroup_9_63 = dataGroup_hi_1593[95:80];
  wire [1023:0] dataGroup_lo_1594 = {dataGroup_lo_hi_1594, dataGroup_lo_lo_1594};
  wire [1023:0] dataGroup_hi_1594 = {dataGroup_hi_hi_1594, dataGroup_hi_lo_1594};
  wire [15:0]   dataGroup_10_63 = dataGroup_hi_1594[207:192];
  wire [1023:0] dataGroup_lo_1595 = {dataGroup_lo_hi_1595, dataGroup_lo_lo_1595};
  wire [1023:0] dataGroup_hi_1595 = {dataGroup_hi_hi_1595, dataGroup_hi_lo_1595};
  wire [15:0]   dataGroup_11_63 = dataGroup_hi_1595[319:304];
  wire [1023:0] dataGroup_lo_1596 = {dataGroup_lo_hi_1596, dataGroup_lo_lo_1596};
  wire [1023:0] dataGroup_hi_1596 = {dataGroup_hi_hi_1596, dataGroup_hi_lo_1596};
  wire [15:0]   dataGroup_12_63 = dataGroup_hi_1596[431:416];
  wire [1023:0] dataGroup_lo_1597 = {dataGroup_lo_hi_1597, dataGroup_lo_lo_1597};
  wire [1023:0] dataGroup_hi_1597 = {dataGroup_hi_hi_1597, dataGroup_hi_lo_1597};
  wire [15:0]   dataGroup_13_63 = dataGroup_hi_1597[543:528];
  wire [1023:0] dataGroup_lo_1598 = {dataGroup_lo_hi_1598, dataGroup_lo_lo_1598};
  wire [1023:0] dataGroup_hi_1598 = {dataGroup_hi_hi_1598, dataGroup_hi_lo_1598};
  wire [15:0]   dataGroup_14_63 = dataGroup_hi_1598[655:640];
  wire [1023:0] dataGroup_lo_1599 = {dataGroup_lo_hi_1599, dataGroup_lo_lo_1599};
  wire [1023:0] dataGroup_hi_1599 = {dataGroup_hi_hi_1599, dataGroup_hi_lo_1599};
  wire [15:0]   dataGroup_15_63 = dataGroup_hi_1599[767:752];
  wire [31:0]   res_lo_lo_lo_63 = {dataGroup_1_63, dataGroup_0_63};
  wire [31:0]   res_lo_lo_hi_63 = {dataGroup_3_63, dataGroup_2_63};
  wire [63:0]   res_lo_lo_63 = {res_lo_lo_hi_63, res_lo_lo_lo_63};
  wire [31:0]   res_lo_hi_lo_63 = {dataGroup_5_63, dataGroup_4_63};
  wire [31:0]   res_lo_hi_hi_63 = {dataGroup_7_63, dataGroup_6_63};
  wire [63:0]   res_lo_hi_63 = {res_lo_hi_hi_63, res_lo_hi_lo_63};
  wire [127:0]  res_lo_63 = {res_lo_hi_63, res_lo_lo_63};
  wire [31:0]   res_hi_lo_lo_63 = {dataGroup_9_63, dataGroup_8_63};
  wire [31:0]   res_hi_lo_hi_63 = {dataGroup_11_63, dataGroup_10_63};
  wire [63:0]   res_hi_lo_63 = {res_hi_lo_hi_63, res_hi_lo_lo_63};
  wire [31:0]   res_hi_hi_lo_63 = {dataGroup_13_63, dataGroup_12_63};
  wire [31:0]   res_hi_hi_hi_63 = {dataGroup_15_63, dataGroup_14_63};
  wire [63:0]   res_hi_hi_63 = {res_hi_hi_hi_63, res_hi_hi_lo_63};
  wire [127:0]  res_hi_63 = {res_hi_hi_63, res_hi_lo_63};
  wire [255:0]  res_118 = {res_hi_63, res_lo_63};
  wire [511:0]  lo_lo_14 = {res_113, res_112};
  wire [511:0]  lo_hi_14 = {res_115, res_114};
  wire [1023:0] lo_14 = {lo_hi_14, lo_lo_14};
  wire [511:0]  hi_lo_14 = {res_117, res_116};
  wire [511:0]  hi_hi_14 = {256'h0, res_118};
  wire [1023:0] hi_14 = {hi_hi_14, hi_lo_14};
  wire [2047:0] regroupLoadData_1_6 = {hi_14, lo_14};
  wire [1023:0] dataGroup_lo_1600 = {dataGroup_lo_hi_1600, dataGroup_lo_lo_1600};
  wire [1023:0] dataGroup_hi_1600 = {dataGroup_hi_hi_1600, dataGroup_hi_lo_1600};
  wire [15:0]   dataGroup_0_64 = dataGroup_lo_1600[15:0];
  wire [1023:0] dataGroup_lo_1601 = {dataGroup_lo_hi_1601, dataGroup_lo_lo_1601};
  wire [1023:0] dataGroup_hi_1601 = {dataGroup_hi_hi_1601, dataGroup_hi_lo_1601};
  wire [15:0]   dataGroup_1_64 = dataGroup_lo_1601[143:128];
  wire [1023:0] dataGroup_lo_1602 = {dataGroup_lo_hi_1602, dataGroup_lo_lo_1602};
  wire [1023:0] dataGroup_hi_1602 = {dataGroup_hi_hi_1602, dataGroup_hi_lo_1602};
  wire [15:0]   dataGroup_2_64 = dataGroup_lo_1602[271:256];
  wire [1023:0] dataGroup_lo_1603 = {dataGroup_lo_hi_1603, dataGroup_lo_lo_1603};
  wire [1023:0] dataGroup_hi_1603 = {dataGroup_hi_hi_1603, dataGroup_hi_lo_1603};
  wire [15:0]   dataGroup_3_64 = dataGroup_lo_1603[399:384];
  wire [1023:0] dataGroup_lo_1604 = {dataGroup_lo_hi_1604, dataGroup_lo_lo_1604};
  wire [1023:0] dataGroup_hi_1604 = {dataGroup_hi_hi_1604, dataGroup_hi_lo_1604};
  wire [15:0]   dataGroup_4_64 = dataGroup_lo_1604[527:512];
  wire [1023:0] dataGroup_lo_1605 = {dataGroup_lo_hi_1605, dataGroup_lo_lo_1605};
  wire [1023:0] dataGroup_hi_1605 = {dataGroup_hi_hi_1605, dataGroup_hi_lo_1605};
  wire [15:0]   dataGroup_5_64 = dataGroup_lo_1605[655:640];
  wire [1023:0] dataGroup_lo_1606 = {dataGroup_lo_hi_1606, dataGroup_lo_lo_1606};
  wire [1023:0] dataGroup_hi_1606 = {dataGroup_hi_hi_1606, dataGroup_hi_lo_1606};
  wire [15:0]   dataGroup_6_64 = dataGroup_lo_1606[783:768];
  wire [1023:0] dataGroup_lo_1607 = {dataGroup_lo_hi_1607, dataGroup_lo_lo_1607};
  wire [1023:0] dataGroup_hi_1607 = {dataGroup_hi_hi_1607, dataGroup_hi_lo_1607};
  wire [15:0]   dataGroup_7_64 = dataGroup_lo_1607[911:896];
  wire [1023:0] dataGroup_lo_1608 = {dataGroup_lo_hi_1608, dataGroup_lo_lo_1608};
  wire [1023:0] dataGroup_hi_1608 = {dataGroup_hi_hi_1608, dataGroup_hi_lo_1608};
  wire [15:0]   dataGroup_8_64 = dataGroup_hi_1608[15:0];
  wire [1023:0] dataGroup_lo_1609 = {dataGroup_lo_hi_1609, dataGroup_lo_lo_1609};
  wire [1023:0] dataGroup_hi_1609 = {dataGroup_hi_hi_1609, dataGroup_hi_lo_1609};
  wire [15:0]   dataGroup_9_64 = dataGroup_hi_1609[143:128];
  wire [1023:0] dataGroup_lo_1610 = {dataGroup_lo_hi_1610, dataGroup_lo_lo_1610};
  wire [1023:0] dataGroup_hi_1610 = {dataGroup_hi_hi_1610, dataGroup_hi_lo_1610};
  wire [15:0]   dataGroup_10_64 = dataGroup_hi_1610[271:256];
  wire [1023:0] dataGroup_lo_1611 = {dataGroup_lo_hi_1611, dataGroup_lo_lo_1611};
  wire [1023:0] dataGroup_hi_1611 = {dataGroup_hi_hi_1611, dataGroup_hi_lo_1611};
  wire [15:0]   dataGroup_11_64 = dataGroup_hi_1611[399:384];
  wire [1023:0] dataGroup_lo_1612 = {dataGroup_lo_hi_1612, dataGroup_lo_lo_1612};
  wire [1023:0] dataGroup_hi_1612 = {dataGroup_hi_hi_1612, dataGroup_hi_lo_1612};
  wire [15:0]   dataGroup_12_64 = dataGroup_hi_1612[527:512];
  wire [1023:0] dataGroup_lo_1613 = {dataGroup_lo_hi_1613, dataGroup_lo_lo_1613};
  wire [1023:0] dataGroup_hi_1613 = {dataGroup_hi_hi_1613, dataGroup_hi_lo_1613};
  wire [15:0]   dataGroup_13_64 = dataGroup_hi_1613[655:640];
  wire [1023:0] dataGroup_lo_1614 = {dataGroup_lo_hi_1614, dataGroup_lo_lo_1614};
  wire [1023:0] dataGroup_hi_1614 = {dataGroup_hi_hi_1614, dataGroup_hi_lo_1614};
  wire [15:0]   dataGroup_14_64 = dataGroup_hi_1614[783:768];
  wire [1023:0] dataGroup_lo_1615 = {dataGroup_lo_hi_1615, dataGroup_lo_lo_1615};
  wire [1023:0] dataGroup_hi_1615 = {dataGroup_hi_hi_1615, dataGroup_hi_lo_1615};
  wire [15:0]   dataGroup_15_64 = dataGroup_hi_1615[911:896];
  wire [31:0]   res_lo_lo_lo_64 = {dataGroup_1_64, dataGroup_0_64};
  wire [31:0]   res_lo_lo_hi_64 = {dataGroup_3_64, dataGroup_2_64};
  wire [63:0]   res_lo_lo_64 = {res_lo_lo_hi_64, res_lo_lo_lo_64};
  wire [31:0]   res_lo_hi_lo_64 = {dataGroup_5_64, dataGroup_4_64};
  wire [31:0]   res_lo_hi_hi_64 = {dataGroup_7_64, dataGroup_6_64};
  wire [63:0]   res_lo_hi_64 = {res_lo_hi_hi_64, res_lo_hi_lo_64};
  wire [127:0]  res_lo_64 = {res_lo_hi_64, res_lo_lo_64};
  wire [31:0]   res_hi_lo_lo_64 = {dataGroup_9_64, dataGroup_8_64};
  wire [31:0]   res_hi_lo_hi_64 = {dataGroup_11_64, dataGroup_10_64};
  wire [63:0]   res_hi_lo_64 = {res_hi_lo_hi_64, res_hi_lo_lo_64};
  wire [31:0]   res_hi_hi_lo_64 = {dataGroup_13_64, dataGroup_12_64};
  wire [31:0]   res_hi_hi_hi_64 = {dataGroup_15_64, dataGroup_14_64};
  wire [63:0]   res_hi_hi_64 = {res_hi_hi_hi_64, res_hi_hi_lo_64};
  wire [127:0]  res_hi_64 = {res_hi_hi_64, res_hi_lo_64};
  wire [255:0]  res_120 = {res_hi_64, res_lo_64};
  wire [1023:0] dataGroup_lo_1616 = {dataGroup_lo_hi_1616, dataGroup_lo_lo_1616};
  wire [1023:0] dataGroup_hi_1616 = {dataGroup_hi_hi_1616, dataGroup_hi_lo_1616};
  wire [15:0]   dataGroup_0_65 = dataGroup_lo_1616[31:16];
  wire [1023:0] dataGroup_lo_1617 = {dataGroup_lo_hi_1617, dataGroup_lo_lo_1617};
  wire [1023:0] dataGroup_hi_1617 = {dataGroup_hi_hi_1617, dataGroup_hi_lo_1617};
  wire [15:0]   dataGroup_1_65 = dataGroup_lo_1617[159:144];
  wire [1023:0] dataGroup_lo_1618 = {dataGroup_lo_hi_1618, dataGroup_lo_lo_1618};
  wire [1023:0] dataGroup_hi_1618 = {dataGroup_hi_hi_1618, dataGroup_hi_lo_1618};
  wire [15:0]   dataGroup_2_65 = dataGroup_lo_1618[287:272];
  wire [1023:0] dataGroup_lo_1619 = {dataGroup_lo_hi_1619, dataGroup_lo_lo_1619};
  wire [1023:0] dataGroup_hi_1619 = {dataGroup_hi_hi_1619, dataGroup_hi_lo_1619};
  wire [15:0]   dataGroup_3_65 = dataGroup_lo_1619[415:400];
  wire [1023:0] dataGroup_lo_1620 = {dataGroup_lo_hi_1620, dataGroup_lo_lo_1620};
  wire [1023:0] dataGroup_hi_1620 = {dataGroup_hi_hi_1620, dataGroup_hi_lo_1620};
  wire [15:0]   dataGroup_4_65 = dataGroup_lo_1620[543:528];
  wire [1023:0] dataGroup_lo_1621 = {dataGroup_lo_hi_1621, dataGroup_lo_lo_1621};
  wire [1023:0] dataGroup_hi_1621 = {dataGroup_hi_hi_1621, dataGroup_hi_lo_1621};
  wire [15:0]   dataGroup_5_65 = dataGroup_lo_1621[671:656];
  wire [1023:0] dataGroup_lo_1622 = {dataGroup_lo_hi_1622, dataGroup_lo_lo_1622};
  wire [1023:0] dataGroup_hi_1622 = {dataGroup_hi_hi_1622, dataGroup_hi_lo_1622};
  wire [15:0]   dataGroup_6_65 = dataGroup_lo_1622[799:784];
  wire [1023:0] dataGroup_lo_1623 = {dataGroup_lo_hi_1623, dataGroup_lo_lo_1623};
  wire [1023:0] dataGroup_hi_1623 = {dataGroup_hi_hi_1623, dataGroup_hi_lo_1623};
  wire [15:0]   dataGroup_7_65 = dataGroup_lo_1623[927:912];
  wire [1023:0] dataGroup_lo_1624 = {dataGroup_lo_hi_1624, dataGroup_lo_lo_1624};
  wire [1023:0] dataGroup_hi_1624 = {dataGroup_hi_hi_1624, dataGroup_hi_lo_1624};
  wire [15:0]   dataGroup_8_65 = dataGroup_hi_1624[31:16];
  wire [1023:0] dataGroup_lo_1625 = {dataGroup_lo_hi_1625, dataGroup_lo_lo_1625};
  wire [1023:0] dataGroup_hi_1625 = {dataGroup_hi_hi_1625, dataGroup_hi_lo_1625};
  wire [15:0]   dataGroup_9_65 = dataGroup_hi_1625[159:144];
  wire [1023:0] dataGroup_lo_1626 = {dataGroup_lo_hi_1626, dataGroup_lo_lo_1626};
  wire [1023:0] dataGroup_hi_1626 = {dataGroup_hi_hi_1626, dataGroup_hi_lo_1626};
  wire [15:0]   dataGroup_10_65 = dataGroup_hi_1626[287:272];
  wire [1023:0] dataGroup_lo_1627 = {dataGroup_lo_hi_1627, dataGroup_lo_lo_1627};
  wire [1023:0] dataGroup_hi_1627 = {dataGroup_hi_hi_1627, dataGroup_hi_lo_1627};
  wire [15:0]   dataGroup_11_65 = dataGroup_hi_1627[415:400];
  wire [1023:0] dataGroup_lo_1628 = {dataGroup_lo_hi_1628, dataGroup_lo_lo_1628};
  wire [1023:0] dataGroup_hi_1628 = {dataGroup_hi_hi_1628, dataGroup_hi_lo_1628};
  wire [15:0]   dataGroup_12_65 = dataGroup_hi_1628[543:528];
  wire [1023:0] dataGroup_lo_1629 = {dataGroup_lo_hi_1629, dataGroup_lo_lo_1629};
  wire [1023:0] dataGroup_hi_1629 = {dataGroup_hi_hi_1629, dataGroup_hi_lo_1629};
  wire [15:0]   dataGroup_13_65 = dataGroup_hi_1629[671:656];
  wire [1023:0] dataGroup_lo_1630 = {dataGroup_lo_hi_1630, dataGroup_lo_lo_1630};
  wire [1023:0] dataGroup_hi_1630 = {dataGroup_hi_hi_1630, dataGroup_hi_lo_1630};
  wire [15:0]   dataGroup_14_65 = dataGroup_hi_1630[799:784];
  wire [1023:0] dataGroup_lo_1631 = {dataGroup_lo_hi_1631, dataGroup_lo_lo_1631};
  wire [1023:0] dataGroup_hi_1631 = {dataGroup_hi_hi_1631, dataGroup_hi_lo_1631};
  wire [15:0]   dataGroup_15_65 = dataGroup_hi_1631[927:912];
  wire [31:0]   res_lo_lo_lo_65 = {dataGroup_1_65, dataGroup_0_65};
  wire [31:0]   res_lo_lo_hi_65 = {dataGroup_3_65, dataGroup_2_65};
  wire [63:0]   res_lo_lo_65 = {res_lo_lo_hi_65, res_lo_lo_lo_65};
  wire [31:0]   res_lo_hi_lo_65 = {dataGroup_5_65, dataGroup_4_65};
  wire [31:0]   res_lo_hi_hi_65 = {dataGroup_7_65, dataGroup_6_65};
  wire [63:0]   res_lo_hi_65 = {res_lo_hi_hi_65, res_lo_hi_lo_65};
  wire [127:0]  res_lo_65 = {res_lo_hi_65, res_lo_lo_65};
  wire [31:0]   res_hi_lo_lo_65 = {dataGroup_9_65, dataGroup_8_65};
  wire [31:0]   res_hi_lo_hi_65 = {dataGroup_11_65, dataGroup_10_65};
  wire [63:0]   res_hi_lo_65 = {res_hi_lo_hi_65, res_hi_lo_lo_65};
  wire [31:0]   res_hi_hi_lo_65 = {dataGroup_13_65, dataGroup_12_65};
  wire [31:0]   res_hi_hi_hi_65 = {dataGroup_15_65, dataGroup_14_65};
  wire [63:0]   res_hi_hi_65 = {res_hi_hi_hi_65, res_hi_hi_lo_65};
  wire [127:0]  res_hi_65 = {res_hi_hi_65, res_hi_lo_65};
  wire [255:0]  res_121 = {res_hi_65, res_lo_65};
  wire [1023:0] dataGroup_lo_1632 = {dataGroup_lo_hi_1632, dataGroup_lo_lo_1632};
  wire [1023:0] dataGroup_hi_1632 = {dataGroup_hi_hi_1632, dataGroup_hi_lo_1632};
  wire [15:0]   dataGroup_0_66 = dataGroup_lo_1632[47:32];
  wire [1023:0] dataGroup_lo_1633 = {dataGroup_lo_hi_1633, dataGroup_lo_lo_1633};
  wire [1023:0] dataGroup_hi_1633 = {dataGroup_hi_hi_1633, dataGroup_hi_lo_1633};
  wire [15:0]   dataGroup_1_66 = dataGroup_lo_1633[175:160];
  wire [1023:0] dataGroup_lo_1634 = {dataGroup_lo_hi_1634, dataGroup_lo_lo_1634};
  wire [1023:0] dataGroup_hi_1634 = {dataGroup_hi_hi_1634, dataGroup_hi_lo_1634};
  wire [15:0]   dataGroup_2_66 = dataGroup_lo_1634[303:288];
  wire [1023:0] dataGroup_lo_1635 = {dataGroup_lo_hi_1635, dataGroup_lo_lo_1635};
  wire [1023:0] dataGroup_hi_1635 = {dataGroup_hi_hi_1635, dataGroup_hi_lo_1635};
  wire [15:0]   dataGroup_3_66 = dataGroup_lo_1635[431:416];
  wire [1023:0] dataGroup_lo_1636 = {dataGroup_lo_hi_1636, dataGroup_lo_lo_1636};
  wire [1023:0] dataGroup_hi_1636 = {dataGroup_hi_hi_1636, dataGroup_hi_lo_1636};
  wire [15:0]   dataGroup_4_66 = dataGroup_lo_1636[559:544];
  wire [1023:0] dataGroup_lo_1637 = {dataGroup_lo_hi_1637, dataGroup_lo_lo_1637};
  wire [1023:0] dataGroup_hi_1637 = {dataGroup_hi_hi_1637, dataGroup_hi_lo_1637};
  wire [15:0]   dataGroup_5_66 = dataGroup_lo_1637[687:672];
  wire [1023:0] dataGroup_lo_1638 = {dataGroup_lo_hi_1638, dataGroup_lo_lo_1638};
  wire [1023:0] dataGroup_hi_1638 = {dataGroup_hi_hi_1638, dataGroup_hi_lo_1638};
  wire [15:0]   dataGroup_6_66 = dataGroup_lo_1638[815:800];
  wire [1023:0] dataGroup_lo_1639 = {dataGroup_lo_hi_1639, dataGroup_lo_lo_1639};
  wire [1023:0] dataGroup_hi_1639 = {dataGroup_hi_hi_1639, dataGroup_hi_lo_1639};
  wire [15:0]   dataGroup_7_66 = dataGroup_lo_1639[943:928];
  wire [1023:0] dataGroup_lo_1640 = {dataGroup_lo_hi_1640, dataGroup_lo_lo_1640};
  wire [1023:0] dataGroup_hi_1640 = {dataGroup_hi_hi_1640, dataGroup_hi_lo_1640};
  wire [15:0]   dataGroup_8_66 = dataGroup_hi_1640[47:32];
  wire [1023:0] dataGroup_lo_1641 = {dataGroup_lo_hi_1641, dataGroup_lo_lo_1641};
  wire [1023:0] dataGroup_hi_1641 = {dataGroup_hi_hi_1641, dataGroup_hi_lo_1641};
  wire [15:0]   dataGroup_9_66 = dataGroup_hi_1641[175:160];
  wire [1023:0] dataGroup_lo_1642 = {dataGroup_lo_hi_1642, dataGroup_lo_lo_1642};
  wire [1023:0] dataGroup_hi_1642 = {dataGroup_hi_hi_1642, dataGroup_hi_lo_1642};
  wire [15:0]   dataGroup_10_66 = dataGroup_hi_1642[303:288];
  wire [1023:0] dataGroup_lo_1643 = {dataGroup_lo_hi_1643, dataGroup_lo_lo_1643};
  wire [1023:0] dataGroup_hi_1643 = {dataGroup_hi_hi_1643, dataGroup_hi_lo_1643};
  wire [15:0]   dataGroup_11_66 = dataGroup_hi_1643[431:416];
  wire [1023:0] dataGroup_lo_1644 = {dataGroup_lo_hi_1644, dataGroup_lo_lo_1644};
  wire [1023:0] dataGroup_hi_1644 = {dataGroup_hi_hi_1644, dataGroup_hi_lo_1644};
  wire [15:0]   dataGroup_12_66 = dataGroup_hi_1644[559:544];
  wire [1023:0] dataGroup_lo_1645 = {dataGroup_lo_hi_1645, dataGroup_lo_lo_1645};
  wire [1023:0] dataGroup_hi_1645 = {dataGroup_hi_hi_1645, dataGroup_hi_lo_1645};
  wire [15:0]   dataGroup_13_66 = dataGroup_hi_1645[687:672];
  wire [1023:0] dataGroup_lo_1646 = {dataGroup_lo_hi_1646, dataGroup_lo_lo_1646};
  wire [1023:0] dataGroup_hi_1646 = {dataGroup_hi_hi_1646, dataGroup_hi_lo_1646};
  wire [15:0]   dataGroup_14_66 = dataGroup_hi_1646[815:800];
  wire [1023:0] dataGroup_lo_1647 = {dataGroup_lo_hi_1647, dataGroup_lo_lo_1647};
  wire [1023:0] dataGroup_hi_1647 = {dataGroup_hi_hi_1647, dataGroup_hi_lo_1647};
  wire [15:0]   dataGroup_15_66 = dataGroup_hi_1647[943:928];
  wire [31:0]   res_lo_lo_lo_66 = {dataGroup_1_66, dataGroup_0_66};
  wire [31:0]   res_lo_lo_hi_66 = {dataGroup_3_66, dataGroup_2_66};
  wire [63:0]   res_lo_lo_66 = {res_lo_lo_hi_66, res_lo_lo_lo_66};
  wire [31:0]   res_lo_hi_lo_66 = {dataGroup_5_66, dataGroup_4_66};
  wire [31:0]   res_lo_hi_hi_66 = {dataGroup_7_66, dataGroup_6_66};
  wire [63:0]   res_lo_hi_66 = {res_lo_hi_hi_66, res_lo_hi_lo_66};
  wire [127:0]  res_lo_66 = {res_lo_hi_66, res_lo_lo_66};
  wire [31:0]   res_hi_lo_lo_66 = {dataGroup_9_66, dataGroup_8_66};
  wire [31:0]   res_hi_lo_hi_66 = {dataGroup_11_66, dataGroup_10_66};
  wire [63:0]   res_hi_lo_66 = {res_hi_lo_hi_66, res_hi_lo_lo_66};
  wire [31:0]   res_hi_hi_lo_66 = {dataGroup_13_66, dataGroup_12_66};
  wire [31:0]   res_hi_hi_hi_66 = {dataGroup_15_66, dataGroup_14_66};
  wire [63:0]   res_hi_hi_66 = {res_hi_hi_hi_66, res_hi_hi_lo_66};
  wire [127:0]  res_hi_66 = {res_hi_hi_66, res_hi_lo_66};
  wire [255:0]  res_122 = {res_hi_66, res_lo_66};
  wire [1023:0] dataGroup_lo_1648 = {dataGroup_lo_hi_1648, dataGroup_lo_lo_1648};
  wire [1023:0] dataGroup_hi_1648 = {dataGroup_hi_hi_1648, dataGroup_hi_lo_1648};
  wire [15:0]   dataGroup_0_67 = dataGroup_lo_1648[63:48];
  wire [1023:0] dataGroup_lo_1649 = {dataGroup_lo_hi_1649, dataGroup_lo_lo_1649};
  wire [1023:0] dataGroup_hi_1649 = {dataGroup_hi_hi_1649, dataGroup_hi_lo_1649};
  wire [15:0]   dataGroup_1_67 = dataGroup_lo_1649[191:176];
  wire [1023:0] dataGroup_lo_1650 = {dataGroup_lo_hi_1650, dataGroup_lo_lo_1650};
  wire [1023:0] dataGroup_hi_1650 = {dataGroup_hi_hi_1650, dataGroup_hi_lo_1650};
  wire [15:0]   dataGroup_2_67 = dataGroup_lo_1650[319:304];
  wire [1023:0] dataGroup_lo_1651 = {dataGroup_lo_hi_1651, dataGroup_lo_lo_1651};
  wire [1023:0] dataGroup_hi_1651 = {dataGroup_hi_hi_1651, dataGroup_hi_lo_1651};
  wire [15:0]   dataGroup_3_67 = dataGroup_lo_1651[447:432];
  wire [1023:0] dataGroup_lo_1652 = {dataGroup_lo_hi_1652, dataGroup_lo_lo_1652};
  wire [1023:0] dataGroup_hi_1652 = {dataGroup_hi_hi_1652, dataGroup_hi_lo_1652};
  wire [15:0]   dataGroup_4_67 = dataGroup_lo_1652[575:560];
  wire [1023:0] dataGroup_lo_1653 = {dataGroup_lo_hi_1653, dataGroup_lo_lo_1653};
  wire [1023:0] dataGroup_hi_1653 = {dataGroup_hi_hi_1653, dataGroup_hi_lo_1653};
  wire [15:0]   dataGroup_5_67 = dataGroup_lo_1653[703:688];
  wire [1023:0] dataGroup_lo_1654 = {dataGroup_lo_hi_1654, dataGroup_lo_lo_1654};
  wire [1023:0] dataGroup_hi_1654 = {dataGroup_hi_hi_1654, dataGroup_hi_lo_1654};
  wire [15:0]   dataGroup_6_67 = dataGroup_lo_1654[831:816];
  wire [1023:0] dataGroup_lo_1655 = {dataGroup_lo_hi_1655, dataGroup_lo_lo_1655};
  wire [1023:0] dataGroup_hi_1655 = {dataGroup_hi_hi_1655, dataGroup_hi_lo_1655};
  wire [15:0]   dataGroup_7_67 = dataGroup_lo_1655[959:944];
  wire [1023:0] dataGroup_lo_1656 = {dataGroup_lo_hi_1656, dataGroup_lo_lo_1656};
  wire [1023:0] dataGroup_hi_1656 = {dataGroup_hi_hi_1656, dataGroup_hi_lo_1656};
  wire [15:0]   dataGroup_8_67 = dataGroup_hi_1656[63:48];
  wire [1023:0] dataGroup_lo_1657 = {dataGroup_lo_hi_1657, dataGroup_lo_lo_1657};
  wire [1023:0] dataGroup_hi_1657 = {dataGroup_hi_hi_1657, dataGroup_hi_lo_1657};
  wire [15:0]   dataGroup_9_67 = dataGroup_hi_1657[191:176];
  wire [1023:0] dataGroup_lo_1658 = {dataGroup_lo_hi_1658, dataGroup_lo_lo_1658};
  wire [1023:0] dataGroup_hi_1658 = {dataGroup_hi_hi_1658, dataGroup_hi_lo_1658};
  wire [15:0]   dataGroup_10_67 = dataGroup_hi_1658[319:304];
  wire [1023:0] dataGroup_lo_1659 = {dataGroup_lo_hi_1659, dataGroup_lo_lo_1659};
  wire [1023:0] dataGroup_hi_1659 = {dataGroup_hi_hi_1659, dataGroup_hi_lo_1659};
  wire [15:0]   dataGroup_11_67 = dataGroup_hi_1659[447:432];
  wire [1023:0] dataGroup_lo_1660 = {dataGroup_lo_hi_1660, dataGroup_lo_lo_1660};
  wire [1023:0] dataGroup_hi_1660 = {dataGroup_hi_hi_1660, dataGroup_hi_lo_1660};
  wire [15:0]   dataGroup_12_67 = dataGroup_hi_1660[575:560];
  wire [1023:0] dataGroup_lo_1661 = {dataGroup_lo_hi_1661, dataGroup_lo_lo_1661};
  wire [1023:0] dataGroup_hi_1661 = {dataGroup_hi_hi_1661, dataGroup_hi_lo_1661};
  wire [15:0]   dataGroup_13_67 = dataGroup_hi_1661[703:688];
  wire [1023:0] dataGroup_lo_1662 = {dataGroup_lo_hi_1662, dataGroup_lo_lo_1662};
  wire [1023:0] dataGroup_hi_1662 = {dataGroup_hi_hi_1662, dataGroup_hi_lo_1662};
  wire [15:0]   dataGroup_14_67 = dataGroup_hi_1662[831:816];
  wire [1023:0] dataGroup_lo_1663 = {dataGroup_lo_hi_1663, dataGroup_lo_lo_1663};
  wire [1023:0] dataGroup_hi_1663 = {dataGroup_hi_hi_1663, dataGroup_hi_lo_1663};
  wire [15:0]   dataGroup_15_67 = dataGroup_hi_1663[959:944];
  wire [31:0]   res_lo_lo_lo_67 = {dataGroup_1_67, dataGroup_0_67};
  wire [31:0]   res_lo_lo_hi_67 = {dataGroup_3_67, dataGroup_2_67};
  wire [63:0]   res_lo_lo_67 = {res_lo_lo_hi_67, res_lo_lo_lo_67};
  wire [31:0]   res_lo_hi_lo_67 = {dataGroup_5_67, dataGroup_4_67};
  wire [31:0]   res_lo_hi_hi_67 = {dataGroup_7_67, dataGroup_6_67};
  wire [63:0]   res_lo_hi_67 = {res_lo_hi_hi_67, res_lo_hi_lo_67};
  wire [127:0]  res_lo_67 = {res_lo_hi_67, res_lo_lo_67};
  wire [31:0]   res_hi_lo_lo_67 = {dataGroup_9_67, dataGroup_8_67};
  wire [31:0]   res_hi_lo_hi_67 = {dataGroup_11_67, dataGroup_10_67};
  wire [63:0]   res_hi_lo_67 = {res_hi_lo_hi_67, res_hi_lo_lo_67};
  wire [31:0]   res_hi_hi_lo_67 = {dataGroup_13_67, dataGroup_12_67};
  wire [31:0]   res_hi_hi_hi_67 = {dataGroup_15_67, dataGroup_14_67};
  wire [63:0]   res_hi_hi_67 = {res_hi_hi_hi_67, res_hi_hi_lo_67};
  wire [127:0]  res_hi_67 = {res_hi_hi_67, res_hi_lo_67};
  wire [255:0]  res_123 = {res_hi_67, res_lo_67};
  wire [1023:0] dataGroup_lo_1664 = {dataGroup_lo_hi_1664, dataGroup_lo_lo_1664};
  wire [1023:0] dataGroup_hi_1664 = {dataGroup_hi_hi_1664, dataGroup_hi_lo_1664};
  wire [15:0]   dataGroup_0_68 = dataGroup_lo_1664[79:64];
  wire [1023:0] dataGroup_lo_1665 = {dataGroup_lo_hi_1665, dataGroup_lo_lo_1665};
  wire [1023:0] dataGroup_hi_1665 = {dataGroup_hi_hi_1665, dataGroup_hi_lo_1665};
  wire [15:0]   dataGroup_1_68 = dataGroup_lo_1665[207:192];
  wire [1023:0] dataGroup_lo_1666 = {dataGroup_lo_hi_1666, dataGroup_lo_lo_1666};
  wire [1023:0] dataGroup_hi_1666 = {dataGroup_hi_hi_1666, dataGroup_hi_lo_1666};
  wire [15:0]   dataGroup_2_68 = dataGroup_lo_1666[335:320];
  wire [1023:0] dataGroup_lo_1667 = {dataGroup_lo_hi_1667, dataGroup_lo_lo_1667};
  wire [1023:0] dataGroup_hi_1667 = {dataGroup_hi_hi_1667, dataGroup_hi_lo_1667};
  wire [15:0]   dataGroup_3_68 = dataGroup_lo_1667[463:448];
  wire [1023:0] dataGroup_lo_1668 = {dataGroup_lo_hi_1668, dataGroup_lo_lo_1668};
  wire [1023:0] dataGroup_hi_1668 = {dataGroup_hi_hi_1668, dataGroup_hi_lo_1668};
  wire [15:0]   dataGroup_4_68 = dataGroup_lo_1668[591:576];
  wire [1023:0] dataGroup_lo_1669 = {dataGroup_lo_hi_1669, dataGroup_lo_lo_1669};
  wire [1023:0] dataGroup_hi_1669 = {dataGroup_hi_hi_1669, dataGroup_hi_lo_1669};
  wire [15:0]   dataGroup_5_68 = dataGroup_lo_1669[719:704];
  wire [1023:0] dataGroup_lo_1670 = {dataGroup_lo_hi_1670, dataGroup_lo_lo_1670};
  wire [1023:0] dataGroup_hi_1670 = {dataGroup_hi_hi_1670, dataGroup_hi_lo_1670};
  wire [15:0]   dataGroup_6_68 = dataGroup_lo_1670[847:832];
  wire [1023:0] dataGroup_lo_1671 = {dataGroup_lo_hi_1671, dataGroup_lo_lo_1671};
  wire [1023:0] dataGroup_hi_1671 = {dataGroup_hi_hi_1671, dataGroup_hi_lo_1671};
  wire [15:0]   dataGroup_7_68 = dataGroup_lo_1671[975:960];
  wire [1023:0] dataGroup_lo_1672 = {dataGroup_lo_hi_1672, dataGroup_lo_lo_1672};
  wire [1023:0] dataGroup_hi_1672 = {dataGroup_hi_hi_1672, dataGroup_hi_lo_1672};
  wire [15:0]   dataGroup_8_68 = dataGroup_hi_1672[79:64];
  wire [1023:0] dataGroup_lo_1673 = {dataGroup_lo_hi_1673, dataGroup_lo_lo_1673};
  wire [1023:0] dataGroup_hi_1673 = {dataGroup_hi_hi_1673, dataGroup_hi_lo_1673};
  wire [15:0]   dataGroup_9_68 = dataGroup_hi_1673[207:192];
  wire [1023:0] dataGroup_lo_1674 = {dataGroup_lo_hi_1674, dataGroup_lo_lo_1674};
  wire [1023:0] dataGroup_hi_1674 = {dataGroup_hi_hi_1674, dataGroup_hi_lo_1674};
  wire [15:0]   dataGroup_10_68 = dataGroup_hi_1674[335:320];
  wire [1023:0] dataGroup_lo_1675 = {dataGroup_lo_hi_1675, dataGroup_lo_lo_1675};
  wire [1023:0] dataGroup_hi_1675 = {dataGroup_hi_hi_1675, dataGroup_hi_lo_1675};
  wire [15:0]   dataGroup_11_68 = dataGroup_hi_1675[463:448];
  wire [1023:0] dataGroup_lo_1676 = {dataGroup_lo_hi_1676, dataGroup_lo_lo_1676};
  wire [1023:0] dataGroup_hi_1676 = {dataGroup_hi_hi_1676, dataGroup_hi_lo_1676};
  wire [15:0]   dataGroup_12_68 = dataGroup_hi_1676[591:576];
  wire [1023:0] dataGroup_lo_1677 = {dataGroup_lo_hi_1677, dataGroup_lo_lo_1677};
  wire [1023:0] dataGroup_hi_1677 = {dataGroup_hi_hi_1677, dataGroup_hi_lo_1677};
  wire [15:0]   dataGroup_13_68 = dataGroup_hi_1677[719:704];
  wire [1023:0] dataGroup_lo_1678 = {dataGroup_lo_hi_1678, dataGroup_lo_lo_1678};
  wire [1023:0] dataGroup_hi_1678 = {dataGroup_hi_hi_1678, dataGroup_hi_lo_1678};
  wire [15:0]   dataGroup_14_68 = dataGroup_hi_1678[847:832];
  wire [1023:0] dataGroup_lo_1679 = {dataGroup_lo_hi_1679, dataGroup_lo_lo_1679};
  wire [1023:0] dataGroup_hi_1679 = {dataGroup_hi_hi_1679, dataGroup_hi_lo_1679};
  wire [15:0]   dataGroup_15_68 = dataGroup_hi_1679[975:960];
  wire [31:0]   res_lo_lo_lo_68 = {dataGroup_1_68, dataGroup_0_68};
  wire [31:0]   res_lo_lo_hi_68 = {dataGroup_3_68, dataGroup_2_68};
  wire [63:0]   res_lo_lo_68 = {res_lo_lo_hi_68, res_lo_lo_lo_68};
  wire [31:0]   res_lo_hi_lo_68 = {dataGroup_5_68, dataGroup_4_68};
  wire [31:0]   res_lo_hi_hi_68 = {dataGroup_7_68, dataGroup_6_68};
  wire [63:0]   res_lo_hi_68 = {res_lo_hi_hi_68, res_lo_hi_lo_68};
  wire [127:0]  res_lo_68 = {res_lo_hi_68, res_lo_lo_68};
  wire [31:0]   res_hi_lo_lo_68 = {dataGroup_9_68, dataGroup_8_68};
  wire [31:0]   res_hi_lo_hi_68 = {dataGroup_11_68, dataGroup_10_68};
  wire [63:0]   res_hi_lo_68 = {res_hi_lo_hi_68, res_hi_lo_lo_68};
  wire [31:0]   res_hi_hi_lo_68 = {dataGroup_13_68, dataGroup_12_68};
  wire [31:0]   res_hi_hi_hi_68 = {dataGroup_15_68, dataGroup_14_68};
  wire [63:0]   res_hi_hi_68 = {res_hi_hi_hi_68, res_hi_hi_lo_68};
  wire [127:0]  res_hi_68 = {res_hi_hi_68, res_hi_lo_68};
  wire [255:0]  res_124 = {res_hi_68, res_lo_68};
  wire [1023:0] dataGroup_lo_1680 = {dataGroup_lo_hi_1680, dataGroup_lo_lo_1680};
  wire [1023:0] dataGroup_hi_1680 = {dataGroup_hi_hi_1680, dataGroup_hi_lo_1680};
  wire [15:0]   dataGroup_0_69 = dataGroup_lo_1680[95:80];
  wire [1023:0] dataGroup_lo_1681 = {dataGroup_lo_hi_1681, dataGroup_lo_lo_1681};
  wire [1023:0] dataGroup_hi_1681 = {dataGroup_hi_hi_1681, dataGroup_hi_lo_1681};
  wire [15:0]   dataGroup_1_69 = dataGroup_lo_1681[223:208];
  wire [1023:0] dataGroup_lo_1682 = {dataGroup_lo_hi_1682, dataGroup_lo_lo_1682};
  wire [1023:0] dataGroup_hi_1682 = {dataGroup_hi_hi_1682, dataGroup_hi_lo_1682};
  wire [15:0]   dataGroup_2_69 = dataGroup_lo_1682[351:336];
  wire [1023:0] dataGroup_lo_1683 = {dataGroup_lo_hi_1683, dataGroup_lo_lo_1683};
  wire [1023:0] dataGroup_hi_1683 = {dataGroup_hi_hi_1683, dataGroup_hi_lo_1683};
  wire [15:0]   dataGroup_3_69 = dataGroup_lo_1683[479:464];
  wire [1023:0] dataGroup_lo_1684 = {dataGroup_lo_hi_1684, dataGroup_lo_lo_1684};
  wire [1023:0] dataGroup_hi_1684 = {dataGroup_hi_hi_1684, dataGroup_hi_lo_1684};
  wire [15:0]   dataGroup_4_69 = dataGroup_lo_1684[607:592];
  wire [1023:0] dataGroup_lo_1685 = {dataGroup_lo_hi_1685, dataGroup_lo_lo_1685};
  wire [1023:0] dataGroup_hi_1685 = {dataGroup_hi_hi_1685, dataGroup_hi_lo_1685};
  wire [15:0]   dataGroup_5_69 = dataGroup_lo_1685[735:720];
  wire [1023:0] dataGroup_lo_1686 = {dataGroup_lo_hi_1686, dataGroup_lo_lo_1686};
  wire [1023:0] dataGroup_hi_1686 = {dataGroup_hi_hi_1686, dataGroup_hi_lo_1686};
  wire [15:0]   dataGroup_6_69 = dataGroup_lo_1686[863:848];
  wire [1023:0] dataGroup_lo_1687 = {dataGroup_lo_hi_1687, dataGroup_lo_lo_1687};
  wire [1023:0] dataGroup_hi_1687 = {dataGroup_hi_hi_1687, dataGroup_hi_lo_1687};
  wire [15:0]   dataGroup_7_69 = dataGroup_lo_1687[991:976];
  wire [1023:0] dataGroup_lo_1688 = {dataGroup_lo_hi_1688, dataGroup_lo_lo_1688};
  wire [1023:0] dataGroup_hi_1688 = {dataGroup_hi_hi_1688, dataGroup_hi_lo_1688};
  wire [15:0]   dataGroup_8_69 = dataGroup_hi_1688[95:80];
  wire [1023:0] dataGroup_lo_1689 = {dataGroup_lo_hi_1689, dataGroup_lo_lo_1689};
  wire [1023:0] dataGroup_hi_1689 = {dataGroup_hi_hi_1689, dataGroup_hi_lo_1689};
  wire [15:0]   dataGroup_9_69 = dataGroup_hi_1689[223:208];
  wire [1023:0] dataGroup_lo_1690 = {dataGroup_lo_hi_1690, dataGroup_lo_lo_1690};
  wire [1023:0] dataGroup_hi_1690 = {dataGroup_hi_hi_1690, dataGroup_hi_lo_1690};
  wire [15:0]   dataGroup_10_69 = dataGroup_hi_1690[351:336];
  wire [1023:0] dataGroup_lo_1691 = {dataGroup_lo_hi_1691, dataGroup_lo_lo_1691};
  wire [1023:0] dataGroup_hi_1691 = {dataGroup_hi_hi_1691, dataGroup_hi_lo_1691};
  wire [15:0]   dataGroup_11_69 = dataGroup_hi_1691[479:464];
  wire [1023:0] dataGroup_lo_1692 = {dataGroup_lo_hi_1692, dataGroup_lo_lo_1692};
  wire [1023:0] dataGroup_hi_1692 = {dataGroup_hi_hi_1692, dataGroup_hi_lo_1692};
  wire [15:0]   dataGroup_12_69 = dataGroup_hi_1692[607:592];
  wire [1023:0] dataGroup_lo_1693 = {dataGroup_lo_hi_1693, dataGroup_lo_lo_1693};
  wire [1023:0] dataGroup_hi_1693 = {dataGroup_hi_hi_1693, dataGroup_hi_lo_1693};
  wire [15:0]   dataGroup_13_69 = dataGroup_hi_1693[735:720];
  wire [1023:0] dataGroup_lo_1694 = {dataGroup_lo_hi_1694, dataGroup_lo_lo_1694};
  wire [1023:0] dataGroup_hi_1694 = {dataGroup_hi_hi_1694, dataGroup_hi_lo_1694};
  wire [15:0]   dataGroup_14_69 = dataGroup_hi_1694[863:848];
  wire [1023:0] dataGroup_lo_1695 = {dataGroup_lo_hi_1695, dataGroup_lo_lo_1695};
  wire [1023:0] dataGroup_hi_1695 = {dataGroup_hi_hi_1695, dataGroup_hi_lo_1695};
  wire [15:0]   dataGroup_15_69 = dataGroup_hi_1695[991:976];
  wire [31:0]   res_lo_lo_lo_69 = {dataGroup_1_69, dataGroup_0_69};
  wire [31:0]   res_lo_lo_hi_69 = {dataGroup_3_69, dataGroup_2_69};
  wire [63:0]   res_lo_lo_69 = {res_lo_lo_hi_69, res_lo_lo_lo_69};
  wire [31:0]   res_lo_hi_lo_69 = {dataGroup_5_69, dataGroup_4_69};
  wire [31:0]   res_lo_hi_hi_69 = {dataGroup_7_69, dataGroup_6_69};
  wire [63:0]   res_lo_hi_69 = {res_lo_hi_hi_69, res_lo_hi_lo_69};
  wire [127:0]  res_lo_69 = {res_lo_hi_69, res_lo_lo_69};
  wire [31:0]   res_hi_lo_lo_69 = {dataGroup_9_69, dataGroup_8_69};
  wire [31:0]   res_hi_lo_hi_69 = {dataGroup_11_69, dataGroup_10_69};
  wire [63:0]   res_hi_lo_69 = {res_hi_lo_hi_69, res_hi_lo_lo_69};
  wire [31:0]   res_hi_hi_lo_69 = {dataGroup_13_69, dataGroup_12_69};
  wire [31:0]   res_hi_hi_hi_69 = {dataGroup_15_69, dataGroup_14_69};
  wire [63:0]   res_hi_hi_69 = {res_hi_hi_hi_69, res_hi_hi_lo_69};
  wire [127:0]  res_hi_69 = {res_hi_hi_69, res_hi_lo_69};
  wire [255:0]  res_125 = {res_hi_69, res_lo_69};
  wire [1023:0] dataGroup_lo_1696 = {dataGroup_lo_hi_1696, dataGroup_lo_lo_1696};
  wire [1023:0] dataGroup_hi_1696 = {dataGroup_hi_hi_1696, dataGroup_hi_lo_1696};
  wire [15:0]   dataGroup_0_70 = dataGroup_lo_1696[111:96];
  wire [1023:0] dataGroup_lo_1697 = {dataGroup_lo_hi_1697, dataGroup_lo_lo_1697};
  wire [1023:0] dataGroup_hi_1697 = {dataGroup_hi_hi_1697, dataGroup_hi_lo_1697};
  wire [15:0]   dataGroup_1_70 = dataGroup_lo_1697[239:224];
  wire [1023:0] dataGroup_lo_1698 = {dataGroup_lo_hi_1698, dataGroup_lo_lo_1698};
  wire [1023:0] dataGroup_hi_1698 = {dataGroup_hi_hi_1698, dataGroup_hi_lo_1698};
  wire [15:0]   dataGroup_2_70 = dataGroup_lo_1698[367:352];
  wire [1023:0] dataGroup_lo_1699 = {dataGroup_lo_hi_1699, dataGroup_lo_lo_1699};
  wire [1023:0] dataGroup_hi_1699 = {dataGroup_hi_hi_1699, dataGroup_hi_lo_1699};
  wire [15:0]   dataGroup_3_70 = dataGroup_lo_1699[495:480];
  wire [1023:0] dataGroup_lo_1700 = {dataGroup_lo_hi_1700, dataGroup_lo_lo_1700};
  wire [1023:0] dataGroup_hi_1700 = {dataGroup_hi_hi_1700, dataGroup_hi_lo_1700};
  wire [15:0]   dataGroup_4_70 = dataGroup_lo_1700[623:608];
  wire [1023:0] dataGroup_lo_1701 = {dataGroup_lo_hi_1701, dataGroup_lo_lo_1701};
  wire [1023:0] dataGroup_hi_1701 = {dataGroup_hi_hi_1701, dataGroup_hi_lo_1701};
  wire [15:0]   dataGroup_5_70 = dataGroup_lo_1701[751:736];
  wire [1023:0] dataGroup_lo_1702 = {dataGroup_lo_hi_1702, dataGroup_lo_lo_1702};
  wire [1023:0] dataGroup_hi_1702 = {dataGroup_hi_hi_1702, dataGroup_hi_lo_1702};
  wire [15:0]   dataGroup_6_70 = dataGroup_lo_1702[879:864];
  wire [1023:0] dataGroup_lo_1703 = {dataGroup_lo_hi_1703, dataGroup_lo_lo_1703};
  wire [1023:0] dataGroup_hi_1703 = {dataGroup_hi_hi_1703, dataGroup_hi_lo_1703};
  wire [15:0]   dataGroup_7_70 = dataGroup_lo_1703[1007:992];
  wire [1023:0] dataGroup_lo_1704 = {dataGroup_lo_hi_1704, dataGroup_lo_lo_1704};
  wire [1023:0] dataGroup_hi_1704 = {dataGroup_hi_hi_1704, dataGroup_hi_lo_1704};
  wire [15:0]   dataGroup_8_70 = dataGroup_hi_1704[111:96];
  wire [1023:0] dataGroup_lo_1705 = {dataGroup_lo_hi_1705, dataGroup_lo_lo_1705};
  wire [1023:0] dataGroup_hi_1705 = {dataGroup_hi_hi_1705, dataGroup_hi_lo_1705};
  wire [15:0]   dataGroup_9_70 = dataGroup_hi_1705[239:224];
  wire [1023:0] dataGroup_lo_1706 = {dataGroup_lo_hi_1706, dataGroup_lo_lo_1706};
  wire [1023:0] dataGroup_hi_1706 = {dataGroup_hi_hi_1706, dataGroup_hi_lo_1706};
  wire [15:0]   dataGroup_10_70 = dataGroup_hi_1706[367:352];
  wire [1023:0] dataGroup_lo_1707 = {dataGroup_lo_hi_1707, dataGroup_lo_lo_1707};
  wire [1023:0] dataGroup_hi_1707 = {dataGroup_hi_hi_1707, dataGroup_hi_lo_1707};
  wire [15:0]   dataGroup_11_70 = dataGroup_hi_1707[495:480];
  wire [1023:0] dataGroup_lo_1708 = {dataGroup_lo_hi_1708, dataGroup_lo_lo_1708};
  wire [1023:0] dataGroup_hi_1708 = {dataGroup_hi_hi_1708, dataGroup_hi_lo_1708};
  wire [15:0]   dataGroup_12_70 = dataGroup_hi_1708[623:608];
  wire [1023:0] dataGroup_lo_1709 = {dataGroup_lo_hi_1709, dataGroup_lo_lo_1709};
  wire [1023:0] dataGroup_hi_1709 = {dataGroup_hi_hi_1709, dataGroup_hi_lo_1709};
  wire [15:0]   dataGroup_13_70 = dataGroup_hi_1709[751:736];
  wire [1023:0] dataGroup_lo_1710 = {dataGroup_lo_hi_1710, dataGroup_lo_lo_1710};
  wire [1023:0] dataGroup_hi_1710 = {dataGroup_hi_hi_1710, dataGroup_hi_lo_1710};
  wire [15:0]   dataGroup_14_70 = dataGroup_hi_1710[879:864];
  wire [1023:0] dataGroup_lo_1711 = {dataGroup_lo_hi_1711, dataGroup_lo_lo_1711};
  wire [1023:0] dataGroup_hi_1711 = {dataGroup_hi_hi_1711, dataGroup_hi_lo_1711};
  wire [15:0]   dataGroup_15_70 = dataGroup_hi_1711[1007:992];
  wire [31:0]   res_lo_lo_lo_70 = {dataGroup_1_70, dataGroup_0_70};
  wire [31:0]   res_lo_lo_hi_70 = {dataGroup_3_70, dataGroup_2_70};
  wire [63:0]   res_lo_lo_70 = {res_lo_lo_hi_70, res_lo_lo_lo_70};
  wire [31:0]   res_lo_hi_lo_70 = {dataGroup_5_70, dataGroup_4_70};
  wire [31:0]   res_lo_hi_hi_70 = {dataGroup_7_70, dataGroup_6_70};
  wire [63:0]   res_lo_hi_70 = {res_lo_hi_hi_70, res_lo_hi_lo_70};
  wire [127:0]  res_lo_70 = {res_lo_hi_70, res_lo_lo_70};
  wire [31:0]   res_hi_lo_lo_70 = {dataGroup_9_70, dataGroup_8_70};
  wire [31:0]   res_hi_lo_hi_70 = {dataGroup_11_70, dataGroup_10_70};
  wire [63:0]   res_hi_lo_70 = {res_hi_lo_hi_70, res_hi_lo_lo_70};
  wire [31:0]   res_hi_hi_lo_70 = {dataGroup_13_70, dataGroup_12_70};
  wire [31:0]   res_hi_hi_hi_70 = {dataGroup_15_70, dataGroup_14_70};
  wire [63:0]   res_hi_hi_70 = {res_hi_hi_hi_70, res_hi_hi_lo_70};
  wire [127:0]  res_hi_70 = {res_hi_hi_70, res_hi_lo_70};
  wire [255:0]  res_126 = {res_hi_70, res_lo_70};
  wire [1023:0] dataGroup_lo_1712 = {dataGroup_lo_hi_1712, dataGroup_lo_lo_1712};
  wire [1023:0] dataGroup_hi_1712 = {dataGroup_hi_hi_1712, dataGroup_hi_lo_1712};
  wire [15:0]   dataGroup_0_71 = dataGroup_lo_1712[127:112];
  wire [1023:0] dataGroup_lo_1713 = {dataGroup_lo_hi_1713, dataGroup_lo_lo_1713};
  wire [1023:0] dataGroup_hi_1713 = {dataGroup_hi_hi_1713, dataGroup_hi_lo_1713};
  wire [15:0]   dataGroup_1_71 = dataGroup_lo_1713[255:240];
  wire [1023:0] dataGroup_lo_1714 = {dataGroup_lo_hi_1714, dataGroup_lo_lo_1714};
  wire [1023:0] dataGroup_hi_1714 = {dataGroup_hi_hi_1714, dataGroup_hi_lo_1714};
  wire [15:0]   dataGroup_2_71 = dataGroup_lo_1714[383:368];
  wire [1023:0] dataGroup_lo_1715 = {dataGroup_lo_hi_1715, dataGroup_lo_lo_1715};
  wire [1023:0] dataGroup_hi_1715 = {dataGroup_hi_hi_1715, dataGroup_hi_lo_1715};
  wire [15:0]   dataGroup_3_71 = dataGroup_lo_1715[511:496];
  wire [1023:0] dataGroup_lo_1716 = {dataGroup_lo_hi_1716, dataGroup_lo_lo_1716};
  wire [1023:0] dataGroup_hi_1716 = {dataGroup_hi_hi_1716, dataGroup_hi_lo_1716};
  wire [15:0]   dataGroup_4_71 = dataGroup_lo_1716[639:624];
  wire [1023:0] dataGroup_lo_1717 = {dataGroup_lo_hi_1717, dataGroup_lo_lo_1717};
  wire [1023:0] dataGroup_hi_1717 = {dataGroup_hi_hi_1717, dataGroup_hi_lo_1717};
  wire [15:0]   dataGroup_5_71 = dataGroup_lo_1717[767:752];
  wire [1023:0] dataGroup_lo_1718 = {dataGroup_lo_hi_1718, dataGroup_lo_lo_1718};
  wire [1023:0] dataGroup_hi_1718 = {dataGroup_hi_hi_1718, dataGroup_hi_lo_1718};
  wire [15:0]   dataGroup_6_71 = dataGroup_lo_1718[895:880];
  wire [1023:0] dataGroup_lo_1719 = {dataGroup_lo_hi_1719, dataGroup_lo_lo_1719};
  wire [1023:0] dataGroup_hi_1719 = {dataGroup_hi_hi_1719, dataGroup_hi_lo_1719};
  wire [15:0]   dataGroup_7_71 = dataGroup_lo_1719[1023:1008];
  wire [1023:0] dataGroup_lo_1720 = {dataGroup_lo_hi_1720, dataGroup_lo_lo_1720};
  wire [1023:0] dataGroup_hi_1720 = {dataGroup_hi_hi_1720, dataGroup_hi_lo_1720};
  wire [15:0]   dataGroup_8_71 = dataGroup_hi_1720[127:112];
  wire [1023:0] dataGroup_lo_1721 = {dataGroup_lo_hi_1721, dataGroup_lo_lo_1721};
  wire [1023:0] dataGroup_hi_1721 = {dataGroup_hi_hi_1721, dataGroup_hi_lo_1721};
  wire [15:0]   dataGroup_9_71 = dataGroup_hi_1721[255:240];
  wire [1023:0] dataGroup_lo_1722 = {dataGroup_lo_hi_1722, dataGroup_lo_lo_1722};
  wire [1023:0] dataGroup_hi_1722 = {dataGroup_hi_hi_1722, dataGroup_hi_lo_1722};
  wire [15:0]   dataGroup_10_71 = dataGroup_hi_1722[383:368];
  wire [1023:0] dataGroup_lo_1723 = {dataGroup_lo_hi_1723, dataGroup_lo_lo_1723};
  wire [1023:0] dataGroup_hi_1723 = {dataGroup_hi_hi_1723, dataGroup_hi_lo_1723};
  wire [15:0]   dataGroup_11_71 = dataGroup_hi_1723[511:496];
  wire [1023:0] dataGroup_lo_1724 = {dataGroup_lo_hi_1724, dataGroup_lo_lo_1724};
  wire [1023:0] dataGroup_hi_1724 = {dataGroup_hi_hi_1724, dataGroup_hi_lo_1724};
  wire [15:0]   dataGroup_12_71 = dataGroup_hi_1724[639:624];
  wire [1023:0] dataGroup_lo_1725 = {dataGroup_lo_hi_1725, dataGroup_lo_lo_1725};
  wire [1023:0] dataGroup_hi_1725 = {dataGroup_hi_hi_1725, dataGroup_hi_lo_1725};
  wire [15:0]   dataGroup_13_71 = dataGroup_hi_1725[767:752];
  wire [1023:0] dataGroup_lo_1726 = {dataGroup_lo_hi_1726, dataGroup_lo_lo_1726};
  wire [1023:0] dataGroup_hi_1726 = {dataGroup_hi_hi_1726, dataGroup_hi_lo_1726};
  wire [15:0]   dataGroup_14_71 = dataGroup_hi_1726[895:880];
  wire [1023:0] dataGroup_lo_1727 = {dataGroup_lo_hi_1727, dataGroup_lo_lo_1727};
  wire [1023:0] dataGroup_hi_1727 = {dataGroup_hi_hi_1727, dataGroup_hi_lo_1727};
  wire [15:0]   dataGroup_15_71 = dataGroup_hi_1727[1023:1008];
  wire [31:0]   res_lo_lo_lo_71 = {dataGroup_1_71, dataGroup_0_71};
  wire [31:0]   res_lo_lo_hi_71 = {dataGroup_3_71, dataGroup_2_71};
  wire [63:0]   res_lo_lo_71 = {res_lo_lo_hi_71, res_lo_lo_lo_71};
  wire [31:0]   res_lo_hi_lo_71 = {dataGroup_5_71, dataGroup_4_71};
  wire [31:0]   res_lo_hi_hi_71 = {dataGroup_7_71, dataGroup_6_71};
  wire [63:0]   res_lo_hi_71 = {res_lo_hi_hi_71, res_lo_hi_lo_71};
  wire [127:0]  res_lo_71 = {res_lo_hi_71, res_lo_lo_71};
  wire [31:0]   res_hi_lo_lo_71 = {dataGroup_9_71, dataGroup_8_71};
  wire [31:0]   res_hi_lo_hi_71 = {dataGroup_11_71, dataGroup_10_71};
  wire [63:0]   res_hi_lo_71 = {res_hi_lo_hi_71, res_hi_lo_lo_71};
  wire [31:0]   res_hi_hi_lo_71 = {dataGroup_13_71, dataGroup_12_71};
  wire [31:0]   res_hi_hi_hi_71 = {dataGroup_15_71, dataGroup_14_71};
  wire [63:0]   res_hi_hi_71 = {res_hi_hi_hi_71, res_hi_hi_lo_71};
  wire [127:0]  res_hi_71 = {res_hi_hi_71, res_hi_lo_71};
  wire [255:0]  res_127 = {res_hi_71, res_lo_71};
  wire [511:0]  lo_lo_15 = {res_121, res_120};
  wire [511:0]  lo_hi_15 = {res_123, res_122};
  wire [1023:0] lo_15 = {lo_hi_15, lo_lo_15};
  wire [511:0]  hi_lo_15 = {res_125, res_124};
  wire [511:0]  hi_hi_15 = {res_127, res_126};
  wire [1023:0] hi_15 = {hi_hi_15, hi_lo_15};
  wire [2047:0] regroupLoadData_1_7 = {hi_15, lo_15};
  wire [1023:0] dataGroup_lo_1728 = {dataGroup_lo_hi_1728, dataGroup_lo_lo_1728};
  wire [1023:0] dataGroup_hi_1728 = {dataGroup_hi_hi_1728, dataGroup_hi_lo_1728};
  wire [31:0]   dataGroup_0_72 = dataGroup_lo_1728[31:0];
  wire [1023:0] dataGroup_lo_1729 = {dataGroup_lo_hi_1729, dataGroup_lo_lo_1729};
  wire [1023:0] dataGroup_hi_1729 = {dataGroup_hi_hi_1729, dataGroup_hi_lo_1729};
  wire [31:0]   dataGroup_1_72 = dataGroup_lo_1729[63:32];
  wire [1023:0] dataGroup_lo_1730 = {dataGroup_lo_hi_1730, dataGroup_lo_lo_1730};
  wire [1023:0] dataGroup_hi_1730 = {dataGroup_hi_hi_1730, dataGroup_hi_lo_1730};
  wire [31:0]   dataGroup_2_72 = dataGroup_lo_1730[95:64];
  wire [1023:0] dataGroup_lo_1731 = {dataGroup_lo_hi_1731, dataGroup_lo_lo_1731};
  wire [1023:0] dataGroup_hi_1731 = {dataGroup_hi_hi_1731, dataGroup_hi_lo_1731};
  wire [31:0]   dataGroup_3_72 = dataGroup_lo_1731[127:96];
  wire [1023:0] dataGroup_lo_1732 = {dataGroup_lo_hi_1732, dataGroup_lo_lo_1732};
  wire [1023:0] dataGroup_hi_1732 = {dataGroup_hi_hi_1732, dataGroup_hi_lo_1732};
  wire [31:0]   dataGroup_4_72 = dataGroup_lo_1732[159:128];
  wire [1023:0] dataGroup_lo_1733 = {dataGroup_lo_hi_1733, dataGroup_lo_lo_1733};
  wire [1023:0] dataGroup_hi_1733 = {dataGroup_hi_hi_1733, dataGroup_hi_lo_1733};
  wire [31:0]   dataGroup_5_72 = dataGroup_lo_1733[191:160];
  wire [1023:0] dataGroup_lo_1734 = {dataGroup_lo_hi_1734, dataGroup_lo_lo_1734};
  wire [1023:0] dataGroup_hi_1734 = {dataGroup_hi_hi_1734, dataGroup_hi_lo_1734};
  wire [31:0]   dataGroup_6_72 = dataGroup_lo_1734[223:192];
  wire [1023:0] dataGroup_lo_1735 = {dataGroup_lo_hi_1735, dataGroup_lo_lo_1735};
  wire [1023:0] dataGroup_hi_1735 = {dataGroup_hi_hi_1735, dataGroup_hi_lo_1735};
  wire [31:0]   dataGroup_7_72 = dataGroup_lo_1735[255:224];
  wire [63:0]   res_lo_lo_72 = {dataGroup_1_72, dataGroup_0_72};
  wire [63:0]   res_lo_hi_72 = {dataGroup_3_72, dataGroup_2_72};
  wire [127:0]  res_lo_72 = {res_lo_hi_72, res_lo_lo_72};
  wire [63:0]   res_hi_lo_72 = {dataGroup_5_72, dataGroup_4_72};
  wire [63:0]   res_hi_hi_72 = {dataGroup_7_72, dataGroup_6_72};
  wire [127:0]  res_hi_72 = {res_hi_hi_72, res_hi_lo_72};
  wire [255:0]  res_128 = {res_hi_72, res_lo_72};
  wire [511:0]  lo_lo_16 = {256'h0, res_128};
  wire [1023:0] lo_16 = {512'h0, lo_lo_16};
  wire [2047:0] regroupLoadData_2_0 = {1024'h0, lo_16};
  wire [1023:0] dataGroup_lo_1736 = {dataGroup_lo_hi_1736, dataGroup_lo_lo_1736};
  wire [1023:0] dataGroup_hi_1736 = {dataGroup_hi_hi_1736, dataGroup_hi_lo_1736};
  wire [31:0]   dataGroup_0_73 = dataGroup_lo_1736[31:0];
  wire [1023:0] dataGroup_lo_1737 = {dataGroup_lo_hi_1737, dataGroup_lo_lo_1737};
  wire [1023:0] dataGroup_hi_1737 = {dataGroup_hi_hi_1737, dataGroup_hi_lo_1737};
  wire [31:0]   dataGroup_1_73 = dataGroup_lo_1737[95:64];
  wire [1023:0] dataGroup_lo_1738 = {dataGroup_lo_hi_1738, dataGroup_lo_lo_1738};
  wire [1023:0] dataGroup_hi_1738 = {dataGroup_hi_hi_1738, dataGroup_hi_lo_1738};
  wire [31:0]   dataGroup_2_73 = dataGroup_lo_1738[159:128];
  wire [1023:0] dataGroup_lo_1739 = {dataGroup_lo_hi_1739, dataGroup_lo_lo_1739};
  wire [1023:0] dataGroup_hi_1739 = {dataGroup_hi_hi_1739, dataGroup_hi_lo_1739};
  wire [31:0]   dataGroup_3_73 = dataGroup_lo_1739[223:192];
  wire [1023:0] dataGroup_lo_1740 = {dataGroup_lo_hi_1740, dataGroup_lo_lo_1740};
  wire [1023:0] dataGroup_hi_1740 = {dataGroup_hi_hi_1740, dataGroup_hi_lo_1740};
  wire [31:0]   dataGroup_4_73 = dataGroup_lo_1740[287:256];
  wire [1023:0] dataGroup_lo_1741 = {dataGroup_lo_hi_1741, dataGroup_lo_lo_1741};
  wire [1023:0] dataGroup_hi_1741 = {dataGroup_hi_hi_1741, dataGroup_hi_lo_1741};
  wire [31:0]   dataGroup_5_73 = dataGroup_lo_1741[351:320];
  wire [1023:0] dataGroup_lo_1742 = {dataGroup_lo_hi_1742, dataGroup_lo_lo_1742};
  wire [1023:0] dataGroup_hi_1742 = {dataGroup_hi_hi_1742, dataGroup_hi_lo_1742};
  wire [31:0]   dataGroup_6_73 = dataGroup_lo_1742[415:384];
  wire [1023:0] dataGroup_lo_1743 = {dataGroup_lo_hi_1743, dataGroup_lo_lo_1743};
  wire [1023:0] dataGroup_hi_1743 = {dataGroup_hi_hi_1743, dataGroup_hi_lo_1743};
  wire [31:0]   dataGroup_7_73 = dataGroup_lo_1743[479:448];
  wire [63:0]   res_lo_lo_73 = {dataGroup_1_73, dataGroup_0_73};
  wire [63:0]   res_lo_hi_73 = {dataGroup_3_73, dataGroup_2_73};
  wire [127:0]  res_lo_73 = {res_lo_hi_73, res_lo_lo_73};
  wire [63:0]   res_hi_lo_73 = {dataGroup_5_73, dataGroup_4_73};
  wire [63:0]   res_hi_hi_73 = {dataGroup_7_73, dataGroup_6_73};
  wire [127:0]  res_hi_73 = {res_hi_hi_73, res_hi_lo_73};
  wire [255:0]  res_136 = {res_hi_73, res_lo_73};
  wire [1023:0] dataGroup_lo_1744 = {dataGroup_lo_hi_1744, dataGroup_lo_lo_1744};
  wire [1023:0] dataGroup_hi_1744 = {dataGroup_hi_hi_1744, dataGroup_hi_lo_1744};
  wire [31:0]   dataGroup_0_74 = dataGroup_lo_1744[63:32];
  wire [1023:0] dataGroup_lo_1745 = {dataGroup_lo_hi_1745, dataGroup_lo_lo_1745};
  wire [1023:0] dataGroup_hi_1745 = {dataGroup_hi_hi_1745, dataGroup_hi_lo_1745};
  wire [31:0]   dataGroup_1_74 = dataGroup_lo_1745[127:96];
  wire [1023:0] dataGroup_lo_1746 = {dataGroup_lo_hi_1746, dataGroup_lo_lo_1746};
  wire [1023:0] dataGroup_hi_1746 = {dataGroup_hi_hi_1746, dataGroup_hi_lo_1746};
  wire [31:0]   dataGroup_2_74 = dataGroup_lo_1746[191:160];
  wire [1023:0] dataGroup_lo_1747 = {dataGroup_lo_hi_1747, dataGroup_lo_lo_1747};
  wire [1023:0] dataGroup_hi_1747 = {dataGroup_hi_hi_1747, dataGroup_hi_lo_1747};
  wire [31:0]   dataGroup_3_74 = dataGroup_lo_1747[255:224];
  wire [1023:0] dataGroup_lo_1748 = {dataGroup_lo_hi_1748, dataGroup_lo_lo_1748};
  wire [1023:0] dataGroup_hi_1748 = {dataGroup_hi_hi_1748, dataGroup_hi_lo_1748};
  wire [31:0]   dataGroup_4_74 = dataGroup_lo_1748[319:288];
  wire [1023:0] dataGroup_lo_1749 = {dataGroup_lo_hi_1749, dataGroup_lo_lo_1749};
  wire [1023:0] dataGroup_hi_1749 = {dataGroup_hi_hi_1749, dataGroup_hi_lo_1749};
  wire [31:0]   dataGroup_5_74 = dataGroup_lo_1749[383:352];
  wire [1023:0] dataGroup_lo_1750 = {dataGroup_lo_hi_1750, dataGroup_lo_lo_1750};
  wire [1023:0] dataGroup_hi_1750 = {dataGroup_hi_hi_1750, dataGroup_hi_lo_1750};
  wire [31:0]   dataGroup_6_74 = dataGroup_lo_1750[447:416];
  wire [1023:0] dataGroup_lo_1751 = {dataGroup_lo_hi_1751, dataGroup_lo_lo_1751};
  wire [1023:0] dataGroup_hi_1751 = {dataGroup_hi_hi_1751, dataGroup_hi_lo_1751};
  wire [31:0]   dataGroup_7_74 = dataGroup_lo_1751[511:480];
  wire [63:0]   res_lo_lo_74 = {dataGroup_1_74, dataGroup_0_74};
  wire [63:0]   res_lo_hi_74 = {dataGroup_3_74, dataGroup_2_74};
  wire [127:0]  res_lo_74 = {res_lo_hi_74, res_lo_lo_74};
  wire [63:0]   res_hi_lo_74 = {dataGroup_5_74, dataGroup_4_74};
  wire [63:0]   res_hi_hi_74 = {dataGroup_7_74, dataGroup_6_74};
  wire [127:0]  res_hi_74 = {res_hi_hi_74, res_hi_lo_74};
  wire [255:0]  res_137 = {res_hi_74, res_lo_74};
  wire [511:0]  lo_lo_17 = {res_137, res_136};
  wire [1023:0] lo_17 = {512'h0, lo_lo_17};
  wire [2047:0] regroupLoadData_2_1 = {1024'h0, lo_17};
  wire [1023:0] dataGroup_lo_1752 = {dataGroup_lo_hi_1752, dataGroup_lo_lo_1752};
  wire [1023:0] dataGroup_hi_1752 = {dataGroup_hi_hi_1752, dataGroup_hi_lo_1752};
  wire [31:0]   dataGroup_0_75 = dataGroup_lo_1752[31:0];
  wire [1023:0] dataGroup_lo_1753 = {dataGroup_lo_hi_1753, dataGroup_lo_lo_1753};
  wire [1023:0] dataGroup_hi_1753 = {dataGroup_hi_hi_1753, dataGroup_hi_lo_1753};
  wire [31:0]   dataGroup_1_75 = dataGroup_lo_1753[127:96];
  wire [1023:0] dataGroup_lo_1754 = {dataGroup_lo_hi_1754, dataGroup_lo_lo_1754};
  wire [1023:0] dataGroup_hi_1754 = {dataGroup_hi_hi_1754, dataGroup_hi_lo_1754};
  wire [31:0]   dataGroup_2_75 = dataGroup_lo_1754[223:192];
  wire [1023:0] dataGroup_lo_1755 = {dataGroup_lo_hi_1755, dataGroup_lo_lo_1755};
  wire [1023:0] dataGroup_hi_1755 = {dataGroup_hi_hi_1755, dataGroup_hi_lo_1755};
  wire [31:0]   dataGroup_3_75 = dataGroup_lo_1755[319:288];
  wire [1023:0] dataGroup_lo_1756 = {dataGroup_lo_hi_1756, dataGroup_lo_lo_1756};
  wire [1023:0] dataGroup_hi_1756 = {dataGroup_hi_hi_1756, dataGroup_hi_lo_1756};
  wire [31:0]   dataGroup_4_75 = dataGroup_lo_1756[415:384];
  wire [1023:0] dataGroup_lo_1757 = {dataGroup_lo_hi_1757, dataGroup_lo_lo_1757};
  wire [1023:0] dataGroup_hi_1757 = {dataGroup_hi_hi_1757, dataGroup_hi_lo_1757};
  wire [31:0]   dataGroup_5_75 = dataGroup_lo_1757[511:480];
  wire [1023:0] dataGroup_lo_1758 = {dataGroup_lo_hi_1758, dataGroup_lo_lo_1758};
  wire [1023:0] dataGroup_hi_1758 = {dataGroup_hi_hi_1758, dataGroup_hi_lo_1758};
  wire [31:0]   dataGroup_6_75 = dataGroup_lo_1758[607:576];
  wire [1023:0] dataGroup_lo_1759 = {dataGroup_lo_hi_1759, dataGroup_lo_lo_1759};
  wire [1023:0] dataGroup_hi_1759 = {dataGroup_hi_hi_1759, dataGroup_hi_lo_1759};
  wire [31:0]   dataGroup_7_75 = dataGroup_lo_1759[703:672];
  wire [63:0]   res_lo_lo_75 = {dataGroup_1_75, dataGroup_0_75};
  wire [63:0]   res_lo_hi_75 = {dataGroup_3_75, dataGroup_2_75};
  wire [127:0]  res_lo_75 = {res_lo_hi_75, res_lo_lo_75};
  wire [63:0]   res_hi_lo_75 = {dataGroup_5_75, dataGroup_4_75};
  wire [63:0]   res_hi_hi_75 = {dataGroup_7_75, dataGroup_6_75};
  wire [127:0]  res_hi_75 = {res_hi_hi_75, res_hi_lo_75};
  wire [255:0]  res_144 = {res_hi_75, res_lo_75};
  wire [1023:0] dataGroup_lo_1760 = {dataGroup_lo_hi_1760, dataGroup_lo_lo_1760};
  wire [1023:0] dataGroup_hi_1760 = {dataGroup_hi_hi_1760, dataGroup_hi_lo_1760};
  wire [31:0]   dataGroup_0_76 = dataGroup_lo_1760[63:32];
  wire [1023:0] dataGroup_lo_1761 = {dataGroup_lo_hi_1761, dataGroup_lo_lo_1761};
  wire [1023:0] dataGroup_hi_1761 = {dataGroup_hi_hi_1761, dataGroup_hi_lo_1761};
  wire [31:0]   dataGroup_1_76 = dataGroup_lo_1761[159:128];
  wire [1023:0] dataGroup_lo_1762 = {dataGroup_lo_hi_1762, dataGroup_lo_lo_1762};
  wire [1023:0] dataGroup_hi_1762 = {dataGroup_hi_hi_1762, dataGroup_hi_lo_1762};
  wire [31:0]   dataGroup_2_76 = dataGroup_lo_1762[255:224];
  wire [1023:0] dataGroup_lo_1763 = {dataGroup_lo_hi_1763, dataGroup_lo_lo_1763};
  wire [1023:0] dataGroup_hi_1763 = {dataGroup_hi_hi_1763, dataGroup_hi_lo_1763};
  wire [31:0]   dataGroup_3_76 = dataGroup_lo_1763[351:320];
  wire [1023:0] dataGroup_lo_1764 = {dataGroup_lo_hi_1764, dataGroup_lo_lo_1764};
  wire [1023:0] dataGroup_hi_1764 = {dataGroup_hi_hi_1764, dataGroup_hi_lo_1764};
  wire [31:0]   dataGroup_4_76 = dataGroup_lo_1764[447:416];
  wire [1023:0] dataGroup_lo_1765 = {dataGroup_lo_hi_1765, dataGroup_lo_lo_1765};
  wire [1023:0] dataGroup_hi_1765 = {dataGroup_hi_hi_1765, dataGroup_hi_lo_1765};
  wire [31:0]   dataGroup_5_76 = dataGroup_lo_1765[543:512];
  wire [1023:0] dataGroup_lo_1766 = {dataGroup_lo_hi_1766, dataGroup_lo_lo_1766};
  wire [1023:0] dataGroup_hi_1766 = {dataGroup_hi_hi_1766, dataGroup_hi_lo_1766};
  wire [31:0]   dataGroup_6_76 = dataGroup_lo_1766[639:608];
  wire [1023:0] dataGroup_lo_1767 = {dataGroup_lo_hi_1767, dataGroup_lo_lo_1767};
  wire [1023:0] dataGroup_hi_1767 = {dataGroup_hi_hi_1767, dataGroup_hi_lo_1767};
  wire [31:0]   dataGroup_7_76 = dataGroup_lo_1767[735:704];
  wire [63:0]   res_lo_lo_76 = {dataGroup_1_76, dataGroup_0_76};
  wire [63:0]   res_lo_hi_76 = {dataGroup_3_76, dataGroup_2_76};
  wire [127:0]  res_lo_76 = {res_lo_hi_76, res_lo_lo_76};
  wire [63:0]   res_hi_lo_76 = {dataGroup_5_76, dataGroup_4_76};
  wire [63:0]   res_hi_hi_76 = {dataGroup_7_76, dataGroup_6_76};
  wire [127:0]  res_hi_76 = {res_hi_hi_76, res_hi_lo_76};
  wire [255:0]  res_145 = {res_hi_76, res_lo_76};
  wire [1023:0] dataGroup_lo_1768 = {dataGroup_lo_hi_1768, dataGroup_lo_lo_1768};
  wire [1023:0] dataGroup_hi_1768 = {dataGroup_hi_hi_1768, dataGroup_hi_lo_1768};
  wire [31:0]   dataGroup_0_77 = dataGroup_lo_1768[95:64];
  wire [1023:0] dataGroup_lo_1769 = {dataGroup_lo_hi_1769, dataGroup_lo_lo_1769};
  wire [1023:0] dataGroup_hi_1769 = {dataGroup_hi_hi_1769, dataGroup_hi_lo_1769};
  wire [31:0]   dataGroup_1_77 = dataGroup_lo_1769[191:160];
  wire [1023:0] dataGroup_lo_1770 = {dataGroup_lo_hi_1770, dataGroup_lo_lo_1770};
  wire [1023:0] dataGroup_hi_1770 = {dataGroup_hi_hi_1770, dataGroup_hi_lo_1770};
  wire [31:0]   dataGroup_2_77 = dataGroup_lo_1770[287:256];
  wire [1023:0] dataGroup_lo_1771 = {dataGroup_lo_hi_1771, dataGroup_lo_lo_1771};
  wire [1023:0] dataGroup_hi_1771 = {dataGroup_hi_hi_1771, dataGroup_hi_lo_1771};
  wire [31:0]   dataGroup_3_77 = dataGroup_lo_1771[383:352];
  wire [1023:0] dataGroup_lo_1772 = {dataGroup_lo_hi_1772, dataGroup_lo_lo_1772};
  wire [1023:0] dataGroup_hi_1772 = {dataGroup_hi_hi_1772, dataGroup_hi_lo_1772};
  wire [31:0]   dataGroup_4_77 = dataGroup_lo_1772[479:448];
  wire [1023:0] dataGroup_lo_1773 = {dataGroup_lo_hi_1773, dataGroup_lo_lo_1773};
  wire [1023:0] dataGroup_hi_1773 = {dataGroup_hi_hi_1773, dataGroup_hi_lo_1773};
  wire [31:0]   dataGroup_5_77 = dataGroup_lo_1773[575:544];
  wire [1023:0] dataGroup_lo_1774 = {dataGroup_lo_hi_1774, dataGroup_lo_lo_1774};
  wire [1023:0] dataGroup_hi_1774 = {dataGroup_hi_hi_1774, dataGroup_hi_lo_1774};
  wire [31:0]   dataGroup_6_77 = dataGroup_lo_1774[671:640];
  wire [1023:0] dataGroup_lo_1775 = {dataGroup_lo_hi_1775, dataGroup_lo_lo_1775};
  wire [1023:0] dataGroup_hi_1775 = {dataGroup_hi_hi_1775, dataGroup_hi_lo_1775};
  wire [31:0]   dataGroup_7_77 = dataGroup_lo_1775[767:736];
  wire [63:0]   res_lo_lo_77 = {dataGroup_1_77, dataGroup_0_77};
  wire [63:0]   res_lo_hi_77 = {dataGroup_3_77, dataGroup_2_77};
  wire [127:0]  res_lo_77 = {res_lo_hi_77, res_lo_lo_77};
  wire [63:0]   res_hi_lo_77 = {dataGroup_5_77, dataGroup_4_77};
  wire [63:0]   res_hi_hi_77 = {dataGroup_7_77, dataGroup_6_77};
  wire [127:0]  res_hi_77 = {res_hi_hi_77, res_hi_lo_77};
  wire [255:0]  res_146 = {res_hi_77, res_lo_77};
  wire [511:0]  lo_lo_18 = {res_145, res_144};
  wire [511:0]  lo_hi_18 = {256'h0, res_146};
  wire [1023:0] lo_18 = {lo_hi_18, lo_lo_18};
  wire [2047:0] regroupLoadData_2_2 = {1024'h0, lo_18};
  wire [1023:0] dataGroup_lo_1776 = {dataGroup_lo_hi_1776, dataGroup_lo_lo_1776};
  wire [1023:0] dataGroup_hi_1776 = {dataGroup_hi_hi_1776, dataGroup_hi_lo_1776};
  wire [31:0]   dataGroup_0_78 = dataGroup_lo_1776[31:0];
  wire [1023:0] dataGroup_lo_1777 = {dataGroup_lo_hi_1777, dataGroup_lo_lo_1777};
  wire [1023:0] dataGroup_hi_1777 = {dataGroup_hi_hi_1777, dataGroup_hi_lo_1777};
  wire [31:0]   dataGroup_1_78 = dataGroup_lo_1777[159:128];
  wire [1023:0] dataGroup_lo_1778 = {dataGroup_lo_hi_1778, dataGroup_lo_lo_1778};
  wire [1023:0] dataGroup_hi_1778 = {dataGroup_hi_hi_1778, dataGroup_hi_lo_1778};
  wire [31:0]   dataGroup_2_78 = dataGroup_lo_1778[287:256];
  wire [1023:0] dataGroup_lo_1779 = {dataGroup_lo_hi_1779, dataGroup_lo_lo_1779};
  wire [1023:0] dataGroup_hi_1779 = {dataGroup_hi_hi_1779, dataGroup_hi_lo_1779};
  wire [31:0]   dataGroup_3_78 = dataGroup_lo_1779[415:384];
  wire [1023:0] dataGroup_lo_1780 = {dataGroup_lo_hi_1780, dataGroup_lo_lo_1780};
  wire [1023:0] dataGroup_hi_1780 = {dataGroup_hi_hi_1780, dataGroup_hi_lo_1780};
  wire [31:0]   dataGroup_4_78 = dataGroup_lo_1780[543:512];
  wire [1023:0] dataGroup_lo_1781 = {dataGroup_lo_hi_1781, dataGroup_lo_lo_1781};
  wire [1023:0] dataGroup_hi_1781 = {dataGroup_hi_hi_1781, dataGroup_hi_lo_1781};
  wire [31:0]   dataGroup_5_78 = dataGroup_lo_1781[671:640];
  wire [1023:0] dataGroup_lo_1782 = {dataGroup_lo_hi_1782, dataGroup_lo_lo_1782};
  wire [1023:0] dataGroup_hi_1782 = {dataGroup_hi_hi_1782, dataGroup_hi_lo_1782};
  wire [31:0]   dataGroup_6_78 = dataGroup_lo_1782[799:768];
  wire [1023:0] dataGroup_lo_1783 = {dataGroup_lo_hi_1783, dataGroup_lo_lo_1783};
  wire [1023:0] dataGroup_hi_1783 = {dataGroup_hi_hi_1783, dataGroup_hi_lo_1783};
  wire [31:0]   dataGroup_7_78 = dataGroup_lo_1783[927:896];
  wire [63:0]   res_lo_lo_78 = {dataGroup_1_78, dataGroup_0_78};
  wire [63:0]   res_lo_hi_78 = {dataGroup_3_78, dataGroup_2_78};
  wire [127:0]  res_lo_78 = {res_lo_hi_78, res_lo_lo_78};
  wire [63:0]   res_hi_lo_78 = {dataGroup_5_78, dataGroup_4_78};
  wire [63:0]   res_hi_hi_78 = {dataGroup_7_78, dataGroup_6_78};
  wire [127:0]  res_hi_78 = {res_hi_hi_78, res_hi_lo_78};
  wire [255:0]  res_152 = {res_hi_78, res_lo_78};
  wire [1023:0] dataGroup_lo_1784 = {dataGroup_lo_hi_1784, dataGroup_lo_lo_1784};
  wire [1023:0] dataGroup_hi_1784 = {dataGroup_hi_hi_1784, dataGroup_hi_lo_1784};
  wire [31:0]   dataGroup_0_79 = dataGroup_lo_1784[63:32];
  wire [1023:0] dataGroup_lo_1785 = {dataGroup_lo_hi_1785, dataGroup_lo_lo_1785};
  wire [1023:0] dataGroup_hi_1785 = {dataGroup_hi_hi_1785, dataGroup_hi_lo_1785};
  wire [31:0]   dataGroup_1_79 = dataGroup_lo_1785[191:160];
  wire [1023:0] dataGroup_lo_1786 = {dataGroup_lo_hi_1786, dataGroup_lo_lo_1786};
  wire [1023:0] dataGroup_hi_1786 = {dataGroup_hi_hi_1786, dataGroup_hi_lo_1786};
  wire [31:0]   dataGroup_2_79 = dataGroup_lo_1786[319:288];
  wire [1023:0] dataGroup_lo_1787 = {dataGroup_lo_hi_1787, dataGroup_lo_lo_1787};
  wire [1023:0] dataGroup_hi_1787 = {dataGroup_hi_hi_1787, dataGroup_hi_lo_1787};
  wire [31:0]   dataGroup_3_79 = dataGroup_lo_1787[447:416];
  wire [1023:0] dataGroup_lo_1788 = {dataGroup_lo_hi_1788, dataGroup_lo_lo_1788};
  wire [1023:0] dataGroup_hi_1788 = {dataGroup_hi_hi_1788, dataGroup_hi_lo_1788};
  wire [31:0]   dataGroup_4_79 = dataGroup_lo_1788[575:544];
  wire [1023:0] dataGroup_lo_1789 = {dataGroup_lo_hi_1789, dataGroup_lo_lo_1789};
  wire [1023:0] dataGroup_hi_1789 = {dataGroup_hi_hi_1789, dataGroup_hi_lo_1789};
  wire [31:0]   dataGroup_5_79 = dataGroup_lo_1789[703:672];
  wire [1023:0] dataGroup_lo_1790 = {dataGroup_lo_hi_1790, dataGroup_lo_lo_1790};
  wire [1023:0] dataGroup_hi_1790 = {dataGroup_hi_hi_1790, dataGroup_hi_lo_1790};
  wire [31:0]   dataGroup_6_79 = dataGroup_lo_1790[831:800];
  wire [1023:0] dataGroup_lo_1791 = {dataGroup_lo_hi_1791, dataGroup_lo_lo_1791};
  wire [1023:0] dataGroup_hi_1791 = {dataGroup_hi_hi_1791, dataGroup_hi_lo_1791};
  wire [31:0]   dataGroup_7_79 = dataGroup_lo_1791[959:928];
  wire [63:0]   res_lo_lo_79 = {dataGroup_1_79, dataGroup_0_79};
  wire [63:0]   res_lo_hi_79 = {dataGroup_3_79, dataGroup_2_79};
  wire [127:0]  res_lo_79 = {res_lo_hi_79, res_lo_lo_79};
  wire [63:0]   res_hi_lo_79 = {dataGroup_5_79, dataGroup_4_79};
  wire [63:0]   res_hi_hi_79 = {dataGroup_7_79, dataGroup_6_79};
  wire [127:0]  res_hi_79 = {res_hi_hi_79, res_hi_lo_79};
  wire [255:0]  res_153 = {res_hi_79, res_lo_79};
  wire [1023:0] dataGroup_lo_1792 = {dataGroup_lo_hi_1792, dataGroup_lo_lo_1792};
  wire [1023:0] dataGroup_hi_1792 = {dataGroup_hi_hi_1792, dataGroup_hi_lo_1792};
  wire [31:0]   dataGroup_0_80 = dataGroup_lo_1792[95:64];
  wire [1023:0] dataGroup_lo_1793 = {dataGroup_lo_hi_1793, dataGroup_lo_lo_1793};
  wire [1023:0] dataGroup_hi_1793 = {dataGroup_hi_hi_1793, dataGroup_hi_lo_1793};
  wire [31:0]   dataGroup_1_80 = dataGroup_lo_1793[223:192];
  wire [1023:0] dataGroup_lo_1794 = {dataGroup_lo_hi_1794, dataGroup_lo_lo_1794};
  wire [1023:0] dataGroup_hi_1794 = {dataGroup_hi_hi_1794, dataGroup_hi_lo_1794};
  wire [31:0]   dataGroup_2_80 = dataGroup_lo_1794[351:320];
  wire [1023:0] dataGroup_lo_1795 = {dataGroup_lo_hi_1795, dataGroup_lo_lo_1795};
  wire [1023:0] dataGroup_hi_1795 = {dataGroup_hi_hi_1795, dataGroup_hi_lo_1795};
  wire [31:0]   dataGroup_3_80 = dataGroup_lo_1795[479:448];
  wire [1023:0] dataGroup_lo_1796 = {dataGroup_lo_hi_1796, dataGroup_lo_lo_1796};
  wire [1023:0] dataGroup_hi_1796 = {dataGroup_hi_hi_1796, dataGroup_hi_lo_1796};
  wire [31:0]   dataGroup_4_80 = dataGroup_lo_1796[607:576];
  wire [1023:0] dataGroup_lo_1797 = {dataGroup_lo_hi_1797, dataGroup_lo_lo_1797};
  wire [1023:0] dataGroup_hi_1797 = {dataGroup_hi_hi_1797, dataGroup_hi_lo_1797};
  wire [31:0]   dataGroup_5_80 = dataGroup_lo_1797[735:704];
  wire [1023:0] dataGroup_lo_1798 = {dataGroup_lo_hi_1798, dataGroup_lo_lo_1798};
  wire [1023:0] dataGroup_hi_1798 = {dataGroup_hi_hi_1798, dataGroup_hi_lo_1798};
  wire [31:0]   dataGroup_6_80 = dataGroup_lo_1798[863:832];
  wire [1023:0] dataGroup_lo_1799 = {dataGroup_lo_hi_1799, dataGroup_lo_lo_1799};
  wire [1023:0] dataGroup_hi_1799 = {dataGroup_hi_hi_1799, dataGroup_hi_lo_1799};
  wire [31:0]   dataGroup_7_80 = dataGroup_lo_1799[991:960];
  wire [63:0]   res_lo_lo_80 = {dataGroup_1_80, dataGroup_0_80};
  wire [63:0]   res_lo_hi_80 = {dataGroup_3_80, dataGroup_2_80};
  wire [127:0]  res_lo_80 = {res_lo_hi_80, res_lo_lo_80};
  wire [63:0]   res_hi_lo_80 = {dataGroup_5_80, dataGroup_4_80};
  wire [63:0]   res_hi_hi_80 = {dataGroup_7_80, dataGroup_6_80};
  wire [127:0]  res_hi_80 = {res_hi_hi_80, res_hi_lo_80};
  wire [255:0]  res_154 = {res_hi_80, res_lo_80};
  wire [1023:0] dataGroup_lo_1800 = {dataGroup_lo_hi_1800, dataGroup_lo_lo_1800};
  wire [1023:0] dataGroup_hi_1800 = {dataGroup_hi_hi_1800, dataGroup_hi_lo_1800};
  wire [31:0]   dataGroup_0_81 = dataGroup_lo_1800[127:96];
  wire [1023:0] dataGroup_lo_1801 = {dataGroup_lo_hi_1801, dataGroup_lo_lo_1801};
  wire [1023:0] dataGroup_hi_1801 = {dataGroup_hi_hi_1801, dataGroup_hi_lo_1801};
  wire [31:0]   dataGroup_1_81 = dataGroup_lo_1801[255:224];
  wire [1023:0] dataGroup_lo_1802 = {dataGroup_lo_hi_1802, dataGroup_lo_lo_1802};
  wire [1023:0] dataGroup_hi_1802 = {dataGroup_hi_hi_1802, dataGroup_hi_lo_1802};
  wire [31:0]   dataGroup_2_81 = dataGroup_lo_1802[383:352];
  wire [1023:0] dataGroup_lo_1803 = {dataGroup_lo_hi_1803, dataGroup_lo_lo_1803};
  wire [1023:0] dataGroup_hi_1803 = {dataGroup_hi_hi_1803, dataGroup_hi_lo_1803};
  wire [31:0]   dataGroup_3_81 = dataGroup_lo_1803[511:480];
  wire [1023:0] dataGroup_lo_1804 = {dataGroup_lo_hi_1804, dataGroup_lo_lo_1804};
  wire [1023:0] dataGroup_hi_1804 = {dataGroup_hi_hi_1804, dataGroup_hi_lo_1804};
  wire [31:0]   dataGroup_4_81 = dataGroup_lo_1804[639:608];
  wire [1023:0] dataGroup_lo_1805 = {dataGroup_lo_hi_1805, dataGroup_lo_lo_1805};
  wire [1023:0] dataGroup_hi_1805 = {dataGroup_hi_hi_1805, dataGroup_hi_lo_1805};
  wire [31:0]   dataGroup_5_81 = dataGroup_lo_1805[767:736];
  wire [1023:0] dataGroup_lo_1806 = {dataGroup_lo_hi_1806, dataGroup_lo_lo_1806};
  wire [1023:0] dataGroup_hi_1806 = {dataGroup_hi_hi_1806, dataGroup_hi_lo_1806};
  wire [31:0]   dataGroup_6_81 = dataGroup_lo_1806[895:864];
  wire [1023:0] dataGroup_lo_1807 = {dataGroup_lo_hi_1807, dataGroup_lo_lo_1807};
  wire [1023:0] dataGroup_hi_1807 = {dataGroup_hi_hi_1807, dataGroup_hi_lo_1807};
  wire [31:0]   dataGroup_7_81 = dataGroup_lo_1807[1023:992];
  wire [63:0]   res_lo_lo_81 = {dataGroup_1_81, dataGroup_0_81};
  wire [63:0]   res_lo_hi_81 = {dataGroup_3_81, dataGroup_2_81};
  wire [127:0]  res_lo_81 = {res_lo_hi_81, res_lo_lo_81};
  wire [63:0]   res_hi_lo_81 = {dataGroup_5_81, dataGroup_4_81};
  wire [63:0]   res_hi_hi_81 = {dataGroup_7_81, dataGroup_6_81};
  wire [127:0]  res_hi_81 = {res_hi_hi_81, res_hi_lo_81};
  wire [255:0]  res_155 = {res_hi_81, res_lo_81};
  wire [511:0]  lo_lo_19 = {res_153, res_152};
  wire [511:0]  lo_hi_19 = {res_155, res_154};
  wire [1023:0] lo_19 = {lo_hi_19, lo_lo_19};
  wire [2047:0] regroupLoadData_2_3 = {1024'h0, lo_19};
  wire [1023:0] dataGroup_lo_1808 = {dataGroup_lo_hi_1808, dataGroup_lo_lo_1808};
  wire [1023:0] dataGroup_hi_1808 = {dataGroup_hi_hi_1808, dataGroup_hi_lo_1808};
  wire [31:0]   dataGroup_0_82 = dataGroup_lo_1808[31:0];
  wire [1023:0] dataGroup_lo_1809 = {dataGroup_lo_hi_1809, dataGroup_lo_lo_1809};
  wire [1023:0] dataGroup_hi_1809 = {dataGroup_hi_hi_1809, dataGroup_hi_lo_1809};
  wire [31:0]   dataGroup_1_82 = dataGroup_lo_1809[191:160];
  wire [1023:0] dataGroup_lo_1810 = {dataGroup_lo_hi_1810, dataGroup_lo_lo_1810};
  wire [1023:0] dataGroup_hi_1810 = {dataGroup_hi_hi_1810, dataGroup_hi_lo_1810};
  wire [31:0]   dataGroup_2_82 = dataGroup_lo_1810[351:320];
  wire [1023:0] dataGroup_lo_1811 = {dataGroup_lo_hi_1811, dataGroup_lo_lo_1811};
  wire [1023:0] dataGroup_hi_1811 = {dataGroup_hi_hi_1811, dataGroup_hi_lo_1811};
  wire [31:0]   dataGroup_3_82 = dataGroup_lo_1811[511:480];
  wire [1023:0] dataGroup_lo_1812 = {dataGroup_lo_hi_1812, dataGroup_lo_lo_1812};
  wire [1023:0] dataGroup_hi_1812 = {dataGroup_hi_hi_1812, dataGroup_hi_lo_1812};
  wire [31:0]   dataGroup_4_82 = dataGroup_lo_1812[671:640];
  wire [1023:0] dataGroup_lo_1813 = {dataGroup_lo_hi_1813, dataGroup_lo_lo_1813};
  wire [1023:0] dataGroup_hi_1813 = {dataGroup_hi_hi_1813, dataGroup_hi_lo_1813};
  wire [31:0]   dataGroup_5_82 = dataGroup_lo_1813[831:800];
  wire [1023:0] dataGroup_lo_1814 = {dataGroup_lo_hi_1814, dataGroup_lo_lo_1814};
  wire [1023:0] dataGroup_hi_1814 = {dataGroup_hi_hi_1814, dataGroup_hi_lo_1814};
  wire [31:0]   dataGroup_6_82 = dataGroup_lo_1814[991:960];
  wire [1023:0] dataGroup_lo_1815 = {dataGroup_lo_hi_1815, dataGroup_lo_lo_1815};
  wire [1023:0] dataGroup_hi_1815 = {dataGroup_hi_hi_1815, dataGroup_hi_lo_1815};
  wire [31:0]   dataGroup_7_82 = dataGroup_hi_1815[127:96];
  wire [63:0]   res_lo_lo_82 = {dataGroup_1_82, dataGroup_0_82};
  wire [63:0]   res_lo_hi_82 = {dataGroup_3_82, dataGroup_2_82};
  wire [127:0]  res_lo_82 = {res_lo_hi_82, res_lo_lo_82};
  wire [63:0]   res_hi_lo_82 = {dataGroup_5_82, dataGroup_4_82};
  wire [63:0]   res_hi_hi_82 = {dataGroup_7_82, dataGroup_6_82};
  wire [127:0]  res_hi_82 = {res_hi_hi_82, res_hi_lo_82};
  wire [255:0]  res_160 = {res_hi_82, res_lo_82};
  wire [1023:0] dataGroup_lo_1816 = {dataGroup_lo_hi_1816, dataGroup_lo_lo_1816};
  wire [1023:0] dataGroup_hi_1816 = {dataGroup_hi_hi_1816, dataGroup_hi_lo_1816};
  wire [31:0]   dataGroup_0_83 = dataGroup_lo_1816[63:32];
  wire [1023:0] dataGroup_lo_1817 = {dataGroup_lo_hi_1817, dataGroup_lo_lo_1817};
  wire [1023:0] dataGroup_hi_1817 = {dataGroup_hi_hi_1817, dataGroup_hi_lo_1817};
  wire [31:0]   dataGroup_1_83 = dataGroup_lo_1817[223:192];
  wire [1023:0] dataGroup_lo_1818 = {dataGroup_lo_hi_1818, dataGroup_lo_lo_1818};
  wire [1023:0] dataGroup_hi_1818 = {dataGroup_hi_hi_1818, dataGroup_hi_lo_1818};
  wire [31:0]   dataGroup_2_83 = dataGroup_lo_1818[383:352];
  wire [1023:0] dataGroup_lo_1819 = {dataGroup_lo_hi_1819, dataGroup_lo_lo_1819};
  wire [1023:0] dataGroup_hi_1819 = {dataGroup_hi_hi_1819, dataGroup_hi_lo_1819};
  wire [31:0]   dataGroup_3_83 = dataGroup_lo_1819[543:512];
  wire [1023:0] dataGroup_lo_1820 = {dataGroup_lo_hi_1820, dataGroup_lo_lo_1820};
  wire [1023:0] dataGroup_hi_1820 = {dataGroup_hi_hi_1820, dataGroup_hi_lo_1820};
  wire [31:0]   dataGroup_4_83 = dataGroup_lo_1820[703:672];
  wire [1023:0] dataGroup_lo_1821 = {dataGroup_lo_hi_1821, dataGroup_lo_lo_1821};
  wire [1023:0] dataGroup_hi_1821 = {dataGroup_hi_hi_1821, dataGroup_hi_lo_1821};
  wire [31:0]   dataGroup_5_83 = dataGroup_lo_1821[863:832];
  wire [1023:0] dataGroup_lo_1822 = {dataGroup_lo_hi_1822, dataGroup_lo_lo_1822};
  wire [1023:0] dataGroup_hi_1822 = {dataGroup_hi_hi_1822, dataGroup_hi_lo_1822};
  wire [31:0]   dataGroup_6_83 = dataGroup_lo_1822[1023:992];
  wire [1023:0] dataGroup_lo_1823 = {dataGroup_lo_hi_1823, dataGroup_lo_lo_1823};
  wire [1023:0] dataGroup_hi_1823 = {dataGroup_hi_hi_1823, dataGroup_hi_lo_1823};
  wire [31:0]   dataGroup_7_83 = dataGroup_hi_1823[159:128];
  wire [63:0]   res_lo_lo_83 = {dataGroup_1_83, dataGroup_0_83};
  wire [63:0]   res_lo_hi_83 = {dataGroup_3_83, dataGroup_2_83};
  wire [127:0]  res_lo_83 = {res_lo_hi_83, res_lo_lo_83};
  wire [63:0]   res_hi_lo_83 = {dataGroup_5_83, dataGroup_4_83};
  wire [63:0]   res_hi_hi_83 = {dataGroup_7_83, dataGroup_6_83};
  wire [127:0]  res_hi_83 = {res_hi_hi_83, res_hi_lo_83};
  wire [255:0]  res_161 = {res_hi_83, res_lo_83};
  wire [1023:0] dataGroup_lo_1824 = {dataGroup_lo_hi_1824, dataGroup_lo_lo_1824};
  wire [1023:0] dataGroup_hi_1824 = {dataGroup_hi_hi_1824, dataGroup_hi_lo_1824};
  wire [31:0]   dataGroup_0_84 = dataGroup_lo_1824[95:64];
  wire [1023:0] dataGroup_lo_1825 = {dataGroup_lo_hi_1825, dataGroup_lo_lo_1825};
  wire [1023:0] dataGroup_hi_1825 = {dataGroup_hi_hi_1825, dataGroup_hi_lo_1825};
  wire [31:0]   dataGroup_1_84 = dataGroup_lo_1825[255:224];
  wire [1023:0] dataGroup_lo_1826 = {dataGroup_lo_hi_1826, dataGroup_lo_lo_1826};
  wire [1023:0] dataGroup_hi_1826 = {dataGroup_hi_hi_1826, dataGroup_hi_lo_1826};
  wire [31:0]   dataGroup_2_84 = dataGroup_lo_1826[415:384];
  wire [1023:0] dataGroup_lo_1827 = {dataGroup_lo_hi_1827, dataGroup_lo_lo_1827};
  wire [1023:0] dataGroup_hi_1827 = {dataGroup_hi_hi_1827, dataGroup_hi_lo_1827};
  wire [31:0]   dataGroup_3_84 = dataGroup_lo_1827[575:544];
  wire [1023:0] dataGroup_lo_1828 = {dataGroup_lo_hi_1828, dataGroup_lo_lo_1828};
  wire [1023:0] dataGroup_hi_1828 = {dataGroup_hi_hi_1828, dataGroup_hi_lo_1828};
  wire [31:0]   dataGroup_4_84 = dataGroup_lo_1828[735:704];
  wire [1023:0] dataGroup_lo_1829 = {dataGroup_lo_hi_1829, dataGroup_lo_lo_1829};
  wire [1023:0] dataGroup_hi_1829 = {dataGroup_hi_hi_1829, dataGroup_hi_lo_1829};
  wire [31:0]   dataGroup_5_84 = dataGroup_lo_1829[895:864];
  wire [1023:0] dataGroup_lo_1830 = {dataGroup_lo_hi_1830, dataGroup_lo_lo_1830};
  wire [1023:0] dataGroup_hi_1830 = {dataGroup_hi_hi_1830, dataGroup_hi_lo_1830};
  wire [31:0]   dataGroup_6_84 = dataGroup_hi_1830[31:0];
  wire [1023:0] dataGroup_lo_1831 = {dataGroup_lo_hi_1831, dataGroup_lo_lo_1831};
  wire [1023:0] dataGroup_hi_1831 = {dataGroup_hi_hi_1831, dataGroup_hi_lo_1831};
  wire [31:0]   dataGroup_7_84 = dataGroup_hi_1831[191:160];
  wire [63:0]   res_lo_lo_84 = {dataGroup_1_84, dataGroup_0_84};
  wire [63:0]   res_lo_hi_84 = {dataGroup_3_84, dataGroup_2_84};
  wire [127:0]  res_lo_84 = {res_lo_hi_84, res_lo_lo_84};
  wire [63:0]   res_hi_lo_84 = {dataGroup_5_84, dataGroup_4_84};
  wire [63:0]   res_hi_hi_84 = {dataGroup_7_84, dataGroup_6_84};
  wire [127:0]  res_hi_84 = {res_hi_hi_84, res_hi_lo_84};
  wire [255:0]  res_162 = {res_hi_84, res_lo_84};
  wire [1023:0] dataGroup_lo_1832 = {dataGroup_lo_hi_1832, dataGroup_lo_lo_1832};
  wire [1023:0] dataGroup_hi_1832 = {dataGroup_hi_hi_1832, dataGroup_hi_lo_1832};
  wire [31:0]   dataGroup_0_85 = dataGroup_lo_1832[127:96];
  wire [1023:0] dataGroup_lo_1833 = {dataGroup_lo_hi_1833, dataGroup_lo_lo_1833};
  wire [1023:0] dataGroup_hi_1833 = {dataGroup_hi_hi_1833, dataGroup_hi_lo_1833};
  wire [31:0]   dataGroup_1_85 = dataGroup_lo_1833[287:256];
  wire [1023:0] dataGroup_lo_1834 = {dataGroup_lo_hi_1834, dataGroup_lo_lo_1834};
  wire [1023:0] dataGroup_hi_1834 = {dataGroup_hi_hi_1834, dataGroup_hi_lo_1834};
  wire [31:0]   dataGroup_2_85 = dataGroup_lo_1834[447:416];
  wire [1023:0] dataGroup_lo_1835 = {dataGroup_lo_hi_1835, dataGroup_lo_lo_1835};
  wire [1023:0] dataGroup_hi_1835 = {dataGroup_hi_hi_1835, dataGroup_hi_lo_1835};
  wire [31:0]   dataGroup_3_85 = dataGroup_lo_1835[607:576];
  wire [1023:0] dataGroup_lo_1836 = {dataGroup_lo_hi_1836, dataGroup_lo_lo_1836};
  wire [1023:0] dataGroup_hi_1836 = {dataGroup_hi_hi_1836, dataGroup_hi_lo_1836};
  wire [31:0]   dataGroup_4_85 = dataGroup_lo_1836[767:736];
  wire [1023:0] dataGroup_lo_1837 = {dataGroup_lo_hi_1837, dataGroup_lo_lo_1837};
  wire [1023:0] dataGroup_hi_1837 = {dataGroup_hi_hi_1837, dataGroup_hi_lo_1837};
  wire [31:0]   dataGroup_5_85 = dataGroup_lo_1837[927:896];
  wire [1023:0] dataGroup_lo_1838 = {dataGroup_lo_hi_1838, dataGroup_lo_lo_1838};
  wire [1023:0] dataGroup_hi_1838 = {dataGroup_hi_hi_1838, dataGroup_hi_lo_1838};
  wire [31:0]   dataGroup_6_85 = dataGroup_hi_1838[63:32];
  wire [1023:0] dataGroup_lo_1839 = {dataGroup_lo_hi_1839, dataGroup_lo_lo_1839};
  wire [1023:0] dataGroup_hi_1839 = {dataGroup_hi_hi_1839, dataGroup_hi_lo_1839};
  wire [31:0]   dataGroup_7_85 = dataGroup_hi_1839[223:192];
  wire [63:0]   res_lo_lo_85 = {dataGroup_1_85, dataGroup_0_85};
  wire [63:0]   res_lo_hi_85 = {dataGroup_3_85, dataGroup_2_85};
  wire [127:0]  res_lo_85 = {res_lo_hi_85, res_lo_lo_85};
  wire [63:0]   res_hi_lo_85 = {dataGroup_5_85, dataGroup_4_85};
  wire [63:0]   res_hi_hi_85 = {dataGroup_7_85, dataGroup_6_85};
  wire [127:0]  res_hi_85 = {res_hi_hi_85, res_hi_lo_85};
  wire [255:0]  res_163 = {res_hi_85, res_lo_85};
  wire [1023:0] dataGroup_lo_1840 = {dataGroup_lo_hi_1840, dataGroup_lo_lo_1840};
  wire [1023:0] dataGroup_hi_1840 = {dataGroup_hi_hi_1840, dataGroup_hi_lo_1840};
  wire [31:0]   dataGroup_0_86 = dataGroup_lo_1840[159:128];
  wire [1023:0] dataGroup_lo_1841 = {dataGroup_lo_hi_1841, dataGroup_lo_lo_1841};
  wire [1023:0] dataGroup_hi_1841 = {dataGroup_hi_hi_1841, dataGroup_hi_lo_1841};
  wire [31:0]   dataGroup_1_86 = dataGroup_lo_1841[319:288];
  wire [1023:0] dataGroup_lo_1842 = {dataGroup_lo_hi_1842, dataGroup_lo_lo_1842};
  wire [1023:0] dataGroup_hi_1842 = {dataGroup_hi_hi_1842, dataGroup_hi_lo_1842};
  wire [31:0]   dataGroup_2_86 = dataGroup_lo_1842[479:448];
  wire [1023:0] dataGroup_lo_1843 = {dataGroup_lo_hi_1843, dataGroup_lo_lo_1843};
  wire [1023:0] dataGroup_hi_1843 = {dataGroup_hi_hi_1843, dataGroup_hi_lo_1843};
  wire [31:0]   dataGroup_3_86 = dataGroup_lo_1843[639:608];
  wire [1023:0] dataGroup_lo_1844 = {dataGroup_lo_hi_1844, dataGroup_lo_lo_1844};
  wire [1023:0] dataGroup_hi_1844 = {dataGroup_hi_hi_1844, dataGroup_hi_lo_1844};
  wire [31:0]   dataGroup_4_86 = dataGroup_lo_1844[799:768];
  wire [1023:0] dataGroup_lo_1845 = {dataGroup_lo_hi_1845, dataGroup_lo_lo_1845};
  wire [1023:0] dataGroup_hi_1845 = {dataGroup_hi_hi_1845, dataGroup_hi_lo_1845};
  wire [31:0]   dataGroup_5_86 = dataGroup_lo_1845[959:928];
  wire [1023:0] dataGroup_lo_1846 = {dataGroup_lo_hi_1846, dataGroup_lo_lo_1846};
  wire [1023:0] dataGroup_hi_1846 = {dataGroup_hi_hi_1846, dataGroup_hi_lo_1846};
  wire [31:0]   dataGroup_6_86 = dataGroup_hi_1846[95:64];
  wire [1023:0] dataGroup_lo_1847 = {dataGroup_lo_hi_1847, dataGroup_lo_lo_1847};
  wire [1023:0] dataGroup_hi_1847 = {dataGroup_hi_hi_1847, dataGroup_hi_lo_1847};
  wire [31:0]   dataGroup_7_86 = dataGroup_hi_1847[255:224];
  wire [63:0]   res_lo_lo_86 = {dataGroup_1_86, dataGroup_0_86};
  wire [63:0]   res_lo_hi_86 = {dataGroup_3_86, dataGroup_2_86};
  wire [127:0]  res_lo_86 = {res_lo_hi_86, res_lo_lo_86};
  wire [63:0]   res_hi_lo_86 = {dataGroup_5_86, dataGroup_4_86};
  wire [63:0]   res_hi_hi_86 = {dataGroup_7_86, dataGroup_6_86};
  wire [127:0]  res_hi_86 = {res_hi_hi_86, res_hi_lo_86};
  wire [255:0]  res_164 = {res_hi_86, res_lo_86};
  wire [511:0]  lo_lo_20 = {res_161, res_160};
  wire [511:0]  lo_hi_20 = {res_163, res_162};
  wire [1023:0] lo_20 = {lo_hi_20, lo_lo_20};
  wire [511:0]  hi_lo_20 = {256'h0, res_164};
  wire [1023:0] hi_20 = {512'h0, hi_lo_20};
  wire [2047:0] regroupLoadData_2_4 = {hi_20, lo_20};
  wire [1023:0] dataGroup_lo_1848 = {dataGroup_lo_hi_1848, dataGroup_lo_lo_1848};
  wire [1023:0] dataGroup_hi_1848 = {dataGroup_hi_hi_1848, dataGroup_hi_lo_1848};
  wire [31:0]   dataGroup_0_87 = dataGroup_lo_1848[31:0];
  wire [1023:0] dataGroup_lo_1849 = {dataGroup_lo_hi_1849, dataGroup_lo_lo_1849};
  wire [1023:0] dataGroup_hi_1849 = {dataGroup_hi_hi_1849, dataGroup_hi_lo_1849};
  wire [31:0]   dataGroup_1_87 = dataGroup_lo_1849[223:192];
  wire [1023:0] dataGroup_lo_1850 = {dataGroup_lo_hi_1850, dataGroup_lo_lo_1850};
  wire [1023:0] dataGroup_hi_1850 = {dataGroup_hi_hi_1850, dataGroup_hi_lo_1850};
  wire [31:0]   dataGroup_2_87 = dataGroup_lo_1850[415:384];
  wire [1023:0] dataGroup_lo_1851 = {dataGroup_lo_hi_1851, dataGroup_lo_lo_1851};
  wire [1023:0] dataGroup_hi_1851 = {dataGroup_hi_hi_1851, dataGroup_hi_lo_1851};
  wire [31:0]   dataGroup_3_87 = dataGroup_lo_1851[607:576];
  wire [1023:0] dataGroup_lo_1852 = {dataGroup_lo_hi_1852, dataGroup_lo_lo_1852};
  wire [1023:0] dataGroup_hi_1852 = {dataGroup_hi_hi_1852, dataGroup_hi_lo_1852};
  wire [31:0]   dataGroup_4_87 = dataGroup_lo_1852[799:768];
  wire [1023:0] dataGroup_lo_1853 = {dataGroup_lo_hi_1853, dataGroup_lo_lo_1853};
  wire [1023:0] dataGroup_hi_1853 = {dataGroup_hi_hi_1853, dataGroup_hi_lo_1853};
  wire [31:0]   dataGroup_5_87 = dataGroup_lo_1853[991:960];
  wire [1023:0] dataGroup_lo_1854 = {dataGroup_lo_hi_1854, dataGroup_lo_lo_1854};
  wire [1023:0] dataGroup_hi_1854 = {dataGroup_hi_hi_1854, dataGroup_hi_lo_1854};
  wire [31:0]   dataGroup_6_87 = dataGroup_hi_1854[159:128];
  wire [1023:0] dataGroup_lo_1855 = {dataGroup_lo_hi_1855, dataGroup_lo_lo_1855};
  wire [1023:0] dataGroup_hi_1855 = {dataGroup_hi_hi_1855, dataGroup_hi_lo_1855};
  wire [31:0]   dataGroup_7_87 = dataGroup_hi_1855[351:320];
  wire [63:0]   res_lo_lo_87 = {dataGroup_1_87, dataGroup_0_87};
  wire [63:0]   res_lo_hi_87 = {dataGroup_3_87, dataGroup_2_87};
  wire [127:0]  res_lo_87 = {res_lo_hi_87, res_lo_lo_87};
  wire [63:0]   res_hi_lo_87 = {dataGroup_5_87, dataGroup_4_87};
  wire [63:0]   res_hi_hi_87 = {dataGroup_7_87, dataGroup_6_87};
  wire [127:0]  res_hi_87 = {res_hi_hi_87, res_hi_lo_87};
  wire [255:0]  res_168 = {res_hi_87, res_lo_87};
  wire [1023:0] dataGroup_lo_1856 = {dataGroup_lo_hi_1856, dataGroup_lo_lo_1856};
  wire [1023:0] dataGroup_hi_1856 = {dataGroup_hi_hi_1856, dataGroup_hi_lo_1856};
  wire [31:0]   dataGroup_0_88 = dataGroup_lo_1856[63:32];
  wire [1023:0] dataGroup_lo_1857 = {dataGroup_lo_hi_1857, dataGroup_lo_lo_1857};
  wire [1023:0] dataGroup_hi_1857 = {dataGroup_hi_hi_1857, dataGroup_hi_lo_1857};
  wire [31:0]   dataGroup_1_88 = dataGroup_lo_1857[255:224];
  wire [1023:0] dataGroup_lo_1858 = {dataGroup_lo_hi_1858, dataGroup_lo_lo_1858};
  wire [1023:0] dataGroup_hi_1858 = {dataGroup_hi_hi_1858, dataGroup_hi_lo_1858};
  wire [31:0]   dataGroup_2_88 = dataGroup_lo_1858[447:416];
  wire [1023:0] dataGroup_lo_1859 = {dataGroup_lo_hi_1859, dataGroup_lo_lo_1859};
  wire [1023:0] dataGroup_hi_1859 = {dataGroup_hi_hi_1859, dataGroup_hi_lo_1859};
  wire [31:0]   dataGroup_3_88 = dataGroup_lo_1859[639:608];
  wire [1023:0] dataGroup_lo_1860 = {dataGroup_lo_hi_1860, dataGroup_lo_lo_1860};
  wire [1023:0] dataGroup_hi_1860 = {dataGroup_hi_hi_1860, dataGroup_hi_lo_1860};
  wire [31:0]   dataGroup_4_88 = dataGroup_lo_1860[831:800];
  wire [1023:0] dataGroup_lo_1861 = {dataGroup_lo_hi_1861, dataGroup_lo_lo_1861};
  wire [1023:0] dataGroup_hi_1861 = {dataGroup_hi_hi_1861, dataGroup_hi_lo_1861};
  wire [31:0]   dataGroup_5_88 = dataGroup_lo_1861[1023:992];
  wire [1023:0] dataGroup_lo_1862 = {dataGroup_lo_hi_1862, dataGroup_lo_lo_1862};
  wire [1023:0] dataGroup_hi_1862 = {dataGroup_hi_hi_1862, dataGroup_hi_lo_1862};
  wire [31:0]   dataGroup_6_88 = dataGroup_hi_1862[191:160];
  wire [1023:0] dataGroup_lo_1863 = {dataGroup_lo_hi_1863, dataGroup_lo_lo_1863};
  wire [1023:0] dataGroup_hi_1863 = {dataGroup_hi_hi_1863, dataGroup_hi_lo_1863};
  wire [31:0]   dataGroup_7_88 = dataGroup_hi_1863[383:352];
  wire [63:0]   res_lo_lo_88 = {dataGroup_1_88, dataGroup_0_88};
  wire [63:0]   res_lo_hi_88 = {dataGroup_3_88, dataGroup_2_88};
  wire [127:0]  res_lo_88 = {res_lo_hi_88, res_lo_lo_88};
  wire [63:0]   res_hi_lo_88 = {dataGroup_5_88, dataGroup_4_88};
  wire [63:0]   res_hi_hi_88 = {dataGroup_7_88, dataGroup_6_88};
  wire [127:0]  res_hi_88 = {res_hi_hi_88, res_hi_lo_88};
  wire [255:0]  res_169 = {res_hi_88, res_lo_88};
  wire [1023:0] dataGroup_lo_1864 = {dataGroup_lo_hi_1864, dataGroup_lo_lo_1864};
  wire [1023:0] dataGroup_hi_1864 = {dataGroup_hi_hi_1864, dataGroup_hi_lo_1864};
  wire [31:0]   dataGroup_0_89 = dataGroup_lo_1864[95:64];
  wire [1023:0] dataGroup_lo_1865 = {dataGroup_lo_hi_1865, dataGroup_lo_lo_1865};
  wire [1023:0] dataGroup_hi_1865 = {dataGroup_hi_hi_1865, dataGroup_hi_lo_1865};
  wire [31:0]   dataGroup_1_89 = dataGroup_lo_1865[287:256];
  wire [1023:0] dataGroup_lo_1866 = {dataGroup_lo_hi_1866, dataGroup_lo_lo_1866};
  wire [1023:0] dataGroup_hi_1866 = {dataGroup_hi_hi_1866, dataGroup_hi_lo_1866};
  wire [31:0]   dataGroup_2_89 = dataGroup_lo_1866[479:448];
  wire [1023:0] dataGroup_lo_1867 = {dataGroup_lo_hi_1867, dataGroup_lo_lo_1867};
  wire [1023:0] dataGroup_hi_1867 = {dataGroup_hi_hi_1867, dataGroup_hi_lo_1867};
  wire [31:0]   dataGroup_3_89 = dataGroup_lo_1867[671:640];
  wire [1023:0] dataGroup_lo_1868 = {dataGroup_lo_hi_1868, dataGroup_lo_lo_1868};
  wire [1023:0] dataGroup_hi_1868 = {dataGroup_hi_hi_1868, dataGroup_hi_lo_1868};
  wire [31:0]   dataGroup_4_89 = dataGroup_lo_1868[863:832];
  wire [1023:0] dataGroup_lo_1869 = {dataGroup_lo_hi_1869, dataGroup_lo_lo_1869};
  wire [1023:0] dataGroup_hi_1869 = {dataGroup_hi_hi_1869, dataGroup_hi_lo_1869};
  wire [31:0]   dataGroup_5_89 = dataGroup_hi_1869[31:0];
  wire [1023:0] dataGroup_lo_1870 = {dataGroup_lo_hi_1870, dataGroup_lo_lo_1870};
  wire [1023:0] dataGroup_hi_1870 = {dataGroup_hi_hi_1870, dataGroup_hi_lo_1870};
  wire [31:0]   dataGroup_6_89 = dataGroup_hi_1870[223:192];
  wire [1023:0] dataGroup_lo_1871 = {dataGroup_lo_hi_1871, dataGroup_lo_lo_1871};
  wire [1023:0] dataGroup_hi_1871 = {dataGroup_hi_hi_1871, dataGroup_hi_lo_1871};
  wire [31:0]   dataGroup_7_89 = dataGroup_hi_1871[415:384];
  wire [63:0]   res_lo_lo_89 = {dataGroup_1_89, dataGroup_0_89};
  wire [63:0]   res_lo_hi_89 = {dataGroup_3_89, dataGroup_2_89};
  wire [127:0]  res_lo_89 = {res_lo_hi_89, res_lo_lo_89};
  wire [63:0]   res_hi_lo_89 = {dataGroup_5_89, dataGroup_4_89};
  wire [63:0]   res_hi_hi_89 = {dataGroup_7_89, dataGroup_6_89};
  wire [127:0]  res_hi_89 = {res_hi_hi_89, res_hi_lo_89};
  wire [255:0]  res_170 = {res_hi_89, res_lo_89};
  wire [1023:0] dataGroup_lo_1872 = {dataGroup_lo_hi_1872, dataGroup_lo_lo_1872};
  wire [1023:0] dataGroup_hi_1872 = {dataGroup_hi_hi_1872, dataGroup_hi_lo_1872};
  wire [31:0]   dataGroup_0_90 = dataGroup_lo_1872[127:96];
  wire [1023:0] dataGroup_lo_1873 = {dataGroup_lo_hi_1873, dataGroup_lo_lo_1873};
  wire [1023:0] dataGroup_hi_1873 = {dataGroup_hi_hi_1873, dataGroup_hi_lo_1873};
  wire [31:0]   dataGroup_1_90 = dataGroup_lo_1873[319:288];
  wire [1023:0] dataGroup_lo_1874 = {dataGroup_lo_hi_1874, dataGroup_lo_lo_1874};
  wire [1023:0] dataGroup_hi_1874 = {dataGroup_hi_hi_1874, dataGroup_hi_lo_1874};
  wire [31:0]   dataGroup_2_90 = dataGroup_lo_1874[511:480];
  wire [1023:0] dataGroup_lo_1875 = {dataGroup_lo_hi_1875, dataGroup_lo_lo_1875};
  wire [1023:0] dataGroup_hi_1875 = {dataGroup_hi_hi_1875, dataGroup_hi_lo_1875};
  wire [31:0]   dataGroup_3_90 = dataGroup_lo_1875[703:672];
  wire [1023:0] dataGroup_lo_1876 = {dataGroup_lo_hi_1876, dataGroup_lo_lo_1876};
  wire [1023:0] dataGroup_hi_1876 = {dataGroup_hi_hi_1876, dataGroup_hi_lo_1876};
  wire [31:0]   dataGroup_4_90 = dataGroup_lo_1876[895:864];
  wire [1023:0] dataGroup_lo_1877 = {dataGroup_lo_hi_1877, dataGroup_lo_lo_1877};
  wire [1023:0] dataGroup_hi_1877 = {dataGroup_hi_hi_1877, dataGroup_hi_lo_1877};
  wire [31:0]   dataGroup_5_90 = dataGroup_hi_1877[63:32];
  wire [1023:0] dataGroup_lo_1878 = {dataGroup_lo_hi_1878, dataGroup_lo_lo_1878};
  wire [1023:0] dataGroup_hi_1878 = {dataGroup_hi_hi_1878, dataGroup_hi_lo_1878};
  wire [31:0]   dataGroup_6_90 = dataGroup_hi_1878[255:224];
  wire [1023:0] dataGroup_lo_1879 = {dataGroup_lo_hi_1879, dataGroup_lo_lo_1879};
  wire [1023:0] dataGroup_hi_1879 = {dataGroup_hi_hi_1879, dataGroup_hi_lo_1879};
  wire [31:0]   dataGroup_7_90 = dataGroup_hi_1879[447:416];
  wire [63:0]   res_lo_lo_90 = {dataGroup_1_90, dataGroup_0_90};
  wire [63:0]   res_lo_hi_90 = {dataGroup_3_90, dataGroup_2_90};
  wire [127:0]  res_lo_90 = {res_lo_hi_90, res_lo_lo_90};
  wire [63:0]   res_hi_lo_90 = {dataGroup_5_90, dataGroup_4_90};
  wire [63:0]   res_hi_hi_90 = {dataGroup_7_90, dataGroup_6_90};
  wire [127:0]  res_hi_90 = {res_hi_hi_90, res_hi_lo_90};
  wire [255:0]  res_171 = {res_hi_90, res_lo_90};
  wire [1023:0] dataGroup_lo_1880 = {dataGroup_lo_hi_1880, dataGroup_lo_lo_1880};
  wire [1023:0] dataGroup_hi_1880 = {dataGroup_hi_hi_1880, dataGroup_hi_lo_1880};
  wire [31:0]   dataGroup_0_91 = dataGroup_lo_1880[159:128];
  wire [1023:0] dataGroup_lo_1881 = {dataGroup_lo_hi_1881, dataGroup_lo_lo_1881};
  wire [1023:0] dataGroup_hi_1881 = {dataGroup_hi_hi_1881, dataGroup_hi_lo_1881};
  wire [31:0]   dataGroup_1_91 = dataGroup_lo_1881[351:320];
  wire [1023:0] dataGroup_lo_1882 = {dataGroup_lo_hi_1882, dataGroup_lo_lo_1882};
  wire [1023:0] dataGroup_hi_1882 = {dataGroup_hi_hi_1882, dataGroup_hi_lo_1882};
  wire [31:0]   dataGroup_2_91 = dataGroup_lo_1882[543:512];
  wire [1023:0] dataGroup_lo_1883 = {dataGroup_lo_hi_1883, dataGroup_lo_lo_1883};
  wire [1023:0] dataGroup_hi_1883 = {dataGroup_hi_hi_1883, dataGroup_hi_lo_1883};
  wire [31:0]   dataGroup_3_91 = dataGroup_lo_1883[735:704];
  wire [1023:0] dataGroup_lo_1884 = {dataGroup_lo_hi_1884, dataGroup_lo_lo_1884};
  wire [1023:0] dataGroup_hi_1884 = {dataGroup_hi_hi_1884, dataGroup_hi_lo_1884};
  wire [31:0]   dataGroup_4_91 = dataGroup_lo_1884[927:896];
  wire [1023:0] dataGroup_lo_1885 = {dataGroup_lo_hi_1885, dataGroup_lo_lo_1885};
  wire [1023:0] dataGroup_hi_1885 = {dataGroup_hi_hi_1885, dataGroup_hi_lo_1885};
  wire [31:0]   dataGroup_5_91 = dataGroup_hi_1885[95:64];
  wire [1023:0] dataGroup_lo_1886 = {dataGroup_lo_hi_1886, dataGroup_lo_lo_1886};
  wire [1023:0] dataGroup_hi_1886 = {dataGroup_hi_hi_1886, dataGroup_hi_lo_1886};
  wire [31:0]   dataGroup_6_91 = dataGroup_hi_1886[287:256];
  wire [1023:0] dataGroup_lo_1887 = {dataGroup_lo_hi_1887, dataGroup_lo_lo_1887};
  wire [1023:0] dataGroup_hi_1887 = {dataGroup_hi_hi_1887, dataGroup_hi_lo_1887};
  wire [31:0]   dataGroup_7_91 = dataGroup_hi_1887[479:448];
  wire [63:0]   res_lo_lo_91 = {dataGroup_1_91, dataGroup_0_91};
  wire [63:0]   res_lo_hi_91 = {dataGroup_3_91, dataGroup_2_91};
  wire [127:0]  res_lo_91 = {res_lo_hi_91, res_lo_lo_91};
  wire [63:0]   res_hi_lo_91 = {dataGroup_5_91, dataGroup_4_91};
  wire [63:0]   res_hi_hi_91 = {dataGroup_7_91, dataGroup_6_91};
  wire [127:0]  res_hi_91 = {res_hi_hi_91, res_hi_lo_91};
  wire [255:0]  res_172 = {res_hi_91, res_lo_91};
  wire [1023:0] dataGroup_lo_1888 = {dataGroup_lo_hi_1888, dataGroup_lo_lo_1888};
  wire [1023:0] dataGroup_hi_1888 = {dataGroup_hi_hi_1888, dataGroup_hi_lo_1888};
  wire [31:0]   dataGroup_0_92 = dataGroup_lo_1888[191:160];
  wire [1023:0] dataGroup_lo_1889 = {dataGroup_lo_hi_1889, dataGroup_lo_lo_1889};
  wire [1023:0] dataGroup_hi_1889 = {dataGroup_hi_hi_1889, dataGroup_hi_lo_1889};
  wire [31:0]   dataGroup_1_92 = dataGroup_lo_1889[383:352];
  wire [1023:0] dataGroup_lo_1890 = {dataGroup_lo_hi_1890, dataGroup_lo_lo_1890};
  wire [1023:0] dataGroup_hi_1890 = {dataGroup_hi_hi_1890, dataGroup_hi_lo_1890};
  wire [31:0]   dataGroup_2_92 = dataGroup_lo_1890[575:544];
  wire [1023:0] dataGroup_lo_1891 = {dataGroup_lo_hi_1891, dataGroup_lo_lo_1891};
  wire [1023:0] dataGroup_hi_1891 = {dataGroup_hi_hi_1891, dataGroup_hi_lo_1891};
  wire [31:0]   dataGroup_3_92 = dataGroup_lo_1891[767:736];
  wire [1023:0] dataGroup_lo_1892 = {dataGroup_lo_hi_1892, dataGroup_lo_lo_1892};
  wire [1023:0] dataGroup_hi_1892 = {dataGroup_hi_hi_1892, dataGroup_hi_lo_1892};
  wire [31:0]   dataGroup_4_92 = dataGroup_lo_1892[959:928];
  wire [1023:0] dataGroup_lo_1893 = {dataGroup_lo_hi_1893, dataGroup_lo_lo_1893};
  wire [1023:0] dataGroup_hi_1893 = {dataGroup_hi_hi_1893, dataGroup_hi_lo_1893};
  wire [31:0]   dataGroup_5_92 = dataGroup_hi_1893[127:96];
  wire [1023:0] dataGroup_lo_1894 = {dataGroup_lo_hi_1894, dataGroup_lo_lo_1894};
  wire [1023:0] dataGroup_hi_1894 = {dataGroup_hi_hi_1894, dataGroup_hi_lo_1894};
  wire [31:0]   dataGroup_6_92 = dataGroup_hi_1894[319:288];
  wire [1023:0] dataGroup_lo_1895 = {dataGroup_lo_hi_1895, dataGroup_lo_lo_1895};
  wire [1023:0] dataGroup_hi_1895 = {dataGroup_hi_hi_1895, dataGroup_hi_lo_1895};
  wire [31:0]   dataGroup_7_92 = dataGroup_hi_1895[511:480];
  wire [63:0]   res_lo_lo_92 = {dataGroup_1_92, dataGroup_0_92};
  wire [63:0]   res_lo_hi_92 = {dataGroup_3_92, dataGroup_2_92};
  wire [127:0]  res_lo_92 = {res_lo_hi_92, res_lo_lo_92};
  wire [63:0]   res_hi_lo_92 = {dataGroup_5_92, dataGroup_4_92};
  wire [63:0]   res_hi_hi_92 = {dataGroup_7_92, dataGroup_6_92};
  wire [127:0]  res_hi_92 = {res_hi_hi_92, res_hi_lo_92};
  wire [255:0]  res_173 = {res_hi_92, res_lo_92};
  wire [511:0]  lo_lo_21 = {res_169, res_168};
  wire [511:0]  lo_hi_21 = {res_171, res_170};
  wire [1023:0] lo_21 = {lo_hi_21, lo_lo_21};
  wire [511:0]  hi_lo_21 = {res_173, res_172};
  wire [1023:0] hi_21 = {512'h0, hi_lo_21};
  wire [2047:0] regroupLoadData_2_5 = {hi_21, lo_21};
  wire [1023:0] dataGroup_lo_1896 = {dataGroup_lo_hi_1896, dataGroup_lo_lo_1896};
  wire [1023:0] dataGroup_hi_1896 = {dataGroup_hi_hi_1896, dataGroup_hi_lo_1896};
  wire [31:0]   dataGroup_0_93 = dataGroup_lo_1896[31:0];
  wire [1023:0] dataGroup_lo_1897 = {dataGroup_lo_hi_1897, dataGroup_lo_lo_1897};
  wire [1023:0] dataGroup_hi_1897 = {dataGroup_hi_hi_1897, dataGroup_hi_lo_1897};
  wire [31:0]   dataGroup_1_93 = dataGroup_lo_1897[255:224];
  wire [1023:0] dataGroup_lo_1898 = {dataGroup_lo_hi_1898, dataGroup_lo_lo_1898};
  wire [1023:0] dataGroup_hi_1898 = {dataGroup_hi_hi_1898, dataGroup_hi_lo_1898};
  wire [31:0]   dataGroup_2_93 = dataGroup_lo_1898[479:448];
  wire [1023:0] dataGroup_lo_1899 = {dataGroup_lo_hi_1899, dataGroup_lo_lo_1899};
  wire [1023:0] dataGroup_hi_1899 = {dataGroup_hi_hi_1899, dataGroup_hi_lo_1899};
  wire [31:0]   dataGroup_3_93 = dataGroup_lo_1899[703:672];
  wire [1023:0] dataGroup_lo_1900 = {dataGroup_lo_hi_1900, dataGroup_lo_lo_1900};
  wire [1023:0] dataGroup_hi_1900 = {dataGroup_hi_hi_1900, dataGroup_hi_lo_1900};
  wire [31:0]   dataGroup_4_93 = dataGroup_lo_1900[927:896];
  wire [1023:0] dataGroup_lo_1901 = {dataGroup_lo_hi_1901, dataGroup_lo_lo_1901};
  wire [1023:0] dataGroup_hi_1901 = {dataGroup_hi_hi_1901, dataGroup_hi_lo_1901};
  wire [31:0]   dataGroup_5_93 = dataGroup_hi_1901[127:96];
  wire [1023:0] dataGroup_lo_1902 = {dataGroup_lo_hi_1902, dataGroup_lo_lo_1902};
  wire [1023:0] dataGroup_hi_1902 = {dataGroup_hi_hi_1902, dataGroup_hi_lo_1902};
  wire [31:0]   dataGroup_6_93 = dataGroup_hi_1902[351:320];
  wire [1023:0] dataGroup_lo_1903 = {dataGroup_lo_hi_1903, dataGroup_lo_lo_1903};
  wire [1023:0] dataGroup_hi_1903 = {dataGroup_hi_hi_1903, dataGroup_hi_lo_1903};
  wire [31:0]   dataGroup_7_93 = dataGroup_hi_1903[575:544];
  wire [63:0]   res_lo_lo_93 = {dataGroup_1_93, dataGroup_0_93};
  wire [63:0]   res_lo_hi_93 = {dataGroup_3_93, dataGroup_2_93};
  wire [127:0]  res_lo_93 = {res_lo_hi_93, res_lo_lo_93};
  wire [63:0]   res_hi_lo_93 = {dataGroup_5_93, dataGroup_4_93};
  wire [63:0]   res_hi_hi_93 = {dataGroup_7_93, dataGroup_6_93};
  wire [127:0]  res_hi_93 = {res_hi_hi_93, res_hi_lo_93};
  wire [255:0]  res_176 = {res_hi_93, res_lo_93};
  wire [1023:0] dataGroup_lo_1904 = {dataGroup_lo_hi_1904, dataGroup_lo_lo_1904};
  wire [1023:0] dataGroup_hi_1904 = {dataGroup_hi_hi_1904, dataGroup_hi_lo_1904};
  wire [31:0]   dataGroup_0_94 = dataGroup_lo_1904[63:32];
  wire [1023:0] dataGroup_lo_1905 = {dataGroup_lo_hi_1905, dataGroup_lo_lo_1905};
  wire [1023:0] dataGroup_hi_1905 = {dataGroup_hi_hi_1905, dataGroup_hi_lo_1905};
  wire [31:0]   dataGroup_1_94 = dataGroup_lo_1905[287:256];
  wire [1023:0] dataGroup_lo_1906 = {dataGroup_lo_hi_1906, dataGroup_lo_lo_1906};
  wire [1023:0] dataGroup_hi_1906 = {dataGroup_hi_hi_1906, dataGroup_hi_lo_1906};
  wire [31:0]   dataGroup_2_94 = dataGroup_lo_1906[511:480];
  wire [1023:0] dataGroup_lo_1907 = {dataGroup_lo_hi_1907, dataGroup_lo_lo_1907};
  wire [1023:0] dataGroup_hi_1907 = {dataGroup_hi_hi_1907, dataGroup_hi_lo_1907};
  wire [31:0]   dataGroup_3_94 = dataGroup_lo_1907[735:704];
  wire [1023:0] dataGroup_lo_1908 = {dataGroup_lo_hi_1908, dataGroup_lo_lo_1908};
  wire [1023:0] dataGroup_hi_1908 = {dataGroup_hi_hi_1908, dataGroup_hi_lo_1908};
  wire [31:0]   dataGroup_4_94 = dataGroup_lo_1908[959:928];
  wire [1023:0] dataGroup_lo_1909 = {dataGroup_lo_hi_1909, dataGroup_lo_lo_1909};
  wire [1023:0] dataGroup_hi_1909 = {dataGroup_hi_hi_1909, dataGroup_hi_lo_1909};
  wire [31:0]   dataGroup_5_94 = dataGroup_hi_1909[159:128];
  wire [1023:0] dataGroup_lo_1910 = {dataGroup_lo_hi_1910, dataGroup_lo_lo_1910};
  wire [1023:0] dataGroup_hi_1910 = {dataGroup_hi_hi_1910, dataGroup_hi_lo_1910};
  wire [31:0]   dataGroup_6_94 = dataGroup_hi_1910[383:352];
  wire [1023:0] dataGroup_lo_1911 = {dataGroup_lo_hi_1911, dataGroup_lo_lo_1911};
  wire [1023:0] dataGroup_hi_1911 = {dataGroup_hi_hi_1911, dataGroup_hi_lo_1911};
  wire [31:0]   dataGroup_7_94 = dataGroup_hi_1911[607:576];
  wire [63:0]   res_lo_lo_94 = {dataGroup_1_94, dataGroup_0_94};
  wire [63:0]   res_lo_hi_94 = {dataGroup_3_94, dataGroup_2_94};
  wire [127:0]  res_lo_94 = {res_lo_hi_94, res_lo_lo_94};
  wire [63:0]   res_hi_lo_94 = {dataGroup_5_94, dataGroup_4_94};
  wire [63:0]   res_hi_hi_94 = {dataGroup_7_94, dataGroup_6_94};
  wire [127:0]  res_hi_94 = {res_hi_hi_94, res_hi_lo_94};
  wire [255:0]  res_177 = {res_hi_94, res_lo_94};
  wire [1023:0] dataGroup_lo_1912 = {dataGroup_lo_hi_1912, dataGroup_lo_lo_1912};
  wire [1023:0] dataGroup_hi_1912 = {dataGroup_hi_hi_1912, dataGroup_hi_lo_1912};
  wire [31:0]   dataGroup_0_95 = dataGroup_lo_1912[95:64];
  wire [1023:0] dataGroup_lo_1913 = {dataGroup_lo_hi_1913, dataGroup_lo_lo_1913};
  wire [1023:0] dataGroup_hi_1913 = {dataGroup_hi_hi_1913, dataGroup_hi_lo_1913};
  wire [31:0]   dataGroup_1_95 = dataGroup_lo_1913[319:288];
  wire [1023:0] dataGroup_lo_1914 = {dataGroup_lo_hi_1914, dataGroup_lo_lo_1914};
  wire [1023:0] dataGroup_hi_1914 = {dataGroup_hi_hi_1914, dataGroup_hi_lo_1914};
  wire [31:0]   dataGroup_2_95 = dataGroup_lo_1914[543:512];
  wire [1023:0] dataGroup_lo_1915 = {dataGroup_lo_hi_1915, dataGroup_lo_lo_1915};
  wire [1023:0] dataGroup_hi_1915 = {dataGroup_hi_hi_1915, dataGroup_hi_lo_1915};
  wire [31:0]   dataGroup_3_95 = dataGroup_lo_1915[767:736];
  wire [1023:0] dataGroup_lo_1916 = {dataGroup_lo_hi_1916, dataGroup_lo_lo_1916};
  wire [1023:0] dataGroup_hi_1916 = {dataGroup_hi_hi_1916, dataGroup_hi_lo_1916};
  wire [31:0]   dataGroup_4_95 = dataGroup_lo_1916[991:960];
  wire [1023:0] dataGroup_lo_1917 = {dataGroup_lo_hi_1917, dataGroup_lo_lo_1917};
  wire [1023:0] dataGroup_hi_1917 = {dataGroup_hi_hi_1917, dataGroup_hi_lo_1917};
  wire [31:0]   dataGroup_5_95 = dataGroup_hi_1917[191:160];
  wire [1023:0] dataGroup_lo_1918 = {dataGroup_lo_hi_1918, dataGroup_lo_lo_1918};
  wire [1023:0] dataGroup_hi_1918 = {dataGroup_hi_hi_1918, dataGroup_hi_lo_1918};
  wire [31:0]   dataGroup_6_95 = dataGroup_hi_1918[415:384];
  wire [1023:0] dataGroup_lo_1919 = {dataGroup_lo_hi_1919, dataGroup_lo_lo_1919};
  wire [1023:0] dataGroup_hi_1919 = {dataGroup_hi_hi_1919, dataGroup_hi_lo_1919};
  wire [31:0]   dataGroup_7_95 = dataGroup_hi_1919[639:608];
  wire [63:0]   res_lo_lo_95 = {dataGroup_1_95, dataGroup_0_95};
  wire [63:0]   res_lo_hi_95 = {dataGroup_3_95, dataGroup_2_95};
  wire [127:0]  res_lo_95 = {res_lo_hi_95, res_lo_lo_95};
  wire [63:0]   res_hi_lo_95 = {dataGroup_5_95, dataGroup_4_95};
  wire [63:0]   res_hi_hi_95 = {dataGroup_7_95, dataGroup_6_95};
  wire [127:0]  res_hi_95 = {res_hi_hi_95, res_hi_lo_95};
  wire [255:0]  res_178 = {res_hi_95, res_lo_95};
  wire [1023:0] dataGroup_lo_1920 = {dataGroup_lo_hi_1920, dataGroup_lo_lo_1920};
  wire [1023:0] dataGroup_hi_1920 = {dataGroup_hi_hi_1920, dataGroup_hi_lo_1920};
  wire [31:0]   dataGroup_0_96 = dataGroup_lo_1920[127:96];
  wire [1023:0] dataGroup_lo_1921 = {dataGroup_lo_hi_1921, dataGroup_lo_lo_1921};
  wire [1023:0] dataGroup_hi_1921 = {dataGroup_hi_hi_1921, dataGroup_hi_lo_1921};
  wire [31:0]   dataGroup_1_96 = dataGroup_lo_1921[351:320];
  wire [1023:0] dataGroup_lo_1922 = {dataGroup_lo_hi_1922, dataGroup_lo_lo_1922};
  wire [1023:0] dataGroup_hi_1922 = {dataGroup_hi_hi_1922, dataGroup_hi_lo_1922};
  wire [31:0]   dataGroup_2_96 = dataGroup_lo_1922[575:544];
  wire [1023:0] dataGroup_lo_1923 = {dataGroup_lo_hi_1923, dataGroup_lo_lo_1923};
  wire [1023:0] dataGroup_hi_1923 = {dataGroup_hi_hi_1923, dataGroup_hi_lo_1923};
  wire [31:0]   dataGroup_3_96 = dataGroup_lo_1923[799:768];
  wire [1023:0] dataGroup_lo_1924 = {dataGroup_lo_hi_1924, dataGroup_lo_lo_1924};
  wire [1023:0] dataGroup_hi_1924 = {dataGroup_hi_hi_1924, dataGroup_hi_lo_1924};
  wire [31:0]   dataGroup_4_96 = dataGroup_lo_1924[1023:992];
  wire [1023:0] dataGroup_lo_1925 = {dataGroup_lo_hi_1925, dataGroup_lo_lo_1925};
  wire [1023:0] dataGroup_hi_1925 = {dataGroup_hi_hi_1925, dataGroup_hi_lo_1925};
  wire [31:0]   dataGroup_5_96 = dataGroup_hi_1925[223:192];
  wire [1023:0] dataGroup_lo_1926 = {dataGroup_lo_hi_1926, dataGroup_lo_lo_1926};
  wire [1023:0] dataGroup_hi_1926 = {dataGroup_hi_hi_1926, dataGroup_hi_lo_1926};
  wire [31:0]   dataGroup_6_96 = dataGroup_hi_1926[447:416];
  wire [1023:0] dataGroup_lo_1927 = {dataGroup_lo_hi_1927, dataGroup_lo_lo_1927};
  wire [1023:0] dataGroup_hi_1927 = {dataGroup_hi_hi_1927, dataGroup_hi_lo_1927};
  wire [31:0]   dataGroup_7_96 = dataGroup_hi_1927[671:640];
  wire [63:0]   res_lo_lo_96 = {dataGroup_1_96, dataGroup_0_96};
  wire [63:0]   res_lo_hi_96 = {dataGroup_3_96, dataGroup_2_96};
  wire [127:0]  res_lo_96 = {res_lo_hi_96, res_lo_lo_96};
  wire [63:0]   res_hi_lo_96 = {dataGroup_5_96, dataGroup_4_96};
  wire [63:0]   res_hi_hi_96 = {dataGroup_7_96, dataGroup_6_96};
  wire [127:0]  res_hi_96 = {res_hi_hi_96, res_hi_lo_96};
  wire [255:0]  res_179 = {res_hi_96, res_lo_96};
  wire [1023:0] dataGroup_lo_1928 = {dataGroup_lo_hi_1928, dataGroup_lo_lo_1928};
  wire [1023:0] dataGroup_hi_1928 = {dataGroup_hi_hi_1928, dataGroup_hi_lo_1928};
  wire [31:0]   dataGroup_0_97 = dataGroup_lo_1928[159:128];
  wire [1023:0] dataGroup_lo_1929 = {dataGroup_lo_hi_1929, dataGroup_lo_lo_1929};
  wire [1023:0] dataGroup_hi_1929 = {dataGroup_hi_hi_1929, dataGroup_hi_lo_1929};
  wire [31:0]   dataGroup_1_97 = dataGroup_lo_1929[383:352];
  wire [1023:0] dataGroup_lo_1930 = {dataGroup_lo_hi_1930, dataGroup_lo_lo_1930};
  wire [1023:0] dataGroup_hi_1930 = {dataGroup_hi_hi_1930, dataGroup_hi_lo_1930};
  wire [31:0]   dataGroup_2_97 = dataGroup_lo_1930[607:576];
  wire [1023:0] dataGroup_lo_1931 = {dataGroup_lo_hi_1931, dataGroup_lo_lo_1931};
  wire [1023:0] dataGroup_hi_1931 = {dataGroup_hi_hi_1931, dataGroup_hi_lo_1931};
  wire [31:0]   dataGroup_3_97 = dataGroup_lo_1931[831:800];
  wire [1023:0] dataGroup_lo_1932 = {dataGroup_lo_hi_1932, dataGroup_lo_lo_1932};
  wire [1023:0] dataGroup_hi_1932 = {dataGroup_hi_hi_1932, dataGroup_hi_lo_1932};
  wire [31:0]   dataGroup_4_97 = dataGroup_hi_1932[31:0];
  wire [1023:0] dataGroup_lo_1933 = {dataGroup_lo_hi_1933, dataGroup_lo_lo_1933};
  wire [1023:0] dataGroup_hi_1933 = {dataGroup_hi_hi_1933, dataGroup_hi_lo_1933};
  wire [31:0]   dataGroup_5_97 = dataGroup_hi_1933[255:224];
  wire [1023:0] dataGroup_lo_1934 = {dataGroup_lo_hi_1934, dataGroup_lo_lo_1934};
  wire [1023:0] dataGroup_hi_1934 = {dataGroup_hi_hi_1934, dataGroup_hi_lo_1934};
  wire [31:0]   dataGroup_6_97 = dataGroup_hi_1934[479:448];
  wire [1023:0] dataGroup_lo_1935 = {dataGroup_lo_hi_1935, dataGroup_lo_lo_1935};
  wire [1023:0] dataGroup_hi_1935 = {dataGroup_hi_hi_1935, dataGroup_hi_lo_1935};
  wire [31:0]   dataGroup_7_97 = dataGroup_hi_1935[703:672];
  wire [63:0]   res_lo_lo_97 = {dataGroup_1_97, dataGroup_0_97};
  wire [63:0]   res_lo_hi_97 = {dataGroup_3_97, dataGroup_2_97};
  wire [127:0]  res_lo_97 = {res_lo_hi_97, res_lo_lo_97};
  wire [63:0]   res_hi_lo_97 = {dataGroup_5_97, dataGroup_4_97};
  wire [63:0]   res_hi_hi_97 = {dataGroup_7_97, dataGroup_6_97};
  wire [127:0]  res_hi_97 = {res_hi_hi_97, res_hi_lo_97};
  wire [255:0]  res_180 = {res_hi_97, res_lo_97};
  wire [1023:0] dataGroup_lo_1936 = {dataGroup_lo_hi_1936, dataGroup_lo_lo_1936};
  wire [1023:0] dataGroup_hi_1936 = {dataGroup_hi_hi_1936, dataGroup_hi_lo_1936};
  wire [31:0]   dataGroup_0_98 = dataGroup_lo_1936[191:160];
  wire [1023:0] dataGroup_lo_1937 = {dataGroup_lo_hi_1937, dataGroup_lo_lo_1937};
  wire [1023:0] dataGroup_hi_1937 = {dataGroup_hi_hi_1937, dataGroup_hi_lo_1937};
  wire [31:0]   dataGroup_1_98 = dataGroup_lo_1937[415:384];
  wire [1023:0] dataGroup_lo_1938 = {dataGroup_lo_hi_1938, dataGroup_lo_lo_1938};
  wire [1023:0] dataGroup_hi_1938 = {dataGroup_hi_hi_1938, dataGroup_hi_lo_1938};
  wire [31:0]   dataGroup_2_98 = dataGroup_lo_1938[639:608];
  wire [1023:0] dataGroup_lo_1939 = {dataGroup_lo_hi_1939, dataGroup_lo_lo_1939};
  wire [1023:0] dataGroup_hi_1939 = {dataGroup_hi_hi_1939, dataGroup_hi_lo_1939};
  wire [31:0]   dataGroup_3_98 = dataGroup_lo_1939[863:832];
  wire [1023:0] dataGroup_lo_1940 = {dataGroup_lo_hi_1940, dataGroup_lo_lo_1940};
  wire [1023:0] dataGroup_hi_1940 = {dataGroup_hi_hi_1940, dataGroup_hi_lo_1940};
  wire [31:0]   dataGroup_4_98 = dataGroup_hi_1940[63:32];
  wire [1023:0] dataGroup_lo_1941 = {dataGroup_lo_hi_1941, dataGroup_lo_lo_1941};
  wire [1023:0] dataGroup_hi_1941 = {dataGroup_hi_hi_1941, dataGroup_hi_lo_1941};
  wire [31:0]   dataGroup_5_98 = dataGroup_hi_1941[287:256];
  wire [1023:0] dataGroup_lo_1942 = {dataGroup_lo_hi_1942, dataGroup_lo_lo_1942};
  wire [1023:0] dataGroup_hi_1942 = {dataGroup_hi_hi_1942, dataGroup_hi_lo_1942};
  wire [31:0]   dataGroup_6_98 = dataGroup_hi_1942[511:480];
  wire [1023:0] dataGroup_lo_1943 = {dataGroup_lo_hi_1943, dataGroup_lo_lo_1943};
  wire [1023:0] dataGroup_hi_1943 = {dataGroup_hi_hi_1943, dataGroup_hi_lo_1943};
  wire [31:0]   dataGroup_7_98 = dataGroup_hi_1943[735:704];
  wire [63:0]   res_lo_lo_98 = {dataGroup_1_98, dataGroup_0_98};
  wire [63:0]   res_lo_hi_98 = {dataGroup_3_98, dataGroup_2_98};
  wire [127:0]  res_lo_98 = {res_lo_hi_98, res_lo_lo_98};
  wire [63:0]   res_hi_lo_98 = {dataGroup_5_98, dataGroup_4_98};
  wire [63:0]   res_hi_hi_98 = {dataGroup_7_98, dataGroup_6_98};
  wire [127:0]  res_hi_98 = {res_hi_hi_98, res_hi_lo_98};
  wire [255:0]  res_181 = {res_hi_98, res_lo_98};
  wire [1023:0] dataGroup_lo_1944 = {dataGroup_lo_hi_1944, dataGroup_lo_lo_1944};
  wire [1023:0] dataGroup_hi_1944 = {dataGroup_hi_hi_1944, dataGroup_hi_lo_1944};
  wire [31:0]   dataGroup_0_99 = dataGroup_lo_1944[223:192];
  wire [1023:0] dataGroup_lo_1945 = {dataGroup_lo_hi_1945, dataGroup_lo_lo_1945};
  wire [1023:0] dataGroup_hi_1945 = {dataGroup_hi_hi_1945, dataGroup_hi_lo_1945};
  wire [31:0]   dataGroup_1_99 = dataGroup_lo_1945[447:416];
  wire [1023:0] dataGroup_lo_1946 = {dataGroup_lo_hi_1946, dataGroup_lo_lo_1946};
  wire [1023:0] dataGroup_hi_1946 = {dataGroup_hi_hi_1946, dataGroup_hi_lo_1946};
  wire [31:0]   dataGroup_2_99 = dataGroup_lo_1946[671:640];
  wire [1023:0] dataGroup_lo_1947 = {dataGroup_lo_hi_1947, dataGroup_lo_lo_1947};
  wire [1023:0] dataGroup_hi_1947 = {dataGroup_hi_hi_1947, dataGroup_hi_lo_1947};
  wire [31:0]   dataGroup_3_99 = dataGroup_lo_1947[895:864];
  wire [1023:0] dataGroup_lo_1948 = {dataGroup_lo_hi_1948, dataGroup_lo_lo_1948};
  wire [1023:0] dataGroup_hi_1948 = {dataGroup_hi_hi_1948, dataGroup_hi_lo_1948};
  wire [31:0]   dataGroup_4_99 = dataGroup_hi_1948[95:64];
  wire [1023:0] dataGroup_lo_1949 = {dataGroup_lo_hi_1949, dataGroup_lo_lo_1949};
  wire [1023:0] dataGroup_hi_1949 = {dataGroup_hi_hi_1949, dataGroup_hi_lo_1949};
  wire [31:0]   dataGroup_5_99 = dataGroup_hi_1949[319:288];
  wire [1023:0] dataGroup_lo_1950 = {dataGroup_lo_hi_1950, dataGroup_lo_lo_1950};
  wire [1023:0] dataGroup_hi_1950 = {dataGroup_hi_hi_1950, dataGroup_hi_lo_1950};
  wire [31:0]   dataGroup_6_99 = dataGroup_hi_1950[543:512];
  wire [1023:0] dataGroup_lo_1951 = {dataGroup_lo_hi_1951, dataGroup_lo_lo_1951};
  wire [1023:0] dataGroup_hi_1951 = {dataGroup_hi_hi_1951, dataGroup_hi_lo_1951};
  wire [31:0]   dataGroup_7_99 = dataGroup_hi_1951[767:736];
  wire [63:0]   res_lo_lo_99 = {dataGroup_1_99, dataGroup_0_99};
  wire [63:0]   res_lo_hi_99 = {dataGroup_3_99, dataGroup_2_99};
  wire [127:0]  res_lo_99 = {res_lo_hi_99, res_lo_lo_99};
  wire [63:0]   res_hi_lo_99 = {dataGroup_5_99, dataGroup_4_99};
  wire [63:0]   res_hi_hi_99 = {dataGroup_7_99, dataGroup_6_99};
  wire [127:0]  res_hi_99 = {res_hi_hi_99, res_hi_lo_99};
  wire [255:0]  res_182 = {res_hi_99, res_lo_99};
  wire [511:0]  lo_lo_22 = {res_177, res_176};
  wire [511:0]  lo_hi_22 = {res_179, res_178};
  wire [1023:0] lo_22 = {lo_hi_22, lo_lo_22};
  wire [511:0]  hi_lo_22 = {res_181, res_180};
  wire [511:0]  hi_hi_22 = {256'h0, res_182};
  wire [1023:0] hi_22 = {hi_hi_22, hi_lo_22};
  wire [2047:0] regroupLoadData_2_6 = {hi_22, lo_22};
  wire [1023:0] dataGroup_lo_1952 = {dataGroup_lo_hi_1952, dataGroup_lo_lo_1952};
  wire [1023:0] dataGroup_hi_1952 = {dataGroup_hi_hi_1952, dataGroup_hi_lo_1952};
  wire [31:0]   dataGroup_0_100 = dataGroup_lo_1952[31:0];
  wire [1023:0] dataGroup_lo_1953 = {dataGroup_lo_hi_1953, dataGroup_lo_lo_1953};
  wire [1023:0] dataGroup_hi_1953 = {dataGroup_hi_hi_1953, dataGroup_hi_lo_1953};
  wire [31:0]   dataGroup_1_100 = dataGroup_lo_1953[287:256];
  wire [1023:0] dataGroup_lo_1954 = {dataGroup_lo_hi_1954, dataGroup_lo_lo_1954};
  wire [1023:0] dataGroup_hi_1954 = {dataGroup_hi_hi_1954, dataGroup_hi_lo_1954};
  wire [31:0]   dataGroup_2_100 = dataGroup_lo_1954[543:512];
  wire [1023:0] dataGroup_lo_1955 = {dataGroup_lo_hi_1955, dataGroup_lo_lo_1955};
  wire [1023:0] dataGroup_hi_1955 = {dataGroup_hi_hi_1955, dataGroup_hi_lo_1955};
  wire [31:0]   dataGroup_3_100 = dataGroup_lo_1955[799:768];
  wire [1023:0] dataGroup_lo_1956 = {dataGroup_lo_hi_1956, dataGroup_lo_lo_1956};
  wire [1023:0] dataGroup_hi_1956 = {dataGroup_hi_hi_1956, dataGroup_hi_lo_1956};
  wire [31:0]   dataGroup_4_100 = dataGroup_hi_1956[31:0];
  wire [1023:0] dataGroup_lo_1957 = {dataGroup_lo_hi_1957, dataGroup_lo_lo_1957};
  wire [1023:0] dataGroup_hi_1957 = {dataGroup_hi_hi_1957, dataGroup_hi_lo_1957};
  wire [31:0]   dataGroup_5_100 = dataGroup_hi_1957[287:256];
  wire [1023:0] dataGroup_lo_1958 = {dataGroup_lo_hi_1958, dataGroup_lo_lo_1958};
  wire [1023:0] dataGroup_hi_1958 = {dataGroup_hi_hi_1958, dataGroup_hi_lo_1958};
  wire [31:0]   dataGroup_6_100 = dataGroup_hi_1958[543:512];
  wire [1023:0] dataGroup_lo_1959 = {dataGroup_lo_hi_1959, dataGroup_lo_lo_1959};
  wire [1023:0] dataGroup_hi_1959 = {dataGroup_hi_hi_1959, dataGroup_hi_lo_1959};
  wire [31:0]   dataGroup_7_100 = dataGroup_hi_1959[799:768];
  wire [63:0]   res_lo_lo_100 = {dataGroup_1_100, dataGroup_0_100};
  wire [63:0]   res_lo_hi_100 = {dataGroup_3_100, dataGroup_2_100};
  wire [127:0]  res_lo_100 = {res_lo_hi_100, res_lo_lo_100};
  wire [63:0]   res_hi_lo_100 = {dataGroup_5_100, dataGroup_4_100};
  wire [63:0]   res_hi_hi_100 = {dataGroup_7_100, dataGroup_6_100};
  wire [127:0]  res_hi_100 = {res_hi_hi_100, res_hi_lo_100};
  wire [255:0]  res_184 = {res_hi_100, res_lo_100};
  wire [1023:0] dataGroup_lo_1960 = {dataGroup_lo_hi_1960, dataGroup_lo_lo_1960};
  wire [1023:0] dataGroup_hi_1960 = {dataGroup_hi_hi_1960, dataGroup_hi_lo_1960};
  wire [31:0]   dataGroup_0_101 = dataGroup_lo_1960[63:32];
  wire [1023:0] dataGroup_lo_1961 = {dataGroup_lo_hi_1961, dataGroup_lo_lo_1961};
  wire [1023:0] dataGroup_hi_1961 = {dataGroup_hi_hi_1961, dataGroup_hi_lo_1961};
  wire [31:0]   dataGroup_1_101 = dataGroup_lo_1961[319:288];
  wire [1023:0] dataGroup_lo_1962 = {dataGroup_lo_hi_1962, dataGroup_lo_lo_1962};
  wire [1023:0] dataGroup_hi_1962 = {dataGroup_hi_hi_1962, dataGroup_hi_lo_1962};
  wire [31:0]   dataGroup_2_101 = dataGroup_lo_1962[575:544];
  wire [1023:0] dataGroup_lo_1963 = {dataGroup_lo_hi_1963, dataGroup_lo_lo_1963};
  wire [1023:0] dataGroup_hi_1963 = {dataGroup_hi_hi_1963, dataGroup_hi_lo_1963};
  wire [31:0]   dataGroup_3_101 = dataGroup_lo_1963[831:800];
  wire [1023:0] dataGroup_lo_1964 = {dataGroup_lo_hi_1964, dataGroup_lo_lo_1964};
  wire [1023:0] dataGroup_hi_1964 = {dataGroup_hi_hi_1964, dataGroup_hi_lo_1964};
  wire [31:0]   dataGroup_4_101 = dataGroup_hi_1964[63:32];
  wire [1023:0] dataGroup_lo_1965 = {dataGroup_lo_hi_1965, dataGroup_lo_lo_1965};
  wire [1023:0] dataGroup_hi_1965 = {dataGroup_hi_hi_1965, dataGroup_hi_lo_1965};
  wire [31:0]   dataGroup_5_101 = dataGroup_hi_1965[319:288];
  wire [1023:0] dataGroup_lo_1966 = {dataGroup_lo_hi_1966, dataGroup_lo_lo_1966};
  wire [1023:0] dataGroup_hi_1966 = {dataGroup_hi_hi_1966, dataGroup_hi_lo_1966};
  wire [31:0]   dataGroup_6_101 = dataGroup_hi_1966[575:544];
  wire [1023:0] dataGroup_lo_1967 = {dataGroup_lo_hi_1967, dataGroup_lo_lo_1967};
  wire [1023:0] dataGroup_hi_1967 = {dataGroup_hi_hi_1967, dataGroup_hi_lo_1967};
  wire [31:0]   dataGroup_7_101 = dataGroup_hi_1967[831:800];
  wire [63:0]   res_lo_lo_101 = {dataGroup_1_101, dataGroup_0_101};
  wire [63:0]   res_lo_hi_101 = {dataGroup_3_101, dataGroup_2_101};
  wire [127:0]  res_lo_101 = {res_lo_hi_101, res_lo_lo_101};
  wire [63:0]   res_hi_lo_101 = {dataGroup_5_101, dataGroup_4_101};
  wire [63:0]   res_hi_hi_101 = {dataGroup_7_101, dataGroup_6_101};
  wire [127:0]  res_hi_101 = {res_hi_hi_101, res_hi_lo_101};
  wire [255:0]  res_185 = {res_hi_101, res_lo_101};
  wire [1023:0] dataGroup_lo_1968 = {dataGroup_lo_hi_1968, dataGroup_lo_lo_1968};
  wire [1023:0] dataGroup_hi_1968 = {dataGroup_hi_hi_1968, dataGroup_hi_lo_1968};
  wire [31:0]   dataGroup_0_102 = dataGroup_lo_1968[95:64];
  wire [1023:0] dataGroup_lo_1969 = {dataGroup_lo_hi_1969, dataGroup_lo_lo_1969};
  wire [1023:0] dataGroup_hi_1969 = {dataGroup_hi_hi_1969, dataGroup_hi_lo_1969};
  wire [31:0]   dataGroup_1_102 = dataGroup_lo_1969[351:320];
  wire [1023:0] dataGroup_lo_1970 = {dataGroup_lo_hi_1970, dataGroup_lo_lo_1970};
  wire [1023:0] dataGroup_hi_1970 = {dataGroup_hi_hi_1970, dataGroup_hi_lo_1970};
  wire [31:0]   dataGroup_2_102 = dataGroup_lo_1970[607:576];
  wire [1023:0] dataGroup_lo_1971 = {dataGroup_lo_hi_1971, dataGroup_lo_lo_1971};
  wire [1023:0] dataGroup_hi_1971 = {dataGroup_hi_hi_1971, dataGroup_hi_lo_1971};
  wire [31:0]   dataGroup_3_102 = dataGroup_lo_1971[863:832];
  wire [1023:0] dataGroup_lo_1972 = {dataGroup_lo_hi_1972, dataGroup_lo_lo_1972};
  wire [1023:0] dataGroup_hi_1972 = {dataGroup_hi_hi_1972, dataGroup_hi_lo_1972};
  wire [31:0]   dataGroup_4_102 = dataGroup_hi_1972[95:64];
  wire [1023:0] dataGroup_lo_1973 = {dataGroup_lo_hi_1973, dataGroup_lo_lo_1973};
  wire [1023:0] dataGroup_hi_1973 = {dataGroup_hi_hi_1973, dataGroup_hi_lo_1973};
  wire [31:0]   dataGroup_5_102 = dataGroup_hi_1973[351:320];
  wire [1023:0] dataGroup_lo_1974 = {dataGroup_lo_hi_1974, dataGroup_lo_lo_1974};
  wire [1023:0] dataGroup_hi_1974 = {dataGroup_hi_hi_1974, dataGroup_hi_lo_1974};
  wire [31:0]   dataGroup_6_102 = dataGroup_hi_1974[607:576];
  wire [1023:0] dataGroup_lo_1975 = {dataGroup_lo_hi_1975, dataGroup_lo_lo_1975};
  wire [1023:0] dataGroup_hi_1975 = {dataGroup_hi_hi_1975, dataGroup_hi_lo_1975};
  wire [31:0]   dataGroup_7_102 = dataGroup_hi_1975[863:832];
  wire [63:0]   res_lo_lo_102 = {dataGroup_1_102, dataGroup_0_102};
  wire [63:0]   res_lo_hi_102 = {dataGroup_3_102, dataGroup_2_102};
  wire [127:0]  res_lo_102 = {res_lo_hi_102, res_lo_lo_102};
  wire [63:0]   res_hi_lo_102 = {dataGroup_5_102, dataGroup_4_102};
  wire [63:0]   res_hi_hi_102 = {dataGroup_7_102, dataGroup_6_102};
  wire [127:0]  res_hi_102 = {res_hi_hi_102, res_hi_lo_102};
  wire [255:0]  res_186 = {res_hi_102, res_lo_102};
  wire [1023:0] dataGroup_lo_1976 = {dataGroup_lo_hi_1976, dataGroup_lo_lo_1976};
  wire [1023:0] dataGroup_hi_1976 = {dataGroup_hi_hi_1976, dataGroup_hi_lo_1976};
  wire [31:0]   dataGroup_0_103 = dataGroup_lo_1976[127:96];
  wire [1023:0] dataGroup_lo_1977 = {dataGroup_lo_hi_1977, dataGroup_lo_lo_1977};
  wire [1023:0] dataGroup_hi_1977 = {dataGroup_hi_hi_1977, dataGroup_hi_lo_1977};
  wire [31:0]   dataGroup_1_103 = dataGroup_lo_1977[383:352];
  wire [1023:0] dataGroup_lo_1978 = {dataGroup_lo_hi_1978, dataGroup_lo_lo_1978};
  wire [1023:0] dataGroup_hi_1978 = {dataGroup_hi_hi_1978, dataGroup_hi_lo_1978};
  wire [31:0]   dataGroup_2_103 = dataGroup_lo_1978[639:608];
  wire [1023:0] dataGroup_lo_1979 = {dataGroup_lo_hi_1979, dataGroup_lo_lo_1979};
  wire [1023:0] dataGroup_hi_1979 = {dataGroup_hi_hi_1979, dataGroup_hi_lo_1979};
  wire [31:0]   dataGroup_3_103 = dataGroup_lo_1979[895:864];
  wire [1023:0] dataGroup_lo_1980 = {dataGroup_lo_hi_1980, dataGroup_lo_lo_1980};
  wire [1023:0] dataGroup_hi_1980 = {dataGroup_hi_hi_1980, dataGroup_hi_lo_1980};
  wire [31:0]   dataGroup_4_103 = dataGroup_hi_1980[127:96];
  wire [1023:0] dataGroup_lo_1981 = {dataGroup_lo_hi_1981, dataGroup_lo_lo_1981};
  wire [1023:0] dataGroup_hi_1981 = {dataGroup_hi_hi_1981, dataGroup_hi_lo_1981};
  wire [31:0]   dataGroup_5_103 = dataGroup_hi_1981[383:352];
  wire [1023:0] dataGroup_lo_1982 = {dataGroup_lo_hi_1982, dataGroup_lo_lo_1982};
  wire [1023:0] dataGroup_hi_1982 = {dataGroup_hi_hi_1982, dataGroup_hi_lo_1982};
  wire [31:0]   dataGroup_6_103 = dataGroup_hi_1982[639:608];
  wire [1023:0] dataGroup_lo_1983 = {dataGroup_lo_hi_1983, dataGroup_lo_lo_1983};
  wire [1023:0] dataGroup_hi_1983 = {dataGroup_hi_hi_1983, dataGroup_hi_lo_1983};
  wire [31:0]   dataGroup_7_103 = dataGroup_hi_1983[895:864];
  wire [63:0]   res_lo_lo_103 = {dataGroup_1_103, dataGroup_0_103};
  wire [63:0]   res_lo_hi_103 = {dataGroup_3_103, dataGroup_2_103};
  wire [127:0]  res_lo_103 = {res_lo_hi_103, res_lo_lo_103};
  wire [63:0]   res_hi_lo_103 = {dataGroup_5_103, dataGroup_4_103};
  wire [63:0]   res_hi_hi_103 = {dataGroup_7_103, dataGroup_6_103};
  wire [127:0]  res_hi_103 = {res_hi_hi_103, res_hi_lo_103};
  wire [255:0]  res_187 = {res_hi_103, res_lo_103};
  wire [1023:0] dataGroup_lo_1984 = {dataGroup_lo_hi_1984, dataGroup_lo_lo_1984};
  wire [1023:0] dataGroup_hi_1984 = {dataGroup_hi_hi_1984, dataGroup_hi_lo_1984};
  wire [31:0]   dataGroup_0_104 = dataGroup_lo_1984[159:128];
  wire [1023:0] dataGroup_lo_1985 = {dataGroup_lo_hi_1985, dataGroup_lo_lo_1985};
  wire [1023:0] dataGroup_hi_1985 = {dataGroup_hi_hi_1985, dataGroup_hi_lo_1985};
  wire [31:0]   dataGroup_1_104 = dataGroup_lo_1985[415:384];
  wire [1023:0] dataGroup_lo_1986 = {dataGroup_lo_hi_1986, dataGroup_lo_lo_1986};
  wire [1023:0] dataGroup_hi_1986 = {dataGroup_hi_hi_1986, dataGroup_hi_lo_1986};
  wire [31:0]   dataGroup_2_104 = dataGroup_lo_1986[671:640];
  wire [1023:0] dataGroup_lo_1987 = {dataGroup_lo_hi_1987, dataGroup_lo_lo_1987};
  wire [1023:0] dataGroup_hi_1987 = {dataGroup_hi_hi_1987, dataGroup_hi_lo_1987};
  wire [31:0]   dataGroup_3_104 = dataGroup_lo_1987[927:896];
  wire [1023:0] dataGroup_lo_1988 = {dataGroup_lo_hi_1988, dataGroup_lo_lo_1988};
  wire [1023:0] dataGroup_hi_1988 = {dataGroup_hi_hi_1988, dataGroup_hi_lo_1988};
  wire [31:0]   dataGroup_4_104 = dataGroup_hi_1988[159:128];
  wire [1023:0] dataGroup_lo_1989 = {dataGroup_lo_hi_1989, dataGroup_lo_lo_1989};
  wire [1023:0] dataGroup_hi_1989 = {dataGroup_hi_hi_1989, dataGroup_hi_lo_1989};
  wire [31:0]   dataGroup_5_104 = dataGroup_hi_1989[415:384];
  wire [1023:0] dataGroup_lo_1990 = {dataGroup_lo_hi_1990, dataGroup_lo_lo_1990};
  wire [1023:0] dataGroup_hi_1990 = {dataGroup_hi_hi_1990, dataGroup_hi_lo_1990};
  wire [31:0]   dataGroup_6_104 = dataGroup_hi_1990[671:640];
  wire [1023:0] dataGroup_lo_1991 = {dataGroup_lo_hi_1991, dataGroup_lo_lo_1991};
  wire [1023:0] dataGroup_hi_1991 = {dataGroup_hi_hi_1991, dataGroup_hi_lo_1991};
  wire [31:0]   dataGroup_7_104 = dataGroup_hi_1991[927:896];
  wire [63:0]   res_lo_lo_104 = {dataGroup_1_104, dataGroup_0_104};
  wire [63:0]   res_lo_hi_104 = {dataGroup_3_104, dataGroup_2_104};
  wire [127:0]  res_lo_104 = {res_lo_hi_104, res_lo_lo_104};
  wire [63:0]   res_hi_lo_104 = {dataGroup_5_104, dataGroup_4_104};
  wire [63:0]   res_hi_hi_104 = {dataGroup_7_104, dataGroup_6_104};
  wire [127:0]  res_hi_104 = {res_hi_hi_104, res_hi_lo_104};
  wire [255:0]  res_188 = {res_hi_104, res_lo_104};
  wire [1023:0] dataGroup_lo_1992 = {dataGroup_lo_hi_1992, dataGroup_lo_lo_1992};
  wire [1023:0] dataGroup_hi_1992 = {dataGroup_hi_hi_1992, dataGroup_hi_lo_1992};
  wire [31:0]   dataGroup_0_105 = dataGroup_lo_1992[191:160];
  wire [1023:0] dataGroup_lo_1993 = {dataGroup_lo_hi_1993, dataGroup_lo_lo_1993};
  wire [1023:0] dataGroup_hi_1993 = {dataGroup_hi_hi_1993, dataGroup_hi_lo_1993};
  wire [31:0]   dataGroup_1_105 = dataGroup_lo_1993[447:416];
  wire [1023:0] dataGroup_lo_1994 = {dataGroup_lo_hi_1994, dataGroup_lo_lo_1994};
  wire [1023:0] dataGroup_hi_1994 = {dataGroup_hi_hi_1994, dataGroup_hi_lo_1994};
  wire [31:0]   dataGroup_2_105 = dataGroup_lo_1994[703:672];
  wire [1023:0] dataGroup_lo_1995 = {dataGroup_lo_hi_1995, dataGroup_lo_lo_1995};
  wire [1023:0] dataGroup_hi_1995 = {dataGroup_hi_hi_1995, dataGroup_hi_lo_1995};
  wire [31:0]   dataGroup_3_105 = dataGroup_lo_1995[959:928];
  wire [1023:0] dataGroup_lo_1996 = {dataGroup_lo_hi_1996, dataGroup_lo_lo_1996};
  wire [1023:0] dataGroup_hi_1996 = {dataGroup_hi_hi_1996, dataGroup_hi_lo_1996};
  wire [31:0]   dataGroup_4_105 = dataGroup_hi_1996[191:160];
  wire [1023:0] dataGroup_lo_1997 = {dataGroup_lo_hi_1997, dataGroup_lo_lo_1997};
  wire [1023:0] dataGroup_hi_1997 = {dataGroup_hi_hi_1997, dataGroup_hi_lo_1997};
  wire [31:0]   dataGroup_5_105 = dataGroup_hi_1997[447:416];
  wire [1023:0] dataGroup_lo_1998 = {dataGroup_lo_hi_1998, dataGroup_lo_lo_1998};
  wire [1023:0] dataGroup_hi_1998 = {dataGroup_hi_hi_1998, dataGroup_hi_lo_1998};
  wire [31:0]   dataGroup_6_105 = dataGroup_hi_1998[703:672];
  wire [1023:0] dataGroup_lo_1999 = {dataGroup_lo_hi_1999, dataGroup_lo_lo_1999};
  wire [1023:0] dataGroup_hi_1999 = {dataGroup_hi_hi_1999, dataGroup_hi_lo_1999};
  wire [31:0]   dataGroup_7_105 = dataGroup_hi_1999[959:928];
  wire [63:0]   res_lo_lo_105 = {dataGroup_1_105, dataGroup_0_105};
  wire [63:0]   res_lo_hi_105 = {dataGroup_3_105, dataGroup_2_105};
  wire [127:0]  res_lo_105 = {res_lo_hi_105, res_lo_lo_105};
  wire [63:0]   res_hi_lo_105 = {dataGroup_5_105, dataGroup_4_105};
  wire [63:0]   res_hi_hi_105 = {dataGroup_7_105, dataGroup_6_105};
  wire [127:0]  res_hi_105 = {res_hi_hi_105, res_hi_lo_105};
  wire [255:0]  res_189 = {res_hi_105, res_lo_105};
  wire [1023:0] dataGroup_lo_2000 = {dataGroup_lo_hi_2000, dataGroup_lo_lo_2000};
  wire [1023:0] dataGroup_hi_2000 = {dataGroup_hi_hi_2000, dataGroup_hi_lo_2000};
  wire [31:0]   dataGroup_0_106 = dataGroup_lo_2000[223:192];
  wire [1023:0] dataGroup_lo_2001 = {dataGroup_lo_hi_2001, dataGroup_lo_lo_2001};
  wire [1023:0] dataGroup_hi_2001 = {dataGroup_hi_hi_2001, dataGroup_hi_lo_2001};
  wire [31:0]   dataGroup_1_106 = dataGroup_lo_2001[479:448];
  wire [1023:0] dataGroup_lo_2002 = {dataGroup_lo_hi_2002, dataGroup_lo_lo_2002};
  wire [1023:0] dataGroup_hi_2002 = {dataGroup_hi_hi_2002, dataGroup_hi_lo_2002};
  wire [31:0]   dataGroup_2_106 = dataGroup_lo_2002[735:704];
  wire [1023:0] dataGroup_lo_2003 = {dataGroup_lo_hi_2003, dataGroup_lo_lo_2003};
  wire [1023:0] dataGroup_hi_2003 = {dataGroup_hi_hi_2003, dataGroup_hi_lo_2003};
  wire [31:0]   dataGroup_3_106 = dataGroup_lo_2003[991:960];
  wire [1023:0] dataGroup_lo_2004 = {dataGroup_lo_hi_2004, dataGroup_lo_lo_2004};
  wire [1023:0] dataGroup_hi_2004 = {dataGroup_hi_hi_2004, dataGroup_hi_lo_2004};
  wire [31:0]   dataGroup_4_106 = dataGroup_hi_2004[223:192];
  wire [1023:0] dataGroup_lo_2005 = {dataGroup_lo_hi_2005, dataGroup_lo_lo_2005};
  wire [1023:0] dataGroup_hi_2005 = {dataGroup_hi_hi_2005, dataGroup_hi_lo_2005};
  wire [31:0]   dataGroup_5_106 = dataGroup_hi_2005[479:448];
  wire [1023:0] dataGroup_lo_2006 = {dataGroup_lo_hi_2006, dataGroup_lo_lo_2006};
  wire [1023:0] dataGroup_hi_2006 = {dataGroup_hi_hi_2006, dataGroup_hi_lo_2006};
  wire [31:0]   dataGroup_6_106 = dataGroup_hi_2006[735:704];
  wire [1023:0] dataGroup_lo_2007 = {dataGroup_lo_hi_2007, dataGroup_lo_lo_2007};
  wire [1023:0] dataGroup_hi_2007 = {dataGroup_hi_hi_2007, dataGroup_hi_lo_2007};
  wire [31:0]   dataGroup_7_106 = dataGroup_hi_2007[991:960];
  wire [63:0]   res_lo_lo_106 = {dataGroup_1_106, dataGroup_0_106};
  wire [63:0]   res_lo_hi_106 = {dataGroup_3_106, dataGroup_2_106};
  wire [127:0]  res_lo_106 = {res_lo_hi_106, res_lo_lo_106};
  wire [63:0]   res_hi_lo_106 = {dataGroup_5_106, dataGroup_4_106};
  wire [63:0]   res_hi_hi_106 = {dataGroup_7_106, dataGroup_6_106};
  wire [127:0]  res_hi_106 = {res_hi_hi_106, res_hi_lo_106};
  wire [255:0]  res_190 = {res_hi_106, res_lo_106};
  wire [1023:0] dataGroup_lo_2008 = {dataGroup_lo_hi_2008, dataGroup_lo_lo_2008};
  wire [1023:0] dataGroup_hi_2008 = {dataGroup_hi_hi_2008, dataGroup_hi_lo_2008};
  wire [31:0]   dataGroup_0_107 = dataGroup_lo_2008[255:224];
  wire [1023:0] dataGroup_lo_2009 = {dataGroup_lo_hi_2009, dataGroup_lo_lo_2009};
  wire [1023:0] dataGroup_hi_2009 = {dataGroup_hi_hi_2009, dataGroup_hi_lo_2009};
  wire [31:0]   dataGroup_1_107 = dataGroup_lo_2009[511:480];
  wire [1023:0] dataGroup_lo_2010 = {dataGroup_lo_hi_2010, dataGroup_lo_lo_2010};
  wire [1023:0] dataGroup_hi_2010 = {dataGroup_hi_hi_2010, dataGroup_hi_lo_2010};
  wire [31:0]   dataGroup_2_107 = dataGroup_lo_2010[767:736];
  wire [1023:0] dataGroup_lo_2011 = {dataGroup_lo_hi_2011, dataGroup_lo_lo_2011};
  wire [1023:0] dataGroup_hi_2011 = {dataGroup_hi_hi_2011, dataGroup_hi_lo_2011};
  wire [31:0]   dataGroup_3_107 = dataGroup_lo_2011[1023:992];
  wire [1023:0] dataGroup_lo_2012 = {dataGroup_lo_hi_2012, dataGroup_lo_lo_2012};
  wire [1023:0] dataGroup_hi_2012 = {dataGroup_hi_hi_2012, dataGroup_hi_lo_2012};
  wire [31:0]   dataGroup_4_107 = dataGroup_hi_2012[255:224];
  wire [1023:0] dataGroup_lo_2013 = {dataGroup_lo_hi_2013, dataGroup_lo_lo_2013};
  wire [1023:0] dataGroup_hi_2013 = {dataGroup_hi_hi_2013, dataGroup_hi_lo_2013};
  wire [31:0]   dataGroup_5_107 = dataGroup_hi_2013[511:480];
  wire [1023:0] dataGroup_lo_2014 = {dataGroup_lo_hi_2014, dataGroup_lo_lo_2014};
  wire [1023:0] dataGroup_hi_2014 = {dataGroup_hi_hi_2014, dataGroup_hi_lo_2014};
  wire [31:0]   dataGroup_6_107 = dataGroup_hi_2014[767:736];
  wire [1023:0] dataGroup_lo_2015 = {dataGroup_lo_hi_2015, dataGroup_lo_lo_2015};
  wire [1023:0] dataGroup_hi_2015 = {dataGroup_hi_hi_2015, dataGroup_hi_lo_2015};
  wire [31:0]   dataGroup_7_107 = dataGroup_hi_2015[1023:992];
  wire [63:0]   res_lo_lo_107 = {dataGroup_1_107, dataGroup_0_107};
  wire [63:0]   res_lo_hi_107 = {dataGroup_3_107, dataGroup_2_107};
  wire [127:0]  res_lo_107 = {res_lo_hi_107, res_lo_lo_107};
  wire [63:0]   res_hi_lo_107 = {dataGroup_5_107, dataGroup_4_107};
  wire [63:0]   res_hi_hi_107 = {dataGroup_7_107, dataGroup_6_107};
  wire [127:0]  res_hi_107 = {res_hi_hi_107, res_hi_lo_107};
  wire [255:0]  res_191 = {res_hi_107, res_lo_107};
  wire [511:0]  lo_lo_23 = {res_185, res_184};
  wire [511:0]  lo_hi_23 = {res_187, res_186};
  wire [1023:0] lo_23 = {lo_hi_23, lo_lo_23};
  wire [511:0]  hi_lo_23 = {res_189, res_188};
  wire [511:0]  hi_hi_23 = {res_191, res_190};
  wire [1023:0] hi_23 = {hi_hi_23, hi_lo_23};
  wire [2047:0] regroupLoadData_2_7 = {hi_23, lo_23};
  wire          vrfWritePort_0_valid_0 = accessState_0 & writeReadyReg;
  wire [3:0]    vrfWritePort_0_bits_mask_0 = maskForGroup[3:0];
  wire [3:0]    vrfWritePort_1_bits_mask_0 = maskForGroup[7:4];
  wire [3:0]    vrfWritePort_2_bits_mask_0 = maskForGroup[11:8];
  wire [3:0]    vrfWritePort_3_bits_mask_0 = maskForGroup[15:12];
  wire [3:0]    vrfWritePort_4_bits_mask_0 = maskForGroup[19:16];
  wire [3:0]    vrfWritePort_5_bits_mask_0 = maskForGroup[23:20];
  wire [3:0]    vrfWritePort_6_bits_mask_0 = maskForGroup[27:24];
  wire [3:0]    vrfWritePort_7_bits_mask_0 = maskForGroup[31:28];
  wire [7:0]    _vrfWritePort_7_bits_data_T = 8'h1 << accessPtr;
  wire [31:0]   vrfWritePort_0_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[31:0] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[31:0] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[31:0] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[31:0] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[31:0] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[31:0] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[31:0] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[31:0] : 32'h0);
  wire [2:0]    vrfWritePort_0_bits_offset_0 = dataGroup[2:0];
  wire [2:0]    vrfWritePort_1_bits_offset_0 = dataGroup[2:0];
  wire [2:0]    vrfWritePort_2_bits_offset_0 = dataGroup[2:0];
  wire [2:0]    vrfWritePort_3_bits_offset_0 = dataGroup[2:0];
  wire [2:0]    vrfWritePort_4_bits_offset_0 = dataGroup[2:0];
  wire [2:0]    vrfWritePort_5_bits_offset_0 = dataGroup[2:0];
  wire [2:0]    vrfWritePort_6_bits_offset_0 = dataGroup[2:0];
  wire [2:0]    vrfWritePort_7_bits_offset_0 = dataGroup[2:0];
  wire [4:0]    _GEN_8 = {2'h0, accessPtr} * {1'h0, segmentInstructionIndexInterval} + {2'h0, dataGroup[5:3]};
  wire [4:0]    vrfWritePort_0_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_0 = ~(vrfWritePort_0_ready_0 & vrfWritePort_0_valid_0) & accessState_0;
  wire          vrfWritePort_1_valid_0 = accessState_1 & writeReadyReg;
  wire [31:0]   vrfWritePort_1_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[63:32] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[63:32] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[63:32] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[63:32] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[63:32] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[63:32] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[63:32] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[63:32] : 32'h0);
  wire [4:0]    vrfWritePort_1_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_1 = ~(vrfWritePort_1_ready_0 & vrfWritePort_1_valid_0) & accessState_1;
  wire          vrfWritePort_2_valid_0 = accessState_2 & writeReadyReg;
  wire [31:0]   vrfWritePort_2_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[95:64] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[95:64] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[95:64] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[95:64] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[95:64] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[95:64] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[95:64] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[95:64] : 32'h0);
  wire [4:0]    vrfWritePort_2_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_2 = ~(vrfWritePort_2_ready_0 & vrfWritePort_2_valid_0) & accessState_2;
  wire          vrfWritePort_3_valid_0 = accessState_3 & writeReadyReg;
  wire [31:0]   vrfWritePort_3_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[127:96] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[127:96] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[127:96] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[127:96] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[127:96] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[127:96] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[127:96] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[127:96] : 32'h0);
  wire [4:0]    vrfWritePort_3_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_3 = ~(vrfWritePort_3_ready_0 & vrfWritePort_3_valid_0) & accessState_3;
  wire          vrfWritePort_4_valid_0 = accessState_4 & writeReadyReg;
  wire [31:0]   vrfWritePort_4_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[159:128] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[159:128] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[159:128] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[159:128] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[159:128] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[159:128] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[159:128] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[159:128] : 32'h0);
  wire [4:0]    vrfWritePort_4_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_4 = ~(vrfWritePort_4_ready_0 & vrfWritePort_4_valid_0) & accessState_4;
  wire          vrfWritePort_5_valid_0 = accessState_5 & writeReadyReg;
  wire [31:0]   vrfWritePort_5_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[191:160] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[191:160] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[191:160] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[191:160] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[191:160] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[191:160] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[191:160] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[191:160] : 32'h0);
  wire [4:0]    vrfWritePort_5_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_5 = ~(vrfWritePort_5_ready_0 & vrfWritePort_5_valid_0) & accessState_5;
  wire          vrfWritePort_6_valid_0 = accessState_6 & writeReadyReg;
  wire [31:0]   vrfWritePort_6_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[223:192] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[223:192] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[223:192] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[223:192] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[223:192] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[223:192] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[223:192] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[223:192] : 32'h0);
  wire [4:0]    vrfWritePort_6_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_6 = ~(vrfWritePort_6_ready_0 & vrfWritePort_6_valid_0) & accessState_6;
  wire          vrfWritePort_7_valid_0 = accessState_7 & writeReadyReg;
  wire [31:0]   vrfWritePort_7_bits_data_0 =
    (_vrfWritePort_7_bits_data_T[0] ? accessData_0[255:224] : 32'h0) | (_vrfWritePort_7_bits_data_T[1] ? accessData_1[255:224] : 32'h0) | (_vrfWritePort_7_bits_data_T[2] ? accessData_2[255:224] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[3] ? accessData_3[255:224] : 32'h0) | (_vrfWritePort_7_bits_data_T[4] ? accessData_4[255:224] : 32'h0) | (_vrfWritePort_7_bits_data_T[5] ? accessData_5[255:224] : 32'h0)
    | (_vrfWritePort_7_bits_data_T[6] ? accessData_6[255:224] : 32'h0) | (_vrfWritePort_7_bits_data_T[7] ? accessData_7[255:224] : 32'h0);
  wire [4:0]    vrfWritePort_7_bits_vd_0 = lsuRequestReg_instructionInformation_vs3 + _GEN_8;
  assign accessStateUpdate_7 = ~(vrfWritePort_7_ready_0 & vrfWritePort_7_valid_0) & accessState_7;
  reg           sendStateReg_0;
  reg           sendStateReg_1;
  reg           sendStateReg_2;
  reg           sendStateReg_3;
  reg           sendStateReg_4;
  reg           sendStateReg_5;
  reg           sendStateReg_6;
  reg           sendStateReg_7;
  wire          lastCacheRequest = lastRequest & _lastCacheRequest_T;
  reg           lastCacheRequestReg;
  reg           lastCacheLineAckReg;
  wire          bufferClear = ~(memResponse_valid_0 | alignedDequeue_valid | bufferFull | ~writeStageReady);
  wire          _status_idle_output = lastCacheRequestReg & lastCacheLineAckReg & bufferClear & ~sendRequest;
  reg           idleNext;
  always @(posedge clock) begin
    if (reset) begin
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 12'h0;
      csrInterfaceReg_vStart <= 12'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      requestFireNext <= 1'h0;
      dataEEW <= 2'h0;
      maskReg <= 32'h0;
      needAmend <= 1'h0;
      lastMaskAmendReg <= 31'h0;
      maskGroupCounter <= 6'h0;
      maskCounterInGroup <= 2'h0;
      maskForGroup <= 32'h0;
      isLastMaskGroup <= 1'h0;
      accessData_0 <= 256'h0;
      accessData_1 <= 256'h0;
      accessData_2 <= 256'h0;
      accessData_3 <= 256'h0;
      accessData_4 <= 256'h0;
      accessData_5 <= 256'h0;
      accessData_6 <= 256'h0;
      accessData_7 <= 256'h0;
      accessPtr <= 3'h0;
      accessState_0 <= 1'h0;
      accessState_1 <= 1'h0;
      accessState_2 <= 1'h0;
      accessState_3 <= 1'h0;
      accessState_4 <= 1'h0;
      accessState_5 <= 1'h0;
      accessState_6 <= 1'h0;
      accessState_7 <= 1'h0;
      dataGroup <= 6'h0;
      dataBuffer_0 <= 256'h0;
      dataBuffer_1 <= 256'h0;
      dataBuffer_2 <= 256'h0;
      dataBuffer_3 <= 256'h0;
      dataBuffer_4 <= 256'h0;
      dataBuffer_5 <= 256'h0;
      dataBuffer_6 <= 256'h0;
      dataBuffer_7 <= 256'h0;
      bufferBaseCacheLineIndex <= 7'h0;
      cacheLineIndexInBuffer <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      lastWriteVrfIndexReg <= 14'h0;
      lastCacheNeedPush <= 1'h0;
      cacheLineNumberReg <= 14'h0;
      sendRequest <= 1'h0;
      writeReadyReg <= 1'h0;
      unalignedCacheLine_valid <= 1'h0;
      unalignedCacheLine_bits_data <= 256'h0;
      unalignedCacheLine_bits_index <= 7'h0;
      bufferFull <= 1'h0;
      waitForFirstDataGroup <= 1'h0;
      sendStateReg_0 <= 1'h0;
      sendStateReg_1 <= 1'h0;
      sendStateReg_2 <= 1'h0;
      sendStateReg_3 <= 1'h0;
      sendStateReg_4 <= 1'h0;
      sendStateReg_5 <= 1'h0;
      sendStateReg_6 <= 1'h0;
      sendStateReg_7 <= 1'h0;
      lastCacheRequestReg <= 1'h1;
      lastCacheLineAckReg <= 1'h1;
      idleNext <= 1'h1;
    end
    else begin
      automatic logic _GEN_9 = bufferDequeueFire | accessStateCheck & ~lastPtr;
      if (lsuRequest_valid) begin
        lsuRequestReg_instructionInformation_nf <= nfCorrection;
        lsuRequestReg_instructionInformation_mew <= ~invalidInstruction & lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataEEW <= lsuRequest_bits_instructionInformation_eew;
        needAmend <= |(csrInterface_vl[4:0]);
        lastMaskAmendReg <= lastMaskAmend;
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
        lastWriteVrfIndexReg <= lastWriteVrfIndex;
        lastCacheNeedPush <= lastCacheLineIndex == lastWriteVrfIndex;
        cacheLineNumberReg <= lastCacheLineIndex;
      end
      requestFireNext <= lsuRequest_valid;
      if (_maskSelect_valid_output | lsuRequest_valid) begin
        maskReg <= maskAmend;
        isLastMaskGroup <= lsuRequest_valid ? csrInterface_vl[11:5] == 7'h0 : {1'h0, _maskSelect_bits_output} == csrInterfaceReg_vl[11:5];
      end
      if (bufferDequeueFire & isLastDataGroup)
        maskGroupCounter <= nextMaskGroup;
      else if (lsuRequest_valid)
        maskGroupCounter <= 6'h0;
      if (lsuRequest_valid | bufferDequeueFire) begin
        maskCounterInGroup <= isLastDataGroup | lsuRequest_valid ? 2'h0 : nextMaskCount;
        waitForFirstDataGroup <= lsuRequest_valid;
      end
      if (bufferDequeueFire) begin
        automatic logic [7:0]    _GEN_10;
        automatic logic [2047:0] _GEN_11;
        _GEN_10 = 8'h1 << lsuRequestReg_instructionInformation_nf;
        _GEN_11 =
          (dataEEWOH[0]
             ? (_GEN_10[0] ? regroupLoadData_0_0 : 2048'h0) | (_GEN_10[1] ? regroupLoadData_0_1 : 2048'h0) | (_GEN_10[2] ? regroupLoadData_0_2 : 2048'h0) | (_GEN_10[3] ? regroupLoadData_0_3 : 2048'h0)
               | (_GEN_10[4] ? regroupLoadData_0_4 : 2048'h0) | (_GEN_10[5] ? regroupLoadData_0_5 : 2048'h0) | (_GEN_10[6] ? regroupLoadData_0_6 : 2048'h0) | (_GEN_10[7] ? regroupLoadData_0_7 : 2048'h0)
             : 2048'h0)
          | (dataEEWOH[1]
               ? (_GEN_10[0] ? regroupLoadData_1_0 : 2048'h0) | (_GEN_10[1] ? regroupLoadData_1_1 : 2048'h0) | (_GEN_10[2] ? regroupLoadData_1_2 : 2048'h0) | (_GEN_10[3] ? regroupLoadData_1_3 : 2048'h0)
                 | (_GEN_10[4] ? regroupLoadData_1_4 : 2048'h0) | (_GEN_10[5] ? regroupLoadData_1_5 : 2048'h0) | (_GEN_10[6] ? regroupLoadData_1_6 : 2048'h0) | (_GEN_10[7] ? regroupLoadData_1_7 : 2048'h0)
               : 2048'h0)
          | (dataEEWOH[2]
               ? (_GEN_10[0] ? regroupLoadData_2_0 : 2048'h0) | (_GEN_10[1] ? regroupLoadData_2_1 : 2048'h0) | (_GEN_10[2] ? regroupLoadData_2_2 : 2048'h0) | (_GEN_10[3] ? regroupLoadData_2_3 : 2048'h0)
                 | (_GEN_10[4] ? regroupLoadData_2_4 : 2048'h0) | (_GEN_10[5] ? regroupLoadData_2_5 : 2048'h0) | (_GEN_10[6] ? regroupLoadData_2_6 : 2048'h0) | (_GEN_10[7] ? regroupLoadData_2_7 : 2048'h0)
               : 2048'h0);
        maskForGroup <= maskForGroupWire;
        accessData_0 <= _GEN_11[255:0];
        accessData_1 <= _GEN_11[511:256];
        accessData_2 <= _GEN_11[767:512];
        accessData_3 <= _GEN_11[1023:768];
        accessData_4 <= _GEN_11[1279:1024];
        accessData_5 <= _GEN_11[1535:1280];
        accessData_6 <= _GEN_11[1791:1536];
        accessData_7 <= _GEN_11[2047:1792];
        dataGroup <= waitForFirstDataGroup ? 6'h0 : dataGroup + 6'h1;
        sendStateReg_0 <= initSendState_0;
        sendStateReg_1 <= initSendState_1;
        sendStateReg_2 <= initSendState_2;
        sendStateReg_3 <= initSendState_3;
        sendStateReg_4 <= initSendState_4;
        sendStateReg_5 <= initSendState_5;
        sendStateReg_6 <= initSendState_6;
        sendStateReg_7 <= initSendState_7;
      end
      if (_GEN_9)
        accessPtr <= bufferDequeueFire ? lsuRequestReg_instructionInformation_nf : accessPtr - 3'h1;
      accessState_0 <= _GEN_9 ? (bufferDequeueFire ? initSendState_0 : sendStateReg_0) : accessStateUpdate_0;
      accessState_1 <= _GEN_9 ? (bufferDequeueFire ? initSendState_1 : sendStateReg_1) : accessStateUpdate_1;
      accessState_2 <= _GEN_9 ? (bufferDequeueFire ? initSendState_2 : sendStateReg_2) : accessStateUpdate_2;
      accessState_3 <= _GEN_9 ? (bufferDequeueFire ? initSendState_3 : sendStateReg_3) : accessStateUpdate_3;
      accessState_4 <= _GEN_9 ? (bufferDequeueFire ? initSendState_4 : sendStateReg_4) : accessStateUpdate_4;
      accessState_5 <= _GEN_9 ? (bufferDequeueFire ? initSendState_5 : sendStateReg_5) : accessStateUpdate_5;
      accessState_6 <= _GEN_9 ? (bufferDequeueFire ? initSendState_6 : sendStateReg_6) : accessStateUpdate_6;
      accessState_7 <= _GEN_9 ? (bufferDequeueFire ? initSendState_7 : sendStateReg_7) : accessStateUpdate_7;
      if (bufferEnqueueSelect[0])
        dataBuffer_0 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[1])
        dataBuffer_1 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[2])
        dataBuffer_2 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[3])
        dataBuffer_3 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[4])
        dataBuffer_4 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[5])
        dataBuffer_5 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[6])
        dataBuffer_6 <= alignedDequeue_bits_data;
      if (bufferEnqueueSelect[7])
        dataBuffer_7 <= alignedDequeue_bits_data;
      if (_bufferTailFire_T & cacheLineIndexInBuffer == 3'h0)
        bufferBaseCacheLineIndex <= alignedDequeue_bits_index;
      if (_bufferTailFire_T | bufferDequeueFire)
        cacheLineIndexInBuffer <= bufferDequeueFire ? 3'h0 : cacheLineIndexInBuffer + 3'h1;
      if (validInstruction | _lastCacheRequest_T & lastRequest)
        sendRequest <= lsuRequest_valid & (|csrInterface_vl);
      writeReadyReg <= ~lsuRequest_valid;
      if (unalignedEnqueueFire ^ _bufferTailFire_T | lsuRequest_valid)
        unalignedCacheLine_valid <= unalignedEnqueueFire;
      if (unalignedEnqueueFire) begin
        unalignedCacheLine_bits_data <= memResponse_bits_data_0;
        unalignedCacheLine_bits_index <= nextIndex;
      end
      if (bufferTailFire | bufferDequeueFire)
        bufferFull <= ~bufferDequeueFire;
      if (lastCacheRequest | validInstruction)
        lastCacheRequestReg <= lastCacheRequest;
      if (anyLastCacheLineAck | validInstruction)
        lastCacheLineAckReg <= anyLastCacheLineAck;
      idleNext <= _status_idle_output;
    end
    invalidInstructionNext <= invalidInstruction & lsuRequest_valid;
    if (_lastCacheRequest_T | lsuRequest_valid)
      cacheLineIndex <= lsuRequest_valid ? 7'h0 : nextCacheLineIndex;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:145];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [7:0] i = 8'h0; i < 8'h92; i += 8'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        lsuRequestReg_instructionInformation_nf = _RANDOM[8'h0][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[8'h0][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[8'h0][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[8'h0][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[8'h0][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[8'h0][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[8'h0][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[8'h0][19];
        lsuRequestReg_rs1Data = {_RANDOM[8'h0][31:20], _RANDOM[8'h1][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[8'h1][31:20], _RANDOM[8'h2][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[8'h2][22:20];
        csrInterfaceReg_vl = {_RANDOM[8'h2][31:23], _RANDOM[8'h3][2:0]};
        csrInterfaceReg_vStart = _RANDOM[8'h3][14:3];
        csrInterfaceReg_vlmul = _RANDOM[8'h3][17:15];
        csrInterfaceReg_vSew = _RANDOM[8'h3][19:18];
        csrInterfaceReg_vxrm = _RANDOM[8'h3][21:20];
        csrInterfaceReg_vta = _RANDOM[8'h3][22];
        csrInterfaceReg_vma = _RANDOM[8'h3][23];
        requestFireNext = _RANDOM[8'h3][24];
        dataEEW = _RANDOM[8'h3][26:25];
        maskReg = {_RANDOM[8'h3][31:27], _RANDOM[8'h4][26:0]};
        needAmend = _RANDOM[8'h4][27];
        lastMaskAmendReg = {_RANDOM[8'h4][31:28], _RANDOM[8'h5][26:0]};
        maskGroupCounter = {_RANDOM[8'h5][31:27], _RANDOM[8'h6][0]};
        maskCounterInGroup = _RANDOM[8'h6][2:1];
        maskForGroup = {_RANDOM[8'h6][31:3], _RANDOM[8'h7][2:0]};
        isLastMaskGroup = _RANDOM[8'h7][3];
        accessData_0 = {_RANDOM[8'h7][31:4], _RANDOM[8'h8], _RANDOM[8'h9], _RANDOM[8'hA], _RANDOM[8'hB], _RANDOM[8'hC], _RANDOM[8'hD], _RANDOM[8'hE], _RANDOM[8'hF][3:0]};
        accessData_1 = {_RANDOM[8'hF][31:4], _RANDOM[8'h10], _RANDOM[8'h11], _RANDOM[8'h12], _RANDOM[8'h13], _RANDOM[8'h14], _RANDOM[8'h15], _RANDOM[8'h16], _RANDOM[8'h17][3:0]};
        accessData_2 = {_RANDOM[8'h17][31:4], _RANDOM[8'h18], _RANDOM[8'h19], _RANDOM[8'h1A], _RANDOM[8'h1B], _RANDOM[8'h1C], _RANDOM[8'h1D], _RANDOM[8'h1E], _RANDOM[8'h1F][3:0]};
        accessData_3 = {_RANDOM[8'h1F][31:4], _RANDOM[8'h20], _RANDOM[8'h21], _RANDOM[8'h22], _RANDOM[8'h23], _RANDOM[8'h24], _RANDOM[8'h25], _RANDOM[8'h26], _RANDOM[8'h27][3:0]};
        accessData_4 = {_RANDOM[8'h27][31:4], _RANDOM[8'h28], _RANDOM[8'h29], _RANDOM[8'h2A], _RANDOM[8'h2B], _RANDOM[8'h2C], _RANDOM[8'h2D], _RANDOM[8'h2E], _RANDOM[8'h2F][3:0]};
        accessData_5 = {_RANDOM[8'h2F][31:4], _RANDOM[8'h30], _RANDOM[8'h31], _RANDOM[8'h32], _RANDOM[8'h33], _RANDOM[8'h34], _RANDOM[8'h35], _RANDOM[8'h36], _RANDOM[8'h37][3:0]};
        accessData_6 = {_RANDOM[8'h37][31:4], _RANDOM[8'h38], _RANDOM[8'h39], _RANDOM[8'h3A], _RANDOM[8'h3B], _RANDOM[8'h3C], _RANDOM[8'h3D], _RANDOM[8'h3E], _RANDOM[8'h3F][3:0]};
        accessData_7 = {_RANDOM[8'h3F][31:4], _RANDOM[8'h40], _RANDOM[8'h41], _RANDOM[8'h42], _RANDOM[8'h43], _RANDOM[8'h44], _RANDOM[8'h45], _RANDOM[8'h46], _RANDOM[8'h47][3:0]};
        accessPtr = _RANDOM[8'h47][6:4];
        accessState_0 = _RANDOM[8'h47][7];
        accessState_1 = _RANDOM[8'h47][8];
        accessState_2 = _RANDOM[8'h47][9];
        accessState_3 = _RANDOM[8'h47][10];
        accessState_4 = _RANDOM[8'h47][11];
        accessState_5 = _RANDOM[8'h47][12];
        accessState_6 = _RANDOM[8'h47][13];
        accessState_7 = _RANDOM[8'h47][14];
        dataGroup = _RANDOM[8'h47][20:15];
        dataBuffer_0 = {_RANDOM[8'h47][31:21], _RANDOM[8'h48], _RANDOM[8'h49], _RANDOM[8'h4A], _RANDOM[8'h4B], _RANDOM[8'h4C], _RANDOM[8'h4D], _RANDOM[8'h4E], _RANDOM[8'h4F][20:0]};
        dataBuffer_1 = {_RANDOM[8'h4F][31:21], _RANDOM[8'h50], _RANDOM[8'h51], _RANDOM[8'h52], _RANDOM[8'h53], _RANDOM[8'h54], _RANDOM[8'h55], _RANDOM[8'h56], _RANDOM[8'h57][20:0]};
        dataBuffer_2 = {_RANDOM[8'h57][31:21], _RANDOM[8'h58], _RANDOM[8'h59], _RANDOM[8'h5A], _RANDOM[8'h5B], _RANDOM[8'h5C], _RANDOM[8'h5D], _RANDOM[8'h5E], _RANDOM[8'h5F][20:0]};
        dataBuffer_3 = {_RANDOM[8'h5F][31:21], _RANDOM[8'h60], _RANDOM[8'h61], _RANDOM[8'h62], _RANDOM[8'h63], _RANDOM[8'h64], _RANDOM[8'h65], _RANDOM[8'h66], _RANDOM[8'h67][20:0]};
        dataBuffer_4 = {_RANDOM[8'h67][31:21], _RANDOM[8'h68], _RANDOM[8'h69], _RANDOM[8'h6A], _RANDOM[8'h6B], _RANDOM[8'h6C], _RANDOM[8'h6D], _RANDOM[8'h6E], _RANDOM[8'h6F][20:0]};
        dataBuffer_5 = {_RANDOM[8'h6F][31:21], _RANDOM[8'h70], _RANDOM[8'h71], _RANDOM[8'h72], _RANDOM[8'h73], _RANDOM[8'h74], _RANDOM[8'h75], _RANDOM[8'h76], _RANDOM[8'h77][20:0]};
        dataBuffer_6 = {_RANDOM[8'h77][31:21], _RANDOM[8'h78], _RANDOM[8'h79], _RANDOM[8'h7A], _RANDOM[8'h7B], _RANDOM[8'h7C], _RANDOM[8'h7D], _RANDOM[8'h7E], _RANDOM[8'h7F][20:0]};
        dataBuffer_7 = {_RANDOM[8'h7F][31:21], _RANDOM[8'h80], _RANDOM[8'h81], _RANDOM[8'h82], _RANDOM[8'h83], _RANDOM[8'h84], _RANDOM[8'h85], _RANDOM[8'h86], _RANDOM[8'h87][20:0]};
        bufferBaseCacheLineIndex = _RANDOM[8'h87][27:21];
        cacheLineIndexInBuffer = _RANDOM[8'h87][30:28];
        invalidInstructionNext = _RANDOM[8'h87][31];
        segmentInstructionIndexInterval = _RANDOM[8'h88][3:0];
        lastWriteVrfIndexReg = _RANDOM[8'h88][17:4];
        lastCacheNeedPush = _RANDOM[8'h88][18];
        cacheLineNumberReg = {_RANDOM[8'h88][31:19], _RANDOM[8'h89][0]};
        cacheLineIndex = _RANDOM[8'h89][7:1];
        sendRequest = _RANDOM[8'h89][8];
        writeReadyReg = _RANDOM[8'h89][9];
        unalignedCacheLine_valid = _RANDOM[8'h89][10];
        unalignedCacheLine_bits_data = {_RANDOM[8'h89][31:11], _RANDOM[8'h8A], _RANDOM[8'h8B], _RANDOM[8'h8C], _RANDOM[8'h8D], _RANDOM[8'h8E], _RANDOM[8'h8F], _RANDOM[8'h90], _RANDOM[8'h91][10:0]};
        unalignedCacheLine_bits_index = _RANDOM[8'h91][17:11];
        bufferFull = _RANDOM[8'h91][18];
        waitForFirstDataGroup = _RANDOM[8'h91][19];
        sendStateReg_0 = _RANDOM[8'h91][20];
        sendStateReg_1 = _RANDOM[8'h91][21];
        sendStateReg_2 = _RANDOM[8'h91][22];
        sendStateReg_3 = _RANDOM[8'h91][23];
        sendStateReg_4 = _RANDOM[8'h91][24];
        sendStateReg_5 = _RANDOM[8'h91][25];
        sendStateReg_6 = _RANDOM[8'h91][26];
        sendStateReg_7 = _RANDOM[8'h91][27];
        lastCacheRequestReg = _RANDOM[8'h91][28];
        lastCacheLineAckReg = _RANDOM[8'h91][29];
        idleNext = _RANDOM[8'h91][30];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign maskSelect_valid = _maskSelect_valid_output;
  assign maskSelect_bits = _maskSelect_bits_output;
  assign memRequest_valid = memRequest_valid_0;
  assign memRequest_bits_src = memRequest_bits_src_0;
  assign memRequest_bits_address = memRequest_bits_address_0;
  assign memResponse_ready = memResponse_ready_0;
  assign status_idle = _status_idle_output;
  assign status_last = ~idleNext & _status_idle_output | invalidInstructionNext;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_changeMaskGroup = _maskSelect_valid_output & ~lsuRequest_valid;
  assign status_startAddress = requestAddress;
  assign status_endAddress = {lsuRequestReg_rs1Data[31:5] + {13'h0, cacheLineNumberReg}, 5'h0};
  assign vrfWritePort_0_valid = vrfWritePort_0_valid_0;
  assign vrfWritePort_0_bits_vd = vrfWritePort_0_bits_vd_0;
  assign vrfWritePort_0_bits_offset = vrfWritePort_0_bits_offset_0;
  assign vrfWritePort_0_bits_mask = vrfWritePort_0_bits_mask_0;
  assign vrfWritePort_0_bits_data = vrfWritePort_0_bits_data_0;
  assign vrfWritePort_0_bits_instructionIndex = vrfWritePort_0_bits_instructionIndex_0;
  assign vrfWritePort_1_valid = vrfWritePort_1_valid_0;
  assign vrfWritePort_1_bits_vd = vrfWritePort_1_bits_vd_0;
  assign vrfWritePort_1_bits_offset = vrfWritePort_1_bits_offset_0;
  assign vrfWritePort_1_bits_mask = vrfWritePort_1_bits_mask_0;
  assign vrfWritePort_1_bits_data = vrfWritePort_1_bits_data_0;
  assign vrfWritePort_1_bits_instructionIndex = vrfWritePort_1_bits_instructionIndex_0;
  assign vrfWritePort_2_valid = vrfWritePort_2_valid_0;
  assign vrfWritePort_2_bits_vd = vrfWritePort_2_bits_vd_0;
  assign vrfWritePort_2_bits_offset = vrfWritePort_2_bits_offset_0;
  assign vrfWritePort_2_bits_mask = vrfWritePort_2_bits_mask_0;
  assign vrfWritePort_2_bits_data = vrfWritePort_2_bits_data_0;
  assign vrfWritePort_2_bits_instructionIndex = vrfWritePort_2_bits_instructionIndex_0;
  assign vrfWritePort_3_valid = vrfWritePort_3_valid_0;
  assign vrfWritePort_3_bits_vd = vrfWritePort_3_bits_vd_0;
  assign vrfWritePort_3_bits_offset = vrfWritePort_3_bits_offset_0;
  assign vrfWritePort_3_bits_mask = vrfWritePort_3_bits_mask_0;
  assign vrfWritePort_3_bits_data = vrfWritePort_3_bits_data_0;
  assign vrfWritePort_3_bits_instructionIndex = vrfWritePort_3_bits_instructionIndex_0;
  assign vrfWritePort_4_valid = vrfWritePort_4_valid_0;
  assign vrfWritePort_4_bits_vd = vrfWritePort_4_bits_vd_0;
  assign vrfWritePort_4_bits_offset = vrfWritePort_4_bits_offset_0;
  assign vrfWritePort_4_bits_mask = vrfWritePort_4_bits_mask_0;
  assign vrfWritePort_4_bits_data = vrfWritePort_4_bits_data_0;
  assign vrfWritePort_4_bits_instructionIndex = vrfWritePort_4_bits_instructionIndex_0;
  assign vrfWritePort_5_valid = vrfWritePort_5_valid_0;
  assign vrfWritePort_5_bits_vd = vrfWritePort_5_bits_vd_0;
  assign vrfWritePort_5_bits_offset = vrfWritePort_5_bits_offset_0;
  assign vrfWritePort_5_bits_mask = vrfWritePort_5_bits_mask_0;
  assign vrfWritePort_5_bits_data = vrfWritePort_5_bits_data_0;
  assign vrfWritePort_5_bits_instructionIndex = vrfWritePort_5_bits_instructionIndex_0;
  assign vrfWritePort_6_valid = vrfWritePort_6_valid_0;
  assign vrfWritePort_6_bits_vd = vrfWritePort_6_bits_vd_0;
  assign vrfWritePort_6_bits_offset = vrfWritePort_6_bits_offset_0;
  assign vrfWritePort_6_bits_mask = vrfWritePort_6_bits_mask_0;
  assign vrfWritePort_6_bits_data = vrfWritePort_6_bits_data_0;
  assign vrfWritePort_6_bits_instructionIndex = vrfWritePort_6_bits_instructionIndex_0;
  assign vrfWritePort_7_valid = vrfWritePort_7_valid_0;
  assign vrfWritePort_7_bits_vd = vrfWritePort_7_bits_vd_0;
  assign vrfWritePort_7_bits_offset = vrfWritePort_7_bits_offset_0;
  assign vrfWritePort_7_bits_mask = vrfWritePort_7_bits_mask_0;
  assign vrfWritePort_7_bits_data = vrfWritePort_7_bits_data_0;
  assign vrfWritePort_7_bits_instructionIndex = vrfWritePort_7_bits_instructionIndex_0;
endmodule

