module LanePopCount(
  input  [31:0] src,
  output [31:0] resp
);

  assign resp =
    {26'h0,
     {1'h0,
      {1'h0, {1'h0, {1'h0, {1'h0, src[0]} + {1'h0, src[1]}} + {1'h0, {1'h0, src[2]} + {1'h0, src[3]}}} + {1'h0, {1'h0, {1'h0, src[4]} + {1'h0, src[5]}} + {1'h0, {1'h0, src[6]} + {1'h0, src[7]}}}}
        + {1'h0, {1'h0, {1'h0, {1'h0, src[8]} + {1'h0, src[9]}} + {1'h0, {1'h0, src[10]} + {1'h0, src[11]}}} + {1'h0, {1'h0, {1'h0, src[12]} + {1'h0, src[13]}} + {1'h0, {1'h0, src[14]} + {1'h0, src[15]}}}}}
       + {1'h0,
          {1'h0, {1'h0, {1'h0, {1'h0, src[16]} + {1'h0, src[17]}} + {1'h0, {1'h0, src[18]} + {1'h0, src[19]}}} + {1'h0, {1'h0, {1'h0, src[20]} + {1'h0, src[21]}} + {1'h0, {1'h0, src[22]} + {1'h0, src[23]}}}}
            + {1'h0, {1'h0, {1'h0, {1'h0, src[24]} + {1'h0, src[25]}} + {1'h0, {1'h0, src[26]} + {1'h0, src[27]}}} + {1'h0, {1'h0, {1'h0, src[28]} + {1'h0, src[29]}} + {1'h0, {1'h0, src[30]} + {1'h0, src[31]}}}}}};
endmodule

