
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module Lane(
  input         clock,
                reset,
  input  [1:0]  laneIndex,
  input         readBusPort_0_enq_valid,
  input  [31:0] readBusPort_0_enq_bits_data,
  output        readBusPort_0_enqRelease,
                readBusPort_0_deq_valid,
  output [31:0] readBusPort_0_deq_bits_data,
  input         readBusPort_0_deqRelease,
                readBusPort_1_enq_valid,
  input  [31:0] readBusPort_1_enq_bits_data,
  output        readBusPort_1_enqRelease,
                readBusPort_1_deq_valid,
  output [31:0] readBusPort_1_deq_bits_data,
  input         readBusPort_1_deqRelease,
                writeBusPort_0_enq_valid,
  input  [31:0] writeBusPort_0_enq_bits_data,
  input  [1:0]  writeBusPort_0_enq_bits_mask,
  input  [2:0]  writeBusPort_0_enq_bits_instructionIndex,
  input  [9:0]  writeBusPort_0_enq_bits_counter,
  output        writeBusPort_0_enqRelease,
                writeBusPort_0_deq_valid,
  output [31:0] writeBusPort_0_deq_bits_data,
  output [1:0]  writeBusPort_0_deq_bits_mask,
  output [2:0]  writeBusPort_0_deq_bits_instructionIndex,
  output [9:0]  writeBusPort_0_deq_bits_counter,
  input         writeBusPort_0_deqRelease,
                writeBusPort_1_enq_valid,
  input  [31:0] writeBusPort_1_enq_bits_data,
  input  [1:0]  writeBusPort_1_enq_bits_mask,
  input  [2:0]  writeBusPort_1_enq_bits_instructionIndex,
  input  [9:0]  writeBusPort_1_enq_bits_counter,
  output        writeBusPort_1_enqRelease,
                writeBusPort_1_deq_valid,
  output [31:0] writeBusPort_1_deq_bits_data,
  output [1:0]  writeBusPort_1_deq_bits_mask,
  output [2:0]  writeBusPort_1_deq_bits_instructionIndex,
  output [9:0]  writeBusPort_1_deq_bits_counter,
  input         writeBusPort_1_deqRelease,
  output        laneRequest_ready,
  input         laneRequest_valid,
  input  [2:0]  laneRequest_bits_instructionIndex,
  input         laneRequest_bits_decodeResult_specialSlot,
  input  [4:0]  laneRequest_bits_decodeResult_topUop,
  input         laneRequest_bits_decodeResult_popCount,
                laneRequest_bits_decodeResult_ffo,
                laneRequest_bits_decodeResult_average,
                laneRequest_bits_decodeResult_reverse,
                laneRequest_bits_decodeResult_dontNeedExecuteInLane,
                laneRequest_bits_decodeResult_scheduler,
                laneRequest_bits_decodeResult_sReadVD,
                laneRequest_bits_decodeResult_vtype,
                laneRequest_bits_decodeResult_sWrite,
                laneRequest_bits_decodeResult_crossRead,
                laneRequest_bits_decodeResult_crossWrite,
                laneRequest_bits_decodeResult_maskUnit,
                laneRequest_bits_decodeResult_special,
                laneRequest_bits_decodeResult_saturate,
                laneRequest_bits_decodeResult_vwmacc,
                laneRequest_bits_decodeResult_readOnly,
                laneRequest_bits_decodeResult_maskSource,
                laneRequest_bits_decodeResult_maskDestination,
                laneRequest_bits_decodeResult_maskLogic,
  input  [3:0]  laneRequest_bits_decodeResult_uop,
  input         laneRequest_bits_decodeResult_iota,
                laneRequest_bits_decodeResult_mv,
                laneRequest_bits_decodeResult_extend,
                laneRequest_bits_decodeResult_unOrderWrite,
                laneRequest_bits_decodeResult_compress,
                laneRequest_bits_decodeResult_gather16,
                laneRequest_bits_decodeResult_gather,
                laneRequest_bits_decodeResult_slid,
                laneRequest_bits_decodeResult_targetRd,
                laneRequest_bits_decodeResult_widenReduce,
                laneRequest_bits_decodeResult_red,
                laneRequest_bits_decodeResult_nr,
                laneRequest_bits_decodeResult_itype,
                laneRequest_bits_decodeResult_unsigned1,
                laneRequest_bits_decodeResult_unsigned0,
                laneRequest_bits_decodeResult_other,
                laneRequest_bits_decodeResult_multiCycle,
                laneRequest_bits_decodeResult_divider,
                laneRequest_bits_decodeResult_multiplier,
                laneRequest_bits_decodeResult_shift,
                laneRequest_bits_decodeResult_adder,
                laneRequest_bits_decodeResult_logic,
                laneRequest_bits_loadStore,
                laneRequest_bits_issueInst,
                laneRequest_bits_store,
                laneRequest_bits_special,
                laneRequest_bits_lsWholeReg,
  input  [4:0]  laneRequest_bits_vs1,
                laneRequest_bits_vs2,
                laneRequest_bits_vd,
  input  [1:0]  laneRequest_bits_loadStoreEEW,
  input         laneRequest_bits_mask,
  input  [2:0]  laneRequest_bits_segment,
  input  [31:0] laneRequest_bits_readFromScalar,
  input  [13:0] laneRequest_bits_csrInterface_vl,
                laneRequest_bits_csrInterface_vStart,
  input  [2:0]  laneRequest_bits_csrInterface_vlmul,
  input  [1:0]  laneRequest_bits_csrInterface_vSew,
                laneRequest_bits_csrInterface_vxrm,
  input         laneRequest_bits_csrInterface_vta,
                laneRequest_bits_csrInterface_vma,
  output        maskUnitRequest_valid,
  output [31:0] maskUnitRequest_bits_source1,
                maskUnitRequest_bits_source2,
  output [2:0]  maskUnitRequest_bits_index,
  output        maskUnitRequest_bits_ffo,
                maskRequestToLSU,
  input         tokenIO_maskRequestRelease,
  output        vrfReadAddressChannel_ready,
  input         vrfReadAddressChannel_valid,
  input  [4:0]  vrfReadAddressChannel_bits_vs,
  input  [1:0]  vrfReadAddressChannel_bits_readSource,
  input  [5:0]  vrfReadAddressChannel_bits_offset,
  input  [2:0]  vrfReadAddressChannel_bits_instructionIndex,
  output [31:0] vrfReadDataChannel,
  output        vrfWriteChannel_ready,
  input         vrfWriteChannel_valid,
  input  [4:0]  vrfWriteChannel_bits_vd,
  input  [5:0]  vrfWriteChannel_bits_offset,
  input  [3:0]  vrfWriteChannel_bits_mask,
  input  [31:0] vrfWriteChannel_bits_data,
  input         vrfWriteChannel_bits_last,
  input  [2:0]  vrfWriteChannel_bits_instructionIndex,
  input         writeFromMask,
  output [7:0]  instructionFinished,
                vxsatReport,
  output        v0Update_valid,
  output [31:0] v0Update_bits_data,
  output [5:0]  v0Update_bits_offset,
  output [3:0]  v0Update_bits_mask,
  input  [31:0] maskInput,
  output [7:0]  maskSelect,
  output [1:0]  maskSelectSew,
  input  [7:0]  lsuLastReport,
                loadDataInLSUWriteQueue,
  input  [9:0]  writeCount,
  output [7:0]  writeQueueValid
);

  wire          _vrfReadArbiter_13_io_out_valid;
  wire [4:0]    _vrfReadArbiter_13_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_13_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_13_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_13_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_12_io_out_valid;
  wire [4:0]    _vrfReadArbiter_12_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_12_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_12_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_12_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_11_io_out_valid;
  wire [4:0]    _vrfReadArbiter_11_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_11_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_11_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_11_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_10_io_out_valid;
  wire [4:0]    _vrfReadArbiter_10_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_10_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_10_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_10_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_9_io_out_valid;
  wire [4:0]    _vrfReadArbiter_9_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_9_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_9_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_9_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_8_io_out_valid;
  wire [4:0]    _vrfReadArbiter_8_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_8_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_8_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_8_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_7_io_out_valid;
  wire [4:0]    _vrfReadArbiter_7_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_7_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_7_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_7_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_6_io_out_valid;
  wire [4:0]    _vrfReadArbiter_6_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_6_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_6_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_6_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_5_io_out_valid;
  wire [4:0]    _vrfReadArbiter_5_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_5_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_5_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_5_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_4_io_out_valid;
  wire [4:0]    _vrfReadArbiter_4_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_4_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_4_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_4_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_3_io_out_valid;
  wire [4:0]    _vrfReadArbiter_3_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_3_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_3_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_3_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_2_io_out_valid;
  wire [4:0]    _vrfReadArbiter_2_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_2_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_2_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_2_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_1_io_out_valid;
  wire [4:0]    _vrfReadArbiter_1_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_1_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_1_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_1_io_out_bits_instructionIndex;
  wire          _vrfReadArbiter_0_io_out_valid;
  wire [4:0]    _vrfReadArbiter_0_io_out_bits_vs;
  wire [1:0]    _vrfReadArbiter_0_io_out_bits_readSource;
  wire [5:0]    _vrfReadArbiter_0_io_out_bits_offset;
  wire [2:0]    _vrfReadArbiter_0_io_out_bits_instructionIndex;
  wire          _vfuResponse_otherArbiter_io_out_valid;
  wire [32:0]   _vfuResponse_otherArbiter_io_out_bits_src_0;
  wire [32:0]   _vfuResponse_otherArbiter_io_out_bits_src_1;
  wire [32:0]   _vfuResponse_otherArbiter_io_out_bits_src_2;
  wire [32:0]   _vfuResponse_otherArbiter_io_out_bits_src_3;
  wire [3:0]    _vfuResponse_otherArbiter_io_out_bits_opcode;
  wire [3:0]    _vfuResponse_otherArbiter_io_out_bits_mask;
  wire [3:0]    _vfuResponse_otherArbiter_io_out_bits_executeMask;
  wire          _vfuResponse_otherArbiter_io_out_bits_sign0;
  wire          _vfuResponse_otherArbiter_io_out_bits_sign;
  wire          _vfuResponse_otherArbiter_io_out_bits_reverse;
  wire          _vfuResponse_otherArbiter_io_out_bits_average;
  wire          _vfuResponse_otherArbiter_io_out_bits_saturate;
  wire [1:0]    _vfuResponse_otherArbiter_io_out_bits_vxrm;
  wire [1:0]    _vfuResponse_otherArbiter_io_out_bits_vSew;
  wire [19:0]   _vfuResponse_otherArbiter_io_out_bits_shifterSize;
  wire          _vfuResponse_otherArbiter_io_out_bits_rem;
  wire [1:0]    _vfuResponse_otherArbiter_io_out_bits_executeIndex;
  wire [13:0]   _vfuResponse_otherArbiter_io_out_bits_popInit;
  wire [9:0]    _vfuResponse_otherArbiter_io_out_bits_groupIndex;
  wire [1:0]    _vfuResponse_otherArbiter_io_out_bits_laneIndex;
  wire          _vfuResponse_otherArbiter_io_out_bits_maskType;
  wire          _vfuResponse_otherArbiter_io_out_bits_narrow;
  wire [1:0]    _vfuResponse_otherArbiter_io_out_bits_tag;
  wire          _vfuResponse_otherDistributor_requestToVfu_valid;
  wire [32:0]   _vfuResponse_otherDistributor_requestToVfu_bits_src_0;
  wire [32:0]   _vfuResponse_otherDistributor_requestToVfu_bits_src_1;
  wire [32:0]   _vfuResponse_otherDistributor_requestToVfu_bits_src_2;
  wire [32:0]   _vfuResponse_otherDistributor_requestToVfu_bits_src_3;
  wire [3:0]    _vfuResponse_otherDistributor_requestToVfu_bits_opcode;
  wire [3:0]    _vfuResponse_otherDistributor_requestToVfu_bits_mask;
  wire          _vfuResponse_otherDistributor_requestToVfu_bits_sign;
  wire [1:0]    _vfuResponse_otherDistributor_requestToVfu_bits_vxrm;
  wire [1:0]    _vfuResponse_otherDistributor_requestToVfu_bits_vSew;
  wire [1:0]    _vfuResponse_otherDistributor_requestToVfu_bits_executeIndex;
  wire [13:0]   _vfuResponse_otherDistributor_requestToVfu_bits_popInit;
  wire [9:0]    _vfuResponse_otherDistributor_requestToVfu_bits_groupIndex;
  wire [1:0]    _vfuResponse_otherDistributor_requestToVfu_bits_laneIndex;
  wire          _vfuResponse_otherDistributor_requestToVfu_bits_maskType;
  wire          _vfuResponse_otherDistributor_requestToVfu_bits_narrow;
  wire [1:0]    _vfuResponse_otherDistributor_requestToVfu_bits_tag;
  wire          _vfuResponse_otherDistributor_requestFromSlot_ready;
  wire          _vfuResponse_otherDistributor_responseToSlot_valid;
  wire [31:0]   _vfuResponse_otherDistributor_responseToSlot_bits_data;
  wire          _vfuResponse_otherDistributor_responseToSlot_bits_ffoSuccess;
  wire [3:0]    _vfuResponse_otherDistributor_responseToSlot_bits_vxsat;
  wire [1:0]    _vfuResponse_otherDistributor_responseToSlot_bits_tag;
  wire          _vfuResponse_dividerArbiter_io_out_valid;
  wire [32:0]   _vfuResponse_dividerArbiter_io_out_bits_src_0;
  wire [32:0]   _vfuResponse_dividerArbiter_io_out_bits_src_1;
  wire [32:0]   _vfuResponse_dividerArbiter_io_out_bits_src_2;
  wire [32:0]   _vfuResponse_dividerArbiter_io_out_bits_src_3;
  wire [3:0]    _vfuResponse_dividerArbiter_io_out_bits_opcode;
  wire [3:0]    _vfuResponse_dividerArbiter_io_out_bits_mask;
  wire [3:0]    _vfuResponse_dividerArbiter_io_out_bits_executeMask;
  wire          _vfuResponse_dividerArbiter_io_out_bits_sign0;
  wire          _vfuResponse_dividerArbiter_io_out_bits_sign;
  wire          _vfuResponse_dividerArbiter_io_out_bits_reverse;
  wire          _vfuResponse_dividerArbiter_io_out_bits_average;
  wire          _vfuResponse_dividerArbiter_io_out_bits_saturate;
  wire [1:0]    _vfuResponse_dividerArbiter_io_out_bits_vxrm;
  wire [1:0]    _vfuResponse_dividerArbiter_io_out_bits_vSew;
  wire [19:0]   _vfuResponse_dividerArbiter_io_out_bits_shifterSize;
  wire          _vfuResponse_dividerArbiter_io_out_bits_rem;
  wire [1:0]    _vfuResponse_dividerArbiter_io_out_bits_executeIndex;
  wire [13:0]   _vfuResponse_dividerArbiter_io_out_bits_popInit;
  wire [9:0]    _vfuResponse_dividerArbiter_io_out_bits_groupIndex;
  wire [1:0]    _vfuResponse_dividerArbiter_io_out_bits_laneIndex;
  wire          _vfuResponse_dividerArbiter_io_out_bits_maskType;
  wire          _vfuResponse_dividerArbiter_io_out_bits_narrow;
  wire [1:0]    _vfuResponse_dividerArbiter_io_out_bits_tag;
  wire          _vfuResponse_dividerDistributor_requestToVfu_valid;
  wire [32:0]   _vfuResponse_dividerDistributor_requestToVfu_bits_src_0;
  wire [32:0]   _vfuResponse_dividerDistributor_requestToVfu_bits_src_1;
  wire [3:0]    _vfuResponse_dividerDistributor_requestToVfu_bits_opcode;
  wire          _vfuResponse_dividerDistributor_requestToVfu_bits_sign;
  wire [1:0]    _vfuResponse_dividerDistributor_requestToVfu_bits_executeIndex;
  wire [1:0]    _vfuResponse_dividerDistributor_requestToVfu_bits_tag;
  wire          _vfuResponse_dividerDistributor_requestFromSlot_ready;
  wire          _vfuResponse_dividerDistributor_responseToSlot_valid;
  wire [31:0]   _vfuResponse_dividerDistributor_responseToSlot_bits_data;
  wire          _vfuResponse_dividerDistributor_responseToSlot_bits_ffoSuccess;
  wire [3:0]    _vfuResponse_dividerDistributor_responseToSlot_bits_vxsat;
  wire [1:0]    _vfuResponse_dividerDistributor_responseToSlot_bits_tag;
  wire          _vfuResponse_multiplierArbiter_io_out_valid;
  wire [32:0]   _vfuResponse_multiplierArbiter_io_out_bits_src_0;
  wire [32:0]   _vfuResponse_multiplierArbiter_io_out_bits_src_1;
  wire [32:0]   _vfuResponse_multiplierArbiter_io_out_bits_src_2;
  wire [3:0]    _vfuResponse_multiplierArbiter_io_out_bits_opcode;
  wire          _vfuResponse_multiplierArbiter_io_out_bits_sign0;
  wire          _vfuResponse_multiplierArbiter_io_out_bits_sign;
  wire          _vfuResponse_multiplierArbiter_io_out_bits_saturate;
  wire [1:0]    _vfuResponse_multiplierArbiter_io_out_bits_vxrm;
  wire [1:0]    _vfuResponse_multiplierArbiter_io_out_bits_vSew;
  wire [1:0]    _vfuResponse_multiplierArbiter_io_out_bits_tag;
  wire          _vfuResponse_shiftArbiter_io_out_valid;
  wire [32:0]   _vfuResponse_shiftArbiter_io_out_bits_src_0;
  wire [32:0]   _vfuResponse_shiftArbiter_io_out_bits_src_1;
  wire [32:0]   _vfuResponse_shiftArbiter_io_out_bits_src_2;
  wire [32:0]   _vfuResponse_shiftArbiter_io_out_bits_src_3;
  wire [3:0]    _vfuResponse_shiftArbiter_io_out_bits_opcode;
  wire [3:0]    _vfuResponse_shiftArbiter_io_out_bits_mask;
  wire [3:0]    _vfuResponse_shiftArbiter_io_out_bits_executeMask;
  wire          _vfuResponse_shiftArbiter_io_out_bits_sign0;
  wire          _vfuResponse_shiftArbiter_io_out_bits_sign;
  wire          _vfuResponse_shiftArbiter_io_out_bits_reverse;
  wire          _vfuResponse_shiftArbiter_io_out_bits_average;
  wire          _vfuResponse_shiftArbiter_io_out_bits_saturate;
  wire [1:0]    _vfuResponse_shiftArbiter_io_out_bits_vxrm;
  wire [1:0]    _vfuResponse_shiftArbiter_io_out_bits_vSew;
  wire [19:0]   _vfuResponse_shiftArbiter_io_out_bits_shifterSize;
  wire          _vfuResponse_shiftArbiter_io_out_bits_rem;
  wire [1:0]    _vfuResponse_shiftArbiter_io_out_bits_executeIndex;
  wire [13:0]   _vfuResponse_shiftArbiter_io_out_bits_popInit;
  wire [9:0]    _vfuResponse_shiftArbiter_io_out_bits_groupIndex;
  wire [1:0]    _vfuResponse_shiftArbiter_io_out_bits_laneIndex;
  wire          _vfuResponse_shiftArbiter_io_out_bits_maskType;
  wire          _vfuResponse_shiftArbiter_io_out_bits_narrow;
  wire [1:0]    _vfuResponse_shiftArbiter_io_out_bits_tag;
  wire          _vfuResponse_shiftDistributor_requestToVfu_valid;
  wire [32:0]   _vfuResponse_shiftDistributor_requestToVfu_bits_src_0;
  wire [32:0]   _vfuResponse_shiftDistributor_requestToVfu_bits_src_1;
  wire [3:0]    _vfuResponse_shiftDistributor_requestToVfu_bits_opcode;
  wire [1:0]    _vfuResponse_shiftDistributor_requestToVfu_bits_vxrm;
  wire [19:0]   _vfuResponse_shiftDistributor_requestToVfu_bits_shifterSize;
  wire [1:0]    _vfuResponse_shiftDistributor_requestToVfu_bits_tag;
  wire          _vfuResponse_shiftDistributor_requestFromSlot_ready;
  wire          _vfuResponse_shiftDistributor_responseToSlot_valid;
  wire [31:0]   _vfuResponse_shiftDistributor_responseToSlot_bits_data;
  wire          _vfuResponse_shiftDistributor_responseToSlot_bits_ffoSuccess;
  wire [3:0]    _vfuResponse_shiftDistributor_responseToSlot_bits_vxsat;
  wire [1:0]    _vfuResponse_shiftDistributor_responseToSlot_bits_tag;
  wire          _vfuResponse_adderArbiter_io_out_valid;
  wire [32:0]   _vfuResponse_adderArbiter_io_out_bits_src_0;
  wire [32:0]   _vfuResponse_adderArbiter_io_out_bits_src_1;
  wire [3:0]    _vfuResponse_adderArbiter_io_out_bits_opcode;
  wire [3:0]    _vfuResponse_adderArbiter_io_out_bits_mask;
  wire          _vfuResponse_adderArbiter_io_out_bits_sign;
  wire          _vfuResponse_adderArbiter_io_out_bits_reverse;
  wire          _vfuResponse_adderArbiter_io_out_bits_average;
  wire          _vfuResponse_adderArbiter_io_out_bits_saturate;
  wire [1:0]    _vfuResponse_adderArbiter_io_out_bits_vxrm;
  wire [1:0]    _vfuResponse_adderArbiter_io_out_bits_vSew;
  wire [1:0]    _vfuResponse_adderArbiter_io_out_bits_executeIndex;
  wire [1:0]    _vfuResponse_adderArbiter_io_out_bits_tag;
  wire          _vfuResponse_logicArbiter_io_out_valid;
  wire [32:0]   _vfuResponse_logicArbiter_io_out_bits_src_0;
  wire [32:0]   _vfuResponse_logicArbiter_io_out_bits_src_1;
  wire [32:0]   _vfuResponse_logicArbiter_io_out_bits_src_2;
  wire [32:0]   _vfuResponse_logicArbiter_io_out_bits_src_3;
  wire [3:0]    _vfuResponse_logicArbiter_io_out_bits_opcode;
  wire [1:0]    _vfuResponse_logicArbiter_io_out_bits_tag;
  wire          _divider_requestIO_ready;
  wire          _multiplier_responseIO_bits_vxsat;
  wire          _stage3_3_vrfWriteRequest_valid;
  wire [3:0]    _stage3_3_vrfWriteRequest_bits_mask;
  wire [2:0]    _stage3_3_vrfWriteRequest_bits_instructionIndex;
  wire          _executionUnit_3_enqueue_ready;
  wire          _executionUnit_3_dequeue_valid;
  wire          _executionUnit_3_vfuRequest_valid;
  wire [2:0]    _executionUnit_3_responseIndex;
  wire          _stage2_3_enqueue_ready;
  wire          _stage2_3_dequeue_valid;
  wire          _stage1_3_enqueue_ready;
  wire          _stage1_3_dequeue_valid;
  wire [3:0]    _stage1_3_dequeue_bits_maskForFilter;
  wire [3:0]    _stage1_3_dequeue_bits_mask;
  wire [9:0]    _stage1_3_dequeue_bits_groupCounter;
  wire [31:0]   _stage1_3_dequeue_bits_src_0;
  wire [31:0]   _stage1_3_dequeue_bits_src_1;
  wire [31:0]   _stage1_3_dequeue_bits_src_2;
  wire          _stage1_3_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage1_3_dequeue_bits_decodeResult_topUop;
  wire          _stage1_3_dequeue_bits_decodeResult_popCount;
  wire          _stage1_3_dequeue_bits_decodeResult_ffo;
  wire          _stage1_3_dequeue_bits_decodeResult_average;
  wire          _stage1_3_dequeue_bits_decodeResult_reverse;
  wire          _stage1_3_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage1_3_dequeue_bits_decodeResult_scheduler;
  wire          _stage1_3_dequeue_bits_decodeResult_sReadVD;
  wire          _stage1_3_dequeue_bits_decodeResult_vtype;
  wire          _stage1_3_dequeue_bits_decodeResult_sWrite;
  wire          _stage1_3_dequeue_bits_decodeResult_crossRead;
  wire          _stage1_3_dequeue_bits_decodeResult_crossWrite;
  wire          _stage1_3_dequeue_bits_decodeResult_maskUnit;
  wire          _stage1_3_dequeue_bits_decodeResult_special;
  wire          _stage1_3_dequeue_bits_decodeResult_saturate;
  wire          _stage1_3_dequeue_bits_decodeResult_vwmacc;
  wire          _stage1_3_dequeue_bits_decodeResult_readOnly;
  wire          _stage1_3_dequeue_bits_decodeResult_maskSource;
  wire          _stage1_3_dequeue_bits_decodeResult_maskDestination;
  wire          _stage1_3_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage1_3_dequeue_bits_decodeResult_uop;
  wire          _stage1_3_dequeue_bits_decodeResult_iota;
  wire          _stage1_3_dequeue_bits_decodeResult_mv;
  wire          _stage1_3_dequeue_bits_decodeResult_extend;
  wire          _stage1_3_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage1_3_dequeue_bits_decodeResult_compress;
  wire          _stage1_3_dequeue_bits_decodeResult_gather16;
  wire          _stage1_3_dequeue_bits_decodeResult_gather;
  wire          _stage1_3_dequeue_bits_decodeResult_slid;
  wire          _stage1_3_dequeue_bits_decodeResult_targetRd;
  wire          _stage1_3_dequeue_bits_decodeResult_widenReduce;
  wire          _stage1_3_dequeue_bits_decodeResult_red;
  wire          _stage1_3_dequeue_bits_decodeResult_nr;
  wire          _stage1_3_dequeue_bits_decodeResult_itype;
  wire          _stage1_3_dequeue_bits_decodeResult_unsigned1;
  wire          _stage1_3_dequeue_bits_decodeResult_unsigned0;
  wire          _stage1_3_dequeue_bits_decodeResult_other;
  wire          _stage1_3_dequeue_bits_decodeResult_multiCycle;
  wire          _stage1_3_dequeue_bits_decodeResult_divider;
  wire          _stage1_3_dequeue_bits_decodeResult_multiplier;
  wire          _stage1_3_dequeue_bits_decodeResult_shift;
  wire          _stage1_3_dequeue_bits_decodeResult_adder;
  wire          _stage1_3_dequeue_bits_decodeResult_logic;
  wire [2:0]    _stage1_3_dequeue_bits_vSew1H;
  wire [13:0]   _stage1_3_dequeue_bits_csr_vl;
  wire [13:0]   _stage1_3_dequeue_bits_csr_vStart;
  wire [2:0]    _stage1_3_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage1_3_dequeue_bits_csr_vSew;
  wire [1:0]    _stage1_3_dequeue_bits_csr_vxrm;
  wire          _stage1_3_dequeue_bits_csr_vta;
  wire          _stage1_3_dequeue_bits_csr_vma;
  wire          _stage1_3_dequeue_bits_maskType;
  wire [1:0]    _stage1_3_dequeue_bits_laneIndex;
  wire [2:0]    _stage1_3_dequeue_bits_instructionIndex;
  wire          _stage1_3_dequeue_bits_loadStore;
  wire [4:0]    _stage1_3_dequeue_bits_vd;
  wire          _stage1_3_dequeue_bits_bordersForMaskLogic;
  wire          _stage0_3_enqueue_ready;
  wire          _stage0_3_dequeue_valid;
  wire [3:0]    _stage0_3_dequeue_bits_maskForMaskInput;
  wire [3:0]    _stage0_3_dequeue_bits_boundaryMaskCorrection;
  wire [9:0]    _stage0_3_dequeue_bits_groupCounter;
  wire [31:0]   _stage0_3_dequeue_bits_readFromScalar;
  wire [2:0]    _stage0_3_dequeue_bits_instructionIndex;
  wire          _stage0_3_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage0_3_dequeue_bits_decodeResult_topUop;
  wire          _stage0_3_dequeue_bits_decodeResult_popCount;
  wire          _stage0_3_dequeue_bits_decodeResult_ffo;
  wire          _stage0_3_dequeue_bits_decodeResult_average;
  wire          _stage0_3_dequeue_bits_decodeResult_reverse;
  wire          _stage0_3_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage0_3_dequeue_bits_decodeResult_scheduler;
  wire          _stage0_3_dequeue_bits_decodeResult_sReadVD;
  wire          _stage0_3_dequeue_bits_decodeResult_vtype;
  wire          _stage0_3_dequeue_bits_decodeResult_sWrite;
  wire          _stage0_3_dequeue_bits_decodeResult_crossRead;
  wire          _stage0_3_dequeue_bits_decodeResult_crossWrite;
  wire          _stage0_3_dequeue_bits_decodeResult_maskUnit;
  wire          _stage0_3_dequeue_bits_decodeResult_special;
  wire          _stage0_3_dequeue_bits_decodeResult_saturate;
  wire          _stage0_3_dequeue_bits_decodeResult_vwmacc;
  wire          _stage0_3_dequeue_bits_decodeResult_readOnly;
  wire          _stage0_3_dequeue_bits_decodeResult_maskSource;
  wire          _stage0_3_dequeue_bits_decodeResult_maskDestination;
  wire          _stage0_3_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage0_3_dequeue_bits_decodeResult_uop;
  wire          _stage0_3_dequeue_bits_decodeResult_iota;
  wire          _stage0_3_dequeue_bits_decodeResult_mv;
  wire          _stage0_3_dequeue_bits_decodeResult_extend;
  wire          _stage0_3_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage0_3_dequeue_bits_decodeResult_compress;
  wire          _stage0_3_dequeue_bits_decodeResult_gather16;
  wire          _stage0_3_dequeue_bits_decodeResult_gather;
  wire          _stage0_3_dequeue_bits_decodeResult_slid;
  wire          _stage0_3_dequeue_bits_decodeResult_targetRd;
  wire          _stage0_3_dequeue_bits_decodeResult_widenReduce;
  wire          _stage0_3_dequeue_bits_decodeResult_red;
  wire          _stage0_3_dequeue_bits_decodeResult_nr;
  wire          _stage0_3_dequeue_bits_decodeResult_itype;
  wire          _stage0_3_dequeue_bits_decodeResult_unsigned1;
  wire          _stage0_3_dequeue_bits_decodeResult_unsigned0;
  wire          _stage0_3_dequeue_bits_decodeResult_other;
  wire          _stage0_3_dequeue_bits_decodeResult_multiCycle;
  wire          _stage0_3_dequeue_bits_decodeResult_divider;
  wire          _stage0_3_dequeue_bits_decodeResult_multiplier;
  wire          _stage0_3_dequeue_bits_decodeResult_shift;
  wire          _stage0_3_dequeue_bits_decodeResult_adder;
  wire          _stage0_3_dequeue_bits_decodeResult_logic;
  wire [1:0]    _stage0_3_dequeue_bits_laneIndex;
  wire          _stage0_3_dequeue_bits_skipRead;
  wire [4:0]    _stage0_3_dequeue_bits_vs1;
  wire [4:0]    _stage0_3_dequeue_bits_vs2;
  wire [4:0]    _stage0_3_dequeue_bits_vd;
  wire [2:0]    _stage0_3_dequeue_bits_vSew1H;
  wire          _stage0_3_dequeue_bits_maskNotMaskedElement;
  wire [13:0]   _stage0_3_dequeue_bits_csr_vl;
  wire [13:0]   _stage0_3_dequeue_bits_csr_vStart;
  wire [2:0]    _stage0_3_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage0_3_dequeue_bits_csr_vSew;
  wire [1:0]    _stage0_3_dequeue_bits_csr_vxrm;
  wire          _stage0_3_dequeue_bits_csr_vta;
  wire          _stage0_3_dequeue_bits_csr_vma;
  wire          _stage0_3_dequeue_bits_maskType;
  wire          _stage0_3_dequeue_bits_loadStore;
  wire          _stage0_3_dequeue_bits_bordersForMaskLogic;
  wire [7:0]    _stage0_3_updateLaneState_maskGroupCount;
  wire [4:0]    _stage0_3_updateLaneState_maskIndex;
  wire          _stage0_3_updateLaneState_outOfExecutionRange;
  wire          _stage0_3_updateLaneState_maskExhausted;
  wire          _stage0_3_tokenReport_valid;
  wire          _stage0_3_tokenReport_bits_decodeResult_sWrite;
  wire          _stage0_3_tokenReport_bits_decodeResult_maskUnit;
  wire [2:0]    _stage0_3_tokenReport_bits_instructionIndex;
  wire          _stage3_2_vrfWriteRequest_valid;
  wire [3:0]    _stage3_2_vrfWriteRequest_bits_mask;
  wire [2:0]    _stage3_2_vrfWriteRequest_bits_instructionIndex;
  wire          _executionUnit_2_enqueue_ready;
  wire          _executionUnit_2_dequeue_valid;
  wire          _executionUnit_2_vfuRequest_valid;
  wire [2:0]    _executionUnit_2_responseIndex;
  wire          _stage2_2_enqueue_ready;
  wire          _stage2_2_dequeue_valid;
  wire          _stage1_2_enqueue_ready;
  wire          _stage1_2_dequeue_valid;
  wire [3:0]    _stage1_2_dequeue_bits_maskForFilter;
  wire [3:0]    _stage1_2_dequeue_bits_mask;
  wire [9:0]    _stage1_2_dequeue_bits_groupCounter;
  wire [31:0]   _stage1_2_dequeue_bits_src_0;
  wire [31:0]   _stage1_2_dequeue_bits_src_1;
  wire [31:0]   _stage1_2_dequeue_bits_src_2;
  wire          _stage1_2_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage1_2_dequeue_bits_decodeResult_topUop;
  wire          _stage1_2_dequeue_bits_decodeResult_popCount;
  wire          _stage1_2_dequeue_bits_decodeResult_ffo;
  wire          _stage1_2_dequeue_bits_decodeResult_average;
  wire          _stage1_2_dequeue_bits_decodeResult_reverse;
  wire          _stage1_2_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage1_2_dequeue_bits_decodeResult_scheduler;
  wire          _stage1_2_dequeue_bits_decodeResult_sReadVD;
  wire          _stage1_2_dequeue_bits_decodeResult_vtype;
  wire          _stage1_2_dequeue_bits_decodeResult_sWrite;
  wire          _stage1_2_dequeue_bits_decodeResult_crossRead;
  wire          _stage1_2_dequeue_bits_decodeResult_crossWrite;
  wire          _stage1_2_dequeue_bits_decodeResult_maskUnit;
  wire          _stage1_2_dequeue_bits_decodeResult_special;
  wire          _stage1_2_dequeue_bits_decodeResult_saturate;
  wire          _stage1_2_dequeue_bits_decodeResult_vwmacc;
  wire          _stage1_2_dequeue_bits_decodeResult_readOnly;
  wire          _stage1_2_dequeue_bits_decodeResult_maskSource;
  wire          _stage1_2_dequeue_bits_decodeResult_maskDestination;
  wire          _stage1_2_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage1_2_dequeue_bits_decodeResult_uop;
  wire          _stage1_2_dequeue_bits_decodeResult_iota;
  wire          _stage1_2_dequeue_bits_decodeResult_mv;
  wire          _stage1_2_dequeue_bits_decodeResult_extend;
  wire          _stage1_2_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage1_2_dequeue_bits_decodeResult_compress;
  wire          _stage1_2_dequeue_bits_decodeResult_gather16;
  wire          _stage1_2_dequeue_bits_decodeResult_gather;
  wire          _stage1_2_dequeue_bits_decodeResult_slid;
  wire          _stage1_2_dequeue_bits_decodeResult_targetRd;
  wire          _stage1_2_dequeue_bits_decodeResult_widenReduce;
  wire          _stage1_2_dequeue_bits_decodeResult_red;
  wire          _stage1_2_dequeue_bits_decodeResult_nr;
  wire          _stage1_2_dequeue_bits_decodeResult_itype;
  wire          _stage1_2_dequeue_bits_decodeResult_unsigned1;
  wire          _stage1_2_dequeue_bits_decodeResult_unsigned0;
  wire          _stage1_2_dequeue_bits_decodeResult_other;
  wire          _stage1_2_dequeue_bits_decodeResult_multiCycle;
  wire          _stage1_2_dequeue_bits_decodeResult_divider;
  wire          _stage1_2_dequeue_bits_decodeResult_multiplier;
  wire          _stage1_2_dequeue_bits_decodeResult_shift;
  wire          _stage1_2_dequeue_bits_decodeResult_adder;
  wire          _stage1_2_dequeue_bits_decodeResult_logic;
  wire [2:0]    _stage1_2_dequeue_bits_vSew1H;
  wire [13:0]   _stage1_2_dequeue_bits_csr_vl;
  wire [13:0]   _stage1_2_dequeue_bits_csr_vStart;
  wire [2:0]    _stage1_2_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage1_2_dequeue_bits_csr_vSew;
  wire [1:0]    _stage1_2_dequeue_bits_csr_vxrm;
  wire          _stage1_2_dequeue_bits_csr_vta;
  wire          _stage1_2_dequeue_bits_csr_vma;
  wire          _stage1_2_dequeue_bits_maskType;
  wire [1:0]    _stage1_2_dequeue_bits_laneIndex;
  wire [2:0]    _stage1_2_dequeue_bits_instructionIndex;
  wire          _stage1_2_dequeue_bits_loadStore;
  wire [4:0]    _stage1_2_dequeue_bits_vd;
  wire          _stage1_2_dequeue_bits_bordersForMaskLogic;
  wire          _stage0_2_enqueue_ready;
  wire          _stage0_2_dequeue_valid;
  wire [3:0]    _stage0_2_dequeue_bits_maskForMaskInput;
  wire [3:0]    _stage0_2_dequeue_bits_boundaryMaskCorrection;
  wire [9:0]    _stage0_2_dequeue_bits_groupCounter;
  wire [31:0]   _stage0_2_dequeue_bits_readFromScalar;
  wire [2:0]    _stage0_2_dequeue_bits_instructionIndex;
  wire          _stage0_2_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage0_2_dequeue_bits_decodeResult_topUop;
  wire          _stage0_2_dequeue_bits_decodeResult_popCount;
  wire          _stage0_2_dequeue_bits_decodeResult_ffo;
  wire          _stage0_2_dequeue_bits_decodeResult_average;
  wire          _stage0_2_dequeue_bits_decodeResult_reverse;
  wire          _stage0_2_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage0_2_dequeue_bits_decodeResult_scheduler;
  wire          _stage0_2_dequeue_bits_decodeResult_sReadVD;
  wire          _stage0_2_dequeue_bits_decodeResult_vtype;
  wire          _stage0_2_dequeue_bits_decodeResult_sWrite;
  wire          _stage0_2_dequeue_bits_decodeResult_crossRead;
  wire          _stage0_2_dequeue_bits_decodeResult_crossWrite;
  wire          _stage0_2_dequeue_bits_decodeResult_maskUnit;
  wire          _stage0_2_dequeue_bits_decodeResult_special;
  wire          _stage0_2_dequeue_bits_decodeResult_saturate;
  wire          _stage0_2_dequeue_bits_decodeResult_vwmacc;
  wire          _stage0_2_dequeue_bits_decodeResult_readOnly;
  wire          _stage0_2_dequeue_bits_decodeResult_maskSource;
  wire          _stage0_2_dequeue_bits_decodeResult_maskDestination;
  wire          _stage0_2_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage0_2_dequeue_bits_decodeResult_uop;
  wire          _stage0_2_dequeue_bits_decodeResult_iota;
  wire          _stage0_2_dequeue_bits_decodeResult_mv;
  wire          _stage0_2_dequeue_bits_decodeResult_extend;
  wire          _stage0_2_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage0_2_dequeue_bits_decodeResult_compress;
  wire          _stage0_2_dequeue_bits_decodeResult_gather16;
  wire          _stage0_2_dequeue_bits_decodeResult_gather;
  wire          _stage0_2_dequeue_bits_decodeResult_slid;
  wire          _stage0_2_dequeue_bits_decodeResult_targetRd;
  wire          _stage0_2_dequeue_bits_decodeResult_widenReduce;
  wire          _stage0_2_dequeue_bits_decodeResult_red;
  wire          _stage0_2_dequeue_bits_decodeResult_nr;
  wire          _stage0_2_dequeue_bits_decodeResult_itype;
  wire          _stage0_2_dequeue_bits_decodeResult_unsigned1;
  wire          _stage0_2_dequeue_bits_decodeResult_unsigned0;
  wire          _stage0_2_dequeue_bits_decodeResult_other;
  wire          _stage0_2_dequeue_bits_decodeResult_multiCycle;
  wire          _stage0_2_dequeue_bits_decodeResult_divider;
  wire          _stage0_2_dequeue_bits_decodeResult_multiplier;
  wire          _stage0_2_dequeue_bits_decodeResult_shift;
  wire          _stage0_2_dequeue_bits_decodeResult_adder;
  wire          _stage0_2_dequeue_bits_decodeResult_logic;
  wire [1:0]    _stage0_2_dequeue_bits_laneIndex;
  wire          _stage0_2_dequeue_bits_skipRead;
  wire [4:0]    _stage0_2_dequeue_bits_vs1;
  wire [4:0]    _stage0_2_dequeue_bits_vs2;
  wire [4:0]    _stage0_2_dequeue_bits_vd;
  wire [2:0]    _stage0_2_dequeue_bits_vSew1H;
  wire          _stage0_2_dequeue_bits_maskNotMaskedElement;
  wire [13:0]   _stage0_2_dequeue_bits_csr_vl;
  wire [13:0]   _stage0_2_dequeue_bits_csr_vStart;
  wire [2:0]    _stage0_2_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage0_2_dequeue_bits_csr_vSew;
  wire [1:0]    _stage0_2_dequeue_bits_csr_vxrm;
  wire          _stage0_2_dequeue_bits_csr_vta;
  wire          _stage0_2_dequeue_bits_csr_vma;
  wire          _stage0_2_dequeue_bits_maskType;
  wire          _stage0_2_dequeue_bits_loadStore;
  wire          _stage0_2_dequeue_bits_bordersForMaskLogic;
  wire [7:0]    _stage0_2_updateLaneState_maskGroupCount;
  wire [4:0]    _stage0_2_updateLaneState_maskIndex;
  wire          _stage0_2_updateLaneState_outOfExecutionRange;
  wire          _stage0_2_updateLaneState_maskExhausted;
  wire          _stage0_2_tokenReport_valid;
  wire          _stage0_2_tokenReport_bits_decodeResult_sWrite;
  wire          _stage0_2_tokenReport_bits_decodeResult_maskUnit;
  wire [2:0]    _stage0_2_tokenReport_bits_instructionIndex;
  wire          _stage3_1_vrfWriteRequest_valid;
  wire [3:0]    _stage3_1_vrfWriteRequest_bits_mask;
  wire [2:0]    _stage3_1_vrfWriteRequest_bits_instructionIndex;
  wire          _executionUnit_1_enqueue_ready;
  wire          _executionUnit_1_dequeue_valid;
  wire          _executionUnit_1_vfuRequest_valid;
  wire [2:0]    _executionUnit_1_responseIndex;
  wire          _stage2_1_enqueue_ready;
  wire          _stage2_1_dequeue_valid;
  wire          _stage1_1_enqueue_ready;
  wire          _stage1_1_dequeue_valid;
  wire [3:0]    _stage1_1_dequeue_bits_maskForFilter;
  wire [3:0]    _stage1_1_dequeue_bits_mask;
  wire [9:0]    _stage1_1_dequeue_bits_groupCounter;
  wire [31:0]   _stage1_1_dequeue_bits_src_0;
  wire [31:0]   _stage1_1_dequeue_bits_src_1;
  wire [31:0]   _stage1_1_dequeue_bits_src_2;
  wire          _stage1_1_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage1_1_dequeue_bits_decodeResult_topUop;
  wire          _stage1_1_dequeue_bits_decodeResult_popCount;
  wire          _stage1_1_dequeue_bits_decodeResult_ffo;
  wire          _stage1_1_dequeue_bits_decodeResult_average;
  wire          _stage1_1_dequeue_bits_decodeResult_reverse;
  wire          _stage1_1_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage1_1_dequeue_bits_decodeResult_scheduler;
  wire          _stage1_1_dequeue_bits_decodeResult_sReadVD;
  wire          _stage1_1_dequeue_bits_decodeResult_vtype;
  wire          _stage1_1_dequeue_bits_decodeResult_sWrite;
  wire          _stage1_1_dequeue_bits_decodeResult_crossRead;
  wire          _stage1_1_dequeue_bits_decodeResult_crossWrite;
  wire          _stage1_1_dequeue_bits_decodeResult_maskUnit;
  wire          _stage1_1_dequeue_bits_decodeResult_special;
  wire          _stage1_1_dequeue_bits_decodeResult_saturate;
  wire          _stage1_1_dequeue_bits_decodeResult_vwmacc;
  wire          _stage1_1_dequeue_bits_decodeResult_readOnly;
  wire          _stage1_1_dequeue_bits_decodeResult_maskSource;
  wire          _stage1_1_dequeue_bits_decodeResult_maskDestination;
  wire          _stage1_1_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage1_1_dequeue_bits_decodeResult_uop;
  wire          _stage1_1_dequeue_bits_decodeResult_iota;
  wire          _stage1_1_dequeue_bits_decodeResult_mv;
  wire          _stage1_1_dequeue_bits_decodeResult_extend;
  wire          _stage1_1_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage1_1_dequeue_bits_decodeResult_compress;
  wire          _stage1_1_dequeue_bits_decodeResult_gather16;
  wire          _stage1_1_dequeue_bits_decodeResult_gather;
  wire          _stage1_1_dequeue_bits_decodeResult_slid;
  wire          _stage1_1_dequeue_bits_decodeResult_targetRd;
  wire          _stage1_1_dequeue_bits_decodeResult_widenReduce;
  wire          _stage1_1_dequeue_bits_decodeResult_red;
  wire          _stage1_1_dequeue_bits_decodeResult_nr;
  wire          _stage1_1_dequeue_bits_decodeResult_itype;
  wire          _stage1_1_dequeue_bits_decodeResult_unsigned1;
  wire          _stage1_1_dequeue_bits_decodeResult_unsigned0;
  wire          _stage1_1_dequeue_bits_decodeResult_other;
  wire          _stage1_1_dequeue_bits_decodeResult_multiCycle;
  wire          _stage1_1_dequeue_bits_decodeResult_divider;
  wire          _stage1_1_dequeue_bits_decodeResult_multiplier;
  wire          _stage1_1_dequeue_bits_decodeResult_shift;
  wire          _stage1_1_dequeue_bits_decodeResult_adder;
  wire          _stage1_1_dequeue_bits_decodeResult_logic;
  wire [2:0]    _stage1_1_dequeue_bits_vSew1H;
  wire [13:0]   _stage1_1_dequeue_bits_csr_vl;
  wire [13:0]   _stage1_1_dequeue_bits_csr_vStart;
  wire [2:0]    _stage1_1_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage1_1_dequeue_bits_csr_vSew;
  wire [1:0]    _stage1_1_dequeue_bits_csr_vxrm;
  wire          _stage1_1_dequeue_bits_csr_vta;
  wire          _stage1_1_dequeue_bits_csr_vma;
  wire          _stage1_1_dequeue_bits_maskType;
  wire [1:0]    _stage1_1_dequeue_bits_laneIndex;
  wire [2:0]    _stage1_1_dequeue_bits_instructionIndex;
  wire          _stage1_1_dequeue_bits_loadStore;
  wire [4:0]    _stage1_1_dequeue_bits_vd;
  wire          _stage1_1_dequeue_bits_bordersForMaskLogic;
  wire          _stage0_1_enqueue_ready;
  wire          _stage0_1_dequeue_valid;
  wire [3:0]    _stage0_1_dequeue_bits_maskForMaskInput;
  wire [3:0]    _stage0_1_dequeue_bits_boundaryMaskCorrection;
  wire [9:0]    _stage0_1_dequeue_bits_groupCounter;
  wire [31:0]   _stage0_1_dequeue_bits_readFromScalar;
  wire [2:0]    _stage0_1_dequeue_bits_instructionIndex;
  wire          _stage0_1_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage0_1_dequeue_bits_decodeResult_topUop;
  wire          _stage0_1_dequeue_bits_decodeResult_popCount;
  wire          _stage0_1_dequeue_bits_decodeResult_ffo;
  wire          _stage0_1_dequeue_bits_decodeResult_average;
  wire          _stage0_1_dequeue_bits_decodeResult_reverse;
  wire          _stage0_1_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage0_1_dequeue_bits_decodeResult_scheduler;
  wire          _stage0_1_dequeue_bits_decodeResult_sReadVD;
  wire          _stage0_1_dequeue_bits_decodeResult_vtype;
  wire          _stage0_1_dequeue_bits_decodeResult_sWrite;
  wire          _stage0_1_dequeue_bits_decodeResult_crossRead;
  wire          _stage0_1_dequeue_bits_decodeResult_crossWrite;
  wire          _stage0_1_dequeue_bits_decodeResult_maskUnit;
  wire          _stage0_1_dequeue_bits_decodeResult_special;
  wire          _stage0_1_dequeue_bits_decodeResult_saturate;
  wire          _stage0_1_dequeue_bits_decodeResult_vwmacc;
  wire          _stage0_1_dequeue_bits_decodeResult_readOnly;
  wire          _stage0_1_dequeue_bits_decodeResult_maskSource;
  wire          _stage0_1_dequeue_bits_decodeResult_maskDestination;
  wire          _stage0_1_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage0_1_dequeue_bits_decodeResult_uop;
  wire          _stage0_1_dequeue_bits_decodeResult_iota;
  wire          _stage0_1_dequeue_bits_decodeResult_mv;
  wire          _stage0_1_dequeue_bits_decodeResult_extend;
  wire          _stage0_1_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage0_1_dequeue_bits_decodeResult_compress;
  wire          _stage0_1_dequeue_bits_decodeResult_gather16;
  wire          _stage0_1_dequeue_bits_decodeResult_gather;
  wire          _stage0_1_dequeue_bits_decodeResult_slid;
  wire          _stage0_1_dequeue_bits_decodeResult_targetRd;
  wire          _stage0_1_dequeue_bits_decodeResult_widenReduce;
  wire          _stage0_1_dequeue_bits_decodeResult_red;
  wire          _stage0_1_dequeue_bits_decodeResult_nr;
  wire          _stage0_1_dequeue_bits_decodeResult_itype;
  wire          _stage0_1_dequeue_bits_decodeResult_unsigned1;
  wire          _stage0_1_dequeue_bits_decodeResult_unsigned0;
  wire          _stage0_1_dequeue_bits_decodeResult_other;
  wire          _stage0_1_dequeue_bits_decodeResult_multiCycle;
  wire          _stage0_1_dequeue_bits_decodeResult_divider;
  wire          _stage0_1_dequeue_bits_decodeResult_multiplier;
  wire          _stage0_1_dequeue_bits_decodeResult_shift;
  wire          _stage0_1_dequeue_bits_decodeResult_adder;
  wire          _stage0_1_dequeue_bits_decodeResult_logic;
  wire [1:0]    _stage0_1_dequeue_bits_laneIndex;
  wire          _stage0_1_dequeue_bits_skipRead;
  wire [4:0]    _stage0_1_dequeue_bits_vs1;
  wire [4:0]    _stage0_1_dequeue_bits_vs2;
  wire [4:0]    _stage0_1_dequeue_bits_vd;
  wire [2:0]    _stage0_1_dequeue_bits_vSew1H;
  wire          _stage0_1_dequeue_bits_maskNotMaskedElement;
  wire [13:0]   _stage0_1_dequeue_bits_csr_vl;
  wire [13:0]   _stage0_1_dequeue_bits_csr_vStart;
  wire [2:0]    _stage0_1_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage0_1_dequeue_bits_csr_vSew;
  wire [1:0]    _stage0_1_dequeue_bits_csr_vxrm;
  wire          _stage0_1_dequeue_bits_csr_vta;
  wire          _stage0_1_dequeue_bits_csr_vma;
  wire          _stage0_1_dequeue_bits_maskType;
  wire          _stage0_1_dequeue_bits_loadStore;
  wire          _stage0_1_dequeue_bits_bordersForMaskLogic;
  wire [7:0]    _stage0_1_updateLaneState_maskGroupCount;
  wire [4:0]    _stage0_1_updateLaneState_maskIndex;
  wire          _stage0_1_updateLaneState_outOfExecutionRange;
  wire          _stage0_1_updateLaneState_maskExhausted;
  wire          _stage0_1_tokenReport_valid;
  wire          _stage0_1_tokenReport_bits_decodeResult_sWrite;
  wire          _stage0_1_tokenReport_bits_decodeResult_maskUnit;
  wire [2:0]    _stage0_1_tokenReport_bits_instructionIndex;
  wire          _queue_fifo_1_empty;
  wire          _queue_fifo_1_full;
  wire          _queue_fifo_1_error;
  wire          _queue_fifo_empty;
  wire          _queue_fifo_full;
  wire          _queue_fifo_error;
  wire          _stage3_enqueue_ready;
  wire          _stage3_vrfWriteRequest_valid;
  wire [3:0]    _stage3_vrfWriteRequest_bits_mask;
  wire [2:0]    _stage3_vrfWriteRequest_bits_instructionIndex;
  wire          _stage3_crossWritePort_0_valid;
  wire          _stage3_crossWritePort_1_valid;
  wire          _maskStage_dequeue_valid;
  wire [9:0]    _maskStage_dequeue_bits_groupCounter;
  wire [31:0]   _maskStage_dequeue_bits_data;
  wire [31:0]   _maskStage_dequeue_bits_pipeData;
  wire [3:0]    _maskStage_dequeue_bits_mask;
  wire [10:0]   _maskStage_dequeue_bits_ffoIndex;
  wire [31:0]   _maskStage_dequeue_bits_crossWriteData_0;
  wire [31:0]   _maskStage_dequeue_bits_crossWriteData_1;
  wire          _maskStage_dequeue_bits_sSendResponse;
  wire          _maskStage_dequeue_bits_ffoSuccess;
  wire          _maskStage_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _maskStage_dequeue_bits_decodeResult_topUop;
  wire          _maskStage_dequeue_bits_decodeResult_popCount;
  wire          _maskStage_dequeue_bits_decodeResult_ffo;
  wire          _maskStage_dequeue_bits_decodeResult_average;
  wire          _maskStage_dequeue_bits_decodeResult_reverse;
  wire          _maskStage_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _maskStage_dequeue_bits_decodeResult_scheduler;
  wire          _maskStage_dequeue_bits_decodeResult_sReadVD;
  wire          _maskStage_dequeue_bits_decodeResult_vtype;
  wire          _maskStage_dequeue_bits_decodeResult_sWrite;
  wire          _maskStage_dequeue_bits_decodeResult_crossRead;
  wire          _maskStage_dequeue_bits_decodeResult_crossWrite;
  wire          _maskStage_dequeue_bits_decodeResult_maskUnit;
  wire          _maskStage_dequeue_bits_decodeResult_special;
  wire          _maskStage_dequeue_bits_decodeResult_saturate;
  wire          _maskStage_dequeue_bits_decodeResult_vwmacc;
  wire          _maskStage_dequeue_bits_decodeResult_readOnly;
  wire          _maskStage_dequeue_bits_decodeResult_maskSource;
  wire          _maskStage_dequeue_bits_decodeResult_maskDestination;
  wire          _maskStage_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _maskStage_dequeue_bits_decodeResult_uop;
  wire          _maskStage_dequeue_bits_decodeResult_iota;
  wire          _maskStage_dequeue_bits_decodeResult_mv;
  wire          _maskStage_dequeue_bits_decodeResult_extend;
  wire          _maskStage_dequeue_bits_decodeResult_unOrderWrite;
  wire          _maskStage_dequeue_bits_decodeResult_compress;
  wire          _maskStage_dequeue_bits_decodeResult_gather16;
  wire          _maskStage_dequeue_bits_decodeResult_gather;
  wire          _maskStage_dequeue_bits_decodeResult_slid;
  wire          _maskStage_dequeue_bits_decodeResult_targetRd;
  wire          _maskStage_dequeue_bits_decodeResult_widenReduce;
  wire          _maskStage_dequeue_bits_decodeResult_red;
  wire          _maskStage_dequeue_bits_decodeResult_nr;
  wire          _maskStage_dequeue_bits_decodeResult_itype;
  wire          _maskStage_dequeue_bits_decodeResult_unsigned1;
  wire          _maskStage_dequeue_bits_decodeResult_unsigned0;
  wire          _maskStage_dequeue_bits_decodeResult_other;
  wire          _maskStage_dequeue_bits_decodeResult_multiCycle;
  wire          _maskStage_dequeue_bits_decodeResult_divider;
  wire          _maskStage_dequeue_bits_decodeResult_multiplier;
  wire          _maskStage_dequeue_bits_decodeResult_shift;
  wire          _maskStage_dequeue_bits_decodeResult_adder;
  wire          _maskStage_dequeue_bits_decodeResult_logic;
  wire [2:0]    _maskStage_dequeue_bits_instructionIndex;
  wire          _maskStage_dequeue_bits_loadStore;
  wire [4:0]    _maskStage_dequeue_bits_vd;
  wire          _maskStage_maskReq_valid;
  wire [2:0]    _maskStage_maskReq_bits_index;
  wire          _executionUnit_enqueue_ready;
  wire          _executionUnit_dequeue_valid;
  wire          _executionUnit_vfuRequest_valid;
  wire [2:0]    _executionUnit_responseIndex;
  wire          _stage2_enqueue_ready;
  wire          _stage2_dequeue_valid;
  wire          _stage1_enqueue_ready;
  wire          _stage1_dequeue_valid;
  wire [3:0]    _stage1_dequeue_bits_maskForFilter;
  wire [3:0]    _stage1_dequeue_bits_mask;
  wire [9:0]    _stage1_dequeue_bits_groupCounter;
  wire          _stage1_dequeue_bits_sSendResponse;
  wire [31:0]   _stage1_dequeue_bits_src_0;
  wire [31:0]   _stage1_dequeue_bits_src_1;
  wire [31:0]   _stage1_dequeue_bits_src_2;
  wire [63:0]   _stage1_dequeue_bits_crossReadSource;
  wire          _stage1_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage1_dequeue_bits_decodeResult_topUop;
  wire          _stage1_dequeue_bits_decodeResult_popCount;
  wire          _stage1_dequeue_bits_decodeResult_ffo;
  wire          _stage1_dequeue_bits_decodeResult_average;
  wire          _stage1_dequeue_bits_decodeResult_reverse;
  wire          _stage1_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage1_dequeue_bits_decodeResult_scheduler;
  wire          _stage1_dequeue_bits_decodeResult_sReadVD;
  wire          _stage1_dequeue_bits_decodeResult_vtype;
  wire          _stage1_dequeue_bits_decodeResult_sWrite;
  wire          _stage1_dequeue_bits_decodeResult_crossRead;
  wire          _stage1_dequeue_bits_decodeResult_crossWrite;
  wire          _stage1_dequeue_bits_decodeResult_maskUnit;
  wire          _stage1_dequeue_bits_decodeResult_special;
  wire          _stage1_dequeue_bits_decodeResult_saturate;
  wire          _stage1_dequeue_bits_decodeResult_vwmacc;
  wire          _stage1_dequeue_bits_decodeResult_readOnly;
  wire          _stage1_dequeue_bits_decodeResult_maskSource;
  wire          _stage1_dequeue_bits_decodeResult_maskDestination;
  wire          _stage1_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage1_dequeue_bits_decodeResult_uop;
  wire          _stage1_dequeue_bits_decodeResult_iota;
  wire          _stage1_dequeue_bits_decodeResult_mv;
  wire          _stage1_dequeue_bits_decodeResult_extend;
  wire          _stage1_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage1_dequeue_bits_decodeResult_compress;
  wire          _stage1_dequeue_bits_decodeResult_gather16;
  wire          _stage1_dequeue_bits_decodeResult_gather;
  wire          _stage1_dequeue_bits_decodeResult_slid;
  wire          _stage1_dequeue_bits_decodeResult_targetRd;
  wire          _stage1_dequeue_bits_decodeResult_widenReduce;
  wire          _stage1_dequeue_bits_decodeResult_red;
  wire          _stage1_dequeue_bits_decodeResult_nr;
  wire          _stage1_dequeue_bits_decodeResult_itype;
  wire          _stage1_dequeue_bits_decodeResult_unsigned1;
  wire          _stage1_dequeue_bits_decodeResult_unsigned0;
  wire          _stage1_dequeue_bits_decodeResult_other;
  wire          _stage1_dequeue_bits_decodeResult_multiCycle;
  wire          _stage1_dequeue_bits_decodeResult_divider;
  wire          _stage1_dequeue_bits_decodeResult_multiplier;
  wire          _stage1_dequeue_bits_decodeResult_shift;
  wire          _stage1_dequeue_bits_decodeResult_adder;
  wire          _stage1_dequeue_bits_decodeResult_logic;
  wire [2:0]    _stage1_dequeue_bits_vSew1H;
  wire [13:0]   _stage1_dequeue_bits_csr_vl;
  wire [13:0]   _stage1_dequeue_bits_csr_vStart;
  wire [2:0]    _stage1_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage1_dequeue_bits_csr_vSew;
  wire [1:0]    _stage1_dequeue_bits_csr_vxrm;
  wire          _stage1_dequeue_bits_csr_vta;
  wire          _stage1_dequeue_bits_csr_vma;
  wire          _stage1_dequeue_bits_maskType;
  wire [1:0]    _stage1_dequeue_bits_laneIndex;
  wire [2:0]    _stage1_dequeue_bits_instructionIndex;
  wire          _stage1_dequeue_bits_loadStore;
  wire [4:0]    _stage1_dequeue_bits_vd;
  wire          _stage1_dequeue_bits_bordersForMaskLogic;
  wire          _stage1_readBusRequest_0_valid;
  wire          _stage1_readBusRequest_1_valid;
  wire          _stage0_enqueue_ready;
  wire          _stage0_dequeue_valid;
  wire [3:0]    _stage0_dequeue_bits_maskForMaskInput;
  wire [3:0]    _stage0_dequeue_bits_boundaryMaskCorrection;
  wire          _stage0_dequeue_bits_sSendResponse;
  wire [9:0]    _stage0_dequeue_bits_groupCounter;
  wire [31:0]   _stage0_dequeue_bits_readFromScalar;
  wire [2:0]    _stage0_dequeue_bits_instructionIndex;
  wire          _stage0_dequeue_bits_decodeResult_specialSlot;
  wire [4:0]    _stage0_dequeue_bits_decodeResult_topUop;
  wire          _stage0_dequeue_bits_decodeResult_popCount;
  wire          _stage0_dequeue_bits_decodeResult_ffo;
  wire          _stage0_dequeue_bits_decodeResult_average;
  wire          _stage0_dequeue_bits_decodeResult_reverse;
  wire          _stage0_dequeue_bits_decodeResult_dontNeedExecuteInLane;
  wire          _stage0_dequeue_bits_decodeResult_scheduler;
  wire          _stage0_dequeue_bits_decodeResult_sReadVD;
  wire          _stage0_dequeue_bits_decodeResult_vtype;
  wire          _stage0_dequeue_bits_decodeResult_sWrite;
  wire          _stage0_dequeue_bits_decodeResult_crossRead;
  wire          _stage0_dequeue_bits_decodeResult_crossWrite;
  wire          _stage0_dequeue_bits_decodeResult_maskUnit;
  wire          _stage0_dequeue_bits_decodeResult_special;
  wire          _stage0_dequeue_bits_decodeResult_saturate;
  wire          _stage0_dequeue_bits_decodeResult_vwmacc;
  wire          _stage0_dequeue_bits_decodeResult_readOnly;
  wire          _stage0_dequeue_bits_decodeResult_maskSource;
  wire          _stage0_dequeue_bits_decodeResult_maskDestination;
  wire          _stage0_dequeue_bits_decodeResult_maskLogic;
  wire [3:0]    _stage0_dequeue_bits_decodeResult_uop;
  wire          _stage0_dequeue_bits_decodeResult_iota;
  wire          _stage0_dequeue_bits_decodeResult_mv;
  wire          _stage0_dequeue_bits_decodeResult_extend;
  wire          _stage0_dequeue_bits_decodeResult_unOrderWrite;
  wire          _stage0_dequeue_bits_decodeResult_compress;
  wire          _stage0_dequeue_bits_decodeResult_gather16;
  wire          _stage0_dequeue_bits_decodeResult_gather;
  wire          _stage0_dequeue_bits_decodeResult_slid;
  wire          _stage0_dequeue_bits_decodeResult_targetRd;
  wire          _stage0_dequeue_bits_decodeResult_widenReduce;
  wire          _stage0_dequeue_bits_decodeResult_red;
  wire          _stage0_dequeue_bits_decodeResult_nr;
  wire          _stage0_dequeue_bits_decodeResult_itype;
  wire          _stage0_dequeue_bits_decodeResult_unsigned1;
  wire          _stage0_dequeue_bits_decodeResult_unsigned0;
  wire          _stage0_dequeue_bits_decodeResult_other;
  wire          _stage0_dequeue_bits_decodeResult_multiCycle;
  wire          _stage0_dequeue_bits_decodeResult_divider;
  wire          _stage0_dequeue_bits_decodeResult_multiplier;
  wire          _stage0_dequeue_bits_decodeResult_shift;
  wire          _stage0_dequeue_bits_decodeResult_adder;
  wire          _stage0_dequeue_bits_decodeResult_logic;
  wire [1:0]    _stage0_dequeue_bits_laneIndex;
  wire          _stage0_dequeue_bits_skipRead;
  wire [4:0]    _stage0_dequeue_bits_vs1;
  wire [4:0]    _stage0_dequeue_bits_vs2;
  wire [4:0]    _stage0_dequeue_bits_vd;
  wire [2:0]    _stage0_dequeue_bits_vSew1H;
  wire          _stage0_dequeue_bits_maskNotMaskedElement;
  wire [13:0]   _stage0_dequeue_bits_csr_vl;
  wire [13:0]   _stage0_dequeue_bits_csr_vStart;
  wire [2:0]    _stage0_dequeue_bits_csr_vlmul;
  wire [1:0]    _stage0_dequeue_bits_csr_vSew;
  wire [1:0]    _stage0_dequeue_bits_csr_vxrm;
  wire          _stage0_dequeue_bits_csr_vta;
  wire          _stage0_dequeue_bits_csr_vma;
  wire          _stage0_dequeue_bits_maskType;
  wire          _stage0_dequeue_bits_loadStore;
  wire          _stage0_dequeue_bits_bordersForMaskLogic;
  wire [7:0]    _stage0_updateLaneState_maskGroupCount;
  wire [4:0]    _stage0_updateLaneState_maskIndex;
  wire          _stage0_updateLaneState_outOfExecutionRange;
  wire          _stage0_updateLaneState_maskExhausted;
  wire          _stage0_tokenReport_valid;
  wire          _stage0_tokenReport_bits_decodeResult_sWrite;
  wire          _stage0_tokenReport_bits_decodeResult_crossWrite;
  wire          _stage0_tokenReport_bits_decodeResult_maskUnit;
  wire [2:0]    _stage0_tokenReport_bits_instructionIndex;
  wire          _stage0_tokenReport_bits_sSendResponse;
  wire [7:0]    _tokenManager_instructionValid;
  wire          _maskedWriteUnit_dequeue_valid;
  wire [4:0]    _maskedWriteUnit_dequeue_bits_vd;
  wire [5:0]    _maskedWriteUnit_dequeue_bits_offset;
  wire [3:0]    _maskedWriteUnit_dequeue_bits_mask;
  wire [31:0]   _maskedWriteUnit_dequeue_bits_data;
  wire          _maskedWriteUnit_dequeue_bits_last;
  wire [2:0]    _maskedWriteUnit_dequeue_bits_instructionIndex;
  wire          _crossLaneWriteQueue_fifo_1_empty;
  wire          _crossLaneWriteQueue_fifo_1_full;
  wire          _crossLaneWriteQueue_fifo_1_error;
  wire [50:0]   _crossLaneWriteQueue_fifo_1_data_out;
  wire          _crossLaneWriteQueue_fifo_empty;
  wire          _crossLaneWriteQueue_fifo_full;
  wire          _crossLaneWriteQueue_fifo_error;
  wire [50:0]   _crossLaneWriteQueue_fifo_data_out;
  wire          _vrf_readRequests_0_ready;
  wire          _vrf_readRequests_1_ready;
  wire          _vrf_readRequests_2_ready;
  wire          _vrf_readRequests_3_ready;
  wire          _vrf_readRequests_4_ready;
  wire          _vrf_readRequests_5_ready;
  wire          _vrf_readRequests_6_ready;
  wire          _vrf_readRequests_7_ready;
  wire          _vrf_readRequests_8_ready;
  wire          _vrf_readRequests_9_ready;
  wire          _vrf_readRequests_10_ready;
  wire          _vrf_readRequests_11_ready;
  wire          _vrf_readRequests_12_ready;
  wire          _vrf_readRequests_13_ready;
  wire [31:0]   _vrf_readResults_0;
  wire          _vrf_write_ready;
  wire          _vrf_writeAllow_0;
  wire          _vrf_writeAllow_1;
  wire          _vrf_writeAllow_2;
  wire          _vrf_writeAllow_3;
  wire          _vrf_writeAllow_4;
  wire          _vrf_writeAllow_5;
  wire          _vrf_writeAllow_6;
  wire [7:0]    _vrf_vrfSlotRelease;
  wire          vrfReadAddressChannel_ready_0;
  wire [1:0]    vfuResponse_responseBundle_2_bits_tag;
  wire          vfuResponse_responseBundle_2_bits_ffoSuccess;
  wire          vfuResponse_responseBundle_2_bits_clipFail;
  wire [31:0]   vfuResponse_responseBundle_2_bits_data;
  wire          vfuResponse_responseBundle_2_valid;
  wire [1:0]    vfuResponse_responseBundle_1_bits_tag;
  wire [1:0]    vfuResponse_responseBundle_1_bits_executeIndex;
  wire [31:0]   vfuResponse_responseBundle_1_bits_data;
  wire          vfuResponse_responseBundle_1_valid;
  wire [1:0]    vfuResponse_responseBundle_bits_tag;
  wire [31:0]   vfuResponse_responseBundle_bits_data;
  wire          vfuResponse_responseBundle_valid;
  wire [10:0]   stage3EnqWire_3_bits_ffoIndex;
  wire [31:0]   stage3EnqWire_3_bits_data;
  wire          responseDecodeVec_3_multiCycle;
  wire          responseDecodeVec_3_unsigned0;
  wire          responseDecodeVec_3_unsigned1;
  wire          responseDecodeVec_3_itype;
  wire          responseDecodeVec_3_nr;
  wire          responseDecodeVec_3_red;
  wire          responseDecodeVec_3_widenReduce;
  wire          responseDecodeVec_3_targetRd;
  wire          responseDecodeVec_3_slid;
  wire          responseDecodeVec_3_gather;
  wire          responseDecodeVec_3_gather16;
  wire          responseDecodeVec_3_compress;
  wire          responseDecodeVec_3_unOrderWrite;
  wire          responseDecodeVec_3_extend;
  wire          responseDecodeVec_3_mv;
  wire          responseDecodeVec_3_iota;
  wire [3:0]    responseDecodeVec_3_uop;
  wire          responseDecodeVec_3_maskLogic;
  wire          responseDecodeVec_3_maskDestination;
  wire          responseDecodeVec_3_maskSource;
  wire          responseDecodeVec_3_readOnly;
  wire          responseDecodeVec_3_vwmacc;
  wire          responseDecodeVec_3_saturate;
  wire          responseDecodeVec_3_special;
  wire          responseDecodeVec_3_maskUnit;
  wire          responseDecodeVec_3_crossWrite;
  wire          responseDecodeVec_3_crossRead;
  wire          responseDecodeVec_3_sWrite;
  wire          responseDecodeVec_3_vtype;
  wire          responseDecodeVec_3_sReadVD;
  wire          responseDecodeVec_3_scheduler;
  wire          responseDecodeVec_3_dontNeedExecuteInLane;
  wire          responseDecodeVec_3_reverse;
  wire          responseDecodeVec_3_average;
  wire          responseDecodeVec_3_ffo;
  wire          responseDecodeVec_3_popCount;
  wire [4:0]    responseDecodeVec_3_topUop;
  wire          responseDecodeVec_3_specialSlot;
  wire          executeDecodeVec_3_multiCycle;
  wire          executeDecodeVec_3_unsigned0;
  wire          executeDecodeVec_3_unsigned1;
  wire          executeDecodeVec_3_itype;
  wire          executeDecodeVec_3_nr;
  wire          executeDecodeVec_3_red;
  wire          executeDecodeVec_3_widenReduce;
  wire          executeDecodeVec_3_targetRd;
  wire          executeDecodeVec_3_slid;
  wire          executeDecodeVec_3_gather;
  wire          executeDecodeVec_3_gather16;
  wire          executeDecodeVec_3_compress;
  wire          executeDecodeVec_3_unOrderWrite;
  wire          executeDecodeVec_3_extend;
  wire          executeDecodeVec_3_mv;
  wire          executeDecodeVec_3_iota;
  wire [3:0]    executeDecodeVec_3_uop;
  wire          executeDecodeVec_3_maskLogic;
  wire          executeDecodeVec_3_maskDestination;
  wire          executeDecodeVec_3_maskSource;
  wire          executeDecodeVec_3_readOnly;
  wire          executeDecodeVec_3_vwmacc;
  wire          executeDecodeVec_3_saturate;
  wire          executeDecodeVec_3_special;
  wire          executeDecodeVec_3_maskUnit;
  wire          executeDecodeVec_3_crossWrite;
  wire          executeDecodeVec_3_crossRead;
  wire          executeDecodeVec_3_sWrite;
  wire          executeDecodeVec_3_vtype;
  wire          executeDecodeVec_3_sReadVD;
  wire          executeDecodeVec_3_scheduler;
  wire          executeDecodeVec_3_dontNeedExecuteInLane;
  wire          executeDecodeVec_3_reverse;
  wire          executeDecodeVec_3_average;
  wire          executeDecodeVec_3_ffo;
  wire          executeDecodeVec_3_popCount;
  wire [4:0]    executeDecodeVec_3_topUop;
  wire          executeDecodeVec_3_specialSlot;
  wire [4:0]    stage3EnqWire_3_bits_vd;
  wire          stage3EnqWire_3_bits_loadStore;
  wire [2:0]    stage3EnqWire_3_bits_instructionIndex;
  wire          stage3EnqWire_3_bits_decodeResult_logic;
  wire          stage3EnqWire_3_bits_decodeResult_adder;
  wire          stage3EnqWire_3_bits_decodeResult_shift;
  wire          stage3EnqWire_3_bits_decodeResult_multiplier;
  wire          stage3EnqWire_3_bits_decodeResult_divider;
  wire          stage3EnqWire_3_bits_decodeResult_multiCycle;
  wire          stage3EnqWire_3_bits_decodeResult_other;
  wire          stage3EnqWire_3_bits_decodeResult_unsigned0;
  wire          stage3EnqWire_3_bits_decodeResult_unsigned1;
  wire          stage3EnqWire_3_bits_decodeResult_itype;
  wire          stage3EnqWire_3_bits_decodeResult_nr;
  wire          stage3EnqWire_3_bits_decodeResult_red;
  wire          stage3EnqWire_3_bits_decodeResult_widenReduce;
  wire          stage3EnqWire_3_bits_decodeResult_targetRd;
  wire          stage3EnqWire_3_bits_decodeResult_slid;
  wire          stage3EnqWire_3_bits_decodeResult_gather;
  wire          stage3EnqWire_3_bits_decodeResult_gather16;
  wire          stage3EnqWire_3_bits_decodeResult_compress;
  wire          stage3EnqWire_3_bits_decodeResult_unOrderWrite;
  wire          stage3EnqWire_3_bits_decodeResult_extend;
  wire          stage3EnqWire_3_bits_decodeResult_mv;
  wire          stage3EnqWire_3_bits_decodeResult_iota;
  wire [3:0]    stage3EnqWire_3_bits_decodeResult_uop;
  wire          stage3EnqWire_3_bits_decodeResult_maskLogic;
  wire          stage3EnqWire_3_bits_decodeResult_maskDestination;
  wire          stage3EnqWire_3_bits_decodeResult_maskSource;
  wire          stage3EnqWire_3_bits_decodeResult_readOnly;
  wire          stage3EnqWire_3_bits_decodeResult_vwmacc;
  wire          stage3EnqWire_3_bits_decodeResult_saturate;
  wire          stage3EnqWire_3_bits_decodeResult_special;
  wire          stage3EnqWire_3_bits_decodeResult_maskUnit;
  wire          stage3EnqWire_3_bits_decodeResult_crossWrite;
  wire          stage3EnqWire_3_bits_decodeResult_crossRead;
  wire          stage3EnqWire_3_bits_decodeResult_sWrite;
  wire          stage3EnqWire_3_bits_decodeResult_vtype;
  wire          stage3EnqWire_3_bits_decodeResult_sReadVD;
  wire          stage3EnqWire_3_bits_decodeResult_scheduler;
  wire          stage3EnqWire_3_bits_decodeResult_dontNeedExecuteInLane;
  wire          stage3EnqWire_3_bits_decodeResult_reverse;
  wire          stage3EnqWire_3_bits_decodeResult_average;
  wire          stage3EnqWire_3_bits_decodeResult_ffo;
  wire          stage3EnqWire_3_bits_decodeResult_popCount;
  wire [4:0]    stage3EnqWire_3_bits_decodeResult_topUop;
  wire          stage3EnqWire_3_bits_decodeResult_specialSlot;
  wire [3:0]    stage3EnqWire_3_bits_mask;
  wire [9:0]    stage3EnqWire_3_bits_groupCounter;
  wire [1:0]    readCheckRequestVec_2_readSource;
  wire [1:0]    readCheckRequestVec_1_readSource;
  wire [1:0]    readCheckRequestVec_0_readSource;
  wire [2:0]    vrfReadRequest_3_2_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_3_2_bits_offset;
  wire [1:0]    vrfReadRequest_3_2_bits_readSource;
  wire [4:0]    vrfReadRequest_3_2_bits_vs;
  wire          vrfReadRequest_3_2_valid;
  wire [2:0]    vrfReadRequest_3_1_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_3_1_bits_offset;
  wire [1:0]    vrfReadRequest_3_1_bits_readSource;
  wire [4:0]    vrfReadRequest_3_1_bits_vs;
  wire          vrfReadRequest_3_1_valid;
  wire [2:0]    vrfReadRequest_3_0_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_3_0_bits_offset;
  wire [1:0]    vrfReadRequest_3_0_bits_readSource;
  wire [4:0]    vrfReadRequest_3_0_bits_vs;
  wire          vrfReadRequest_3_0_valid;
  wire [10:0]   stage3EnqWire_2_bits_ffoIndex;
  wire [31:0]   stage3EnqWire_2_bits_data;
  wire          responseDecodeVec_2_multiCycle;
  wire          responseDecodeVec_2_unsigned0;
  wire          responseDecodeVec_2_unsigned1;
  wire          responseDecodeVec_2_itype;
  wire          responseDecodeVec_2_nr;
  wire          responseDecodeVec_2_red;
  wire          responseDecodeVec_2_widenReduce;
  wire          responseDecodeVec_2_targetRd;
  wire          responseDecodeVec_2_slid;
  wire          responseDecodeVec_2_gather;
  wire          responseDecodeVec_2_gather16;
  wire          responseDecodeVec_2_compress;
  wire          responseDecodeVec_2_unOrderWrite;
  wire          responseDecodeVec_2_extend;
  wire          responseDecodeVec_2_mv;
  wire          responseDecodeVec_2_iota;
  wire [3:0]    responseDecodeVec_2_uop;
  wire          responseDecodeVec_2_maskLogic;
  wire          responseDecodeVec_2_maskDestination;
  wire          responseDecodeVec_2_maskSource;
  wire          responseDecodeVec_2_readOnly;
  wire          responseDecodeVec_2_vwmacc;
  wire          responseDecodeVec_2_saturate;
  wire          responseDecodeVec_2_special;
  wire          responseDecodeVec_2_maskUnit;
  wire          responseDecodeVec_2_crossWrite;
  wire          responseDecodeVec_2_crossRead;
  wire          responseDecodeVec_2_sWrite;
  wire          responseDecodeVec_2_vtype;
  wire          responseDecodeVec_2_sReadVD;
  wire          responseDecodeVec_2_scheduler;
  wire          responseDecodeVec_2_dontNeedExecuteInLane;
  wire          responseDecodeVec_2_reverse;
  wire          responseDecodeVec_2_average;
  wire          responseDecodeVec_2_ffo;
  wire          responseDecodeVec_2_popCount;
  wire [4:0]    responseDecodeVec_2_topUop;
  wire          responseDecodeVec_2_specialSlot;
  wire          executeDecodeVec_2_multiCycle;
  wire          executeDecodeVec_2_unsigned0;
  wire          executeDecodeVec_2_unsigned1;
  wire          executeDecodeVec_2_itype;
  wire          executeDecodeVec_2_nr;
  wire          executeDecodeVec_2_red;
  wire          executeDecodeVec_2_widenReduce;
  wire          executeDecodeVec_2_targetRd;
  wire          executeDecodeVec_2_slid;
  wire          executeDecodeVec_2_gather;
  wire          executeDecodeVec_2_gather16;
  wire          executeDecodeVec_2_compress;
  wire          executeDecodeVec_2_unOrderWrite;
  wire          executeDecodeVec_2_extend;
  wire          executeDecodeVec_2_mv;
  wire          executeDecodeVec_2_iota;
  wire [3:0]    executeDecodeVec_2_uop;
  wire          executeDecodeVec_2_maskLogic;
  wire          executeDecodeVec_2_maskDestination;
  wire          executeDecodeVec_2_maskSource;
  wire          executeDecodeVec_2_readOnly;
  wire          executeDecodeVec_2_vwmacc;
  wire          executeDecodeVec_2_saturate;
  wire          executeDecodeVec_2_special;
  wire          executeDecodeVec_2_maskUnit;
  wire          executeDecodeVec_2_crossWrite;
  wire          executeDecodeVec_2_crossRead;
  wire          executeDecodeVec_2_sWrite;
  wire          executeDecodeVec_2_vtype;
  wire          executeDecodeVec_2_sReadVD;
  wire          executeDecodeVec_2_scheduler;
  wire          executeDecodeVec_2_dontNeedExecuteInLane;
  wire          executeDecodeVec_2_reverse;
  wire          executeDecodeVec_2_average;
  wire          executeDecodeVec_2_ffo;
  wire          executeDecodeVec_2_popCount;
  wire [4:0]    executeDecodeVec_2_topUop;
  wire          executeDecodeVec_2_specialSlot;
  wire [4:0]    stage3EnqWire_2_bits_vd;
  wire          stage3EnqWire_2_bits_loadStore;
  wire [2:0]    stage3EnqWire_2_bits_instructionIndex;
  wire          stage3EnqWire_2_bits_decodeResult_logic;
  wire          stage3EnqWire_2_bits_decodeResult_adder;
  wire          stage3EnqWire_2_bits_decodeResult_shift;
  wire          stage3EnqWire_2_bits_decodeResult_multiplier;
  wire          stage3EnqWire_2_bits_decodeResult_divider;
  wire          stage3EnqWire_2_bits_decodeResult_multiCycle;
  wire          stage3EnqWire_2_bits_decodeResult_other;
  wire          stage3EnqWire_2_bits_decodeResult_unsigned0;
  wire          stage3EnqWire_2_bits_decodeResult_unsigned1;
  wire          stage3EnqWire_2_bits_decodeResult_itype;
  wire          stage3EnqWire_2_bits_decodeResult_nr;
  wire          stage3EnqWire_2_bits_decodeResult_red;
  wire          stage3EnqWire_2_bits_decodeResult_widenReduce;
  wire          stage3EnqWire_2_bits_decodeResult_targetRd;
  wire          stage3EnqWire_2_bits_decodeResult_slid;
  wire          stage3EnqWire_2_bits_decodeResult_gather;
  wire          stage3EnqWire_2_bits_decodeResult_gather16;
  wire          stage3EnqWire_2_bits_decodeResult_compress;
  wire          stage3EnqWire_2_bits_decodeResult_unOrderWrite;
  wire          stage3EnqWire_2_bits_decodeResult_extend;
  wire          stage3EnqWire_2_bits_decodeResult_mv;
  wire          stage3EnqWire_2_bits_decodeResult_iota;
  wire [3:0]    stage3EnqWire_2_bits_decodeResult_uop;
  wire          stage3EnqWire_2_bits_decodeResult_maskLogic;
  wire          stage3EnqWire_2_bits_decodeResult_maskDestination;
  wire          stage3EnqWire_2_bits_decodeResult_maskSource;
  wire          stage3EnqWire_2_bits_decodeResult_readOnly;
  wire          stage3EnqWire_2_bits_decodeResult_vwmacc;
  wire          stage3EnqWire_2_bits_decodeResult_saturate;
  wire          stage3EnqWire_2_bits_decodeResult_special;
  wire          stage3EnqWire_2_bits_decodeResult_maskUnit;
  wire          stage3EnqWire_2_bits_decodeResult_crossWrite;
  wire          stage3EnqWire_2_bits_decodeResult_crossRead;
  wire          stage3EnqWire_2_bits_decodeResult_sWrite;
  wire          stage3EnqWire_2_bits_decodeResult_vtype;
  wire          stage3EnqWire_2_bits_decodeResult_sReadVD;
  wire          stage3EnqWire_2_bits_decodeResult_scheduler;
  wire          stage3EnqWire_2_bits_decodeResult_dontNeedExecuteInLane;
  wire          stage3EnqWire_2_bits_decodeResult_reverse;
  wire          stage3EnqWire_2_bits_decodeResult_average;
  wire          stage3EnqWire_2_bits_decodeResult_ffo;
  wire          stage3EnqWire_2_bits_decodeResult_popCount;
  wire [4:0]    stage3EnqWire_2_bits_decodeResult_topUop;
  wire          stage3EnqWire_2_bits_decodeResult_specialSlot;
  wire [3:0]    stage3EnqWire_2_bits_mask;
  wire [9:0]    stage3EnqWire_2_bits_groupCounter;
  wire [1:0]    readCheckRequestVec_5_readSource;
  wire [1:0]    readCheckRequestVec_4_readSource;
  wire [1:0]    readCheckRequestVec_3_readSource;
  wire [2:0]    vrfReadRequest_2_2_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_2_2_bits_offset;
  wire [1:0]    vrfReadRequest_2_2_bits_readSource;
  wire [4:0]    vrfReadRequest_2_2_bits_vs;
  wire          vrfReadRequest_2_2_valid;
  wire [2:0]    vrfReadRequest_2_1_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_2_1_bits_offset;
  wire [1:0]    vrfReadRequest_2_1_bits_readSource;
  wire [4:0]    vrfReadRequest_2_1_bits_vs;
  wire          vrfReadRequest_2_1_valid;
  wire [2:0]    vrfReadRequest_2_0_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_2_0_bits_offset;
  wire [1:0]    vrfReadRequest_2_0_bits_readSource;
  wire [4:0]    vrfReadRequest_2_0_bits_vs;
  wire          vrfReadRequest_2_0_valid;
  wire [10:0]   stage3EnqWire_1_bits_ffoIndex;
  wire [31:0]   stage3EnqWire_1_bits_data;
  wire          responseDecodeVec_1_multiCycle;
  wire          responseDecodeVec_1_unsigned0;
  wire          responseDecodeVec_1_unsigned1;
  wire          responseDecodeVec_1_itype;
  wire          responseDecodeVec_1_nr;
  wire          responseDecodeVec_1_red;
  wire          responseDecodeVec_1_widenReduce;
  wire          responseDecodeVec_1_targetRd;
  wire          responseDecodeVec_1_slid;
  wire          responseDecodeVec_1_gather;
  wire          responseDecodeVec_1_gather16;
  wire          responseDecodeVec_1_compress;
  wire          responseDecodeVec_1_unOrderWrite;
  wire          responseDecodeVec_1_extend;
  wire          responseDecodeVec_1_mv;
  wire          responseDecodeVec_1_iota;
  wire [3:0]    responseDecodeVec_1_uop;
  wire          responseDecodeVec_1_maskLogic;
  wire          responseDecodeVec_1_maskDestination;
  wire          responseDecodeVec_1_maskSource;
  wire          responseDecodeVec_1_readOnly;
  wire          responseDecodeVec_1_vwmacc;
  wire          responseDecodeVec_1_saturate;
  wire          responseDecodeVec_1_special;
  wire          responseDecodeVec_1_maskUnit;
  wire          responseDecodeVec_1_crossWrite;
  wire          responseDecodeVec_1_crossRead;
  wire          responseDecodeVec_1_sWrite;
  wire          responseDecodeVec_1_vtype;
  wire          responseDecodeVec_1_sReadVD;
  wire          responseDecodeVec_1_scheduler;
  wire          responseDecodeVec_1_dontNeedExecuteInLane;
  wire          responseDecodeVec_1_reverse;
  wire          responseDecodeVec_1_average;
  wire          responseDecodeVec_1_ffo;
  wire          responseDecodeVec_1_popCount;
  wire [4:0]    responseDecodeVec_1_topUop;
  wire          responseDecodeVec_1_specialSlot;
  wire          executeDecodeVec_1_multiCycle;
  wire          executeDecodeVec_1_unsigned0;
  wire          executeDecodeVec_1_unsigned1;
  wire          executeDecodeVec_1_itype;
  wire          executeDecodeVec_1_nr;
  wire          executeDecodeVec_1_red;
  wire          executeDecodeVec_1_widenReduce;
  wire          executeDecodeVec_1_targetRd;
  wire          executeDecodeVec_1_slid;
  wire          executeDecodeVec_1_gather;
  wire          executeDecodeVec_1_gather16;
  wire          executeDecodeVec_1_compress;
  wire          executeDecodeVec_1_unOrderWrite;
  wire          executeDecodeVec_1_extend;
  wire          executeDecodeVec_1_mv;
  wire          executeDecodeVec_1_iota;
  wire [3:0]    executeDecodeVec_1_uop;
  wire          executeDecodeVec_1_maskLogic;
  wire          executeDecodeVec_1_maskDestination;
  wire          executeDecodeVec_1_maskSource;
  wire          executeDecodeVec_1_readOnly;
  wire          executeDecodeVec_1_vwmacc;
  wire          executeDecodeVec_1_saturate;
  wire          executeDecodeVec_1_special;
  wire          executeDecodeVec_1_maskUnit;
  wire          executeDecodeVec_1_crossWrite;
  wire          executeDecodeVec_1_crossRead;
  wire          executeDecodeVec_1_sWrite;
  wire          executeDecodeVec_1_vtype;
  wire          executeDecodeVec_1_sReadVD;
  wire          executeDecodeVec_1_scheduler;
  wire          executeDecodeVec_1_dontNeedExecuteInLane;
  wire          executeDecodeVec_1_reverse;
  wire          executeDecodeVec_1_average;
  wire          executeDecodeVec_1_ffo;
  wire          executeDecodeVec_1_popCount;
  wire [4:0]    executeDecodeVec_1_topUop;
  wire          executeDecodeVec_1_specialSlot;
  wire [4:0]    stage3EnqWire_1_bits_vd;
  wire          stage3EnqWire_1_bits_loadStore;
  wire [2:0]    stage3EnqWire_1_bits_instructionIndex;
  wire          stage3EnqWire_1_bits_decodeResult_logic;
  wire          stage3EnqWire_1_bits_decodeResult_adder;
  wire          stage3EnqWire_1_bits_decodeResult_shift;
  wire          stage3EnqWire_1_bits_decodeResult_multiplier;
  wire          stage3EnqWire_1_bits_decodeResult_divider;
  wire          stage3EnqWire_1_bits_decodeResult_multiCycle;
  wire          stage3EnqWire_1_bits_decodeResult_other;
  wire          stage3EnqWire_1_bits_decodeResult_unsigned0;
  wire          stage3EnqWire_1_bits_decodeResult_unsigned1;
  wire          stage3EnqWire_1_bits_decodeResult_itype;
  wire          stage3EnqWire_1_bits_decodeResult_nr;
  wire          stage3EnqWire_1_bits_decodeResult_red;
  wire          stage3EnqWire_1_bits_decodeResult_widenReduce;
  wire          stage3EnqWire_1_bits_decodeResult_targetRd;
  wire          stage3EnqWire_1_bits_decodeResult_slid;
  wire          stage3EnqWire_1_bits_decodeResult_gather;
  wire          stage3EnqWire_1_bits_decodeResult_gather16;
  wire          stage3EnqWire_1_bits_decodeResult_compress;
  wire          stage3EnqWire_1_bits_decodeResult_unOrderWrite;
  wire          stage3EnqWire_1_bits_decodeResult_extend;
  wire          stage3EnqWire_1_bits_decodeResult_mv;
  wire          stage3EnqWire_1_bits_decodeResult_iota;
  wire [3:0]    stage3EnqWire_1_bits_decodeResult_uop;
  wire          stage3EnqWire_1_bits_decodeResult_maskLogic;
  wire          stage3EnqWire_1_bits_decodeResult_maskDestination;
  wire          stage3EnqWire_1_bits_decodeResult_maskSource;
  wire          stage3EnqWire_1_bits_decodeResult_readOnly;
  wire          stage3EnqWire_1_bits_decodeResult_vwmacc;
  wire          stage3EnqWire_1_bits_decodeResult_saturate;
  wire          stage3EnqWire_1_bits_decodeResult_special;
  wire          stage3EnqWire_1_bits_decodeResult_maskUnit;
  wire          stage3EnqWire_1_bits_decodeResult_crossWrite;
  wire          stage3EnqWire_1_bits_decodeResult_crossRead;
  wire          stage3EnqWire_1_bits_decodeResult_sWrite;
  wire          stage3EnqWire_1_bits_decodeResult_vtype;
  wire          stage3EnqWire_1_bits_decodeResult_sReadVD;
  wire          stage3EnqWire_1_bits_decodeResult_scheduler;
  wire          stage3EnqWire_1_bits_decodeResult_dontNeedExecuteInLane;
  wire          stage3EnqWire_1_bits_decodeResult_reverse;
  wire          stage3EnqWire_1_bits_decodeResult_average;
  wire          stage3EnqWire_1_bits_decodeResult_ffo;
  wire          stage3EnqWire_1_bits_decodeResult_popCount;
  wire [4:0]    stage3EnqWire_1_bits_decodeResult_topUop;
  wire          stage3EnqWire_1_bits_decodeResult_specialSlot;
  wire [3:0]    stage3EnqWire_1_bits_mask;
  wire [9:0]    stage3EnqWire_1_bits_groupCounter;
  wire [1:0]    readCheckRequestVec_8_readSource;
  wire [1:0]    readCheckRequestVec_7_readSource;
  wire [1:0]    readCheckRequestVec_6_readSource;
  wire [2:0]    vrfReadRequest_1_2_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_1_2_bits_offset;
  wire [1:0]    vrfReadRequest_1_2_bits_readSource;
  wire [4:0]    vrfReadRequest_1_2_bits_vs;
  wire          vrfReadRequest_1_2_valid;
  wire [2:0]    vrfReadRequest_1_1_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_1_1_bits_offset;
  wire [1:0]    vrfReadRequest_1_1_bits_readSource;
  wire [4:0]    vrfReadRequest_1_1_bits_vs;
  wire          vrfReadRequest_1_1_valid;
  wire [2:0]    vrfReadRequest_1_0_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_1_0_bits_offset;
  wire [1:0]    vrfReadRequest_1_0_bits_readSource;
  wire [4:0]    vrfReadRequest_1_0_bits_vs;
  wire          vrfReadRequest_1_0_valid;
  wire          queue_1_almostFull;
  wire          queue_1_almostEmpty;
  wire          queue_almostFull;
  wire          queue_almostEmpty;
  wire [9:0]    writeBusPort_1_deq_bits_counter_0;
  wire [2:0]    writeBusPort_1_deq_bits_instructionIndex_0;
  wire [1:0]    writeBusPort_1_deq_bits_mask_0;
  wire [31:0]   writeBusPort_1_deq_bits_data_0;
  wire [9:0]    writeBusPort_0_deq_bits_counter_0;
  wire [2:0]    writeBusPort_0_deq_bits_instructionIndex_0;
  wire [1:0]    writeBusPort_0_deq_bits_mask_0;
  wire [31:0]   writeBusPort_0_deq_bits_data_0;
  wire          stage3EnqWire_bits_ffoSuccess;
  wire [31:0]   stage3EnqWire_bits_crossWriteData_1;
  wire [31:0]   stage3EnqWire_bits_crossWriteData_0;
  wire [10:0]   stage3EnqWire_bits_ffoIndex;
  wire [31:0]   stage3EnqWire_bits_data;
  wire          responseDecodeVec_0_multiCycle;
  wire          responseDecodeVec_0_unsigned0;
  wire          responseDecodeVec_0_unsigned1;
  wire          responseDecodeVec_0_itype;
  wire          responseDecodeVec_0_nr;
  wire          responseDecodeVec_0_red;
  wire          responseDecodeVec_0_widenReduce;
  wire          responseDecodeVec_0_targetRd;
  wire          responseDecodeVec_0_slid;
  wire          responseDecodeVec_0_gather;
  wire          responseDecodeVec_0_gather16;
  wire          responseDecodeVec_0_compress;
  wire          responseDecodeVec_0_unOrderWrite;
  wire          responseDecodeVec_0_extend;
  wire          responseDecodeVec_0_mv;
  wire          responseDecodeVec_0_iota;
  wire [3:0]    responseDecodeVec_0_uop;
  wire          responseDecodeVec_0_maskLogic;
  wire          responseDecodeVec_0_maskDestination;
  wire          responseDecodeVec_0_maskSource;
  wire          responseDecodeVec_0_readOnly;
  wire          responseDecodeVec_0_vwmacc;
  wire          responseDecodeVec_0_saturate;
  wire          responseDecodeVec_0_special;
  wire          responseDecodeVec_0_maskUnit;
  wire          responseDecodeVec_0_crossWrite;
  wire          responseDecodeVec_0_crossRead;
  wire          responseDecodeVec_0_sWrite;
  wire          responseDecodeVec_0_vtype;
  wire          responseDecodeVec_0_sReadVD;
  wire          responseDecodeVec_0_scheduler;
  wire          responseDecodeVec_0_dontNeedExecuteInLane;
  wire          responseDecodeVec_0_reverse;
  wire          responseDecodeVec_0_average;
  wire          responseDecodeVec_0_ffo;
  wire          responseDecodeVec_0_popCount;
  wire [4:0]    responseDecodeVec_0_topUop;
  wire          responseDecodeVec_0_specialSlot;
  wire          executeDecodeVec_0_multiCycle;
  wire          executeDecodeVec_0_unsigned0;
  wire          executeDecodeVec_0_unsigned1;
  wire          executeDecodeVec_0_itype;
  wire          executeDecodeVec_0_nr;
  wire          executeDecodeVec_0_red;
  wire          executeDecodeVec_0_widenReduce;
  wire          executeDecodeVec_0_targetRd;
  wire          executeDecodeVec_0_slid;
  wire          executeDecodeVec_0_gather;
  wire          executeDecodeVec_0_gather16;
  wire          executeDecodeVec_0_compress;
  wire          executeDecodeVec_0_unOrderWrite;
  wire          executeDecodeVec_0_extend;
  wire          executeDecodeVec_0_mv;
  wire          executeDecodeVec_0_iota;
  wire [3:0]    executeDecodeVec_0_uop;
  wire          executeDecodeVec_0_maskLogic;
  wire          executeDecodeVec_0_maskDestination;
  wire          executeDecodeVec_0_maskSource;
  wire          executeDecodeVec_0_readOnly;
  wire          executeDecodeVec_0_vwmacc;
  wire          executeDecodeVec_0_saturate;
  wire          executeDecodeVec_0_special;
  wire          executeDecodeVec_0_maskUnit;
  wire          executeDecodeVec_0_crossWrite;
  wire          executeDecodeVec_0_crossRead;
  wire          executeDecodeVec_0_sWrite;
  wire          executeDecodeVec_0_vtype;
  wire          executeDecodeVec_0_sReadVD;
  wire          executeDecodeVec_0_scheduler;
  wire          executeDecodeVec_0_dontNeedExecuteInLane;
  wire          executeDecodeVec_0_reverse;
  wire          executeDecodeVec_0_average;
  wire          executeDecodeVec_0_ffo;
  wire          executeDecodeVec_0_popCount;
  wire [4:0]    executeDecodeVec_0_topUop;
  wire          executeDecodeVec_0_specialSlot;
  wire [4:0]    stage3EnqWire_bits_vd;
  wire          stage3EnqWire_bits_loadStore;
  wire [2:0]    stage3EnqWire_bits_instructionIndex;
  wire          stage3EnqWire_bits_decodeResult_logic;
  wire          stage3EnqWire_bits_decodeResult_adder;
  wire          stage3EnqWire_bits_decodeResult_shift;
  wire          stage3EnqWire_bits_decodeResult_multiplier;
  wire          stage3EnqWire_bits_decodeResult_divider;
  wire          stage3EnqWire_bits_decodeResult_multiCycle;
  wire          stage3EnqWire_bits_decodeResult_other;
  wire          stage3EnqWire_bits_decodeResult_unsigned0;
  wire          stage3EnqWire_bits_decodeResult_unsigned1;
  wire          stage3EnqWire_bits_decodeResult_itype;
  wire          stage3EnqWire_bits_decodeResult_nr;
  wire          stage3EnqWire_bits_decodeResult_red;
  wire          stage3EnqWire_bits_decodeResult_widenReduce;
  wire          stage3EnqWire_bits_decodeResult_targetRd;
  wire          stage3EnqWire_bits_decodeResult_slid;
  wire          stage3EnqWire_bits_decodeResult_gather;
  wire          stage3EnqWire_bits_decodeResult_gather16;
  wire          stage3EnqWire_bits_decodeResult_compress;
  wire          stage3EnqWire_bits_decodeResult_unOrderWrite;
  wire          stage3EnqWire_bits_decodeResult_extend;
  wire          stage3EnqWire_bits_decodeResult_mv;
  wire          stage3EnqWire_bits_decodeResult_iota;
  wire [3:0]    stage3EnqWire_bits_decodeResult_uop;
  wire          stage3EnqWire_bits_decodeResult_maskLogic;
  wire          stage3EnqWire_bits_decodeResult_maskDestination;
  wire          stage3EnqWire_bits_decodeResult_maskSource;
  wire          stage3EnqWire_bits_decodeResult_readOnly;
  wire          stage3EnqWire_bits_decodeResult_vwmacc;
  wire          stage3EnqWire_bits_decodeResult_saturate;
  wire          stage3EnqWire_bits_decodeResult_special;
  wire          stage3EnqWire_bits_decodeResult_maskUnit;
  wire          stage3EnqWire_bits_decodeResult_crossWrite;
  wire          stage3EnqWire_bits_decodeResult_crossRead;
  wire          stage3EnqWire_bits_decodeResult_sWrite;
  wire          stage3EnqWire_bits_decodeResult_vtype;
  wire          stage3EnqWire_bits_decodeResult_sReadVD;
  wire          stage3EnqWire_bits_decodeResult_scheduler;
  wire          stage3EnqWire_bits_decodeResult_dontNeedExecuteInLane;
  wire          stage3EnqWire_bits_decodeResult_reverse;
  wire          stage3EnqWire_bits_decodeResult_average;
  wire          stage3EnqWire_bits_decodeResult_ffo;
  wire          stage3EnqWire_bits_decodeResult_popCount;
  wire [4:0]    stage3EnqWire_bits_decodeResult_topUop;
  wire          stage3EnqWire_bits_decodeResult_specialSlot;
  wire          stage3EnqWire_bits_sSendResponse;
  wire [3:0]    stage3EnqWire_bits_mask;
  wire [31:0]   stage3EnqWire_bits_pipeData;
  wire [9:0]    stage3EnqWire_bits_groupCounter;
  wire [9:0]    readBusDequeueGroup;
  wire [1:0]    readCheckRequestVec_13_readSource;
  wire [1:0]    readCheckRequestVec_12_readSource;
  wire [1:0]    readCheckRequestVec_11_readSource;
  wire [1:0]    readCheckRequestVec_10_readSource;
  wire [1:0]    readCheckRequestVec_9_readSource;
  wire [2:0]    vrfReadRequest_0_2_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_0_2_bits_offset;
  wire [1:0]    vrfReadRequest_0_2_bits_readSource;
  wire [4:0]    vrfReadRequest_0_2_bits_vs;
  wire          vrfReadRequest_0_2_valid;
  wire [2:0]    vrfReadRequest_0_1_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_0_1_bits_offset;
  wire [1:0]    vrfReadRequest_0_1_bits_readSource;
  wire [4:0]    vrfReadRequest_0_1_bits_vs;
  wire          vrfReadRequest_0_1_valid;
  wire [2:0]    vrfReadRequest_0_0_bits_instructionIndex;
  wire [5:0]    vrfReadRequest_0_0_bits_offset;
  wire [1:0]    vrfReadRequest_0_0_bits_readSource;
  wire [4:0]    vrfReadRequest_0_0_bits_vs;
  wire          vrfReadRequest_0_0_valid;
  wire [31:0]   readBusPort_1_deq_bits_data_0;
  wire [31:0]   readBusPort_0_deq_bits_data_0;
  wire [2:0]    readBeforeMaskedWrite_bits_instructionIndex;
  wire [5:0]    readBeforeMaskedWrite_bits_offset;
  wire [4:0]    readBeforeMaskedWrite_bits_vs;
  wire          readBeforeMaskedWrite_valid;
  wire          crossLaneWriteQueue_1_almostFull;
  wire          crossLaneWriteQueue_1_almostEmpty;
  wire          crossLaneWriteQueue_0_almostFull;
  wire          crossLaneWriteQueue_0_almostEmpty;
  wire          readCheckResult_13;
  wire          readCheckResult_12;
  wire          readCheckResult_11;
  wire          readCheckResult_10;
  wire          readCheckResult_9;
  wire          readCheckResult_8;
  wire          readCheckResult_7;
  wire          readCheckResult_6;
  wire          readCheckResult_5;
  wire          readCheckResult_4;
  wire          readCheckResult_3;
  wire          readCheckResult_2;
  wire          readCheckResult_1;
  wire          readCheckResult_0;
  wire [31:0]   vrfReadResult_3_2;
  wire [31:0]   vrfReadResult_3_1;
  wire [31:0]   vrfReadResult_3_0;
  wire [31:0]   vrfReadResult_2_2;
  wire [31:0]   vrfReadResult_2_1;
  wire [31:0]   vrfReadResult_2_0;
  wire [31:0]   vrfReadResult_1_2;
  wire [31:0]   vrfReadResult_1_1;
  wire [31:0]   vrfReadResult_1_0;
  wire [31:0]   vrfReadResult_0_2;
  wire [31:0]   vrfReadResult_0_1;
  wire [31:0]   vrfReadResult_0_0;
  wire          requestVec_3_narrow;
  wire          requestVec_3_maskType;
  wire [1:0]    requestVec_3_laneIndex;
  wire [9:0]    requestVec_3_groupIndex;
  wire          requestVec_3_rem;
  wire [19:0]   requestVec_3_shifterSize;
  wire [1:0]    requestVec_3_vSew;
  wire [1:0]    requestVec_3_vxrm;
  wire          requestVec_3_saturate;
  wire          requestVec_3_average;
  wire          requestVec_3_reverse;
  wire          requestVec_3_sign;
  wire          requestVec_3_sign0;
  wire [3:0]    requestVec_3_executeMask;
  wire [3:0]    requestVec_3_mask;
  wire [3:0]    requestVec_3_opcode;
  wire [32:0]   requestVec_3_src_3;
  wire [32:0]   requestVec_3_src_2;
  wire [32:0]   requestVec_3_src_1;
  wire [32:0]   requestVec_3_src_0;
  wire          requestVec_2_narrow;
  wire          requestVec_2_maskType;
  wire [1:0]    requestVec_2_laneIndex;
  wire [9:0]    requestVec_2_groupIndex;
  wire          requestVec_2_rem;
  wire [19:0]   requestVec_2_shifterSize;
  wire [1:0]    requestVec_2_vSew;
  wire [1:0]    requestVec_2_vxrm;
  wire          requestVec_2_saturate;
  wire          requestVec_2_average;
  wire          requestVec_2_reverse;
  wire          requestVec_2_sign;
  wire          requestVec_2_sign0;
  wire [3:0]    requestVec_2_executeMask;
  wire [3:0]    requestVec_2_mask;
  wire [3:0]    requestVec_2_opcode;
  wire [32:0]   requestVec_2_src_3;
  wire [32:0]   requestVec_2_src_2;
  wire [32:0]   requestVec_2_src_1;
  wire [32:0]   requestVec_2_src_0;
  wire          requestVec_1_narrow;
  wire          requestVec_1_maskType;
  wire [1:0]    requestVec_1_laneIndex;
  wire [9:0]    requestVec_1_groupIndex;
  wire          requestVec_1_rem;
  wire [19:0]   requestVec_1_shifterSize;
  wire [1:0]    requestVec_1_vSew;
  wire [1:0]    requestVec_1_vxrm;
  wire          requestVec_1_saturate;
  wire          requestVec_1_average;
  wire          requestVec_1_reverse;
  wire          requestVec_1_sign;
  wire          requestVec_1_sign0;
  wire [3:0]    requestVec_1_executeMask;
  wire [3:0]    requestVec_1_mask;
  wire [3:0]    requestVec_1_opcode;
  wire [32:0]   requestVec_1_src_3;
  wire [32:0]   requestVec_1_src_2;
  wire [32:0]   requestVec_1_src_1;
  wire [32:0]   requestVec_1_src_0;
  wire          requestVec_0_narrow;
  wire          requestVec_0_maskType;
  wire [1:0]    requestVec_0_laneIndex;
  wire [9:0]    requestVec_0_groupIndex;
  wire [13:0]   requestVec_0_popInit;
  wire [1:0]    requestVec_0_executeIndex;
  wire          requestVec_0_rem;
  wire [19:0]   requestVec_0_shifterSize;
  wire [1:0]    requestVec_0_vSew;
  wire [1:0]    requestVec_0_vxrm;
  wire          requestVec_0_saturate;
  wire          requestVec_0_average;
  wire          requestVec_0_reverse;
  wire          requestVec_0_sign;
  wire          requestVec_0_sign0;
  wire [3:0]    requestVec_0_executeMask;
  wire [3:0]    requestVec_0_mask;
  wire [3:0]    requestVec_0_opcode;
  wire [32:0]   requestVec_0_src_3;
  wire [32:0]   requestVec_0_src_2;
  wire [32:0]   requestVec_0_src_1;
  wire [32:0]   requestVec_0_src_0;
  wire          slotShiftValid_3;
  wire          slotShiftValid_2;
  wire          slotShiftValid_1;
  wire          readBusPort_0_enq_valid_0 = readBusPort_0_enq_valid;
  wire [31:0]   readBusPort_0_enq_bits_data_0 = readBusPort_0_enq_bits_data;
  wire          readBusPort_0_deqRelease_0 = readBusPort_0_deqRelease;
  wire          readBusPort_1_enq_valid_0 = readBusPort_1_enq_valid;
  wire [31:0]   readBusPort_1_enq_bits_data_0 = readBusPort_1_enq_bits_data;
  wire          readBusPort_1_deqRelease_0 = readBusPort_1_deqRelease;
  wire          writeBusPort_0_enq_valid_0 = writeBusPort_0_enq_valid;
  wire [31:0]   writeBusPort_0_enq_bits_data_0 = writeBusPort_0_enq_bits_data;
  wire [1:0]    writeBusPort_0_enq_bits_mask_0 = writeBusPort_0_enq_bits_mask;
  wire [2:0]    writeBusPort_0_enq_bits_instructionIndex_0 = writeBusPort_0_enq_bits_instructionIndex;
  wire [9:0]    writeBusPort_0_enq_bits_counter_0 = writeBusPort_0_enq_bits_counter;
  wire          writeBusPort_0_deqRelease_0 = writeBusPort_0_deqRelease;
  wire          writeBusPort_1_enq_valid_0 = writeBusPort_1_enq_valid;
  wire [31:0]   writeBusPort_1_enq_bits_data_0 = writeBusPort_1_enq_bits_data;
  wire [1:0]    writeBusPort_1_enq_bits_mask_0 = writeBusPort_1_enq_bits_mask;
  wire [2:0]    writeBusPort_1_enq_bits_instructionIndex_0 = writeBusPort_1_enq_bits_instructionIndex;
  wire [9:0]    writeBusPort_1_enq_bits_counter_0 = writeBusPort_1_enq_bits_counter;
  wire          writeBusPort_1_deqRelease_0 = writeBusPort_1_deqRelease;
  wire          laneRequest_valid_0 = laneRequest_valid;
  wire [2:0]    laneRequest_bits_instructionIndex_0 = laneRequest_bits_instructionIndex;
  wire          laneRequest_bits_decodeResult_specialSlot_0 = laneRequest_bits_decodeResult_specialSlot;
  wire [4:0]    laneRequest_bits_decodeResult_topUop_0 = laneRequest_bits_decodeResult_topUop;
  wire          laneRequest_bits_decodeResult_popCount_0 = laneRequest_bits_decodeResult_popCount;
  wire          laneRequest_bits_decodeResult_ffo_0 = laneRequest_bits_decodeResult_ffo;
  wire          laneRequest_bits_decodeResult_average_0 = laneRequest_bits_decodeResult_average;
  wire          laneRequest_bits_decodeResult_reverse_0 = laneRequest_bits_decodeResult_reverse;
  wire          laneRequest_bits_decodeResult_dontNeedExecuteInLane_0 = laneRequest_bits_decodeResult_dontNeedExecuteInLane;
  wire          laneRequest_bits_decodeResult_scheduler_0 = laneRequest_bits_decodeResult_scheduler;
  wire          laneRequest_bits_decodeResult_sReadVD_0 = laneRequest_bits_decodeResult_sReadVD;
  wire          laneRequest_bits_decodeResult_vtype_0 = laneRequest_bits_decodeResult_vtype;
  wire          laneRequest_bits_decodeResult_sWrite_0 = laneRequest_bits_decodeResult_sWrite;
  wire          laneRequest_bits_decodeResult_crossRead_0 = laneRequest_bits_decodeResult_crossRead;
  wire          laneRequest_bits_decodeResult_crossWrite_0 = laneRequest_bits_decodeResult_crossWrite;
  wire          laneRequest_bits_decodeResult_maskUnit_0 = laneRequest_bits_decodeResult_maskUnit;
  wire          laneRequest_bits_decodeResult_special_0 = laneRequest_bits_decodeResult_special;
  wire          laneRequest_bits_decodeResult_saturate_0 = laneRequest_bits_decodeResult_saturate;
  wire          laneRequest_bits_decodeResult_vwmacc_0 = laneRequest_bits_decodeResult_vwmacc;
  wire          laneRequest_bits_decodeResult_readOnly_0 = laneRequest_bits_decodeResult_readOnly;
  wire          laneRequest_bits_decodeResult_maskSource_0 = laneRequest_bits_decodeResult_maskSource;
  wire          laneRequest_bits_decodeResult_maskDestination_0 = laneRequest_bits_decodeResult_maskDestination;
  wire          laneRequest_bits_decodeResult_maskLogic_0 = laneRequest_bits_decodeResult_maskLogic;
  wire [3:0]    laneRequest_bits_decodeResult_uop_0 = laneRequest_bits_decodeResult_uop;
  wire          laneRequest_bits_decodeResult_iota_0 = laneRequest_bits_decodeResult_iota;
  wire          laneRequest_bits_decodeResult_mv_0 = laneRequest_bits_decodeResult_mv;
  wire          laneRequest_bits_decodeResult_extend_0 = laneRequest_bits_decodeResult_extend;
  wire          laneRequest_bits_decodeResult_unOrderWrite_0 = laneRequest_bits_decodeResult_unOrderWrite;
  wire          laneRequest_bits_decodeResult_compress_0 = laneRequest_bits_decodeResult_compress;
  wire          laneRequest_bits_decodeResult_gather16_0 = laneRequest_bits_decodeResult_gather16;
  wire          laneRequest_bits_decodeResult_gather_0 = laneRequest_bits_decodeResult_gather;
  wire          laneRequest_bits_decodeResult_slid_0 = laneRequest_bits_decodeResult_slid;
  wire          laneRequest_bits_decodeResult_targetRd_0 = laneRequest_bits_decodeResult_targetRd;
  wire          laneRequest_bits_decodeResult_widenReduce_0 = laneRequest_bits_decodeResult_widenReduce;
  wire          laneRequest_bits_decodeResult_red_0 = laneRequest_bits_decodeResult_red;
  wire          laneRequest_bits_decodeResult_nr_0 = laneRequest_bits_decodeResult_nr;
  wire          laneRequest_bits_decodeResult_itype_0 = laneRequest_bits_decodeResult_itype;
  wire          laneRequest_bits_decodeResult_unsigned1_0 = laneRequest_bits_decodeResult_unsigned1;
  wire          laneRequest_bits_decodeResult_unsigned0_0 = laneRequest_bits_decodeResult_unsigned0;
  wire          laneRequest_bits_decodeResult_other_0 = laneRequest_bits_decodeResult_other;
  wire          laneRequest_bits_decodeResult_multiCycle_0 = laneRequest_bits_decodeResult_multiCycle;
  wire          laneRequest_bits_decodeResult_divider_0 = laneRequest_bits_decodeResult_divider;
  wire          laneRequest_bits_decodeResult_multiplier_0 = laneRequest_bits_decodeResult_multiplier;
  wire          laneRequest_bits_decodeResult_shift_0 = laneRequest_bits_decodeResult_shift;
  wire          laneRequest_bits_decodeResult_adder_0 = laneRequest_bits_decodeResult_adder;
  wire          laneRequest_bits_decodeResult_logic_0 = laneRequest_bits_decodeResult_logic;
  wire          laneRequest_bits_loadStore_0 = laneRequest_bits_loadStore;
  wire          laneRequest_bits_issueInst_0 = laneRequest_bits_issueInst;
  wire          laneRequest_bits_store_0 = laneRequest_bits_store;
  wire          laneRequest_bits_special_0 = laneRequest_bits_special;
  wire          laneRequest_bits_lsWholeReg_0 = laneRequest_bits_lsWholeReg;
  wire [4:0]    laneRequest_bits_vs1_0 = laneRequest_bits_vs1;
  wire [4:0]    laneRequest_bits_vs2_0 = laneRequest_bits_vs2;
  wire [4:0]    laneRequest_bits_vd_0 = laneRequest_bits_vd;
  wire [1:0]    laneRequest_bits_loadStoreEEW_0 = laneRequest_bits_loadStoreEEW;
  wire          laneRequest_bits_mask_0 = laneRequest_bits_mask;
  wire [2:0]    laneRequest_bits_segment_0 = laneRequest_bits_segment;
  wire [31:0]   laneRequest_bits_readFromScalar_0 = laneRequest_bits_readFromScalar;
  wire [13:0]   laneRequest_bits_csrInterface_vl_0 = laneRequest_bits_csrInterface_vl;
  wire [13:0]   laneRequest_bits_csrInterface_vStart_0 = laneRequest_bits_csrInterface_vStart;
  wire [2:0]    laneRequest_bits_csrInterface_vlmul_0 = laneRequest_bits_csrInterface_vlmul;
  wire [1:0]    laneRequest_bits_csrInterface_vSew_0 = laneRequest_bits_csrInterface_vSew;
  wire [1:0]    laneRequest_bits_csrInterface_vxrm_0 = laneRequest_bits_csrInterface_vxrm;
  wire          laneRequest_bits_csrInterface_vta_0 = laneRequest_bits_csrInterface_vta;
  wire          laneRequest_bits_csrInterface_vma_0 = laneRequest_bits_csrInterface_vma;
  wire          tokenIO_maskRequestRelease_0 = tokenIO_maskRequestRelease;
  wire          vrfReadAddressChannel_valid_0 = vrfReadAddressChannel_valid;
  wire [4:0]    vrfReadAddressChannel_bits_vs_0 = vrfReadAddressChannel_bits_vs;
  wire [1:0]    vrfReadAddressChannel_bits_readSource_0 = vrfReadAddressChannel_bits_readSource;
  wire [5:0]    vrfReadAddressChannel_bits_offset_0 = vrfReadAddressChannel_bits_offset;
  wire [2:0]    vrfReadAddressChannel_bits_instructionIndex_0 = vrfReadAddressChannel_bits_instructionIndex;
  wire          vrfWriteChannel_valid_0 = vrfWriteChannel_valid;
  wire [4:0]    vrfWriteChannel_bits_vd_0 = vrfWriteChannel_bits_vd;
  wire [5:0]    vrfWriteChannel_bits_offset_0 = vrfWriteChannel_bits_offset;
  wire [3:0]    vrfWriteChannel_bits_mask_0 = vrfWriteChannel_bits_mask;
  wire [31:0]   vrfWriteChannel_bits_data_0 = vrfWriteChannel_bits_data;
  wire          vrfWriteChannel_bits_last_0 = vrfWriteChannel_bits_last;
  wire [2:0]    vrfWriteChannel_bits_instructionIndex_0 = vrfWriteChannel_bits_instructionIndex;
  wire [1:0]    laneState_laneIndex = laneIndex;
  wire [1:0]    laneState_1_laneIndex = laneIndex;
  wire [1:0]    laneState_2_laneIndex = laneIndex;
  wire [1:0]    laneState_3_laneIndex = laneIndex;
  wire [1:0]    requestVec_1_tag = 2'h1;
  wire [1:0]    requestVecFromSlot_1_other_bits_tag = 2'h1;
  wire [1:0]    requestVecFromSlot_1_divider_bits_tag = 2'h1;
  wire [1:0]    requestVecFromSlot_1_multiplier_bits_tag = 2'h1;
  wire [1:0]    requestVecFromSlot_1_shift_bits_tag = 2'h1;
  wire [1:0]    requestVecFromSlot_1_adder_bits_tag = 2'h1;
  wire [1:0]    requestVecFromSlot_1_logic_bits_tag = 2'h1;
  wire [13:0]   requestVec_1_popInit = 14'h0;
  wire [13:0]   requestVec_2_popInit = 14'h0;
  wire [13:0]   requestVec_3_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_1_other_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_1_divider_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_1_multiplier_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_1_shift_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_1_adder_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_1_logic_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_2_other_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_2_divider_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_2_multiplier_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_2_shift_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_2_adder_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_2_logic_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_3_other_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_3_divider_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_3_multiplier_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_3_shift_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_3_adder_bits_popInit = 14'h0;
  wire [13:0]   requestVecFromSlot_3_logic_bits_popInit = 14'h0;
  wire [1:0]    requestVec_3_tag = 2'h3;
  wire [1:0]    requestVecFromSlot_3_other_bits_tag = 2'h3;
  wire [1:0]    requestVecFromSlot_3_divider_bits_tag = 2'h3;
  wire [1:0]    requestVecFromSlot_3_multiplier_bits_tag = 2'h3;
  wire [1:0]    requestVecFromSlot_3_shift_bits_tag = 2'h3;
  wire [1:0]    requestVecFromSlot_3_adder_bits_tag = 2'h3;
  wire [1:0]    requestVecFromSlot_3_logic_bits_tag = 2'h3;
  wire [2:0]    vfuResponse_VFUNotClear_lo = 3'h0;
  wire [2:0]    vfuResponse_VFUNotClear_lo_1 = 3'h0;
  wire [2:0]    vfuResponse_VFUNotClear_lo_2 = 3'h0;
  wire [2:0]    vfuResponse_VFUNotClear_lo_3 = 3'h0;
  wire [2:0]    vfuResponse_VFUNotClear_lo_4 = 3'h0;
  wire [2:0]    vfuResponse_VFUNotClear_lo_5 = 3'h0;
  wire [1:0]    requestVec_2_tag = 2'h2;
  wire [1:0]    requestVecFromSlot_2_other_bits_tag = 2'h2;
  wire [1:0]    requestVecFromSlot_2_divider_bits_tag = 2'h2;
  wire [1:0]    requestVecFromSlot_2_multiplier_bits_tag = 2'h2;
  wire [1:0]    requestVecFromSlot_2_shift_bits_tag = 2'h2;
  wire [1:0]    requestVecFromSlot_2_adder_bits_tag = 2'h2;
  wire [1:0]    requestVecFromSlot_2_logic_bits_tag = 2'h2;
  wire [1:0]    readBeforeMaskedWrite_bits_readSource = 2'h2;
  wire [31:0]   stage3EnqWire_1_bits_pipeData = 32'h0;
  wire [31:0]   stage3EnqWire_1_bits_crossWriteData_0 = 32'h0;
  wire [31:0]   stage3EnqWire_1_bits_crossWriteData_1 = 32'h0;
  wire [31:0]   stage3EnqWire_2_bits_pipeData = 32'h0;
  wire [31:0]   stage3EnqWire_2_bits_crossWriteData_0 = 32'h0;
  wire [31:0]   stage3EnqWire_2_bits_crossWriteData_1 = 32'h0;
  wire [31:0]   stage3EnqWire_3_bits_pipeData = 32'h0;
  wire [31:0]   stage3EnqWire_3_bits_crossWriteData_0 = 32'h0;
  wire [31:0]   stage3EnqWire_3_bits_crossWriteData_1 = 32'h0;
  wire [31:0]   entranceControl_mask_bits = 32'h0;
  wire [63:0]   segmentMask_notAccessForRegister = 64'hFFFFFFFFFFFFFFFF;
  wire          slotCanShift_1 = 1'h1;
  wire          slotCanShift_2 = 1'h1;
  wire          slotCanShift_3 = 1'h1;
  wire [4:0]    responseVec_0_bits_exceptionFlags = 5'h0;
  wire [4:0]    responseVec_1_bits_exceptionFlags = 5'h0;
  wire [4:0]    responseVec_2_bits_exceptionFlags = 5'h0;
  wire [4:0]    responseVec_3_bits_exceptionFlags = 5'h0;
  wire [4:0]    vfuResponse_0_bits_exceptionFlags = 5'h0;
  wire [4:0]    vfuResponse_1_bits_exceptionFlags = 5'h0;
  wire [4:0]    vfuResponse_responseBundle_bits_exceptionFlags = 5'h0;
  wire [4:0]    vfuResponse_3_bits_exceptionFlags = 5'h0;
  wire [4:0]    vfuResponse_responseBundle_1_bits_exceptionFlags = 5'h0;
  wire [4:0]    vfuResponse_responseBundle_2_bits_exceptionFlags = 5'h0;
  wire [4:0]    selectResponse_bits_exceptionFlags = 5'h0;
  wire [4:0]    selectResponse_1_bits_exceptionFlags = 5'h0;
  wire [4:0]    selectResponse_2_bits_exceptionFlags = 5'h0;
  wire [4:0]    selectResponse_3_bits_exceptionFlags = 5'h0;
  wire [1:0]    requestVec_0_tag = 2'h0;
  wire [1:0]    requestVec_1_executeIndex = 2'h0;
  wire [1:0]    requestVec_2_executeIndex = 2'h0;
  wire [1:0]    requestVec_3_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_0_other_bits_tag = 2'h0;
  wire [1:0]    requestVecFromSlot_0_divider_bits_tag = 2'h0;
  wire [1:0]    requestVecFromSlot_0_multiplier_bits_tag = 2'h0;
  wire [1:0]    requestVecFromSlot_0_shift_bits_tag = 2'h0;
  wire [1:0]    requestVecFromSlot_0_adder_bits_tag = 2'h0;
  wire [1:0]    requestVecFromSlot_0_logic_bits_tag = 2'h0;
  wire [1:0]    requestVecFromSlot_1_other_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_1_divider_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_1_multiplier_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_1_shift_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_1_adder_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_1_logic_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_2_other_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_2_divider_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_2_multiplier_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_2_shift_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_2_adder_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_2_logic_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_3_other_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_3_divider_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_3_multiplier_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_3_shift_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_3_adder_bits_executeIndex = 2'h0;
  wire [1:0]    requestVecFromSlot_3_logic_bits_executeIndex = 2'h0;
  wire [1:0]    vfuResponse_0_bits_executeIndex = 2'h0;
  wire [1:0]    vfuResponse_VFUNotClear_lo_hi = 2'h0;
  wire [1:0]    vfuResponse_VFUNotClear_lo_hi_1 = 2'h0;
  wire [1:0]    vfuResponse_responseBundle_bits_executeIndex = 2'h0;
  wire [1:0]    vfuResponse_VFUNotClear_lo_hi_2 = 2'h0;
  wire [1:0]    vfuResponse_3_bits_executeIndex = 2'h0;
  wire [1:0]    vfuResponse_VFUNotClear_lo_hi_3 = 2'h0;
  wire [1:0]    vfuResponse_VFUNotClear_lo_hi_4 = 2'h0;
  wire [1:0]    vfuResponse_responseBundle_2_bits_executeIndex = 2'h0;
  wire [1:0]    vfuResponse_VFUNotClear_lo_hi_5 = 2'h0;
  wire [1:0]    entranceControl_executeIndex = 2'h0;
  wire          requestVec_0_complete = 1'h0;
  wire          requestVec_1_complete = 1'h0;
  wire          requestVec_2_complete = 1'h0;
  wire          requestVec_3_complete = 1'h0;
  wire          responseVec_0_bits_clipFail = 1'h0;
  wire          responseVec_0_bits_divBusy = 1'h0;
  wire          responseVec_1_bits_clipFail = 1'h0;
  wire          responseVec_1_bits_divBusy = 1'h0;
  wire          responseVec_2_bits_clipFail = 1'h0;
  wire          responseVec_2_bits_divBusy = 1'h0;
  wire          responseVec_3_bits_clipFail = 1'h0;
  wire          responseVec_3_bits_divBusy = 1'h0;
  wire          crossLaneWriteQueue_0_enq_bits_last = 1'h0;
  wire          crossLaneWriteQueue_1_enq_bits_last = 1'h0;
  wire          stage3EnqWire_bits_ffoByOtherLanes = 1'h0;
  wire          stage3EnqWire_1_bits_sSendResponse = 1'h0;
  wire          stage3EnqWire_1_bits_ffoSuccess = 1'h0;
  wire          stage3EnqWire_1_bits_ffoByOtherLanes = 1'h0;
  wire          stage3EnqWire_2_bits_sSendResponse = 1'h0;
  wire          stage3EnqWire_2_bits_ffoSuccess = 1'h0;
  wire          stage3EnqWire_2_bits_ffoByOtherLanes = 1'h0;
  wire          stage3EnqWire_3_bits_sSendResponse = 1'h0;
  wire          stage3EnqWire_3_bits_ffoSuccess = 1'h0;
  wire          stage3EnqWire_3_bits_ffoByOtherLanes = 1'h0;
  wire          requestVecFromSlot_0_other_bits_complete = 1'h0;
  wire          requestVecFromSlot_0_divider_bits_complete = 1'h0;
  wire          requestVecFromSlot_0_multiplier_bits_complete = 1'h0;
  wire          requestVecFromSlot_0_shift_bits_complete = 1'h0;
  wire          requestVecFromSlot_0_adder_bits_complete = 1'h0;
  wire          requestVecFromSlot_0_logic_bits_complete = 1'h0;
  wire          requestVecFromSlot_1_other_bits_complete = 1'h0;
  wire          requestVecFromSlot_1_divider_bits_complete = 1'h0;
  wire          requestVecFromSlot_1_multiplier_bits_complete = 1'h0;
  wire          requestVecFromSlot_1_shift_bits_complete = 1'h0;
  wire          requestVecFromSlot_1_adder_bits_complete = 1'h0;
  wire          requestVecFromSlot_1_logic_bits_complete = 1'h0;
  wire          requestVecFromSlot_2_other_bits_complete = 1'h0;
  wire          requestVecFromSlot_2_divider_bits_complete = 1'h0;
  wire          requestVecFromSlot_2_multiplier_bits_complete = 1'h0;
  wire          requestVecFromSlot_2_shift_bits_complete = 1'h0;
  wire          requestVecFromSlot_2_adder_bits_complete = 1'h0;
  wire          requestVecFromSlot_2_logic_bits_complete = 1'h0;
  wire          requestVecFromSlot_3_other_bits_complete = 1'h0;
  wire          requestVecFromSlot_3_divider_bits_complete = 1'h0;
  wire          requestVecFromSlot_3_multiplier_bits_complete = 1'h0;
  wire          requestVecFromSlot_3_shift_bits_complete = 1'h0;
  wire          requestVecFromSlot_3_adder_bits_complete = 1'h0;
  wire          requestVecFromSlot_3_logic_bits_complete = 1'h0;
  wire          vrfIsBusy_0 = 1'h0;
  wire          vrfIsBusy_1 = 1'h0;
  wire          vrfIsBusy_2 = 1'h0;
  wire          vrfIsBusy_3 = 1'h0;
  wire          vrfIsBusy_5 = 1'h0;
  wire          vfuResponse_0_bits_clipFail = 1'h0;
  wire          vfuResponse_0_bits_ffoSuccess = 1'h0;
  wire          vfuResponse_0_bits_divBusy = 1'h0;
  wire          vfuResponse_1_bits_clipFail = 1'h0;
  wire          vfuResponse_1_bits_ffoSuccess = 1'h0;
  wire          vfuResponse_1_bits_divBusy = 1'h0;
  wire          vfuResponse_responseBundle_bits_clipFail = 1'h0;
  wire          vfuResponse_responseBundle_bits_ffoSuccess = 1'h0;
  wire          vfuResponse_responseBundle_bits_divBusy = 1'h0;
  wire          vfuResponse_3_bits_clipFail = 1'h0;
  wire          vfuResponse_3_bits_ffoSuccess = 1'h0;
  wire          vfuResponse_3_bits_divBusy = 1'h0;
  wire          vfuResponse_responseBundle_1_bits_clipFail = 1'h0;
  wire          vfuResponse_responseBundle_1_bits_ffoSuccess = 1'h0;
  wire          vfuResponse_responseBundle_1_bits_divBusy = 1'h0;
  wire          vfuResponse_responseBundle_2_bits_divBusy = 1'h0;
  wire          selectResponse_bits_clipFail = 1'h0;
  wire          selectResponse_bits_divBusy = 1'h0;
  wire          selectResponse_1_bits_clipFail = 1'h0;
  wire          selectResponse_1_bits_divBusy = 1'h0;
  wire          selectResponse_2_bits_clipFail = 1'h0;
  wire          selectResponse_2_bits_divBusy = 1'h0;
  wire          selectResponse_3_bits_clipFail = 1'h0;
  wire          selectResponse_3_bits_divBusy = 1'h0;
  wire          entranceControl_mask_valid = 1'h0;
  wire [3:0]    vfuResponse_0_bits_adderMaskResp = 4'h0;
  wire [3:0]    vfuResponse_0_bits_vxsat = 4'h0;
  wire [3:0]    vfuResponse_responseBundle_bits_adderMaskResp = 4'h0;
  wire [3:0]    vfuResponse_responseBundle_bits_vxsat = 4'h0;
  wire [3:0]    vfuResponse_3_bits_adderMaskResp = 4'h0;
  wire [3:0]    vfuResponse_responseBundle_1_bits_adderMaskResp = 4'h0;
  wire [3:0]    vfuResponse_responseBundle_1_bits_vxsat = 4'h0;
  wire [3:0]    vfuResponse_responseBundle_2_bits_adderMaskResp = 4'h0;
  wire [3:0]    vfuResponse_responseBundle_2_bits_vxsat = 4'h0;
  wire [3:0]    entranceControl_vrfWriteMask = 4'h0;
  wire          queue_enq_valid = readBusPort_0_enq_valid_0;
  wire [31:0]   queue_enq_bits_data = readBusPort_0_enq_bits_data_0;
  wire          queue_1_enq_valid = readBusPort_1_enq_valid_0;
  wire [31:0]   queue_1_enq_bits_data = readBusPort_1_enq_bits_data_0;
  wire          crossLaneWriteQueue_0_enq_valid = writeBusPort_0_enq_valid_0;
  wire [31:0]   crossLaneWriteQueue_0_enq_bits_data = writeBusPort_0_enq_bits_data_0;
  wire [2:0]    crossLaneWriteQueue_0_enq_bits_instructionIndex = writeBusPort_0_enq_bits_instructionIndex_0;
  wire          crossLaneWriteQueue_1_enq_valid = writeBusPort_1_enq_valid_0;
  wire [31:0]   crossLaneWriteQueue_1_enq_bits_data = writeBusPort_1_enq_bits_data_0;
  wire [2:0]    crossLaneWriteQueue_1_enq_bits_instructionIndex = writeBusPort_1_enq_bits_instructionIndex_0;
  wire          slotFree;
  wire          enqueueValid_3 = laneRequest_valid_0;
  wire [2:0]    entranceControl_laneRequest_instructionIndex = laneRequest_bits_instructionIndex_0;
  wire          entranceControl_laneRequest_decodeResult_specialSlot = laneRequest_bits_decodeResult_specialSlot_0;
  wire [4:0]    entranceControl_laneRequest_decodeResult_topUop = laneRequest_bits_decodeResult_topUop_0;
  wire          entranceControl_laneRequest_decodeResult_popCount = laneRequest_bits_decodeResult_popCount_0;
  wire          entranceControl_laneRequest_decodeResult_ffo = laneRequest_bits_decodeResult_ffo_0;
  wire          entranceControl_laneRequest_decodeResult_average = laneRequest_bits_decodeResult_average_0;
  wire          entranceControl_laneRequest_decodeResult_reverse = laneRequest_bits_decodeResult_reverse_0;
  wire          entranceControl_laneRequest_decodeResult_dontNeedExecuteInLane = laneRequest_bits_decodeResult_dontNeedExecuteInLane_0;
  wire          entranceControl_laneRequest_decodeResult_scheduler = laneRequest_bits_decodeResult_scheduler_0;
  wire          entranceControl_laneRequest_decodeResult_sReadVD = laneRequest_bits_decodeResult_sReadVD_0;
  wire          entranceControl_laneRequest_decodeResult_vtype = laneRequest_bits_decodeResult_vtype_0;
  wire          entranceControl_laneRequest_decodeResult_sWrite = laneRequest_bits_decodeResult_sWrite_0;
  wire          entranceControl_laneRequest_decodeResult_crossRead = laneRequest_bits_decodeResult_crossRead_0;
  wire          entranceControl_laneRequest_decodeResult_crossWrite = laneRequest_bits_decodeResult_crossWrite_0;
  wire          entranceControl_laneRequest_decodeResult_maskUnit = laneRequest_bits_decodeResult_maskUnit_0;
  wire          entranceControl_laneRequest_decodeResult_special = laneRequest_bits_decodeResult_special_0;
  wire          entranceControl_laneRequest_decodeResult_saturate = laneRequest_bits_decodeResult_saturate_0;
  wire          entranceControl_laneRequest_decodeResult_vwmacc = laneRequest_bits_decodeResult_vwmacc_0;
  wire          entranceControl_laneRequest_decodeResult_readOnly = laneRequest_bits_decodeResult_readOnly_0;
  wire          entranceControl_laneRequest_decodeResult_maskSource = laneRequest_bits_decodeResult_maskSource_0;
  wire          entranceControl_laneRequest_decodeResult_maskDestination = laneRequest_bits_decodeResult_maskDestination_0;
  wire          entranceControl_laneRequest_decodeResult_maskLogic = laneRequest_bits_decodeResult_maskLogic_0;
  wire [3:0]    entranceControl_laneRequest_decodeResult_uop = laneRequest_bits_decodeResult_uop_0;
  wire          entranceControl_laneRequest_decodeResult_iota = laneRequest_bits_decodeResult_iota_0;
  wire          entranceControl_laneRequest_decodeResult_mv = laneRequest_bits_decodeResult_mv_0;
  wire          entranceControl_laneRequest_decodeResult_extend = laneRequest_bits_decodeResult_extend_0;
  wire          entranceControl_laneRequest_decodeResult_unOrderWrite = laneRequest_bits_decodeResult_unOrderWrite_0;
  wire          entranceControl_laneRequest_decodeResult_compress = laneRequest_bits_decodeResult_compress_0;
  wire          entranceControl_laneRequest_decodeResult_gather16 = laneRequest_bits_decodeResult_gather16_0;
  wire          entranceControl_laneRequest_decodeResult_gather = laneRequest_bits_decodeResult_gather_0;
  wire          entranceControl_laneRequest_decodeResult_slid = laneRequest_bits_decodeResult_slid_0;
  wire          entranceControl_laneRequest_decodeResult_targetRd = laneRequest_bits_decodeResult_targetRd_0;
  wire          entranceControl_laneRequest_decodeResult_widenReduce = laneRequest_bits_decodeResult_widenReduce_0;
  wire          entranceControl_laneRequest_decodeResult_red = laneRequest_bits_decodeResult_red_0;
  wire          entranceControl_laneRequest_decodeResult_nr = laneRequest_bits_decodeResult_nr_0;
  wire          entranceControl_laneRequest_decodeResult_itype = laneRequest_bits_decodeResult_itype_0;
  wire          entranceControl_laneRequest_decodeResult_unsigned1 = laneRequest_bits_decodeResult_unsigned1_0;
  wire          entranceControl_laneRequest_decodeResult_unsigned0 = laneRequest_bits_decodeResult_unsigned0_0;
  wire          entranceControl_laneRequest_decodeResult_other = laneRequest_bits_decodeResult_other_0;
  wire          entranceControl_laneRequest_decodeResult_multiCycle = laneRequest_bits_decodeResult_multiCycle_0;
  wire          entranceControl_laneRequest_decodeResult_divider = laneRequest_bits_decodeResult_divider_0;
  wire          entranceControl_laneRequest_decodeResult_multiplier = laneRequest_bits_decodeResult_multiplier_0;
  wire          entranceControl_laneRequest_decodeResult_shift = laneRequest_bits_decodeResult_shift_0;
  wire          entranceControl_laneRequest_decodeResult_adder = laneRequest_bits_decodeResult_adder_0;
  wire          entranceControl_laneRequest_decodeResult_logic = laneRequest_bits_decodeResult_logic_0;
  wire          entranceControl_laneRequest_loadStore = laneRequest_bits_loadStore_0;
  wire          entranceControl_laneRequest_issueInst = laneRequest_bits_issueInst_0;
  wire          entranceControl_laneRequest_store = laneRequest_bits_store_0;
  wire          entranceControl_laneRequest_special = laneRequest_bits_special_0;
  wire          entranceControl_laneRequest_lsWholeReg = laneRequest_bits_lsWholeReg_0;
  wire [4:0]    entranceControl_laneRequest_vs1 = laneRequest_bits_vs1_0;
  wire [4:0]    entranceControl_laneRequest_vs2 = laneRequest_bits_vs2_0;
  wire [4:0]    entranceControl_laneRequest_vd = laneRequest_bits_vd_0;
  wire [1:0]    entranceControl_laneRequest_loadStoreEEW = laneRequest_bits_loadStoreEEW_0;
  wire          entranceControl_laneRequest_mask = laneRequest_bits_mask_0;
  wire [2:0]    entranceControl_laneRequest_segment = laneRequest_bits_segment_0;
  wire [31:0]   entranceControl_laneRequest_readFromScalar = laneRequest_bits_readFromScalar_0;
  wire [13:0]   entranceControl_laneRequest_csrInterface_vl = laneRequest_bits_csrInterface_vl_0;
  wire [13:0]   entranceControl_laneRequest_csrInterface_vStart = laneRequest_bits_csrInterface_vStart_0;
  wire [2:0]    entranceControl_laneRequest_csrInterface_vlmul = laneRequest_bits_csrInterface_vlmul_0;
  wire [1:0]    entranceControl_laneRequest_csrInterface_vSew = laneRequest_bits_csrInterface_vSew_0;
  wire [1:0]    entranceControl_laneRequest_csrInterface_vxrm = laneRequest_bits_csrInterface_vxrm_0;
  wire          entranceControl_laneRequest_csrInterface_vta = laneRequest_bits_csrInterface_vta_0;
  wire          entranceControl_laneRequest_csrInterface_vma = laneRequest_bits_csrInterface_vma_0;
  wire          vrfWriteArbiter_4_ready;
  wire          vrfWriteArbiter_4_valid = vrfWriteChannel_valid_0;
  wire [4:0]    vrfWriteArbiter_4_bits_vd = vrfWriteChannel_bits_vd_0;
  wire [5:0]    vrfWriteArbiter_4_bits_offset = vrfWriteChannel_bits_offset_0;
  wire [3:0]    vrfWriteArbiter_4_bits_mask = vrfWriteChannel_bits_mask_0;
  wire [31:0]   vrfWriteArbiter_4_bits_data = vrfWriteChannel_bits_data_0;
  wire          vrfWriteArbiter_4_bits_last = vrfWriteChannel_bits_last_0;
  wire [2:0]    vrfWriteArbiter_4_bits_instructionIndex = vrfWriteChannel_bits_instructionIndex_0;
  reg           slotOccupied_0;
  wire          slotActive_0 = slotOccupied_0;
  reg           slotOccupied_1;
  wire          enqueueValid = slotOccupied_1;
  reg           slotOccupied_2;
  wire          enqueueValid_1 = slotOccupied_2;
  reg           slotOccupied_3;
  wire          enqueueValid_2 = slotOccupied_3;
  reg  [7:0]    maskGroupCountVec_0;
  reg  [7:0]    maskGroupCountVec_1;
  reg  [7:0]    maskGroupCountVec_2;
  reg  [7:0]    maskGroupCountVec_3;
  reg  [4:0]    maskIndexVec_0;
  reg  [4:0]    maskIndexVec_1;
  reg  [4:0]    maskIndexVec_2;
  reg  [4:0]    maskIndexVec_3;
  wire          enqReady;
  wire          enqReady_1;
  wire          enqReady_2;
  wire          enqReady_3;
  wire          enqReady_4;
  wire          vrfWriteChannel_ready_0 = vrfWriteArbiter_4_ready;
  reg  [4:0]    allVrfWriteAfterCheck_0_vd;
  reg  [5:0]    allVrfWriteAfterCheck_0_offset;
  reg  [3:0]    allVrfWriteAfterCheck_0_mask;
  reg  [31:0]   allVrfWriteAfterCheck_0_data;
  reg           allVrfWriteAfterCheck_0_last;
  reg  [2:0]    allVrfWriteAfterCheck_0_instructionIndex;
  reg  [4:0]    allVrfWriteAfterCheck_1_vd;
  reg  [5:0]    allVrfWriteAfterCheck_1_offset;
  reg  [3:0]    allVrfWriteAfterCheck_1_mask;
  reg  [31:0]   allVrfWriteAfterCheck_1_data;
  reg           allVrfWriteAfterCheck_1_last;
  reg  [2:0]    allVrfWriteAfterCheck_1_instructionIndex;
  reg  [4:0]    allVrfWriteAfterCheck_2_vd;
  reg  [5:0]    allVrfWriteAfterCheck_2_offset;
  reg  [3:0]    allVrfWriteAfterCheck_2_mask;
  reg  [31:0]   allVrfWriteAfterCheck_2_data;
  reg           allVrfWriteAfterCheck_2_last;
  reg  [2:0]    allVrfWriteAfterCheck_2_instructionIndex;
  reg  [4:0]    allVrfWriteAfterCheck_3_vd;
  reg  [5:0]    allVrfWriteAfterCheck_3_offset;
  reg  [3:0]    allVrfWriteAfterCheck_3_mask;
  reg  [31:0]   allVrfWriteAfterCheck_3_data;
  reg           allVrfWriteAfterCheck_3_last;
  reg  [2:0]    allVrfWriteAfterCheck_3_instructionIndex;
  reg  [4:0]    allVrfWriteAfterCheck_4_vd;
  reg  [5:0]    allVrfWriteAfterCheck_4_offset;
  reg  [3:0]    allVrfWriteAfterCheck_4_mask;
  reg  [31:0]   allVrfWriteAfterCheck_4_data;
  reg           allVrfWriteAfterCheck_4_last;
  reg  [2:0]    allVrfWriteAfterCheck_4_instructionIndex;
  reg  [4:0]    allVrfWriteAfterCheck_5_vd;
  reg  [5:0]    allVrfWriteAfterCheck_5_offset;
  reg  [3:0]    allVrfWriteAfterCheck_5_mask;
  reg  [31:0]   allVrfWriteAfterCheck_5_data;
  reg           allVrfWriteAfterCheck_5_last;
  reg  [2:0]    allVrfWriteAfterCheck_5_instructionIndex;
  reg  [4:0]    allVrfWriteAfterCheck_6_vd;
  reg  [5:0]    allVrfWriteAfterCheck_6_offset;
  reg  [3:0]    allVrfWriteAfterCheck_6_mask;
  reg  [31:0]   allVrfWriteAfterCheck_6_data;
  reg           allVrfWriteAfterCheck_6_last;
  reg  [2:0]    allVrfWriteAfterCheck_6_instructionIndex;
  reg           afterCheckValid_0;
  reg           afterCheckValid_1;
  reg           afterCheckValid_2;
  reg           afterCheckValid_3;
  reg           afterCheckValid_4;
  reg           afterCheckValid_5;
  reg           afterCheckValid_6;
  wire          afterCheckDequeueReady_0;
  wire          afterCheckDequeueFire_0 = afterCheckValid_0 & afterCheckDequeueReady_0;
  wire          afterCheckDequeueReady_1;
  wire          afterCheckDequeueFire_1 = afterCheckValid_1 & afterCheckDequeueReady_1;
  wire          afterCheckDequeueReady_2;
  wire          afterCheckDequeueFire_2 = afterCheckValid_2 & afterCheckDequeueReady_2;
  wire          afterCheckDequeueReady_3;
  wire          afterCheckDequeueFire_3 = afterCheckValid_3 & afterCheckDequeueReady_3;
  wire          afterCheckDequeueReady_4;
  wire          afterCheckDequeueFire_4 = afterCheckValid_4 & afterCheckDequeueReady_4;
  wire          afterCheckDequeueReady_5;
  wire          afterCheckDequeueFire_5 = afterCheckValid_5 & afterCheckDequeueReady_5;
  wire          afterCheckDequeueReady_6;
  wire          afterCheckDequeueFire_6 = afterCheckValid_6 & afterCheckDequeueReady_6;
  wire          maskControlReq_0;
  wire          maskControlReq_1;
  wire [1:0]    maskControlReqSelect_lo = {maskControlReq_1, maskControlReq_0};
  wire          maskControlReq_2;
  wire          maskControlReq_3;
  wire [1:0]    maskControlReqSelect_hi = {maskControlReq_3, maskControlReq_2};
  wire [2:0]    _maskControlReqSelect_T_3 = {maskControlReqSelect_hi[0], maskControlReqSelect_lo} | {maskControlReqSelect_lo, 1'h0};
  wire [3:0]    maskControlReqSelect = {~(_maskControlReqSelect_T_3 | {_maskControlReqSelect_T_3[0], 2'h0}), 1'h1} & {maskControlReqSelect_hi, maskControlReqSelect_lo};
  reg  [2:0]    maskControlVec_0_index;
  reg  [1:0]    maskControlVec_0_sew;
  reg  [31:0]   maskControlVec_0_maskData;
  reg  [7:0]    maskControlVec_0_group;
  reg           maskControlVec_0_dataValid;
  reg           maskControlVec_0_waiteResponse;
  reg           maskControlVec_0_controlValid;
  wire [2:0]    maskControlRelease_0_bits;
  wire          maskControlRelease_0_valid;
  wire [2:0]    maskControlRelease_1_bits;
  wire          maskControlRelease_1_valid;
  wire [2:0]    maskControlRelease_2_bits;
  wire          maskControlRelease_2_valid;
  wire [2:0]    maskControlRelease_3_bits;
  wire          maskControlRelease_3_valid;
  wire          maskControlVec_releaseHit =
    maskControlRelease_0_valid & maskControlRelease_0_bits == maskControlVec_0_index | maskControlRelease_1_valid & maskControlRelease_1_bits == maskControlVec_0_index | maskControlRelease_2_valid
    & maskControlRelease_2_bits == maskControlVec_0_index | maskControlRelease_3_valid & maskControlRelease_3_bits == maskControlVec_0_index;
  reg           maskControlVec_responseFire_pipe_v;
  reg           maskControlVec_responseFire_pipe_pipe_v;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_v;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_pipe_v;
  wire          maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_valid = maskControlVec_responseFire_pipe_pipe_pipe_pipe_v;
  assign maskControlReq_0 = maskControlVec_0_controlValid & ~maskControlVec_0_dataValid & ~maskControlVec_0_waiteResponse;
  reg  [2:0]    maskControlVec_1_index;
  reg  [1:0]    maskControlVec_1_sew;
  reg  [31:0]   maskControlVec_1_maskData;
  reg  [7:0]    maskControlVec_1_group;
  reg           maskControlVec_1_dataValid;
  reg           maskControlVec_1_waiteResponse;
  reg           maskControlVec_1_controlValid;
  wire          maskControlVec_releaseHit_1 =
    maskControlRelease_0_valid & maskControlRelease_0_bits == maskControlVec_1_index | maskControlRelease_1_valid & maskControlRelease_1_bits == maskControlVec_1_index | maskControlRelease_2_valid
    & maskControlRelease_2_bits == maskControlVec_1_index | maskControlRelease_3_valid & maskControlRelease_3_bits == maskControlVec_1_index;
  reg           maskControlVec_responseFire_pipe_v_1;
  reg           maskControlVec_responseFire_pipe_pipe_v_1;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_v_1;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_1;
  wire          maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_1_valid = maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_1;
  assign maskControlReq_1 = maskControlVec_1_controlValid & ~maskControlVec_1_dataValid & ~maskControlVec_1_waiteResponse;
  reg  [2:0]    maskControlVec_2_index;
  reg  [1:0]    maskControlVec_2_sew;
  reg  [31:0]   maskControlVec_2_maskData;
  reg  [7:0]    maskControlVec_2_group;
  reg           maskControlVec_2_dataValid;
  reg           maskControlVec_2_waiteResponse;
  reg           maskControlVec_2_controlValid;
  wire          maskControlVec_releaseHit_2 =
    maskControlRelease_0_valid & maskControlRelease_0_bits == maskControlVec_2_index | maskControlRelease_1_valid & maskControlRelease_1_bits == maskControlVec_2_index | maskControlRelease_2_valid
    & maskControlRelease_2_bits == maskControlVec_2_index | maskControlRelease_3_valid & maskControlRelease_3_bits == maskControlVec_2_index;
  reg           maskControlVec_responseFire_pipe_v_2;
  reg           maskControlVec_responseFire_pipe_pipe_v_2;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_v_2;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_2;
  wire          maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_2_valid = maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_2;
  assign maskControlReq_2 = maskControlVec_2_controlValid & ~maskControlVec_2_dataValid & ~maskControlVec_2_waiteResponse;
  reg  [2:0]    maskControlVec_3_index;
  reg  [1:0]    maskControlVec_3_sew;
  reg  [31:0]   maskControlVec_3_maskData;
  reg  [7:0]    maskControlVec_3_group;
  reg           maskControlVec_3_dataValid;
  reg           maskControlVec_3_waiteResponse;
  reg           maskControlVec_3_controlValid;
  wire          maskControlVec_releaseHit_3 =
    maskControlRelease_0_valid & maskControlRelease_0_bits == maskControlVec_3_index | maskControlRelease_1_valid & maskControlRelease_1_bits == maskControlVec_3_index | maskControlRelease_2_valid
    & maskControlRelease_2_bits == maskControlVec_3_index | maskControlRelease_3_valid & maskControlRelease_3_bits == maskControlVec_3_index;
  reg           maskControlVec_responseFire_pipe_v_3;
  reg           maskControlVec_responseFire_pipe_pipe_v_3;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_v_3;
  reg           maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_3;
  wire          maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_3_valid = maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_3;
  assign maskControlReq_3 = maskControlVec_3_controlValid & ~maskControlVec_3_dataValid & ~maskControlVec_3_waiteResponse;
  wire          maskControlFree_0 = ~maskControlVec_0_controlValid & ~maskControlVec_0_waiteResponse;
  wire          maskControlFree_1 = ~maskControlVec_1_controlValid & ~maskControlVec_1_waiteResponse;
  wire          maskControlFree_2 = ~maskControlVec_2_controlValid & ~maskControlVec_2_waiteResponse;
  wire          maskControlFree_3 = ~maskControlVec_3_controlValid & ~maskControlVec_3_waiteResponse;
  wire [1:0]    freeSelect_lo = {maskControlFree_1, maskControlFree_0};
  wire [1:0]    freeSelect_hi = {maskControlFree_3, maskControlFree_2};
  wire [2:0]    _freeSelect_T_3 = {freeSelect_hi[0], freeSelect_lo} | {freeSelect_lo, 1'h0};
  wire [3:0]    freeSelect = {~(_freeSelect_T_3 | {_freeSelect_T_3[0], 2'h0}), 1'h1} & {freeSelect_hi, freeSelect_lo};
  wire          laneRequest_ready_0;
  wire [3:0]    maskControlEnq = laneRequest_ready_0 & laneRequest_valid_0 & laneRequest_bits_mask_0 ? freeSelect : 4'h0;
  wire          maskControlDataDeq_maskRequestFire;
  wire          maskControlDataDeq_maskRequestFire_1;
  wire          maskControlDataDeq_maskRequestFire_2;
  wire          maskControlDataDeq_maskRequestFire_3;
  wire [31:0]   maskControlDataDeq_data;
  wire [31:0]   maskControlDataDeq_data_1;
  wire [31:0]   maskControlDataDeq_data_2;
  wire [31:0]   maskControlDataDeq_data_3;
  reg  [2:0]    slotControl_0_laneRequest_instructionIndex;
  assign maskControlRelease_0_bits = slotControl_0_laneRequest_instructionIndex;
  wire [2:0]    laneState_instructionIndex = slotControl_0_laneRequest_instructionIndex;
  reg           slotControl_0_laneRequest_decodeResult_specialSlot;
  wire          laneState_decodeResult_specialSlot = slotControl_0_laneRequest_decodeResult_specialSlot;
  reg  [4:0]    slotControl_0_laneRequest_decodeResult_topUop;
  wire [4:0]    laneState_decodeResult_topUop = slotControl_0_laneRequest_decodeResult_topUop;
  reg           slotControl_0_laneRequest_decodeResult_popCount;
  wire          laneState_decodeResult_popCount = slotControl_0_laneRequest_decodeResult_popCount;
  reg           slotControl_0_laneRequest_decodeResult_ffo;
  wire          laneState_decodeResult_ffo = slotControl_0_laneRequest_decodeResult_ffo;
  reg           slotControl_0_laneRequest_decodeResult_average;
  wire          laneState_decodeResult_average = slotControl_0_laneRequest_decodeResult_average;
  reg           slotControl_0_laneRequest_decodeResult_reverse;
  wire          laneState_decodeResult_reverse = slotControl_0_laneRequest_decodeResult_reverse;
  reg           slotControl_0_laneRequest_decodeResult_dontNeedExecuteInLane;
  wire          laneState_decodeResult_dontNeedExecuteInLane = slotControl_0_laneRequest_decodeResult_dontNeedExecuteInLane;
  reg           slotControl_0_laneRequest_decodeResult_scheduler;
  wire          laneState_decodeResult_scheduler = slotControl_0_laneRequest_decodeResult_scheduler;
  reg           slotControl_0_laneRequest_decodeResult_sReadVD;
  wire          laneState_decodeResult_sReadVD = slotControl_0_laneRequest_decodeResult_sReadVD;
  reg           slotControl_0_laneRequest_decodeResult_vtype;
  wire          laneState_decodeResult_vtype = slotControl_0_laneRequest_decodeResult_vtype;
  reg           slotControl_0_laneRequest_decodeResult_sWrite;
  wire          laneState_decodeResult_sWrite = slotControl_0_laneRequest_decodeResult_sWrite;
  reg           slotControl_0_laneRequest_decodeResult_crossRead;
  wire          laneState_decodeResult_crossRead = slotControl_0_laneRequest_decodeResult_crossRead;
  reg           slotControl_0_laneRequest_decodeResult_crossWrite;
  wire          laneState_decodeResult_crossWrite = slotControl_0_laneRequest_decodeResult_crossWrite;
  reg           slotControl_0_laneRequest_decodeResult_maskUnit;
  wire          laneState_decodeResult_maskUnit = slotControl_0_laneRequest_decodeResult_maskUnit;
  reg           slotControl_0_laneRequest_decodeResult_special;
  wire          laneState_decodeResult_special = slotControl_0_laneRequest_decodeResult_special;
  reg           slotControl_0_laneRequest_decodeResult_saturate;
  wire          laneState_decodeResult_saturate = slotControl_0_laneRequest_decodeResult_saturate;
  reg           slotControl_0_laneRequest_decodeResult_vwmacc;
  wire          laneState_decodeResult_vwmacc = slotControl_0_laneRequest_decodeResult_vwmacc;
  reg           slotControl_0_laneRequest_decodeResult_readOnly;
  wire          laneState_decodeResult_readOnly = slotControl_0_laneRequest_decodeResult_readOnly;
  reg           slotControl_0_laneRequest_decodeResult_maskSource;
  wire          laneState_decodeResult_maskSource = slotControl_0_laneRequest_decodeResult_maskSource;
  reg           slotControl_0_laneRequest_decodeResult_maskDestination;
  wire          laneState_decodeResult_maskDestination = slotControl_0_laneRequest_decodeResult_maskDestination;
  reg           slotControl_0_laneRequest_decodeResult_maskLogic;
  wire          laneState_decodeResult_maskLogic = slotControl_0_laneRequest_decodeResult_maskLogic;
  reg  [3:0]    slotControl_0_laneRequest_decodeResult_uop;
  wire [3:0]    laneState_decodeResult_uop = slotControl_0_laneRequest_decodeResult_uop;
  reg           slotControl_0_laneRequest_decodeResult_iota;
  wire          laneState_decodeResult_iota = slotControl_0_laneRequest_decodeResult_iota;
  reg           slotControl_0_laneRequest_decodeResult_mv;
  wire          laneState_decodeResult_mv = slotControl_0_laneRequest_decodeResult_mv;
  reg           slotControl_0_laneRequest_decodeResult_extend;
  wire          laneState_decodeResult_extend = slotControl_0_laneRequest_decodeResult_extend;
  reg           slotControl_0_laneRequest_decodeResult_unOrderWrite;
  wire          laneState_decodeResult_unOrderWrite = slotControl_0_laneRequest_decodeResult_unOrderWrite;
  reg           slotControl_0_laneRequest_decodeResult_compress;
  wire          laneState_decodeResult_compress = slotControl_0_laneRequest_decodeResult_compress;
  reg           slotControl_0_laneRequest_decodeResult_gather16;
  wire          laneState_decodeResult_gather16 = slotControl_0_laneRequest_decodeResult_gather16;
  reg           slotControl_0_laneRequest_decodeResult_gather;
  wire          laneState_decodeResult_gather = slotControl_0_laneRequest_decodeResult_gather;
  reg           slotControl_0_laneRequest_decodeResult_slid;
  wire          laneState_decodeResult_slid = slotControl_0_laneRequest_decodeResult_slid;
  reg           slotControl_0_laneRequest_decodeResult_targetRd;
  wire          laneState_decodeResult_targetRd = slotControl_0_laneRequest_decodeResult_targetRd;
  reg           slotControl_0_laneRequest_decodeResult_widenReduce;
  wire          laneState_decodeResult_widenReduce = slotControl_0_laneRequest_decodeResult_widenReduce;
  reg           slotControl_0_laneRequest_decodeResult_red;
  wire          laneState_decodeResult_red = slotControl_0_laneRequest_decodeResult_red;
  reg           slotControl_0_laneRequest_decodeResult_nr;
  wire          laneState_decodeResult_nr = slotControl_0_laneRequest_decodeResult_nr;
  reg           slotControl_0_laneRequest_decodeResult_itype;
  wire          laneState_decodeResult_itype = slotControl_0_laneRequest_decodeResult_itype;
  reg           slotControl_0_laneRequest_decodeResult_unsigned1;
  wire          laneState_decodeResult_unsigned1 = slotControl_0_laneRequest_decodeResult_unsigned1;
  reg           slotControl_0_laneRequest_decodeResult_unsigned0;
  wire          laneState_decodeResult_unsigned0 = slotControl_0_laneRequest_decodeResult_unsigned0;
  reg           slotControl_0_laneRequest_decodeResult_other;
  wire          laneState_decodeResult_other = slotControl_0_laneRequest_decodeResult_other;
  reg           slotControl_0_laneRequest_decodeResult_multiCycle;
  wire          laneState_decodeResult_multiCycle = slotControl_0_laneRequest_decodeResult_multiCycle;
  reg           slotControl_0_laneRequest_decodeResult_divider;
  wire          laneState_decodeResult_divider = slotControl_0_laneRequest_decodeResult_divider;
  reg           slotControl_0_laneRequest_decodeResult_multiplier;
  wire          laneState_decodeResult_multiplier = slotControl_0_laneRequest_decodeResult_multiplier;
  reg           slotControl_0_laneRequest_decodeResult_shift;
  wire          laneState_decodeResult_shift = slotControl_0_laneRequest_decodeResult_shift;
  reg           slotControl_0_laneRequest_decodeResult_adder;
  wire          laneState_decodeResult_adder = slotControl_0_laneRequest_decodeResult_adder;
  reg           slotControl_0_laneRequest_decodeResult_logic;
  wire          laneState_decodeResult_logic = slotControl_0_laneRequest_decodeResult_logic;
  reg           slotControl_0_laneRequest_loadStore;
  wire          laneState_loadStore = slotControl_0_laneRequest_loadStore;
  reg           slotControl_0_laneRequest_issueInst;
  reg           slotControl_0_laneRequest_store;
  reg           slotControl_0_laneRequest_special;
  reg           slotControl_0_laneRequest_lsWholeReg;
  reg  [4:0]    slotControl_0_laneRequest_vs1;
  wire [4:0]    laneState_vs1 = slotControl_0_laneRequest_vs1;
  reg  [4:0]    slotControl_0_laneRequest_vs2;
  wire [4:0]    laneState_vs2 = slotControl_0_laneRequest_vs2;
  reg  [4:0]    slotControl_0_laneRequest_vd;
  wire [4:0]    laneState_vd = slotControl_0_laneRequest_vd;
  reg  [1:0]    slotControl_0_laneRequest_loadStoreEEW;
  reg           slotControl_0_laneRequest_mask;
  wire          laneState_maskType = slotControl_0_laneRequest_mask;
  reg  [2:0]    slotControl_0_laneRequest_segment;
  reg  [31:0]   slotControl_0_laneRequest_readFromScalar;
  reg  [13:0]   slotControl_0_laneRequest_csrInterface_vl;
  wire [13:0]   laneState_csr_vl = slotControl_0_laneRequest_csrInterface_vl;
  reg  [13:0]   slotControl_0_laneRequest_csrInterface_vStart;
  wire [13:0]   laneState_csr_vStart = slotControl_0_laneRequest_csrInterface_vStart;
  reg  [2:0]    slotControl_0_laneRequest_csrInterface_vlmul;
  wire [2:0]    laneState_csr_vlmul = slotControl_0_laneRequest_csrInterface_vlmul;
  reg  [1:0]    slotControl_0_laneRequest_csrInterface_vSew;
  wire [1:0]    laneState_csr_vSew = slotControl_0_laneRequest_csrInterface_vSew;
  reg  [1:0]    slotControl_0_laneRequest_csrInterface_vxrm;
  wire [1:0]    laneState_csr_vxrm = slotControl_0_laneRequest_csrInterface_vxrm;
  reg           slotControl_0_laneRequest_csrInterface_vta;
  wire          laneState_csr_vta = slotControl_0_laneRequest_csrInterface_vta;
  reg           slotControl_0_laneRequest_csrInterface_vma;
  wire          laneState_csr_vma = slotControl_0_laneRequest_csrInterface_vma;
  reg  [9:0]    slotControl_0_lastGroupForInstruction;
  wire [9:0]    laneState_lastGroupForInstruction = slotControl_0_lastGroupForInstruction;
  reg           slotControl_0_isLastLaneForInstruction;
  wire          laneState_isLastLaneForInstruction = slotControl_0_isLastLaneForInstruction;
  reg           slotControl_0_additionalRW;
  wire          laneState_additionalRW = slotControl_0_additionalRW;
  reg           slotControl_0_instructionFinished;
  wire          laneState_instructionFinished = slotControl_0_instructionFinished;
  reg           slotControl_0_mask_valid;
  reg  [31:0]   slotControl_0_mask_bits;
  reg  [2:0]    slotControl_1_laneRequest_instructionIndex;
  assign maskControlRelease_1_bits = slotControl_1_laneRequest_instructionIndex;
  wire [2:0]    laneState_1_instructionIndex = slotControl_1_laneRequest_instructionIndex;
  reg           slotControl_1_laneRequest_decodeResult_specialSlot;
  wire          laneState_1_decodeResult_specialSlot = slotControl_1_laneRequest_decodeResult_specialSlot;
  reg  [4:0]    slotControl_1_laneRequest_decodeResult_topUop;
  wire [4:0]    laneState_1_decodeResult_topUop = slotControl_1_laneRequest_decodeResult_topUop;
  reg           slotControl_1_laneRequest_decodeResult_popCount;
  wire          laneState_1_decodeResult_popCount = slotControl_1_laneRequest_decodeResult_popCount;
  reg           slotControl_1_laneRequest_decodeResult_ffo;
  wire          laneState_1_decodeResult_ffo = slotControl_1_laneRequest_decodeResult_ffo;
  reg           slotControl_1_laneRequest_decodeResult_average;
  wire          laneState_1_decodeResult_average = slotControl_1_laneRequest_decodeResult_average;
  reg           slotControl_1_laneRequest_decodeResult_reverse;
  wire          laneState_1_decodeResult_reverse = slotControl_1_laneRequest_decodeResult_reverse;
  reg           slotControl_1_laneRequest_decodeResult_dontNeedExecuteInLane;
  wire          laneState_1_decodeResult_dontNeedExecuteInLane = slotControl_1_laneRequest_decodeResult_dontNeedExecuteInLane;
  reg           slotControl_1_laneRequest_decodeResult_scheduler;
  wire          laneState_1_decodeResult_scheduler = slotControl_1_laneRequest_decodeResult_scheduler;
  reg           slotControl_1_laneRequest_decodeResult_sReadVD;
  wire          laneState_1_decodeResult_sReadVD = slotControl_1_laneRequest_decodeResult_sReadVD;
  reg           slotControl_1_laneRequest_decodeResult_vtype;
  wire          laneState_1_decodeResult_vtype = slotControl_1_laneRequest_decodeResult_vtype;
  reg           slotControl_1_laneRequest_decodeResult_sWrite;
  wire          laneState_1_decodeResult_sWrite = slotControl_1_laneRequest_decodeResult_sWrite;
  reg           slotControl_1_laneRequest_decodeResult_crossRead;
  wire          laneState_1_decodeResult_crossRead = slotControl_1_laneRequest_decodeResult_crossRead;
  reg           slotControl_1_laneRequest_decodeResult_crossWrite;
  wire          laneState_1_decodeResult_crossWrite = slotControl_1_laneRequest_decodeResult_crossWrite;
  reg           slotControl_1_laneRequest_decodeResult_maskUnit;
  wire          laneState_1_decodeResult_maskUnit = slotControl_1_laneRequest_decodeResult_maskUnit;
  reg           slotControl_1_laneRequest_decodeResult_special;
  wire          laneState_1_decodeResult_special = slotControl_1_laneRequest_decodeResult_special;
  reg           slotControl_1_laneRequest_decodeResult_saturate;
  wire          laneState_1_decodeResult_saturate = slotControl_1_laneRequest_decodeResult_saturate;
  reg           slotControl_1_laneRequest_decodeResult_vwmacc;
  wire          laneState_1_decodeResult_vwmacc = slotControl_1_laneRequest_decodeResult_vwmacc;
  reg           slotControl_1_laneRequest_decodeResult_readOnly;
  wire          laneState_1_decodeResult_readOnly = slotControl_1_laneRequest_decodeResult_readOnly;
  reg           slotControl_1_laneRequest_decodeResult_maskSource;
  wire          laneState_1_decodeResult_maskSource = slotControl_1_laneRequest_decodeResult_maskSource;
  reg           slotControl_1_laneRequest_decodeResult_maskDestination;
  wire          laneState_1_decodeResult_maskDestination = slotControl_1_laneRequest_decodeResult_maskDestination;
  reg           slotControl_1_laneRequest_decodeResult_maskLogic;
  wire          laneState_1_decodeResult_maskLogic = slotControl_1_laneRequest_decodeResult_maskLogic;
  reg  [3:0]    slotControl_1_laneRequest_decodeResult_uop;
  wire [3:0]    laneState_1_decodeResult_uop = slotControl_1_laneRequest_decodeResult_uop;
  reg           slotControl_1_laneRequest_decodeResult_iota;
  wire          laneState_1_decodeResult_iota = slotControl_1_laneRequest_decodeResult_iota;
  reg           slotControl_1_laneRequest_decodeResult_mv;
  wire          laneState_1_decodeResult_mv = slotControl_1_laneRequest_decodeResult_mv;
  reg           slotControl_1_laneRequest_decodeResult_extend;
  wire          laneState_1_decodeResult_extend = slotControl_1_laneRequest_decodeResult_extend;
  reg           slotControl_1_laneRequest_decodeResult_unOrderWrite;
  wire          laneState_1_decodeResult_unOrderWrite = slotControl_1_laneRequest_decodeResult_unOrderWrite;
  reg           slotControl_1_laneRequest_decodeResult_compress;
  wire          laneState_1_decodeResult_compress = slotControl_1_laneRequest_decodeResult_compress;
  reg           slotControl_1_laneRequest_decodeResult_gather16;
  wire          laneState_1_decodeResult_gather16 = slotControl_1_laneRequest_decodeResult_gather16;
  reg           slotControl_1_laneRequest_decodeResult_gather;
  wire          laneState_1_decodeResult_gather = slotControl_1_laneRequest_decodeResult_gather;
  reg           slotControl_1_laneRequest_decodeResult_slid;
  wire          laneState_1_decodeResult_slid = slotControl_1_laneRequest_decodeResult_slid;
  reg           slotControl_1_laneRequest_decodeResult_targetRd;
  wire          laneState_1_decodeResult_targetRd = slotControl_1_laneRequest_decodeResult_targetRd;
  reg           slotControl_1_laneRequest_decodeResult_widenReduce;
  wire          laneState_1_decodeResult_widenReduce = slotControl_1_laneRequest_decodeResult_widenReduce;
  reg           slotControl_1_laneRequest_decodeResult_red;
  wire          laneState_1_decodeResult_red = slotControl_1_laneRequest_decodeResult_red;
  reg           slotControl_1_laneRequest_decodeResult_nr;
  wire          laneState_1_decodeResult_nr = slotControl_1_laneRequest_decodeResult_nr;
  reg           slotControl_1_laneRequest_decodeResult_itype;
  wire          laneState_1_decodeResult_itype = slotControl_1_laneRequest_decodeResult_itype;
  reg           slotControl_1_laneRequest_decodeResult_unsigned1;
  wire          laneState_1_decodeResult_unsigned1 = slotControl_1_laneRequest_decodeResult_unsigned1;
  reg           slotControl_1_laneRequest_decodeResult_unsigned0;
  wire          laneState_1_decodeResult_unsigned0 = slotControl_1_laneRequest_decodeResult_unsigned0;
  reg           slotControl_1_laneRequest_decodeResult_other;
  wire          laneState_1_decodeResult_other = slotControl_1_laneRequest_decodeResult_other;
  reg           slotControl_1_laneRequest_decodeResult_multiCycle;
  wire          laneState_1_decodeResult_multiCycle = slotControl_1_laneRequest_decodeResult_multiCycle;
  reg           slotControl_1_laneRequest_decodeResult_divider;
  wire          laneState_1_decodeResult_divider = slotControl_1_laneRequest_decodeResult_divider;
  reg           slotControl_1_laneRequest_decodeResult_multiplier;
  wire          laneState_1_decodeResult_multiplier = slotControl_1_laneRequest_decodeResult_multiplier;
  reg           slotControl_1_laneRequest_decodeResult_shift;
  wire          laneState_1_decodeResult_shift = slotControl_1_laneRequest_decodeResult_shift;
  reg           slotControl_1_laneRequest_decodeResult_adder;
  wire          laneState_1_decodeResult_adder = slotControl_1_laneRequest_decodeResult_adder;
  reg           slotControl_1_laneRequest_decodeResult_logic;
  wire          laneState_1_decodeResult_logic = slotControl_1_laneRequest_decodeResult_logic;
  reg           slotControl_1_laneRequest_loadStore;
  wire          laneState_1_loadStore = slotControl_1_laneRequest_loadStore;
  reg           slotControl_1_laneRequest_issueInst;
  reg           slotControl_1_laneRequest_store;
  reg           slotControl_1_laneRequest_special;
  reg           slotControl_1_laneRequest_lsWholeReg;
  reg  [4:0]    slotControl_1_laneRequest_vs1;
  wire [4:0]    laneState_1_vs1 = slotControl_1_laneRequest_vs1;
  reg  [4:0]    slotControl_1_laneRequest_vs2;
  wire [4:0]    laneState_1_vs2 = slotControl_1_laneRequest_vs2;
  reg  [4:0]    slotControl_1_laneRequest_vd;
  wire [4:0]    laneState_1_vd = slotControl_1_laneRequest_vd;
  reg  [1:0]    slotControl_1_laneRequest_loadStoreEEW;
  reg           slotControl_1_laneRequest_mask;
  wire          laneState_1_maskType = slotControl_1_laneRequest_mask;
  reg  [2:0]    slotControl_1_laneRequest_segment;
  reg  [31:0]   slotControl_1_laneRequest_readFromScalar;
  reg  [13:0]   slotControl_1_laneRequest_csrInterface_vl;
  wire [13:0]   laneState_1_csr_vl = slotControl_1_laneRequest_csrInterface_vl;
  reg  [13:0]   slotControl_1_laneRequest_csrInterface_vStart;
  wire [13:0]   laneState_1_csr_vStart = slotControl_1_laneRequest_csrInterface_vStart;
  reg  [2:0]    slotControl_1_laneRequest_csrInterface_vlmul;
  wire [2:0]    laneState_1_csr_vlmul = slotControl_1_laneRequest_csrInterface_vlmul;
  reg  [1:0]    slotControl_1_laneRequest_csrInterface_vSew;
  wire [1:0]    laneState_1_csr_vSew = slotControl_1_laneRequest_csrInterface_vSew;
  reg  [1:0]    slotControl_1_laneRequest_csrInterface_vxrm;
  wire [1:0]    laneState_1_csr_vxrm = slotControl_1_laneRequest_csrInterface_vxrm;
  reg           slotControl_1_laneRequest_csrInterface_vta;
  wire          laneState_1_csr_vta = slotControl_1_laneRequest_csrInterface_vta;
  reg           slotControl_1_laneRequest_csrInterface_vma;
  wire          laneState_1_csr_vma = slotControl_1_laneRequest_csrInterface_vma;
  reg  [9:0]    slotControl_1_lastGroupForInstruction;
  wire [9:0]    laneState_1_lastGroupForInstruction = slotControl_1_lastGroupForInstruction;
  reg           slotControl_1_isLastLaneForInstruction;
  wire          laneState_1_isLastLaneForInstruction = slotControl_1_isLastLaneForInstruction;
  reg           slotControl_1_additionalRW;
  wire          laneState_1_additionalRW = slotControl_1_additionalRW;
  reg           slotControl_1_instructionFinished;
  wire          laneState_1_instructionFinished = slotControl_1_instructionFinished;
  reg           slotControl_1_mask_valid;
  reg  [31:0]   slotControl_1_mask_bits;
  reg  [2:0]    slotControl_2_laneRequest_instructionIndex;
  assign maskControlRelease_2_bits = slotControl_2_laneRequest_instructionIndex;
  wire [2:0]    laneState_2_instructionIndex = slotControl_2_laneRequest_instructionIndex;
  reg           slotControl_2_laneRequest_decodeResult_specialSlot;
  wire          laneState_2_decodeResult_specialSlot = slotControl_2_laneRequest_decodeResult_specialSlot;
  reg  [4:0]    slotControl_2_laneRequest_decodeResult_topUop;
  wire [4:0]    laneState_2_decodeResult_topUop = slotControl_2_laneRequest_decodeResult_topUop;
  reg           slotControl_2_laneRequest_decodeResult_popCount;
  wire          laneState_2_decodeResult_popCount = slotControl_2_laneRequest_decodeResult_popCount;
  reg           slotControl_2_laneRequest_decodeResult_ffo;
  wire          laneState_2_decodeResult_ffo = slotControl_2_laneRequest_decodeResult_ffo;
  reg           slotControl_2_laneRequest_decodeResult_average;
  wire          laneState_2_decodeResult_average = slotControl_2_laneRequest_decodeResult_average;
  reg           slotControl_2_laneRequest_decodeResult_reverse;
  wire          laneState_2_decodeResult_reverse = slotControl_2_laneRequest_decodeResult_reverse;
  reg           slotControl_2_laneRequest_decodeResult_dontNeedExecuteInLane;
  wire          laneState_2_decodeResult_dontNeedExecuteInLane = slotControl_2_laneRequest_decodeResult_dontNeedExecuteInLane;
  reg           slotControl_2_laneRequest_decodeResult_scheduler;
  wire          laneState_2_decodeResult_scheduler = slotControl_2_laneRequest_decodeResult_scheduler;
  reg           slotControl_2_laneRequest_decodeResult_sReadVD;
  wire          laneState_2_decodeResult_sReadVD = slotControl_2_laneRequest_decodeResult_sReadVD;
  reg           slotControl_2_laneRequest_decodeResult_vtype;
  wire          laneState_2_decodeResult_vtype = slotControl_2_laneRequest_decodeResult_vtype;
  reg           slotControl_2_laneRequest_decodeResult_sWrite;
  wire          laneState_2_decodeResult_sWrite = slotControl_2_laneRequest_decodeResult_sWrite;
  reg           slotControl_2_laneRequest_decodeResult_crossRead;
  wire          laneState_2_decodeResult_crossRead = slotControl_2_laneRequest_decodeResult_crossRead;
  reg           slotControl_2_laneRequest_decodeResult_crossWrite;
  wire          laneState_2_decodeResult_crossWrite = slotControl_2_laneRequest_decodeResult_crossWrite;
  reg           slotControl_2_laneRequest_decodeResult_maskUnit;
  wire          laneState_2_decodeResult_maskUnit = slotControl_2_laneRequest_decodeResult_maskUnit;
  reg           slotControl_2_laneRequest_decodeResult_special;
  wire          laneState_2_decodeResult_special = slotControl_2_laneRequest_decodeResult_special;
  reg           slotControl_2_laneRequest_decodeResult_saturate;
  wire          laneState_2_decodeResult_saturate = slotControl_2_laneRequest_decodeResult_saturate;
  reg           slotControl_2_laneRequest_decodeResult_vwmacc;
  wire          laneState_2_decodeResult_vwmacc = slotControl_2_laneRequest_decodeResult_vwmacc;
  reg           slotControl_2_laneRequest_decodeResult_readOnly;
  wire          laneState_2_decodeResult_readOnly = slotControl_2_laneRequest_decodeResult_readOnly;
  reg           slotControl_2_laneRequest_decodeResult_maskSource;
  wire          laneState_2_decodeResult_maskSource = slotControl_2_laneRequest_decodeResult_maskSource;
  reg           slotControl_2_laneRequest_decodeResult_maskDestination;
  wire          laneState_2_decodeResult_maskDestination = slotControl_2_laneRequest_decodeResult_maskDestination;
  reg           slotControl_2_laneRequest_decodeResult_maskLogic;
  wire          laneState_2_decodeResult_maskLogic = slotControl_2_laneRequest_decodeResult_maskLogic;
  reg  [3:0]    slotControl_2_laneRequest_decodeResult_uop;
  wire [3:0]    laneState_2_decodeResult_uop = slotControl_2_laneRequest_decodeResult_uop;
  reg           slotControl_2_laneRequest_decodeResult_iota;
  wire          laneState_2_decodeResult_iota = slotControl_2_laneRequest_decodeResult_iota;
  reg           slotControl_2_laneRequest_decodeResult_mv;
  wire          laneState_2_decodeResult_mv = slotControl_2_laneRequest_decodeResult_mv;
  reg           slotControl_2_laneRequest_decodeResult_extend;
  wire          laneState_2_decodeResult_extend = slotControl_2_laneRequest_decodeResult_extend;
  reg           slotControl_2_laneRequest_decodeResult_unOrderWrite;
  wire          laneState_2_decodeResult_unOrderWrite = slotControl_2_laneRequest_decodeResult_unOrderWrite;
  reg           slotControl_2_laneRequest_decodeResult_compress;
  wire          laneState_2_decodeResult_compress = slotControl_2_laneRequest_decodeResult_compress;
  reg           slotControl_2_laneRequest_decodeResult_gather16;
  wire          laneState_2_decodeResult_gather16 = slotControl_2_laneRequest_decodeResult_gather16;
  reg           slotControl_2_laneRequest_decodeResult_gather;
  wire          laneState_2_decodeResult_gather = slotControl_2_laneRequest_decodeResult_gather;
  reg           slotControl_2_laneRequest_decodeResult_slid;
  wire          laneState_2_decodeResult_slid = slotControl_2_laneRequest_decodeResult_slid;
  reg           slotControl_2_laneRequest_decodeResult_targetRd;
  wire          laneState_2_decodeResult_targetRd = slotControl_2_laneRequest_decodeResult_targetRd;
  reg           slotControl_2_laneRequest_decodeResult_widenReduce;
  wire          laneState_2_decodeResult_widenReduce = slotControl_2_laneRequest_decodeResult_widenReduce;
  reg           slotControl_2_laneRequest_decodeResult_red;
  wire          laneState_2_decodeResult_red = slotControl_2_laneRequest_decodeResult_red;
  reg           slotControl_2_laneRequest_decodeResult_nr;
  wire          laneState_2_decodeResult_nr = slotControl_2_laneRequest_decodeResult_nr;
  reg           slotControl_2_laneRequest_decodeResult_itype;
  wire          laneState_2_decodeResult_itype = slotControl_2_laneRequest_decodeResult_itype;
  reg           slotControl_2_laneRequest_decodeResult_unsigned1;
  wire          laneState_2_decodeResult_unsigned1 = slotControl_2_laneRequest_decodeResult_unsigned1;
  reg           slotControl_2_laneRequest_decodeResult_unsigned0;
  wire          laneState_2_decodeResult_unsigned0 = slotControl_2_laneRequest_decodeResult_unsigned0;
  reg           slotControl_2_laneRequest_decodeResult_other;
  wire          laneState_2_decodeResult_other = slotControl_2_laneRequest_decodeResult_other;
  reg           slotControl_2_laneRequest_decodeResult_multiCycle;
  wire          laneState_2_decodeResult_multiCycle = slotControl_2_laneRequest_decodeResult_multiCycle;
  reg           slotControl_2_laneRequest_decodeResult_divider;
  wire          laneState_2_decodeResult_divider = slotControl_2_laneRequest_decodeResult_divider;
  reg           slotControl_2_laneRequest_decodeResult_multiplier;
  wire          laneState_2_decodeResult_multiplier = slotControl_2_laneRequest_decodeResult_multiplier;
  reg           slotControl_2_laneRequest_decodeResult_shift;
  wire          laneState_2_decodeResult_shift = slotControl_2_laneRequest_decodeResult_shift;
  reg           slotControl_2_laneRequest_decodeResult_adder;
  wire          laneState_2_decodeResult_adder = slotControl_2_laneRequest_decodeResult_adder;
  reg           slotControl_2_laneRequest_decodeResult_logic;
  wire          laneState_2_decodeResult_logic = slotControl_2_laneRequest_decodeResult_logic;
  reg           slotControl_2_laneRequest_loadStore;
  wire          laneState_2_loadStore = slotControl_2_laneRequest_loadStore;
  reg           slotControl_2_laneRequest_issueInst;
  reg           slotControl_2_laneRequest_store;
  reg           slotControl_2_laneRequest_special;
  reg           slotControl_2_laneRequest_lsWholeReg;
  reg  [4:0]    slotControl_2_laneRequest_vs1;
  wire [4:0]    laneState_2_vs1 = slotControl_2_laneRequest_vs1;
  reg  [4:0]    slotControl_2_laneRequest_vs2;
  wire [4:0]    laneState_2_vs2 = slotControl_2_laneRequest_vs2;
  reg  [4:0]    slotControl_2_laneRequest_vd;
  wire [4:0]    laneState_2_vd = slotControl_2_laneRequest_vd;
  reg  [1:0]    slotControl_2_laneRequest_loadStoreEEW;
  reg           slotControl_2_laneRequest_mask;
  wire          laneState_2_maskType = slotControl_2_laneRequest_mask;
  reg  [2:0]    slotControl_2_laneRequest_segment;
  reg  [31:0]   slotControl_2_laneRequest_readFromScalar;
  reg  [13:0]   slotControl_2_laneRequest_csrInterface_vl;
  wire [13:0]   laneState_2_csr_vl = slotControl_2_laneRequest_csrInterface_vl;
  reg  [13:0]   slotControl_2_laneRequest_csrInterface_vStart;
  wire [13:0]   laneState_2_csr_vStart = slotControl_2_laneRequest_csrInterface_vStart;
  reg  [2:0]    slotControl_2_laneRequest_csrInterface_vlmul;
  wire [2:0]    laneState_2_csr_vlmul = slotControl_2_laneRequest_csrInterface_vlmul;
  reg  [1:0]    slotControl_2_laneRequest_csrInterface_vSew;
  wire [1:0]    laneState_2_csr_vSew = slotControl_2_laneRequest_csrInterface_vSew;
  reg  [1:0]    slotControl_2_laneRequest_csrInterface_vxrm;
  wire [1:0]    laneState_2_csr_vxrm = slotControl_2_laneRequest_csrInterface_vxrm;
  reg           slotControl_2_laneRequest_csrInterface_vta;
  wire          laneState_2_csr_vta = slotControl_2_laneRequest_csrInterface_vta;
  reg           slotControl_2_laneRequest_csrInterface_vma;
  wire          laneState_2_csr_vma = slotControl_2_laneRequest_csrInterface_vma;
  reg  [9:0]    slotControl_2_lastGroupForInstruction;
  wire [9:0]    laneState_2_lastGroupForInstruction = slotControl_2_lastGroupForInstruction;
  reg           slotControl_2_isLastLaneForInstruction;
  wire          laneState_2_isLastLaneForInstruction = slotControl_2_isLastLaneForInstruction;
  reg           slotControl_2_additionalRW;
  wire          laneState_2_additionalRW = slotControl_2_additionalRW;
  reg           slotControl_2_instructionFinished;
  wire          laneState_2_instructionFinished = slotControl_2_instructionFinished;
  reg           slotControl_2_mask_valid;
  reg  [31:0]   slotControl_2_mask_bits;
  reg  [2:0]    slotControl_3_laneRequest_instructionIndex;
  assign maskControlRelease_3_bits = slotControl_3_laneRequest_instructionIndex;
  wire [2:0]    laneState_3_instructionIndex = slotControl_3_laneRequest_instructionIndex;
  reg           slotControl_3_laneRequest_decodeResult_specialSlot;
  wire          laneState_3_decodeResult_specialSlot = slotControl_3_laneRequest_decodeResult_specialSlot;
  reg  [4:0]    slotControl_3_laneRequest_decodeResult_topUop;
  wire [4:0]    laneState_3_decodeResult_topUop = slotControl_3_laneRequest_decodeResult_topUop;
  reg           slotControl_3_laneRequest_decodeResult_popCount;
  wire          laneState_3_decodeResult_popCount = slotControl_3_laneRequest_decodeResult_popCount;
  reg           slotControl_3_laneRequest_decodeResult_ffo;
  wire          laneState_3_decodeResult_ffo = slotControl_3_laneRequest_decodeResult_ffo;
  reg           slotControl_3_laneRequest_decodeResult_average;
  wire          laneState_3_decodeResult_average = slotControl_3_laneRequest_decodeResult_average;
  reg           slotControl_3_laneRequest_decodeResult_reverse;
  wire          laneState_3_decodeResult_reverse = slotControl_3_laneRequest_decodeResult_reverse;
  reg           slotControl_3_laneRequest_decodeResult_dontNeedExecuteInLane;
  wire          laneState_3_decodeResult_dontNeedExecuteInLane = slotControl_3_laneRequest_decodeResult_dontNeedExecuteInLane;
  reg           slotControl_3_laneRequest_decodeResult_scheduler;
  wire          laneState_3_decodeResult_scheduler = slotControl_3_laneRequest_decodeResult_scheduler;
  reg           slotControl_3_laneRequest_decodeResult_sReadVD;
  wire          laneState_3_decodeResult_sReadVD = slotControl_3_laneRequest_decodeResult_sReadVD;
  reg           slotControl_3_laneRequest_decodeResult_vtype;
  wire          laneState_3_decodeResult_vtype = slotControl_3_laneRequest_decodeResult_vtype;
  reg           slotControl_3_laneRequest_decodeResult_sWrite;
  wire          laneState_3_decodeResult_sWrite = slotControl_3_laneRequest_decodeResult_sWrite;
  reg           slotControl_3_laneRequest_decodeResult_crossRead;
  wire          laneState_3_decodeResult_crossRead = slotControl_3_laneRequest_decodeResult_crossRead;
  reg           slotControl_3_laneRequest_decodeResult_crossWrite;
  wire          laneState_3_decodeResult_crossWrite = slotControl_3_laneRequest_decodeResult_crossWrite;
  reg           slotControl_3_laneRequest_decodeResult_maskUnit;
  wire          laneState_3_decodeResult_maskUnit = slotControl_3_laneRequest_decodeResult_maskUnit;
  reg           slotControl_3_laneRequest_decodeResult_special;
  wire          laneState_3_decodeResult_special = slotControl_3_laneRequest_decodeResult_special;
  reg           slotControl_3_laneRequest_decodeResult_saturate;
  wire          laneState_3_decodeResult_saturate = slotControl_3_laneRequest_decodeResult_saturate;
  reg           slotControl_3_laneRequest_decodeResult_vwmacc;
  wire          laneState_3_decodeResult_vwmacc = slotControl_3_laneRequest_decodeResult_vwmacc;
  reg           slotControl_3_laneRequest_decodeResult_readOnly;
  wire          laneState_3_decodeResult_readOnly = slotControl_3_laneRequest_decodeResult_readOnly;
  reg           slotControl_3_laneRequest_decodeResult_maskSource;
  wire          laneState_3_decodeResult_maskSource = slotControl_3_laneRequest_decodeResult_maskSource;
  reg           slotControl_3_laneRequest_decodeResult_maskDestination;
  wire          laneState_3_decodeResult_maskDestination = slotControl_3_laneRequest_decodeResult_maskDestination;
  reg           slotControl_3_laneRequest_decodeResult_maskLogic;
  wire          laneState_3_decodeResult_maskLogic = slotControl_3_laneRequest_decodeResult_maskLogic;
  reg  [3:0]    slotControl_3_laneRequest_decodeResult_uop;
  wire [3:0]    laneState_3_decodeResult_uop = slotControl_3_laneRequest_decodeResult_uop;
  reg           slotControl_3_laneRequest_decodeResult_iota;
  wire          laneState_3_decodeResult_iota = slotControl_3_laneRequest_decodeResult_iota;
  reg           slotControl_3_laneRequest_decodeResult_mv;
  wire          laneState_3_decodeResult_mv = slotControl_3_laneRequest_decodeResult_mv;
  reg           slotControl_3_laneRequest_decodeResult_extend;
  wire          laneState_3_decodeResult_extend = slotControl_3_laneRequest_decodeResult_extend;
  reg           slotControl_3_laneRequest_decodeResult_unOrderWrite;
  wire          laneState_3_decodeResult_unOrderWrite = slotControl_3_laneRequest_decodeResult_unOrderWrite;
  reg           slotControl_3_laneRequest_decodeResult_compress;
  wire          laneState_3_decodeResult_compress = slotControl_3_laneRequest_decodeResult_compress;
  reg           slotControl_3_laneRequest_decodeResult_gather16;
  wire          laneState_3_decodeResult_gather16 = slotControl_3_laneRequest_decodeResult_gather16;
  reg           slotControl_3_laneRequest_decodeResult_gather;
  wire          laneState_3_decodeResult_gather = slotControl_3_laneRequest_decodeResult_gather;
  reg           slotControl_3_laneRequest_decodeResult_slid;
  wire          laneState_3_decodeResult_slid = slotControl_3_laneRequest_decodeResult_slid;
  reg           slotControl_3_laneRequest_decodeResult_targetRd;
  wire          laneState_3_decodeResult_targetRd = slotControl_3_laneRequest_decodeResult_targetRd;
  reg           slotControl_3_laneRequest_decodeResult_widenReduce;
  wire          laneState_3_decodeResult_widenReduce = slotControl_3_laneRequest_decodeResult_widenReduce;
  reg           slotControl_3_laneRequest_decodeResult_red;
  wire          laneState_3_decodeResult_red = slotControl_3_laneRequest_decodeResult_red;
  reg           slotControl_3_laneRequest_decodeResult_nr;
  wire          laneState_3_decodeResult_nr = slotControl_3_laneRequest_decodeResult_nr;
  reg           slotControl_3_laneRequest_decodeResult_itype;
  wire          laneState_3_decodeResult_itype = slotControl_3_laneRequest_decodeResult_itype;
  reg           slotControl_3_laneRequest_decodeResult_unsigned1;
  wire          laneState_3_decodeResult_unsigned1 = slotControl_3_laneRequest_decodeResult_unsigned1;
  reg           slotControl_3_laneRequest_decodeResult_unsigned0;
  wire          laneState_3_decodeResult_unsigned0 = slotControl_3_laneRequest_decodeResult_unsigned0;
  reg           slotControl_3_laneRequest_decodeResult_other;
  wire          laneState_3_decodeResult_other = slotControl_3_laneRequest_decodeResult_other;
  reg           slotControl_3_laneRequest_decodeResult_multiCycle;
  wire          laneState_3_decodeResult_multiCycle = slotControl_3_laneRequest_decodeResult_multiCycle;
  reg           slotControl_3_laneRequest_decodeResult_divider;
  wire          laneState_3_decodeResult_divider = slotControl_3_laneRequest_decodeResult_divider;
  reg           slotControl_3_laneRequest_decodeResult_multiplier;
  wire          laneState_3_decodeResult_multiplier = slotControl_3_laneRequest_decodeResult_multiplier;
  reg           slotControl_3_laneRequest_decodeResult_shift;
  wire          laneState_3_decodeResult_shift = slotControl_3_laneRequest_decodeResult_shift;
  reg           slotControl_3_laneRequest_decodeResult_adder;
  wire          laneState_3_decodeResult_adder = slotControl_3_laneRequest_decodeResult_adder;
  reg           slotControl_3_laneRequest_decodeResult_logic;
  wire          laneState_3_decodeResult_logic = slotControl_3_laneRequest_decodeResult_logic;
  reg           slotControl_3_laneRequest_loadStore;
  wire          laneState_3_loadStore = slotControl_3_laneRequest_loadStore;
  reg           slotControl_3_laneRequest_issueInst;
  reg           slotControl_3_laneRequest_store;
  reg           slotControl_3_laneRequest_special;
  reg           slotControl_3_laneRequest_lsWholeReg;
  reg  [4:0]    slotControl_3_laneRequest_vs1;
  wire [4:0]    laneState_3_vs1 = slotControl_3_laneRequest_vs1;
  reg  [4:0]    slotControl_3_laneRequest_vs2;
  wire [4:0]    laneState_3_vs2 = slotControl_3_laneRequest_vs2;
  reg  [4:0]    slotControl_3_laneRequest_vd;
  wire [4:0]    laneState_3_vd = slotControl_3_laneRequest_vd;
  reg  [1:0]    slotControl_3_laneRequest_loadStoreEEW;
  reg           slotControl_3_laneRequest_mask;
  wire          laneState_3_maskType = slotControl_3_laneRequest_mask;
  reg  [2:0]    slotControl_3_laneRequest_segment;
  reg  [31:0]   slotControl_3_laneRequest_readFromScalar;
  reg  [13:0]   slotControl_3_laneRequest_csrInterface_vl;
  wire [13:0]   laneState_3_csr_vl = slotControl_3_laneRequest_csrInterface_vl;
  reg  [13:0]   slotControl_3_laneRequest_csrInterface_vStart;
  wire [13:0]   laneState_3_csr_vStart = slotControl_3_laneRequest_csrInterface_vStart;
  reg  [2:0]    slotControl_3_laneRequest_csrInterface_vlmul;
  wire [2:0]    laneState_3_csr_vlmul = slotControl_3_laneRequest_csrInterface_vlmul;
  reg  [1:0]    slotControl_3_laneRequest_csrInterface_vSew;
  wire [1:0]    laneState_3_csr_vSew = slotControl_3_laneRequest_csrInterface_vSew;
  reg  [1:0]    slotControl_3_laneRequest_csrInterface_vxrm;
  wire [1:0]    laneState_3_csr_vxrm = slotControl_3_laneRequest_csrInterface_vxrm;
  reg           slotControl_3_laneRequest_csrInterface_vta;
  wire          laneState_3_csr_vta = slotControl_3_laneRequest_csrInterface_vta;
  reg           slotControl_3_laneRequest_csrInterface_vma;
  wire          laneState_3_csr_vma = slotControl_3_laneRequest_csrInterface_vma;
  reg  [9:0]    slotControl_3_lastGroupForInstruction;
  wire [9:0]    laneState_3_lastGroupForInstruction = slotControl_3_lastGroupForInstruction;
  reg           slotControl_3_isLastLaneForInstruction;
  wire          laneState_3_isLastLaneForInstruction = slotControl_3_isLastLaneForInstruction;
  reg           slotControl_3_additionalRW;
  wire          laneState_3_additionalRW = slotControl_3_additionalRW;
  reg           slotControl_3_instructionFinished;
  wire          laneState_3_instructionFinished = slotControl_3_instructionFinished;
  reg           slotControl_3_mask_valid;
  reg  [31:0]   slotControl_3_mask_bits;
  wire          slotShiftValid_0;
  assign slotShiftValid_0 = ~slotOccupied_0;
  wire          enqueueReady = slotShiftValid_0;
  wire          enqueueReady_1 = slotShiftValid_1;
  wire          enqueueReady_2 = slotShiftValid_2;
  wire          enqueueReady_3 = slotShiftValid_3;
  wire          slotCanShift_0;
  assign slotCanShift_0 = ~slotOccupied_0;
  wire [32:0]   requestVecFromSlot_0_other_bits_src_0 = requestVec_0_src_0;
  wire [32:0]   requestVecFromSlot_0_divider_bits_src_0 = requestVec_0_src_0;
  wire [32:0]   requestVecFromSlot_0_multiplier_bits_src_0 = requestVec_0_src_0;
  wire [32:0]   requestVecFromSlot_0_shift_bits_src_0 = requestVec_0_src_0;
  wire [32:0]   requestVecFromSlot_0_adder_bits_src_0 = requestVec_0_src_0;
  wire [32:0]   requestVecFromSlot_0_logic_bits_src_0 = requestVec_0_src_0;
  wire [32:0]   requestVecFromSlot_0_other_bits_src_1 = requestVec_0_src_1;
  wire [32:0]   requestVecFromSlot_0_divider_bits_src_1 = requestVec_0_src_1;
  wire [32:0]   requestVecFromSlot_0_multiplier_bits_src_1 = requestVec_0_src_1;
  wire [32:0]   requestVecFromSlot_0_shift_bits_src_1 = requestVec_0_src_1;
  wire [32:0]   requestVecFromSlot_0_adder_bits_src_1 = requestVec_0_src_1;
  wire [32:0]   requestVecFromSlot_0_logic_bits_src_1 = requestVec_0_src_1;
  wire [32:0]   requestVecFromSlot_0_other_bits_src_2 = requestVec_0_src_2;
  wire [32:0]   requestVecFromSlot_0_divider_bits_src_2 = requestVec_0_src_2;
  wire [32:0]   requestVecFromSlot_0_multiplier_bits_src_2 = requestVec_0_src_2;
  wire [32:0]   requestVecFromSlot_0_shift_bits_src_2 = requestVec_0_src_2;
  wire [32:0]   requestVecFromSlot_0_adder_bits_src_2 = requestVec_0_src_2;
  wire [32:0]   requestVecFromSlot_0_logic_bits_src_2 = requestVec_0_src_2;
  wire [32:0]   requestVecFromSlot_0_other_bits_src_3 = requestVec_0_src_3;
  wire [32:0]   requestVecFromSlot_0_divider_bits_src_3 = requestVec_0_src_3;
  wire [32:0]   requestVecFromSlot_0_multiplier_bits_src_3 = requestVec_0_src_3;
  wire [32:0]   requestVecFromSlot_0_shift_bits_src_3 = requestVec_0_src_3;
  wire [32:0]   requestVecFromSlot_0_adder_bits_src_3 = requestVec_0_src_3;
  wire [32:0]   requestVecFromSlot_0_logic_bits_src_3 = requestVec_0_src_3;
  wire [3:0]    requestVecFromSlot_0_other_bits_opcode = requestVec_0_opcode;
  wire [3:0]    requestVecFromSlot_0_divider_bits_opcode = requestVec_0_opcode;
  wire [3:0]    requestVecFromSlot_0_multiplier_bits_opcode = requestVec_0_opcode;
  wire [3:0]    requestVecFromSlot_0_shift_bits_opcode = requestVec_0_opcode;
  wire [3:0]    requestVecFromSlot_0_adder_bits_opcode = requestVec_0_opcode;
  wire [3:0]    requestVecFromSlot_0_logic_bits_opcode = requestVec_0_opcode;
  wire [3:0]    requestVecFromSlot_0_other_bits_mask = requestVec_0_mask;
  wire [3:0]    requestVecFromSlot_0_divider_bits_mask = requestVec_0_mask;
  wire [3:0]    requestVecFromSlot_0_multiplier_bits_mask = requestVec_0_mask;
  wire [3:0]    requestVecFromSlot_0_shift_bits_mask = requestVec_0_mask;
  wire [3:0]    requestVecFromSlot_0_adder_bits_mask = requestVec_0_mask;
  wire [3:0]    requestVecFromSlot_0_logic_bits_mask = requestVec_0_mask;
  wire [3:0]    requestVecFromSlot_0_other_bits_executeMask = requestVec_0_executeMask;
  wire [3:0]    requestVecFromSlot_0_divider_bits_executeMask = requestVec_0_executeMask;
  wire [3:0]    requestVecFromSlot_0_multiplier_bits_executeMask = requestVec_0_executeMask;
  wire [3:0]    requestVecFromSlot_0_shift_bits_executeMask = requestVec_0_executeMask;
  wire [3:0]    requestVecFromSlot_0_adder_bits_executeMask = requestVec_0_executeMask;
  wire [3:0]    requestVecFromSlot_0_logic_bits_executeMask = requestVec_0_executeMask;
  wire          requestVecFromSlot_0_other_bits_sign0 = requestVec_0_sign0;
  wire          requestVecFromSlot_0_divider_bits_sign0 = requestVec_0_sign0;
  wire          requestVecFromSlot_0_multiplier_bits_sign0 = requestVec_0_sign0;
  wire          requestVecFromSlot_0_shift_bits_sign0 = requestVec_0_sign0;
  wire          requestVecFromSlot_0_adder_bits_sign0 = requestVec_0_sign0;
  wire          requestVecFromSlot_0_logic_bits_sign0 = requestVec_0_sign0;
  wire          requestVecFromSlot_0_other_bits_sign = requestVec_0_sign;
  wire          requestVecFromSlot_0_divider_bits_sign = requestVec_0_sign;
  wire          requestVecFromSlot_0_multiplier_bits_sign = requestVec_0_sign;
  wire          requestVecFromSlot_0_shift_bits_sign = requestVec_0_sign;
  wire          requestVecFromSlot_0_adder_bits_sign = requestVec_0_sign;
  wire          requestVecFromSlot_0_logic_bits_sign = requestVec_0_sign;
  wire          requestVecFromSlot_0_other_bits_reverse = requestVec_0_reverse;
  wire          requestVecFromSlot_0_divider_bits_reverse = requestVec_0_reverse;
  wire          requestVecFromSlot_0_multiplier_bits_reverse = requestVec_0_reverse;
  wire          requestVecFromSlot_0_shift_bits_reverse = requestVec_0_reverse;
  wire          requestVecFromSlot_0_adder_bits_reverse = requestVec_0_reverse;
  wire          requestVecFromSlot_0_logic_bits_reverse = requestVec_0_reverse;
  wire          requestVecFromSlot_0_other_bits_average = requestVec_0_average;
  wire          requestVecFromSlot_0_divider_bits_average = requestVec_0_average;
  wire          requestVecFromSlot_0_multiplier_bits_average = requestVec_0_average;
  wire          requestVecFromSlot_0_shift_bits_average = requestVec_0_average;
  wire          requestVecFromSlot_0_adder_bits_average = requestVec_0_average;
  wire          requestVecFromSlot_0_logic_bits_average = requestVec_0_average;
  wire          requestVecFromSlot_0_other_bits_saturate = requestVec_0_saturate;
  wire          requestVecFromSlot_0_divider_bits_saturate = requestVec_0_saturate;
  wire          requestVecFromSlot_0_multiplier_bits_saturate = requestVec_0_saturate;
  wire          requestVecFromSlot_0_shift_bits_saturate = requestVec_0_saturate;
  wire          requestVecFromSlot_0_adder_bits_saturate = requestVec_0_saturate;
  wire          requestVecFromSlot_0_logic_bits_saturate = requestVec_0_saturate;
  wire [1:0]    requestVecFromSlot_0_other_bits_vxrm = requestVec_0_vxrm;
  wire [1:0]    requestVecFromSlot_0_divider_bits_vxrm = requestVec_0_vxrm;
  wire [1:0]    requestVecFromSlot_0_multiplier_bits_vxrm = requestVec_0_vxrm;
  wire [1:0]    requestVecFromSlot_0_shift_bits_vxrm = requestVec_0_vxrm;
  wire [1:0]    requestVecFromSlot_0_adder_bits_vxrm = requestVec_0_vxrm;
  wire [1:0]    requestVecFromSlot_0_logic_bits_vxrm = requestVec_0_vxrm;
  wire [1:0]    requestVecFromSlot_0_other_bits_vSew = requestVec_0_vSew;
  wire [1:0]    requestVecFromSlot_0_divider_bits_vSew = requestVec_0_vSew;
  wire [1:0]    requestVecFromSlot_0_multiplier_bits_vSew = requestVec_0_vSew;
  wire [1:0]    requestVecFromSlot_0_shift_bits_vSew = requestVec_0_vSew;
  wire [1:0]    requestVecFromSlot_0_adder_bits_vSew = requestVec_0_vSew;
  wire [1:0]    requestVecFromSlot_0_logic_bits_vSew = requestVec_0_vSew;
  wire [19:0]   requestVecFromSlot_0_other_bits_shifterSize = requestVec_0_shifterSize;
  wire [19:0]   requestVecFromSlot_0_divider_bits_shifterSize = requestVec_0_shifterSize;
  wire [19:0]   requestVecFromSlot_0_multiplier_bits_shifterSize = requestVec_0_shifterSize;
  wire [19:0]   requestVecFromSlot_0_shift_bits_shifterSize = requestVec_0_shifterSize;
  wire [19:0]   requestVecFromSlot_0_adder_bits_shifterSize = requestVec_0_shifterSize;
  wire [19:0]   requestVecFromSlot_0_logic_bits_shifterSize = requestVec_0_shifterSize;
  wire          requestVecFromSlot_0_other_bits_rem = requestVec_0_rem;
  wire          requestVecFromSlot_0_divider_bits_rem = requestVec_0_rem;
  wire          requestVecFromSlot_0_multiplier_bits_rem = requestVec_0_rem;
  wire          requestVecFromSlot_0_shift_bits_rem = requestVec_0_rem;
  wire          requestVecFromSlot_0_adder_bits_rem = requestVec_0_rem;
  wire          requestVecFromSlot_0_logic_bits_rem = requestVec_0_rem;
  wire [1:0]    requestVecFromSlot_0_other_bits_executeIndex = requestVec_0_executeIndex;
  wire [1:0]    requestVecFromSlot_0_divider_bits_executeIndex = requestVec_0_executeIndex;
  wire [1:0]    requestVecFromSlot_0_multiplier_bits_executeIndex = requestVec_0_executeIndex;
  wire [1:0]    requestVecFromSlot_0_shift_bits_executeIndex = requestVec_0_executeIndex;
  wire [1:0]    requestVecFromSlot_0_adder_bits_executeIndex = requestVec_0_executeIndex;
  wire [1:0]    requestVecFromSlot_0_logic_bits_executeIndex = requestVec_0_executeIndex;
  wire [13:0]   requestVecFromSlot_0_other_bits_popInit = requestVec_0_popInit;
  wire [13:0]   requestVecFromSlot_0_divider_bits_popInit = requestVec_0_popInit;
  wire [13:0]   requestVecFromSlot_0_multiplier_bits_popInit = requestVec_0_popInit;
  wire [13:0]   requestVecFromSlot_0_shift_bits_popInit = requestVec_0_popInit;
  wire [13:0]   requestVecFromSlot_0_adder_bits_popInit = requestVec_0_popInit;
  wire [13:0]   requestVecFromSlot_0_logic_bits_popInit = requestVec_0_popInit;
  wire [9:0]    requestVecFromSlot_0_other_bits_groupIndex = requestVec_0_groupIndex;
  wire [9:0]    requestVecFromSlot_0_divider_bits_groupIndex = requestVec_0_groupIndex;
  wire [9:0]    requestVecFromSlot_0_multiplier_bits_groupIndex = requestVec_0_groupIndex;
  wire [9:0]    requestVecFromSlot_0_shift_bits_groupIndex = requestVec_0_groupIndex;
  wire [9:0]    requestVecFromSlot_0_adder_bits_groupIndex = requestVec_0_groupIndex;
  wire [9:0]    requestVecFromSlot_0_logic_bits_groupIndex = requestVec_0_groupIndex;
  wire [1:0]    requestVecFromSlot_0_other_bits_laneIndex = requestVec_0_laneIndex;
  wire [1:0]    requestVecFromSlot_0_divider_bits_laneIndex = requestVec_0_laneIndex;
  wire [1:0]    requestVecFromSlot_0_multiplier_bits_laneIndex = requestVec_0_laneIndex;
  wire [1:0]    requestVecFromSlot_0_shift_bits_laneIndex = requestVec_0_laneIndex;
  wire [1:0]    requestVecFromSlot_0_adder_bits_laneIndex = requestVec_0_laneIndex;
  wire [1:0]    requestVecFromSlot_0_logic_bits_laneIndex = requestVec_0_laneIndex;
  wire          requestVecFromSlot_0_other_bits_maskType = requestVec_0_maskType;
  wire          requestVecFromSlot_0_divider_bits_maskType = requestVec_0_maskType;
  wire          requestVecFromSlot_0_multiplier_bits_maskType = requestVec_0_maskType;
  wire          requestVecFromSlot_0_shift_bits_maskType = requestVec_0_maskType;
  wire          requestVecFromSlot_0_adder_bits_maskType = requestVec_0_maskType;
  wire          requestVecFromSlot_0_logic_bits_maskType = requestVec_0_maskType;
  wire          requestVecFromSlot_0_other_bits_narrow = requestVec_0_narrow;
  wire          requestVecFromSlot_0_divider_bits_narrow = requestVec_0_narrow;
  wire          requestVecFromSlot_0_multiplier_bits_narrow = requestVec_0_narrow;
  wire          requestVecFromSlot_0_shift_bits_narrow = requestVec_0_narrow;
  wire          requestVecFromSlot_0_adder_bits_narrow = requestVec_0_narrow;
  wire          requestVecFromSlot_0_logic_bits_narrow = requestVec_0_narrow;
  wire [32:0]   requestVecFromSlot_1_other_bits_src_0 = requestVec_1_src_0;
  wire [32:0]   requestVecFromSlot_1_divider_bits_src_0 = requestVec_1_src_0;
  wire [32:0]   requestVecFromSlot_1_multiplier_bits_src_0 = requestVec_1_src_0;
  wire [32:0]   requestVecFromSlot_1_shift_bits_src_0 = requestVec_1_src_0;
  wire [32:0]   requestVecFromSlot_1_adder_bits_src_0 = requestVec_1_src_0;
  wire [32:0]   requestVecFromSlot_1_logic_bits_src_0 = requestVec_1_src_0;
  wire [32:0]   requestVecFromSlot_1_other_bits_src_1 = requestVec_1_src_1;
  wire [32:0]   requestVecFromSlot_1_divider_bits_src_1 = requestVec_1_src_1;
  wire [32:0]   requestVecFromSlot_1_multiplier_bits_src_1 = requestVec_1_src_1;
  wire [32:0]   requestVecFromSlot_1_shift_bits_src_1 = requestVec_1_src_1;
  wire [32:0]   requestVecFromSlot_1_adder_bits_src_1 = requestVec_1_src_1;
  wire [32:0]   requestVecFromSlot_1_logic_bits_src_1 = requestVec_1_src_1;
  wire [32:0]   requestVecFromSlot_1_other_bits_src_2 = requestVec_1_src_2;
  wire [32:0]   requestVecFromSlot_1_divider_bits_src_2 = requestVec_1_src_2;
  wire [32:0]   requestVecFromSlot_1_multiplier_bits_src_2 = requestVec_1_src_2;
  wire [32:0]   requestVecFromSlot_1_shift_bits_src_2 = requestVec_1_src_2;
  wire [32:0]   requestVecFromSlot_1_adder_bits_src_2 = requestVec_1_src_2;
  wire [32:0]   requestVecFromSlot_1_logic_bits_src_2 = requestVec_1_src_2;
  wire [32:0]   requestVecFromSlot_1_other_bits_src_3 = requestVec_1_src_3;
  wire [32:0]   requestVecFromSlot_1_divider_bits_src_3 = requestVec_1_src_3;
  wire [32:0]   requestVecFromSlot_1_multiplier_bits_src_3 = requestVec_1_src_3;
  wire [32:0]   requestVecFromSlot_1_shift_bits_src_3 = requestVec_1_src_3;
  wire [32:0]   requestVecFromSlot_1_adder_bits_src_3 = requestVec_1_src_3;
  wire [32:0]   requestVecFromSlot_1_logic_bits_src_3 = requestVec_1_src_3;
  wire [3:0]    requestVecFromSlot_1_other_bits_opcode = requestVec_1_opcode;
  wire [3:0]    requestVecFromSlot_1_divider_bits_opcode = requestVec_1_opcode;
  wire [3:0]    requestVecFromSlot_1_multiplier_bits_opcode = requestVec_1_opcode;
  wire [3:0]    requestVecFromSlot_1_shift_bits_opcode = requestVec_1_opcode;
  wire [3:0]    requestVecFromSlot_1_adder_bits_opcode = requestVec_1_opcode;
  wire [3:0]    requestVecFromSlot_1_logic_bits_opcode = requestVec_1_opcode;
  wire [3:0]    requestVecFromSlot_1_other_bits_mask = requestVec_1_mask;
  wire [3:0]    requestVecFromSlot_1_divider_bits_mask = requestVec_1_mask;
  wire [3:0]    requestVecFromSlot_1_multiplier_bits_mask = requestVec_1_mask;
  wire [3:0]    requestVecFromSlot_1_shift_bits_mask = requestVec_1_mask;
  wire [3:0]    requestVecFromSlot_1_adder_bits_mask = requestVec_1_mask;
  wire [3:0]    requestVecFromSlot_1_logic_bits_mask = requestVec_1_mask;
  wire [3:0]    requestVecFromSlot_1_other_bits_executeMask = requestVec_1_executeMask;
  wire [3:0]    requestVecFromSlot_1_divider_bits_executeMask = requestVec_1_executeMask;
  wire [3:0]    requestVecFromSlot_1_multiplier_bits_executeMask = requestVec_1_executeMask;
  wire [3:0]    requestVecFromSlot_1_shift_bits_executeMask = requestVec_1_executeMask;
  wire [3:0]    requestVecFromSlot_1_adder_bits_executeMask = requestVec_1_executeMask;
  wire [3:0]    requestVecFromSlot_1_logic_bits_executeMask = requestVec_1_executeMask;
  wire          requestVecFromSlot_1_other_bits_sign0 = requestVec_1_sign0;
  wire          requestVecFromSlot_1_divider_bits_sign0 = requestVec_1_sign0;
  wire          requestVecFromSlot_1_multiplier_bits_sign0 = requestVec_1_sign0;
  wire          requestVecFromSlot_1_shift_bits_sign0 = requestVec_1_sign0;
  wire          requestVecFromSlot_1_adder_bits_sign0 = requestVec_1_sign0;
  wire          requestVecFromSlot_1_logic_bits_sign0 = requestVec_1_sign0;
  wire          requestVecFromSlot_1_other_bits_sign = requestVec_1_sign;
  wire          requestVecFromSlot_1_divider_bits_sign = requestVec_1_sign;
  wire          requestVecFromSlot_1_multiplier_bits_sign = requestVec_1_sign;
  wire          requestVecFromSlot_1_shift_bits_sign = requestVec_1_sign;
  wire          requestVecFromSlot_1_adder_bits_sign = requestVec_1_sign;
  wire          requestVecFromSlot_1_logic_bits_sign = requestVec_1_sign;
  wire          requestVecFromSlot_1_other_bits_reverse = requestVec_1_reverse;
  wire          requestVecFromSlot_1_divider_bits_reverse = requestVec_1_reverse;
  wire          requestVecFromSlot_1_multiplier_bits_reverse = requestVec_1_reverse;
  wire          requestVecFromSlot_1_shift_bits_reverse = requestVec_1_reverse;
  wire          requestVecFromSlot_1_adder_bits_reverse = requestVec_1_reverse;
  wire          requestVecFromSlot_1_logic_bits_reverse = requestVec_1_reverse;
  wire          requestVecFromSlot_1_other_bits_average = requestVec_1_average;
  wire          requestVecFromSlot_1_divider_bits_average = requestVec_1_average;
  wire          requestVecFromSlot_1_multiplier_bits_average = requestVec_1_average;
  wire          requestVecFromSlot_1_shift_bits_average = requestVec_1_average;
  wire          requestVecFromSlot_1_adder_bits_average = requestVec_1_average;
  wire          requestVecFromSlot_1_logic_bits_average = requestVec_1_average;
  wire          requestVecFromSlot_1_other_bits_saturate = requestVec_1_saturate;
  wire          requestVecFromSlot_1_divider_bits_saturate = requestVec_1_saturate;
  wire          requestVecFromSlot_1_multiplier_bits_saturate = requestVec_1_saturate;
  wire          requestVecFromSlot_1_shift_bits_saturate = requestVec_1_saturate;
  wire          requestVecFromSlot_1_adder_bits_saturate = requestVec_1_saturate;
  wire          requestVecFromSlot_1_logic_bits_saturate = requestVec_1_saturate;
  wire [1:0]    requestVecFromSlot_1_other_bits_vxrm = requestVec_1_vxrm;
  wire [1:0]    requestVecFromSlot_1_divider_bits_vxrm = requestVec_1_vxrm;
  wire [1:0]    requestVecFromSlot_1_multiplier_bits_vxrm = requestVec_1_vxrm;
  wire [1:0]    requestVecFromSlot_1_shift_bits_vxrm = requestVec_1_vxrm;
  wire [1:0]    requestVecFromSlot_1_adder_bits_vxrm = requestVec_1_vxrm;
  wire [1:0]    requestVecFromSlot_1_logic_bits_vxrm = requestVec_1_vxrm;
  wire [1:0]    requestVecFromSlot_1_other_bits_vSew = requestVec_1_vSew;
  wire [1:0]    requestVecFromSlot_1_divider_bits_vSew = requestVec_1_vSew;
  wire [1:0]    requestVecFromSlot_1_multiplier_bits_vSew = requestVec_1_vSew;
  wire [1:0]    requestVecFromSlot_1_shift_bits_vSew = requestVec_1_vSew;
  wire [1:0]    requestVecFromSlot_1_adder_bits_vSew = requestVec_1_vSew;
  wire [1:0]    requestVecFromSlot_1_logic_bits_vSew = requestVec_1_vSew;
  wire [19:0]   requestVecFromSlot_1_other_bits_shifterSize = requestVec_1_shifterSize;
  wire [19:0]   requestVecFromSlot_1_divider_bits_shifterSize = requestVec_1_shifterSize;
  wire [19:0]   requestVecFromSlot_1_multiplier_bits_shifterSize = requestVec_1_shifterSize;
  wire [19:0]   requestVecFromSlot_1_shift_bits_shifterSize = requestVec_1_shifterSize;
  wire [19:0]   requestVecFromSlot_1_adder_bits_shifterSize = requestVec_1_shifterSize;
  wire [19:0]   requestVecFromSlot_1_logic_bits_shifterSize = requestVec_1_shifterSize;
  wire          requestVecFromSlot_1_other_bits_rem = requestVec_1_rem;
  wire          requestVecFromSlot_1_divider_bits_rem = requestVec_1_rem;
  wire          requestVecFromSlot_1_multiplier_bits_rem = requestVec_1_rem;
  wire          requestVecFromSlot_1_shift_bits_rem = requestVec_1_rem;
  wire          requestVecFromSlot_1_adder_bits_rem = requestVec_1_rem;
  wire          requestVecFromSlot_1_logic_bits_rem = requestVec_1_rem;
  wire [9:0]    requestVecFromSlot_1_other_bits_groupIndex = requestVec_1_groupIndex;
  wire [9:0]    requestVecFromSlot_1_divider_bits_groupIndex = requestVec_1_groupIndex;
  wire [9:0]    requestVecFromSlot_1_multiplier_bits_groupIndex = requestVec_1_groupIndex;
  wire [9:0]    requestVecFromSlot_1_shift_bits_groupIndex = requestVec_1_groupIndex;
  wire [9:0]    requestVecFromSlot_1_adder_bits_groupIndex = requestVec_1_groupIndex;
  wire [9:0]    requestVecFromSlot_1_logic_bits_groupIndex = requestVec_1_groupIndex;
  wire [1:0]    requestVecFromSlot_1_other_bits_laneIndex = requestVec_1_laneIndex;
  wire [1:0]    requestVecFromSlot_1_divider_bits_laneIndex = requestVec_1_laneIndex;
  wire [1:0]    requestVecFromSlot_1_multiplier_bits_laneIndex = requestVec_1_laneIndex;
  wire [1:0]    requestVecFromSlot_1_shift_bits_laneIndex = requestVec_1_laneIndex;
  wire [1:0]    requestVecFromSlot_1_adder_bits_laneIndex = requestVec_1_laneIndex;
  wire [1:0]    requestVecFromSlot_1_logic_bits_laneIndex = requestVec_1_laneIndex;
  wire          requestVecFromSlot_1_other_bits_maskType = requestVec_1_maskType;
  wire          requestVecFromSlot_1_divider_bits_maskType = requestVec_1_maskType;
  wire          requestVecFromSlot_1_multiplier_bits_maskType = requestVec_1_maskType;
  wire          requestVecFromSlot_1_shift_bits_maskType = requestVec_1_maskType;
  wire          requestVecFromSlot_1_adder_bits_maskType = requestVec_1_maskType;
  wire          requestVecFromSlot_1_logic_bits_maskType = requestVec_1_maskType;
  wire          requestVecFromSlot_1_other_bits_narrow = requestVec_1_narrow;
  wire          requestVecFromSlot_1_divider_bits_narrow = requestVec_1_narrow;
  wire          requestVecFromSlot_1_multiplier_bits_narrow = requestVec_1_narrow;
  wire          requestVecFromSlot_1_shift_bits_narrow = requestVec_1_narrow;
  wire          requestVecFromSlot_1_adder_bits_narrow = requestVec_1_narrow;
  wire          requestVecFromSlot_1_logic_bits_narrow = requestVec_1_narrow;
  wire [32:0]   requestVecFromSlot_2_other_bits_src_0 = requestVec_2_src_0;
  wire [32:0]   requestVecFromSlot_2_divider_bits_src_0 = requestVec_2_src_0;
  wire [32:0]   requestVecFromSlot_2_multiplier_bits_src_0 = requestVec_2_src_0;
  wire [32:0]   requestVecFromSlot_2_shift_bits_src_0 = requestVec_2_src_0;
  wire [32:0]   requestVecFromSlot_2_adder_bits_src_0 = requestVec_2_src_0;
  wire [32:0]   requestVecFromSlot_2_logic_bits_src_0 = requestVec_2_src_0;
  wire [32:0]   requestVecFromSlot_2_other_bits_src_1 = requestVec_2_src_1;
  wire [32:0]   requestVecFromSlot_2_divider_bits_src_1 = requestVec_2_src_1;
  wire [32:0]   requestVecFromSlot_2_multiplier_bits_src_1 = requestVec_2_src_1;
  wire [32:0]   requestVecFromSlot_2_shift_bits_src_1 = requestVec_2_src_1;
  wire [32:0]   requestVecFromSlot_2_adder_bits_src_1 = requestVec_2_src_1;
  wire [32:0]   requestVecFromSlot_2_logic_bits_src_1 = requestVec_2_src_1;
  wire [32:0]   requestVecFromSlot_2_other_bits_src_2 = requestVec_2_src_2;
  wire [32:0]   requestVecFromSlot_2_divider_bits_src_2 = requestVec_2_src_2;
  wire [32:0]   requestVecFromSlot_2_multiplier_bits_src_2 = requestVec_2_src_2;
  wire [32:0]   requestVecFromSlot_2_shift_bits_src_2 = requestVec_2_src_2;
  wire [32:0]   requestVecFromSlot_2_adder_bits_src_2 = requestVec_2_src_2;
  wire [32:0]   requestVecFromSlot_2_logic_bits_src_2 = requestVec_2_src_2;
  wire [32:0]   requestVecFromSlot_2_other_bits_src_3 = requestVec_2_src_3;
  wire [32:0]   requestVecFromSlot_2_divider_bits_src_3 = requestVec_2_src_3;
  wire [32:0]   requestVecFromSlot_2_multiplier_bits_src_3 = requestVec_2_src_3;
  wire [32:0]   requestVecFromSlot_2_shift_bits_src_3 = requestVec_2_src_3;
  wire [32:0]   requestVecFromSlot_2_adder_bits_src_3 = requestVec_2_src_3;
  wire [32:0]   requestVecFromSlot_2_logic_bits_src_3 = requestVec_2_src_3;
  wire [3:0]    requestVecFromSlot_2_other_bits_opcode = requestVec_2_opcode;
  wire [3:0]    requestVecFromSlot_2_divider_bits_opcode = requestVec_2_opcode;
  wire [3:0]    requestVecFromSlot_2_multiplier_bits_opcode = requestVec_2_opcode;
  wire [3:0]    requestVecFromSlot_2_shift_bits_opcode = requestVec_2_opcode;
  wire [3:0]    requestVecFromSlot_2_adder_bits_opcode = requestVec_2_opcode;
  wire [3:0]    requestVecFromSlot_2_logic_bits_opcode = requestVec_2_opcode;
  wire [3:0]    requestVecFromSlot_2_other_bits_mask = requestVec_2_mask;
  wire [3:0]    requestVecFromSlot_2_divider_bits_mask = requestVec_2_mask;
  wire [3:0]    requestVecFromSlot_2_multiplier_bits_mask = requestVec_2_mask;
  wire [3:0]    requestVecFromSlot_2_shift_bits_mask = requestVec_2_mask;
  wire [3:0]    requestVecFromSlot_2_adder_bits_mask = requestVec_2_mask;
  wire [3:0]    requestVecFromSlot_2_logic_bits_mask = requestVec_2_mask;
  wire [3:0]    requestVecFromSlot_2_other_bits_executeMask = requestVec_2_executeMask;
  wire [3:0]    requestVecFromSlot_2_divider_bits_executeMask = requestVec_2_executeMask;
  wire [3:0]    requestVecFromSlot_2_multiplier_bits_executeMask = requestVec_2_executeMask;
  wire [3:0]    requestVecFromSlot_2_shift_bits_executeMask = requestVec_2_executeMask;
  wire [3:0]    requestVecFromSlot_2_adder_bits_executeMask = requestVec_2_executeMask;
  wire [3:0]    requestVecFromSlot_2_logic_bits_executeMask = requestVec_2_executeMask;
  wire          requestVecFromSlot_2_other_bits_sign0 = requestVec_2_sign0;
  wire          requestVecFromSlot_2_divider_bits_sign0 = requestVec_2_sign0;
  wire          requestVecFromSlot_2_multiplier_bits_sign0 = requestVec_2_sign0;
  wire          requestVecFromSlot_2_shift_bits_sign0 = requestVec_2_sign0;
  wire          requestVecFromSlot_2_adder_bits_sign0 = requestVec_2_sign0;
  wire          requestVecFromSlot_2_logic_bits_sign0 = requestVec_2_sign0;
  wire          requestVecFromSlot_2_other_bits_sign = requestVec_2_sign;
  wire          requestVecFromSlot_2_divider_bits_sign = requestVec_2_sign;
  wire          requestVecFromSlot_2_multiplier_bits_sign = requestVec_2_sign;
  wire          requestVecFromSlot_2_shift_bits_sign = requestVec_2_sign;
  wire          requestVecFromSlot_2_adder_bits_sign = requestVec_2_sign;
  wire          requestVecFromSlot_2_logic_bits_sign = requestVec_2_sign;
  wire          requestVecFromSlot_2_other_bits_reverse = requestVec_2_reverse;
  wire          requestVecFromSlot_2_divider_bits_reverse = requestVec_2_reverse;
  wire          requestVecFromSlot_2_multiplier_bits_reverse = requestVec_2_reverse;
  wire          requestVecFromSlot_2_shift_bits_reverse = requestVec_2_reverse;
  wire          requestVecFromSlot_2_adder_bits_reverse = requestVec_2_reverse;
  wire          requestVecFromSlot_2_logic_bits_reverse = requestVec_2_reverse;
  wire          requestVecFromSlot_2_other_bits_average = requestVec_2_average;
  wire          requestVecFromSlot_2_divider_bits_average = requestVec_2_average;
  wire          requestVecFromSlot_2_multiplier_bits_average = requestVec_2_average;
  wire          requestVecFromSlot_2_shift_bits_average = requestVec_2_average;
  wire          requestVecFromSlot_2_adder_bits_average = requestVec_2_average;
  wire          requestVecFromSlot_2_logic_bits_average = requestVec_2_average;
  wire          requestVecFromSlot_2_other_bits_saturate = requestVec_2_saturate;
  wire          requestVecFromSlot_2_divider_bits_saturate = requestVec_2_saturate;
  wire          requestVecFromSlot_2_multiplier_bits_saturate = requestVec_2_saturate;
  wire          requestVecFromSlot_2_shift_bits_saturate = requestVec_2_saturate;
  wire          requestVecFromSlot_2_adder_bits_saturate = requestVec_2_saturate;
  wire          requestVecFromSlot_2_logic_bits_saturate = requestVec_2_saturate;
  wire [1:0]    requestVecFromSlot_2_other_bits_vxrm = requestVec_2_vxrm;
  wire [1:0]    requestVecFromSlot_2_divider_bits_vxrm = requestVec_2_vxrm;
  wire [1:0]    requestVecFromSlot_2_multiplier_bits_vxrm = requestVec_2_vxrm;
  wire [1:0]    requestVecFromSlot_2_shift_bits_vxrm = requestVec_2_vxrm;
  wire [1:0]    requestVecFromSlot_2_adder_bits_vxrm = requestVec_2_vxrm;
  wire [1:0]    requestVecFromSlot_2_logic_bits_vxrm = requestVec_2_vxrm;
  wire [1:0]    requestVecFromSlot_2_other_bits_vSew = requestVec_2_vSew;
  wire [1:0]    requestVecFromSlot_2_divider_bits_vSew = requestVec_2_vSew;
  wire [1:0]    requestVecFromSlot_2_multiplier_bits_vSew = requestVec_2_vSew;
  wire [1:0]    requestVecFromSlot_2_shift_bits_vSew = requestVec_2_vSew;
  wire [1:0]    requestVecFromSlot_2_adder_bits_vSew = requestVec_2_vSew;
  wire [1:0]    requestVecFromSlot_2_logic_bits_vSew = requestVec_2_vSew;
  wire [19:0]   requestVecFromSlot_2_other_bits_shifterSize = requestVec_2_shifterSize;
  wire [19:0]   requestVecFromSlot_2_divider_bits_shifterSize = requestVec_2_shifterSize;
  wire [19:0]   requestVecFromSlot_2_multiplier_bits_shifterSize = requestVec_2_shifterSize;
  wire [19:0]   requestVecFromSlot_2_shift_bits_shifterSize = requestVec_2_shifterSize;
  wire [19:0]   requestVecFromSlot_2_adder_bits_shifterSize = requestVec_2_shifterSize;
  wire [19:0]   requestVecFromSlot_2_logic_bits_shifterSize = requestVec_2_shifterSize;
  wire          requestVecFromSlot_2_other_bits_rem = requestVec_2_rem;
  wire          requestVecFromSlot_2_divider_bits_rem = requestVec_2_rem;
  wire          requestVecFromSlot_2_multiplier_bits_rem = requestVec_2_rem;
  wire          requestVecFromSlot_2_shift_bits_rem = requestVec_2_rem;
  wire          requestVecFromSlot_2_adder_bits_rem = requestVec_2_rem;
  wire          requestVecFromSlot_2_logic_bits_rem = requestVec_2_rem;
  wire [9:0]    requestVecFromSlot_2_other_bits_groupIndex = requestVec_2_groupIndex;
  wire [9:0]    requestVecFromSlot_2_divider_bits_groupIndex = requestVec_2_groupIndex;
  wire [9:0]    requestVecFromSlot_2_multiplier_bits_groupIndex = requestVec_2_groupIndex;
  wire [9:0]    requestVecFromSlot_2_shift_bits_groupIndex = requestVec_2_groupIndex;
  wire [9:0]    requestVecFromSlot_2_adder_bits_groupIndex = requestVec_2_groupIndex;
  wire [9:0]    requestVecFromSlot_2_logic_bits_groupIndex = requestVec_2_groupIndex;
  wire [1:0]    requestVecFromSlot_2_other_bits_laneIndex = requestVec_2_laneIndex;
  wire [1:0]    requestVecFromSlot_2_divider_bits_laneIndex = requestVec_2_laneIndex;
  wire [1:0]    requestVecFromSlot_2_multiplier_bits_laneIndex = requestVec_2_laneIndex;
  wire [1:0]    requestVecFromSlot_2_shift_bits_laneIndex = requestVec_2_laneIndex;
  wire [1:0]    requestVecFromSlot_2_adder_bits_laneIndex = requestVec_2_laneIndex;
  wire [1:0]    requestVecFromSlot_2_logic_bits_laneIndex = requestVec_2_laneIndex;
  wire          requestVecFromSlot_2_other_bits_maskType = requestVec_2_maskType;
  wire          requestVecFromSlot_2_divider_bits_maskType = requestVec_2_maskType;
  wire          requestVecFromSlot_2_multiplier_bits_maskType = requestVec_2_maskType;
  wire          requestVecFromSlot_2_shift_bits_maskType = requestVec_2_maskType;
  wire          requestVecFromSlot_2_adder_bits_maskType = requestVec_2_maskType;
  wire          requestVecFromSlot_2_logic_bits_maskType = requestVec_2_maskType;
  wire          requestVecFromSlot_2_other_bits_narrow = requestVec_2_narrow;
  wire          requestVecFromSlot_2_divider_bits_narrow = requestVec_2_narrow;
  wire          requestVecFromSlot_2_multiplier_bits_narrow = requestVec_2_narrow;
  wire          requestVecFromSlot_2_shift_bits_narrow = requestVec_2_narrow;
  wire          requestVecFromSlot_2_adder_bits_narrow = requestVec_2_narrow;
  wire          requestVecFromSlot_2_logic_bits_narrow = requestVec_2_narrow;
  wire [32:0]   requestVecFromSlot_3_other_bits_src_0 = requestVec_3_src_0;
  wire [32:0]   requestVecFromSlot_3_divider_bits_src_0 = requestVec_3_src_0;
  wire [32:0]   requestVecFromSlot_3_multiplier_bits_src_0 = requestVec_3_src_0;
  wire [32:0]   requestVecFromSlot_3_shift_bits_src_0 = requestVec_3_src_0;
  wire [32:0]   requestVecFromSlot_3_adder_bits_src_0 = requestVec_3_src_0;
  wire [32:0]   requestVecFromSlot_3_logic_bits_src_0 = requestVec_3_src_0;
  wire [32:0]   requestVecFromSlot_3_other_bits_src_1 = requestVec_3_src_1;
  wire [32:0]   requestVecFromSlot_3_divider_bits_src_1 = requestVec_3_src_1;
  wire [32:0]   requestVecFromSlot_3_multiplier_bits_src_1 = requestVec_3_src_1;
  wire [32:0]   requestVecFromSlot_3_shift_bits_src_1 = requestVec_3_src_1;
  wire [32:0]   requestVecFromSlot_3_adder_bits_src_1 = requestVec_3_src_1;
  wire [32:0]   requestVecFromSlot_3_logic_bits_src_1 = requestVec_3_src_1;
  wire [32:0]   requestVecFromSlot_3_other_bits_src_2 = requestVec_3_src_2;
  wire [32:0]   requestVecFromSlot_3_divider_bits_src_2 = requestVec_3_src_2;
  wire [32:0]   requestVecFromSlot_3_multiplier_bits_src_2 = requestVec_3_src_2;
  wire [32:0]   requestVecFromSlot_3_shift_bits_src_2 = requestVec_3_src_2;
  wire [32:0]   requestVecFromSlot_3_adder_bits_src_2 = requestVec_3_src_2;
  wire [32:0]   requestVecFromSlot_3_logic_bits_src_2 = requestVec_3_src_2;
  wire [32:0]   requestVecFromSlot_3_other_bits_src_3 = requestVec_3_src_3;
  wire [32:0]   requestVecFromSlot_3_divider_bits_src_3 = requestVec_3_src_3;
  wire [32:0]   requestVecFromSlot_3_multiplier_bits_src_3 = requestVec_3_src_3;
  wire [32:0]   requestVecFromSlot_3_shift_bits_src_3 = requestVec_3_src_3;
  wire [32:0]   requestVecFromSlot_3_adder_bits_src_3 = requestVec_3_src_3;
  wire [32:0]   requestVecFromSlot_3_logic_bits_src_3 = requestVec_3_src_3;
  wire [3:0]    requestVecFromSlot_3_other_bits_opcode = requestVec_3_opcode;
  wire [3:0]    requestVecFromSlot_3_divider_bits_opcode = requestVec_3_opcode;
  wire [3:0]    requestVecFromSlot_3_multiplier_bits_opcode = requestVec_3_opcode;
  wire [3:0]    requestVecFromSlot_3_shift_bits_opcode = requestVec_3_opcode;
  wire [3:0]    requestVecFromSlot_3_adder_bits_opcode = requestVec_3_opcode;
  wire [3:0]    requestVecFromSlot_3_logic_bits_opcode = requestVec_3_opcode;
  wire [3:0]    requestVecFromSlot_3_other_bits_mask = requestVec_3_mask;
  wire [3:0]    requestVecFromSlot_3_divider_bits_mask = requestVec_3_mask;
  wire [3:0]    requestVecFromSlot_3_multiplier_bits_mask = requestVec_3_mask;
  wire [3:0]    requestVecFromSlot_3_shift_bits_mask = requestVec_3_mask;
  wire [3:0]    requestVecFromSlot_3_adder_bits_mask = requestVec_3_mask;
  wire [3:0]    requestVecFromSlot_3_logic_bits_mask = requestVec_3_mask;
  wire [3:0]    requestVecFromSlot_3_other_bits_executeMask = requestVec_3_executeMask;
  wire [3:0]    requestVecFromSlot_3_divider_bits_executeMask = requestVec_3_executeMask;
  wire [3:0]    requestVecFromSlot_3_multiplier_bits_executeMask = requestVec_3_executeMask;
  wire [3:0]    requestVecFromSlot_3_shift_bits_executeMask = requestVec_3_executeMask;
  wire [3:0]    requestVecFromSlot_3_adder_bits_executeMask = requestVec_3_executeMask;
  wire [3:0]    requestVecFromSlot_3_logic_bits_executeMask = requestVec_3_executeMask;
  wire          requestVecFromSlot_3_other_bits_sign0 = requestVec_3_sign0;
  wire          requestVecFromSlot_3_divider_bits_sign0 = requestVec_3_sign0;
  wire          requestVecFromSlot_3_multiplier_bits_sign0 = requestVec_3_sign0;
  wire          requestVecFromSlot_3_shift_bits_sign0 = requestVec_3_sign0;
  wire          requestVecFromSlot_3_adder_bits_sign0 = requestVec_3_sign0;
  wire          requestVecFromSlot_3_logic_bits_sign0 = requestVec_3_sign0;
  wire          requestVecFromSlot_3_other_bits_sign = requestVec_3_sign;
  wire          requestVecFromSlot_3_divider_bits_sign = requestVec_3_sign;
  wire          requestVecFromSlot_3_multiplier_bits_sign = requestVec_3_sign;
  wire          requestVecFromSlot_3_shift_bits_sign = requestVec_3_sign;
  wire          requestVecFromSlot_3_adder_bits_sign = requestVec_3_sign;
  wire          requestVecFromSlot_3_logic_bits_sign = requestVec_3_sign;
  wire          requestVecFromSlot_3_other_bits_reverse = requestVec_3_reverse;
  wire          requestVecFromSlot_3_divider_bits_reverse = requestVec_3_reverse;
  wire          requestVecFromSlot_3_multiplier_bits_reverse = requestVec_3_reverse;
  wire          requestVecFromSlot_3_shift_bits_reverse = requestVec_3_reverse;
  wire          requestVecFromSlot_3_adder_bits_reverse = requestVec_3_reverse;
  wire          requestVecFromSlot_3_logic_bits_reverse = requestVec_3_reverse;
  wire          requestVecFromSlot_3_other_bits_average = requestVec_3_average;
  wire          requestVecFromSlot_3_divider_bits_average = requestVec_3_average;
  wire          requestVecFromSlot_3_multiplier_bits_average = requestVec_3_average;
  wire          requestVecFromSlot_3_shift_bits_average = requestVec_3_average;
  wire          requestVecFromSlot_3_adder_bits_average = requestVec_3_average;
  wire          requestVecFromSlot_3_logic_bits_average = requestVec_3_average;
  wire          requestVecFromSlot_3_other_bits_saturate = requestVec_3_saturate;
  wire          requestVecFromSlot_3_divider_bits_saturate = requestVec_3_saturate;
  wire          requestVecFromSlot_3_multiplier_bits_saturate = requestVec_3_saturate;
  wire          requestVecFromSlot_3_shift_bits_saturate = requestVec_3_saturate;
  wire          requestVecFromSlot_3_adder_bits_saturate = requestVec_3_saturate;
  wire          requestVecFromSlot_3_logic_bits_saturate = requestVec_3_saturate;
  wire [1:0]    requestVecFromSlot_3_other_bits_vxrm = requestVec_3_vxrm;
  wire [1:0]    requestVecFromSlot_3_divider_bits_vxrm = requestVec_3_vxrm;
  wire [1:0]    requestVecFromSlot_3_multiplier_bits_vxrm = requestVec_3_vxrm;
  wire [1:0]    requestVecFromSlot_3_shift_bits_vxrm = requestVec_3_vxrm;
  wire [1:0]    requestVecFromSlot_3_adder_bits_vxrm = requestVec_3_vxrm;
  wire [1:0]    requestVecFromSlot_3_logic_bits_vxrm = requestVec_3_vxrm;
  wire [1:0]    requestVecFromSlot_3_other_bits_vSew = requestVec_3_vSew;
  wire [1:0]    requestVecFromSlot_3_divider_bits_vSew = requestVec_3_vSew;
  wire [1:0]    requestVecFromSlot_3_multiplier_bits_vSew = requestVec_3_vSew;
  wire [1:0]    requestVecFromSlot_3_shift_bits_vSew = requestVec_3_vSew;
  wire [1:0]    requestVecFromSlot_3_adder_bits_vSew = requestVec_3_vSew;
  wire [1:0]    requestVecFromSlot_3_logic_bits_vSew = requestVec_3_vSew;
  wire [19:0]   requestVecFromSlot_3_other_bits_shifterSize = requestVec_3_shifterSize;
  wire [19:0]   requestVecFromSlot_3_divider_bits_shifterSize = requestVec_3_shifterSize;
  wire [19:0]   requestVecFromSlot_3_multiplier_bits_shifterSize = requestVec_3_shifterSize;
  wire [19:0]   requestVecFromSlot_3_shift_bits_shifterSize = requestVec_3_shifterSize;
  wire [19:0]   requestVecFromSlot_3_adder_bits_shifterSize = requestVec_3_shifterSize;
  wire [19:0]   requestVecFromSlot_3_logic_bits_shifterSize = requestVec_3_shifterSize;
  wire          requestVecFromSlot_3_other_bits_rem = requestVec_3_rem;
  wire          requestVecFromSlot_3_divider_bits_rem = requestVec_3_rem;
  wire          requestVecFromSlot_3_multiplier_bits_rem = requestVec_3_rem;
  wire          requestVecFromSlot_3_shift_bits_rem = requestVec_3_rem;
  wire          requestVecFromSlot_3_adder_bits_rem = requestVec_3_rem;
  wire          requestVecFromSlot_3_logic_bits_rem = requestVec_3_rem;
  wire [9:0]    requestVecFromSlot_3_other_bits_groupIndex = requestVec_3_groupIndex;
  wire [9:0]    requestVecFromSlot_3_divider_bits_groupIndex = requestVec_3_groupIndex;
  wire [9:0]    requestVecFromSlot_3_multiplier_bits_groupIndex = requestVec_3_groupIndex;
  wire [9:0]    requestVecFromSlot_3_shift_bits_groupIndex = requestVec_3_groupIndex;
  wire [9:0]    requestVecFromSlot_3_adder_bits_groupIndex = requestVec_3_groupIndex;
  wire [9:0]    requestVecFromSlot_3_logic_bits_groupIndex = requestVec_3_groupIndex;
  wire [1:0]    requestVecFromSlot_3_other_bits_laneIndex = requestVec_3_laneIndex;
  wire [1:0]    requestVecFromSlot_3_divider_bits_laneIndex = requestVec_3_laneIndex;
  wire [1:0]    requestVecFromSlot_3_multiplier_bits_laneIndex = requestVec_3_laneIndex;
  wire [1:0]    requestVecFromSlot_3_shift_bits_laneIndex = requestVec_3_laneIndex;
  wire [1:0]    requestVecFromSlot_3_adder_bits_laneIndex = requestVec_3_laneIndex;
  wire [1:0]    requestVecFromSlot_3_logic_bits_laneIndex = requestVec_3_laneIndex;
  wire          requestVecFromSlot_3_other_bits_maskType = requestVec_3_maskType;
  wire          requestVecFromSlot_3_divider_bits_maskType = requestVec_3_maskType;
  wire          requestVecFromSlot_3_multiplier_bits_maskType = requestVec_3_maskType;
  wire          requestVecFromSlot_3_shift_bits_maskType = requestVec_3_maskType;
  wire          requestVecFromSlot_3_adder_bits_maskType = requestVec_3_maskType;
  wire          requestVecFromSlot_3_logic_bits_maskType = requestVec_3_maskType;
  wire          requestVecFromSlot_3_other_bits_narrow = requestVec_3_narrow;
  wire          requestVecFromSlot_3_divider_bits_narrow = requestVec_3_narrow;
  wire          requestVecFromSlot_3_multiplier_bits_narrow = requestVec_3_narrow;
  wire          requestVecFromSlot_3_shift_bits_narrow = requestVec_3_narrow;
  wire          requestVecFromSlot_3_adder_bits_narrow = requestVec_3_narrow;
  wire          requestVecFromSlot_3_logic_bits_narrow = requestVec_3_narrow;
  wire [31:0]   selectResponse_bits_data;
  wire [1:0]    selectResponse_bits_executeIndex;
  wire          selectResponse_bits_ffoSuccess;
  wire [3:0]    selectResponse_bits_adderMaskResp;
  wire [3:0]    selectResponse_bits_vxsat;
  wire [1:0]    selectResponse_bits_tag;
  wire [31:0]   selectResponse_1_bits_data;
  wire [1:0]    selectResponse_1_bits_executeIndex;
  wire          selectResponse_1_bits_ffoSuccess;
  wire [3:0]    selectResponse_1_bits_adderMaskResp;
  wire [3:0]    selectResponse_1_bits_vxsat;
  wire [1:0]    selectResponse_1_bits_tag;
  wire [31:0]   selectResponse_2_bits_data;
  wire [1:0]    selectResponse_2_bits_executeIndex;
  wire          selectResponse_2_bits_ffoSuccess;
  wire [3:0]    selectResponse_2_bits_adderMaskResp;
  wire [3:0]    selectResponse_2_bits_vxsat;
  wire [1:0]    selectResponse_2_bits_tag;
  wire [31:0]   selectResponse_3_bits_data;
  wire [1:0]    selectResponse_3_bits_executeIndex;
  wire          selectResponse_3_bits_ffoSuccess;
  wire [3:0]    selectResponse_3_bits_adderMaskResp;
  wire [3:0]    selectResponse_3_bits_vxsat;
  wire [1:0]    selectResponse_3_bits_tag;
  wire          requestFire;
  wire          requestFire_1;
  wire          requestFire_2;
  wire          requestFire_3;
  wire          slotEnqueueFire_0;
  reg  [7:0]    instructionValidNext;
  reg  [7:0]    vxsatResult;
  wire          enqReady_5;
  wire          crossLaneWriteQueue_0_deq_valid;
  assign crossLaneWriteQueue_0_deq_valid = ~_crossLaneWriteQueue_fifo_empty;
  wire [4:0]    crossLaneWriteQueue_dataOut_vd;
  wire [5:0]    crossLaneWriteQueue_dataOut_offset;
  wire [3:0]    crossLaneWriteQueue_dataOut_mask;
  wire [31:0]   crossLaneWriteQueue_dataOut_data;
  wire          crossLaneWriteQueue_dataOut_last;
  wire [2:0]    crossLaneWriteQueue_dataOut_instructionIndex;
  wire [32:0]   crossLaneWriteQueue_dataIn_lo_hi = {crossLaneWriteQueue_0_enq_bits_data, 1'h0};
  wire [35:0]   crossLaneWriteQueue_dataIn_lo = {crossLaneWriteQueue_dataIn_lo_hi, crossLaneWriteQueue_0_enq_bits_instructionIndex};
  wire [4:0]    crossLaneWriteQueue_0_enq_bits_vd;
  wire [5:0]    crossLaneWriteQueue_0_enq_bits_offset;
  wire [10:0]   crossLaneWriteQueue_dataIn_hi_hi = {crossLaneWriteQueue_0_enq_bits_vd, crossLaneWriteQueue_0_enq_bits_offset};
  wire [3:0]    crossLaneWriteQueue_0_enq_bits_mask;
  wire [14:0]   crossLaneWriteQueue_dataIn_hi = {crossLaneWriteQueue_dataIn_hi_hi, crossLaneWriteQueue_0_enq_bits_mask};
  wire [50:0]   crossLaneWriteQueue_dataIn = {crossLaneWriteQueue_dataIn_hi, crossLaneWriteQueue_dataIn_lo};
  assign crossLaneWriteQueue_dataOut_instructionIndex = _crossLaneWriteQueue_fifo_data_out[2:0];
  assign crossLaneWriteQueue_dataOut_last = _crossLaneWriteQueue_fifo_data_out[3];
  assign crossLaneWriteQueue_dataOut_data = _crossLaneWriteQueue_fifo_data_out[35:4];
  assign crossLaneWriteQueue_dataOut_mask = _crossLaneWriteQueue_fifo_data_out[39:36];
  assign crossLaneWriteQueue_dataOut_offset = _crossLaneWriteQueue_fifo_data_out[45:40];
  assign crossLaneWriteQueue_dataOut_vd = _crossLaneWriteQueue_fifo_data_out[50:46];
  wire [4:0]    crossLaneWriteQueue_0_deq_bits_vd = crossLaneWriteQueue_dataOut_vd;
  wire [5:0]    crossLaneWriteQueue_0_deq_bits_offset = crossLaneWriteQueue_dataOut_offset;
  wire [3:0]    crossLaneWriteQueue_0_deq_bits_mask = crossLaneWriteQueue_dataOut_mask;
  wire [31:0]   crossLaneWriteQueue_0_deq_bits_data = crossLaneWriteQueue_dataOut_data;
  wire          crossLaneWriteQueue_0_deq_bits_last = crossLaneWriteQueue_dataOut_last;
  wire [2:0]    crossLaneWriteQueue_0_deq_bits_instructionIndex = crossLaneWriteQueue_dataOut_instructionIndex;
  wire          crossLaneWriteQueue_0_deq_ready;
  wire          crossLaneWriteQueue_0_enq_ready = ~_crossLaneWriteQueue_fifo_full | crossLaneWriteQueue_0_deq_ready;
  wire          enqReady_6;
  wire          crossLaneWriteQueue_1_deq_valid;
  assign crossLaneWriteQueue_1_deq_valid = ~_crossLaneWriteQueue_fifo_1_empty;
  wire [4:0]    crossLaneWriteQueue_dataOut_1_vd;
  wire [5:0]    crossLaneWriteQueue_dataOut_1_offset;
  wire [3:0]    crossLaneWriteQueue_dataOut_1_mask;
  wire [31:0]   crossLaneWriteQueue_dataOut_1_data;
  wire          crossLaneWriteQueue_dataOut_1_last;
  wire [2:0]    crossLaneWriteQueue_dataOut_1_instructionIndex;
  wire [32:0]   crossLaneWriteQueue_dataIn_lo_hi_1 = {crossLaneWriteQueue_1_enq_bits_data, 1'h0};
  wire [35:0]   crossLaneWriteQueue_dataIn_lo_1 = {crossLaneWriteQueue_dataIn_lo_hi_1, crossLaneWriteQueue_1_enq_bits_instructionIndex};
  wire [4:0]    crossLaneWriteQueue_1_enq_bits_vd;
  wire [5:0]    crossLaneWriteQueue_1_enq_bits_offset;
  wire [10:0]   crossLaneWriteQueue_dataIn_hi_hi_1 = {crossLaneWriteQueue_1_enq_bits_vd, crossLaneWriteQueue_1_enq_bits_offset};
  wire [3:0]    crossLaneWriteQueue_1_enq_bits_mask;
  wire [14:0]   crossLaneWriteQueue_dataIn_hi_1 = {crossLaneWriteQueue_dataIn_hi_hi_1, crossLaneWriteQueue_1_enq_bits_mask};
  wire [50:0]   crossLaneWriteQueue_dataIn_1 = {crossLaneWriteQueue_dataIn_hi_1, crossLaneWriteQueue_dataIn_lo_1};
  assign crossLaneWriteQueue_dataOut_1_instructionIndex = _crossLaneWriteQueue_fifo_1_data_out[2:0];
  assign crossLaneWriteQueue_dataOut_1_last = _crossLaneWriteQueue_fifo_1_data_out[3];
  assign crossLaneWriteQueue_dataOut_1_data = _crossLaneWriteQueue_fifo_1_data_out[35:4];
  assign crossLaneWriteQueue_dataOut_1_mask = _crossLaneWriteQueue_fifo_1_data_out[39:36];
  assign crossLaneWriteQueue_dataOut_1_offset = _crossLaneWriteQueue_fifo_1_data_out[45:40];
  assign crossLaneWriteQueue_dataOut_1_vd = _crossLaneWriteQueue_fifo_1_data_out[50:46];
  wire [4:0]    crossLaneWriteQueue_1_deq_bits_vd = crossLaneWriteQueue_dataOut_1_vd;
  wire [5:0]    crossLaneWriteQueue_1_deq_bits_offset = crossLaneWriteQueue_dataOut_1_offset;
  wire [3:0]    crossLaneWriteQueue_1_deq_bits_mask = crossLaneWriteQueue_dataOut_1_mask;
  wire [31:0]   crossLaneWriteQueue_1_deq_bits_data = crossLaneWriteQueue_dataOut_1_data;
  wire          crossLaneWriteQueue_1_deq_bits_last = crossLaneWriteQueue_dataOut_1_last;
  wire [2:0]    crossLaneWriteQueue_1_deq_bits_instructionIndex = crossLaneWriteQueue_dataOut_1_instructionIndex;
  wire          crossLaneWriteQueue_1_deq_ready;
  wire          crossLaneWriteQueue_1_enq_ready = ~_crossLaneWriteQueue_fifo_1_full | crossLaneWriteQueue_1_deq_ready;
  wire          _probeWire_slots_0_decodeResultIsCrossReadOrWrite_T_3 = slotControl_0_laneRequest_decodeResult_crossRead | slotControl_0_laneRequest_decodeResult_crossWrite;
  wire          alwaysNextGroup = _probeWire_slots_0_decodeResultIsCrossReadOrWrite_T_3 | slotControl_0_laneRequest_decodeResult_nr | ~slotControl_0_laneRequest_decodeResult_scheduler | slotControl_0_laneRequest_loadStore;
  wire          _GEN = slotControl_0_laneRequest_decodeResult_maskSource | slotControl_0_laneRequest_decodeResult_maskLogic;
  wire          maskNotMaskedElement = ~slotControl_0_laneRequest_mask | _GEN;
  wire [3:0]    _vSew1H_T = 4'h1 << slotControl_0_laneRequest_csrInterface_vSew;
  wire [2:0]    vSew1H = _vSew1H_T[2:0];
  wire [2:0]    laneState_vSew1H = vSew1H;
  wire          skipEnable = slotControl_0_laneRequest_mask & ~slotControl_0_laneRequest_decodeResult_maskSource & ~slotControl_0_laneRequest_decodeResult_maskLogic & ~alwaysNextGroup;
  wire          laneState_skipEnable = skipEnable;
  wire          laneState_maskNotMaskedElement = ~slotControl_0_laneRequest_mask | _GEN;
  wire          laneState_skipRead = slotControl_0_laneRequest_decodeResult_other & slotControl_0_laneRequest_decodeResult_uop == 4'h9;
  wire          stage0_enqueue_valid = slotActive_0 & (slotControl_0_mask_valid | ~slotControl_0_laneRequest_mask);
  wire          _maskFailure_T = _stage0_enqueue_ready & stage0_enqueue_valid;
  assign maskControlRelease_0_valid = _maskFailure_T & _stage0_updateLaneState_outOfExecutionRange;
  wire          slotMaskRequestVec_0_valid = slotControl_0_laneRequest_mask & slotOccupied_0 & (_maskFailure_T & _stage0_updateLaneState_maskExhausted | ~slotControl_0_mask_valid);
  wire          maskRequestFireOH_0;
  wire          maskUpdateFire = slotMaskRequestVec_0_valid & maskRequestFireOH_0;
  wire          maskFailure = _stage0_updateLaneState_maskExhausted & _maskFailure_T;
  wire [3:0]    instructionIndex1H = 4'h1 << slotControl_0_laneRequest_instructionIndex[1:0];
  wire [3:0]    instructionUnrelatedMaskUnitVec_0 = slotControl_0_laneRequest_decodeResult_maskUnit & slotControl_0_laneRequest_decodeResult_readOnly ? 4'h0 : instructionIndex1H;
  reg  [2:0]    tokenReg;
  wire          tokenReady = tokenReg != 3'h4;
  wire          readBusPort_0_deq_valid_0 = _stage1_readBusRequest_0_valid & tokenReady;
  wire [2:0]    tokenUpdate = readBusPort_0_deq_valid_0 ? 3'h1 : 3'h7;
  wire          queue_deq_valid;
  assign queue_deq_valid = ~_queue_fifo_empty;
  wire [31:0]   queue_dataOut_data;
  wire [31:0]   queue_deq_bits_data = queue_dataOut_data;
  wire          queue_deq_ready;
  wire          queue_enq_ready = ~_queue_fifo_full | queue_deq_ready;
  wire          readBusPort_0_enqRelease_0 = queue_deq_ready & queue_deq_valid;
  reg  [2:0]    tokenReg_1;
  wire          tokenReady_1 = tokenReg_1 != 3'h4;
  wire          readBusPort_1_deq_valid_0 = _stage1_readBusRequest_1_valid & tokenReady_1;
  wire [2:0]    tokenUpdate_1 = readBusPort_1_deq_valid_0 ? 3'h1 : 3'h7;
  wire          queue_1_deq_valid;
  assign queue_1_deq_valid = ~_queue_fifo_1_empty;
  wire [31:0]   queue_dataOut_1_data;
  wire [31:0]   queue_1_deq_bits_data = queue_dataOut_1_data;
  wire          queue_1_deq_ready;
  wire          queue_1_enq_ready = ~_queue_fifo_1_full | queue_1_deq_ready;
  wire          readBusPort_1_enqRelease_0 = queue_1_deq_ready & queue_1_deq_valid;
  reg  [2:0]    tokenReg_2;
  wire          tokenReady_2 = tokenReg_2 != 3'h4;
  wire          writeBusPort_0_deq_valid_0 = _stage3_crossWritePort_0_valid & tokenReady_2;
  wire [2:0]    tokenUpdate_2 = writeBusPort_0_deq_valid_0 ? 3'h1 : 3'h7;
  reg  [2:0]    tokenReg_3;
  wire          tokenReady_3 = tokenReg_3 != 3'h4;
  wire          writeBusPort_1_deq_valid_0 = _stage3_crossWritePort_1_valid & tokenReady_3;
  wire [2:0]    tokenUpdate_3 = writeBusPort_1_deq_valid_0 ? 3'h1 : 3'h7;
  wire [3:0]    responseVec_0_bits_vxsat;
  wire          responseVec_0_valid;
  wire [7:0]    vxsatEnq_0 = responseVec_0_valid & (|responseVec_0_bits_vxsat) ? 8'h1 << _executionUnit_responseIndex : 8'h0;
  wire          stage3EnqWire_ready;
  wire          _probeWire_slots_1_decodeResultIsCrossReadOrWrite_T_3 = slotControl_1_laneRequest_decodeResult_crossRead | slotControl_1_laneRequest_decodeResult_crossWrite;
  wire          alwaysNextGroup_1 = _probeWire_slots_1_decodeResultIsCrossReadOrWrite_T_3 | slotControl_1_laneRequest_decodeResult_nr | ~slotControl_1_laneRequest_decodeResult_scheduler | slotControl_1_laneRequest_loadStore;
  wire          _GEN_0 = slotControl_1_laneRequest_decodeResult_maskSource | slotControl_1_laneRequest_decodeResult_maskLogic;
  wire          maskNotMaskedElement_1 = ~slotControl_1_laneRequest_mask | _GEN_0;
  wire [3:0]    _vSew1H_T_1 = 4'h1 << slotControl_1_laneRequest_csrInterface_vSew;
  wire [2:0]    vSew1H_1 = _vSew1H_T_1[2:0];
  wire [2:0]    laneState_1_vSew1H = vSew1H_1;
  wire          skipEnable_1 = slotControl_1_laneRequest_mask & ~slotControl_1_laneRequest_decodeResult_maskSource & ~slotControl_1_laneRequest_decodeResult_maskLogic & ~alwaysNextGroup_1;
  wire          laneState_1_skipEnable = skipEnable_1;
  wire          slotActive_1 = slotOccupied_1 & ~slotShiftValid_1 & ~(_probeWire_slots_1_decodeResultIsCrossReadOrWrite_T_3 | slotControl_1_laneRequest_decodeResult_widenReduce) & slotControl_1_laneRequest_decodeResult_scheduler;
  wire          laneState_1_maskNotMaskedElement = ~slotControl_1_laneRequest_mask | _GEN_0;
  wire          laneState_1_skipRead = slotControl_1_laneRequest_decodeResult_other & slotControl_1_laneRequest_decodeResult_uop == 4'h9;
  wire          stage0_1_enqueue_valid = slotActive_1 & (slotControl_1_mask_valid | ~slotControl_1_laneRequest_mask);
  wire          _maskFailure_T_1 = _stage0_1_enqueue_ready & stage0_1_enqueue_valid;
  assign maskControlRelease_1_valid = _maskFailure_T_1 & _stage0_1_updateLaneState_outOfExecutionRange;
  wire          slotMaskRequestVec_1_valid = slotControl_1_laneRequest_mask & slotOccupied_1 & (_maskFailure_T_1 & _stage0_1_updateLaneState_maskExhausted | ~slotControl_1_mask_valid);
  wire          maskRequestFireOH_1;
  wire          maskUpdateFire_1 = slotMaskRequestVec_1_valid & maskRequestFireOH_1;
  wire          maskFailure_1 = _stage0_1_updateLaneState_maskExhausted & _maskFailure_T_1;
  wire [3:0]    instructionIndex1H_1 = 4'h1 << slotControl_1_laneRequest_instructionIndex[1:0];
  wire [3:0]    instructionUnrelatedMaskUnitVec_1 = slotControl_1_laneRequest_decodeResult_maskUnit & slotControl_1_laneRequest_decodeResult_readOnly ? 4'h0 : instructionIndex1H_1;
  wire [3:0]    responseVec_1_bits_vxsat;
  wire          responseVec_1_valid;
  wire [7:0]    vxsatEnq_1 = responseVec_1_valid & (|responseVec_1_bits_vxsat) ? 8'h1 << _executionUnit_1_responseIndex : 8'h0;
  wire          stage3EnqWire_1_ready;
  wire          _probeWire_slots_2_decodeResultIsCrossReadOrWrite_T_3 = slotControl_2_laneRequest_decodeResult_crossRead | slotControl_2_laneRequest_decodeResult_crossWrite;
  wire          alwaysNextGroup_2 = _probeWire_slots_2_decodeResultIsCrossReadOrWrite_T_3 | slotControl_2_laneRequest_decodeResult_nr | ~slotControl_2_laneRequest_decodeResult_scheduler | slotControl_2_laneRequest_loadStore;
  wire          _GEN_1 = slotControl_2_laneRequest_decodeResult_maskSource | slotControl_2_laneRequest_decodeResult_maskLogic;
  wire          maskNotMaskedElement_2 = ~slotControl_2_laneRequest_mask | _GEN_1;
  wire [3:0]    _vSew1H_T_2 = 4'h1 << slotControl_2_laneRequest_csrInterface_vSew;
  wire [2:0]    vSew1H_2 = _vSew1H_T_2[2:0];
  wire [2:0]    laneState_2_vSew1H = vSew1H_2;
  wire          skipEnable_2 = slotControl_2_laneRequest_mask & ~slotControl_2_laneRequest_decodeResult_maskSource & ~slotControl_2_laneRequest_decodeResult_maskLogic & ~alwaysNextGroup_2;
  wire          laneState_2_skipEnable = skipEnable_2;
  wire          slotActive_2 = slotOccupied_2 & ~slotShiftValid_2 & ~(_probeWire_slots_2_decodeResultIsCrossReadOrWrite_T_3 | slotControl_2_laneRequest_decodeResult_widenReduce) & slotControl_2_laneRequest_decodeResult_scheduler;
  wire          laneState_2_maskNotMaskedElement = ~slotControl_2_laneRequest_mask | _GEN_1;
  wire          laneState_2_skipRead = slotControl_2_laneRequest_decodeResult_other & slotControl_2_laneRequest_decodeResult_uop == 4'h9;
  wire          stage0_2_enqueue_valid = slotActive_2 & (slotControl_2_mask_valid | ~slotControl_2_laneRequest_mask);
  wire          _maskFailure_T_2 = _stage0_2_enqueue_ready & stage0_2_enqueue_valid;
  assign maskControlRelease_2_valid = _maskFailure_T_2 & _stage0_2_updateLaneState_outOfExecutionRange;
  wire          slotMaskRequestVec_2_valid = slotControl_2_laneRequest_mask & slotOccupied_2 & (_maskFailure_T_2 & _stage0_2_updateLaneState_maskExhausted | ~slotControl_2_mask_valid);
  wire          maskRequestFireOH_2;
  wire          maskUpdateFire_2 = slotMaskRequestVec_2_valid & maskRequestFireOH_2;
  wire          maskFailure_2 = _stage0_2_updateLaneState_maskExhausted & _maskFailure_T_2;
  wire [3:0]    instructionIndex1H_2 = 4'h1 << slotControl_2_laneRequest_instructionIndex[1:0];
  wire [3:0]    instructionUnrelatedMaskUnitVec_2 = slotControl_2_laneRequest_decodeResult_maskUnit & slotControl_2_laneRequest_decodeResult_readOnly ? 4'h0 : instructionIndex1H_2;
  wire [3:0]    responseVec_2_bits_vxsat;
  wire          responseVec_2_valid;
  wire [7:0]    vxsatEnq_2 = responseVec_2_valid & (|responseVec_2_bits_vxsat) ? 8'h1 << _executionUnit_2_responseIndex : 8'h0;
  wire          stage3EnqWire_2_ready;
  wire          _probeWire_slots_3_decodeResultIsCrossReadOrWrite_T_3 = slotControl_3_laneRequest_decodeResult_crossRead | slotControl_3_laneRequest_decodeResult_crossWrite;
  wire          alwaysNextGroup_3 = _probeWire_slots_3_decodeResultIsCrossReadOrWrite_T_3 | slotControl_3_laneRequest_decodeResult_nr | ~slotControl_3_laneRequest_decodeResult_scheduler | slotControl_3_laneRequest_loadStore;
  wire          _GEN_2 = slotControl_3_laneRequest_decodeResult_maskSource | slotControl_3_laneRequest_decodeResult_maskLogic;
  wire          maskNotMaskedElement_3 = ~slotControl_3_laneRequest_mask | _GEN_2;
  wire [3:0]    _vSew1H_T_3 = 4'h1 << slotControl_3_laneRequest_csrInterface_vSew;
  wire [2:0]    vSew1H_3 = _vSew1H_T_3[2:0];
  wire [2:0]    laneState_3_vSew1H = vSew1H_3;
  wire          skipEnable_3 = slotControl_3_laneRequest_mask & ~slotControl_3_laneRequest_decodeResult_maskSource & ~slotControl_3_laneRequest_decodeResult_maskLogic & ~alwaysNextGroup_3;
  wire          laneState_3_skipEnable = skipEnable_3;
  wire          slotActive_3 = slotOccupied_3 & ~slotShiftValid_3 & ~(_probeWire_slots_3_decodeResultIsCrossReadOrWrite_T_3 | slotControl_3_laneRequest_decodeResult_widenReduce) & slotControl_3_laneRequest_decodeResult_scheduler;
  wire          laneState_3_maskNotMaskedElement = ~slotControl_3_laneRequest_mask | _GEN_2;
  wire          laneState_3_skipRead = slotControl_3_laneRequest_decodeResult_other & slotControl_3_laneRequest_decodeResult_uop == 4'h9;
  wire          stage0_3_enqueue_valid = slotActive_3 & (slotControl_3_mask_valid | ~slotControl_3_laneRequest_mask);
  wire          _maskFailure_T_3 = _stage0_3_enqueue_ready & stage0_3_enqueue_valid;
  assign maskControlRelease_3_valid = _maskFailure_T_3 & _stage0_3_updateLaneState_outOfExecutionRange;
  wire          slotMaskRequestVec_3_valid = slotControl_3_laneRequest_mask & slotOccupied_3 & (_maskFailure_T_3 & _stage0_3_updateLaneState_maskExhausted | ~slotControl_3_mask_valid);
  wire          maskRequestFireOH_3;
  wire          maskUpdateFire_3 = slotMaskRequestVec_3_valid & maskRequestFireOH_3;
  wire          maskFailure_3 = _stage0_3_updateLaneState_maskExhausted & _maskFailure_T_3;
  wire [3:0]    instructionIndex1H_3 = 4'h1 << slotControl_3_laneRequest_instructionIndex[1:0];
  wire [3:0]    instructionUnrelatedMaskUnitVec_3 = slotControl_3_laneRequest_decodeResult_maskUnit & slotControl_3_laneRequest_decodeResult_readOnly ? 4'h0 : instructionIndex1H_3;
  wire [3:0]    responseVec_3_bits_vxsat;
  wire          responseVec_3_valid;
  wire [7:0]    vxsatEnq_3 = responseVec_3_valid & (|responseVec_3_bits_vxsat) ? 8'h1 << _executionUnit_3_responseIndex : 8'h0;
  wire          stage3EnqWire_3_ready;
  wire [10:0]   _GEN_3 = {slotControl_0_laneRequest_vd, 6'h0};
  wire [10:0]   baseIndex;
  assign baseIndex = _GEN_3;
  wire [10:0]   baseIndex_1;
  assign baseIndex_1 = _GEN_3;
  wire [9:0]    indexGrowth = {writeBusPort_0_enq_bits_counter_0[8:0], 1'h0};
  wire [10:0]   finalIndex = baseIndex + {1'h0, indexGrowth};
  assign crossLaneWriteQueue_0_enq_bits_vd = finalIndex[10:6];
  assign crossLaneWriteQueue_0_enq_bits_offset = finalIndex[5:0];
  assign crossLaneWriteQueue_0_enq_bits_mask = {{2{writeBusPort_0_enq_bits_mask_0[1]}}, {2{writeBusPort_0_enq_bits_mask_0[0]}}};
  wire          writeBusPort_0_enqRelease_0 = crossLaneWriteQueue_0_deq_ready & crossLaneWriteQueue_0_deq_valid;
  wire [9:0]    indexGrowth_1 = {writeBusPort_1_enq_bits_counter_0[8:0], 1'h1};
  wire [10:0]   finalIndex_1 = baseIndex_1 + {1'h0, indexGrowth_1};
  assign crossLaneWriteQueue_1_enq_bits_vd = finalIndex_1[10:6];
  assign crossLaneWriteQueue_1_enq_bits_offset = finalIndex_1[5:0];
  assign crossLaneWriteQueue_1_enq_bits_mask = {{2{writeBusPort_1_enq_bits_mask_0[1]}}, {2{writeBusPort_1_enq_bits_mask_0[0]}}};
  wire          writeBusPort_1_enqRelease_0 = crossLaneWriteQueue_1_deq_ready & crossLaneWriteQueue_1_deq_valid;
  wire          executeEnqueueValid_0;
  wire          executeDecodeVec_0_logic;
  wire          requestVecFromSlot_0_logic_ready;
  wire          requestVecFromSlot_0_logic_valid = executeEnqueueValid_0 & executeDecodeVec_0_logic;
  wire          executeDecodeVec_0_adder;
  wire          requestVecFromSlot_0_adder_ready;
  wire          requestVecFromSlot_0_adder_valid = executeEnqueueValid_0 & executeDecodeVec_0_adder;
  wire          executeDecodeVec_0_shift;
  wire          requestVecFromSlot_0_shift_ready;
  wire          requestVecFromSlot_0_shift_valid = executeEnqueueValid_0 & executeDecodeVec_0_shift;
  wire          executeDecodeVec_0_multiplier;
  wire          requestVecFromSlot_0_multiplier_ready;
  wire          requestVecFromSlot_0_multiplier_valid = executeEnqueueValid_0 & executeDecodeVec_0_multiplier;
  wire          executeDecodeVec_0_divider;
  wire          requestVecFromSlot_0_divider_ready;
  wire          requestVecFromSlot_0_divider_valid = executeEnqueueValid_0 & executeDecodeVec_0_divider;
  wire          executeDecodeVec_0_other;
  wire          requestVecFromSlot_0_other_ready;
  wire          requestVecFromSlot_0_other_valid = executeEnqueueValid_0 & executeDecodeVec_0_other;
  assign requestFire =
    requestVecFromSlot_0_logic_ready & requestVecFromSlot_0_logic_valid | requestVecFromSlot_0_adder_ready & requestVecFromSlot_0_adder_valid | requestVecFromSlot_0_shift_ready & requestVecFromSlot_0_shift_valid
    | requestVecFromSlot_0_multiplier_ready & requestVecFromSlot_0_multiplier_valid | requestVecFromSlot_0_divider_ready & requestVecFromSlot_0_divider_valid | requestVecFromSlot_0_other_ready & requestVecFromSlot_0_other_valid;
  wire          executeEnqueueValid_1;
  wire          executeDecodeVec_1_logic;
  wire          executeEnqueueFire_0 = requestFire;
  wire          requestVecFromSlot_1_logic_ready;
  wire          requestVecFromSlot_1_logic_valid = executeEnqueueValid_1 & executeDecodeVec_1_logic;
  wire          executeDecodeVec_1_adder;
  wire          requestVecFromSlot_1_adder_ready;
  wire          requestVecFromSlot_1_adder_valid = executeEnqueueValid_1 & executeDecodeVec_1_adder;
  wire          executeDecodeVec_1_shift;
  wire          requestVecFromSlot_1_shift_ready;
  wire          requestVecFromSlot_1_shift_valid = executeEnqueueValid_1 & executeDecodeVec_1_shift;
  wire          executeDecodeVec_1_multiplier;
  wire          requestVecFromSlot_1_multiplier_ready;
  wire          requestVecFromSlot_1_multiplier_valid = executeEnqueueValid_1 & executeDecodeVec_1_multiplier;
  wire          executeDecodeVec_1_divider;
  wire          requestVecFromSlot_1_divider_ready;
  wire          requestVecFromSlot_1_divider_valid = executeEnqueueValid_1 & executeDecodeVec_1_divider;
  wire          executeDecodeVec_1_other;
  wire          requestVecFromSlot_1_other_ready;
  wire          requestVecFromSlot_1_other_valid = executeEnqueueValid_1 & executeDecodeVec_1_other;
  assign requestFire_1 =
    requestVecFromSlot_1_logic_ready & requestVecFromSlot_1_logic_valid | requestVecFromSlot_1_adder_ready & requestVecFromSlot_1_adder_valid | requestVecFromSlot_1_shift_ready & requestVecFromSlot_1_shift_valid
    | requestVecFromSlot_1_multiplier_ready & requestVecFromSlot_1_multiplier_valid | requestVecFromSlot_1_divider_ready & requestVecFromSlot_1_divider_valid | requestVecFromSlot_1_other_ready & requestVecFromSlot_1_other_valid;
  wire          executeEnqueueValid_2;
  wire          executeDecodeVec_2_logic;
  wire          executeEnqueueFire_1 = requestFire_1;
  wire          requestVecFromSlot_2_logic_ready;
  wire          requestVecFromSlot_2_logic_valid = executeEnqueueValid_2 & executeDecodeVec_2_logic;
  wire          executeDecodeVec_2_adder;
  wire          requestVecFromSlot_2_adder_ready;
  wire          requestVecFromSlot_2_adder_valid = executeEnqueueValid_2 & executeDecodeVec_2_adder;
  wire          executeDecodeVec_2_shift;
  wire          requestVecFromSlot_2_shift_ready;
  wire          requestVecFromSlot_2_shift_valid = executeEnqueueValid_2 & executeDecodeVec_2_shift;
  wire          executeDecodeVec_2_multiplier;
  wire          requestVecFromSlot_2_multiplier_ready;
  wire          requestVecFromSlot_2_multiplier_valid = executeEnqueueValid_2 & executeDecodeVec_2_multiplier;
  wire          executeDecodeVec_2_divider;
  wire          requestVecFromSlot_2_divider_ready;
  wire          requestVecFromSlot_2_divider_valid = executeEnqueueValid_2 & executeDecodeVec_2_divider;
  wire          executeDecodeVec_2_other;
  wire          requestVecFromSlot_2_other_ready;
  wire          requestVecFromSlot_2_other_valid = executeEnqueueValid_2 & executeDecodeVec_2_other;
  assign requestFire_2 =
    requestVecFromSlot_2_logic_ready & requestVecFromSlot_2_logic_valid | requestVecFromSlot_2_adder_ready & requestVecFromSlot_2_adder_valid | requestVecFromSlot_2_shift_ready & requestVecFromSlot_2_shift_valid
    | requestVecFromSlot_2_multiplier_ready & requestVecFromSlot_2_multiplier_valid | requestVecFromSlot_2_divider_ready & requestVecFromSlot_2_divider_valid | requestVecFromSlot_2_other_ready & requestVecFromSlot_2_other_valid;
  wire          executeEnqueueValid_3;
  wire          executeDecodeVec_3_logic;
  wire          executeEnqueueFire_2 = requestFire_2;
  wire          requestVecFromSlot_3_logic_ready;
  wire          requestVecFromSlot_3_logic_valid = executeEnqueueValid_3 & executeDecodeVec_3_logic;
  wire          executeDecodeVec_3_adder;
  wire          requestVecFromSlot_3_adder_ready;
  wire          requestVecFromSlot_3_adder_valid = executeEnqueueValid_3 & executeDecodeVec_3_adder;
  wire          executeDecodeVec_3_shift;
  wire          requestVecFromSlot_3_shift_ready;
  wire          requestVecFromSlot_3_shift_valid = executeEnqueueValid_3 & executeDecodeVec_3_shift;
  wire          executeDecodeVec_3_multiplier;
  wire          requestVecFromSlot_3_multiplier_ready;
  wire          requestVecFromSlot_3_multiplier_valid = executeEnqueueValid_3 & executeDecodeVec_3_multiplier;
  wire          executeDecodeVec_3_divider;
  wire          requestVecFromSlot_3_divider_ready;
  wire          requestVecFromSlot_3_divider_valid = executeEnqueueValid_3 & executeDecodeVec_3_divider;
  wire          executeDecodeVec_3_other;
  wire          requestVecFromSlot_3_other_ready;
  wire          requestVecFromSlot_3_other_valid = executeEnqueueValid_3 & executeDecodeVec_3_other;
  assign requestFire_3 =
    requestVecFromSlot_3_logic_ready & requestVecFromSlot_3_logic_valid | requestVecFromSlot_3_adder_ready & requestVecFromSlot_3_adder_valid | requestVecFromSlot_3_shift_ready & requestVecFromSlot_3_shift_valid
    | requestVecFromSlot_3_multiplier_ready & requestVecFromSlot_3_multiplier_valid | requestVecFromSlot_3_divider_ready & requestVecFromSlot_3_divider_valid | requestVecFromSlot_3_other_ready & requestVecFromSlot_3_other_valid;
  wire          executeEnqueueFire_3 = requestFire_3;
  wire          vrfIsBusy_4;
  wire [1:0]    _GEN_4 = {1'h0, vrfIsBusy_4};
  wire [1:0]    vfuResponse_VFUNotClear_hi_hi;
  assign vfuResponse_VFUNotClear_hi_hi = _GEN_4;
  wire [1:0]    vfuResponse_VFUNotClear_hi_hi_1;
  assign vfuResponse_VFUNotClear_hi_hi_1 = _GEN_4;
  wire [1:0]    vfuResponse_VFUNotClear_hi_hi_2;
  assign vfuResponse_VFUNotClear_hi_hi_2 = _GEN_4;
  wire [1:0]    vfuResponse_VFUNotClear_hi_hi_3;
  assign vfuResponse_VFUNotClear_hi_hi_3 = _GEN_4;
  wire [1:0]    vfuResponse_VFUNotClear_hi_hi_4;
  assign vfuResponse_VFUNotClear_hi_hi_4 = _GEN_4;
  wire [1:0]    vfuResponse_VFUNotClear_hi_hi_5;
  assign vfuResponse_VFUNotClear_hi_hi_5 = _GEN_4;
  wire [2:0]    vfuResponse_VFUNotClear_hi = {vfuResponse_VFUNotClear_hi_hi, 1'h0};
  wire [2:0]    vfuResponse_VFUNotClear_hi_1 = {vfuResponse_VFUNotClear_hi_hi_1, 1'h0};
  wire [2:0]    vfuResponse_VFUNotClear_hi_2 = {vfuResponse_VFUNotClear_hi_hi_2, 1'h0};
  wire [3:0]    vfuResponse_3_bits_vxsat = {3'h0, _multiplier_responseIO_bits_vxsat};
  wire [2:0]    vfuResponse_VFUNotClear_hi_3 = {vfuResponse_VFUNotClear_hi_hi_3, 1'h0};
  wire          executeOccupied_4 = _divider_requestIO_ready & _vfuResponse_dividerDistributor_requestToVfu_valid;
  wire [2:0]    vfuResponse_VFUNotClear_hi_4 = {vfuResponse_VFUNotClear_hi_hi_4, 1'h0};
  wire [2:0]    vfuResponse_VFUNotClear_hi_5 = {vfuResponse_VFUNotClear_hi_hi_5, 1'h0};
  wire          VFUNotClear = |vfuResponse_VFUNotClear_hi_5;
  wire [31:0]   responseVec_0_bits_data = selectResponse_bits_data;
  wire [1:0]    responseVec_0_bits_executeIndex = selectResponse_bits_executeIndex;
  wire          responseVec_0_bits_ffoSuccess = selectResponse_bits_ffoSuccess;
  wire [3:0]    responseVec_0_bits_adderMaskResp = selectResponse_bits_adderMaskResp;
  assign responseVec_0_bits_vxsat = selectResponse_bits_vxsat;
  wire          responseDecodeVec_0_logic;
  wire [1:0]    responseVec_0_bits_tag = selectResponse_bits_tag;
  wire [1:0]    vfuResponse_0_bits_tag;
  wire          responseDecodeVec_0_adder;
  wire [1:0]    vfuResponse_1_bits_tag;
  wire          responseDecodeVec_0_shift;
  wire          responseDecodeVec_0_multiplier;
  wire [1:0]    vfuResponse_3_bits_tag;
  wire          responseDecodeVec_0_divider;
  wire          responseDecodeVec_0_other;
  wire [3:0]    vfuResponse_1_bits_vxsat;
  assign selectResponse_bits_tag =
    (responseDecodeVec_0_logic ? vfuResponse_0_bits_tag : 2'h0) | (responseDecodeVec_0_adder ? vfuResponse_1_bits_tag : 2'h0) | (responseDecodeVec_0_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_0_multiplier ? vfuResponse_3_bits_tag : 2'h0) | (responseDecodeVec_0_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_0_other ? _vfuResponse_otherDistributor_responseToSlot_bits_tag : 2'h0);
  wire [3:0]    vfuResponse_1_bits_adderMaskResp;
  assign selectResponse_bits_vxsat =
    (responseDecodeVec_0_adder ? vfuResponse_1_bits_vxsat : 4'h0) | (responseDecodeVec_0_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_0_multiplier ? vfuResponse_3_bits_vxsat : 4'h0)
    | (responseDecodeVec_0_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_0_other ? _vfuResponse_otherDistributor_responseToSlot_bits_vxsat : 4'h0);
  assign selectResponse_bits_adderMaskResp = responseDecodeVec_0_adder ? vfuResponse_1_bits_adderMaskResp : 4'h0;
  wire [1:0]    vfuResponse_1_bits_executeIndex;
  assign selectResponse_bits_ffoSuccess =
    responseDecodeVec_0_shift & _vfuResponse_shiftDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_0_divider & _vfuResponse_dividerDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_0_other
    & _vfuResponse_otherDistributor_responseToSlot_bits_ffoSuccess;
  wire [31:0]   vfuResponse_0_bits_data;
  assign selectResponse_bits_executeIndex = responseDecodeVec_0_adder ? vfuResponse_1_bits_executeIndex : 2'h0;
  wire [31:0]   vfuResponse_1_bits_data;
  wire [31:0]   vfuResponse_3_bits_data;
  wire          vfuResponse_0_valid;
  assign selectResponse_bits_data =
    (responseDecodeVec_0_logic ? vfuResponse_0_bits_data : 32'h0) | (responseDecodeVec_0_adder ? vfuResponse_1_bits_data : 32'h0) | (responseDecodeVec_0_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_0_multiplier ? vfuResponse_3_bits_data : 32'h0) | (responseDecodeVec_0_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_0_other ? _vfuResponse_otherDistributor_responseToSlot_bits_data : 32'h0);
  wire          vfuResponse_1_valid;
  wire          vfuResponse_3_valid;
  wire          selectResponse_valid =
    responseDecodeVec_0_logic & vfuResponse_0_valid | responseDecodeVec_0_adder & vfuResponse_1_valid | responseDecodeVec_0_shift & _vfuResponse_shiftDistributor_responseToSlot_valid | responseDecodeVec_0_multiplier & vfuResponse_3_valid
    | responseDecodeVec_0_divider & _vfuResponse_dividerDistributor_responseToSlot_valid | responseDecodeVec_0_other & _vfuResponse_otherDistributor_responseToSlot_valid;
  assign responseVec_0_valid = selectResponse_valid & selectResponse_bits_tag == 2'h0;
  wire [31:0]   responseVec_1_bits_data = selectResponse_1_bits_data;
  wire [1:0]    responseVec_1_bits_executeIndex = selectResponse_1_bits_executeIndex;
  wire          responseVec_1_bits_ffoSuccess = selectResponse_1_bits_ffoSuccess;
  wire [3:0]    responseVec_1_bits_adderMaskResp = selectResponse_1_bits_adderMaskResp;
  assign responseVec_1_bits_vxsat = selectResponse_1_bits_vxsat;
  wire          responseDecodeVec_1_logic;
  wire [1:0]    responseVec_1_bits_tag = selectResponse_1_bits_tag;
  wire          responseDecodeVec_1_adder;
  wire          responseDecodeVec_1_shift;
  wire          responseDecodeVec_1_multiplier;
  wire          responseDecodeVec_1_divider;
  wire          responseDecodeVec_1_other;
  assign selectResponse_1_bits_tag =
    (responseDecodeVec_1_logic ? vfuResponse_0_bits_tag : 2'h0) | (responseDecodeVec_1_adder ? vfuResponse_1_bits_tag : 2'h0) | (responseDecodeVec_1_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_1_multiplier ? vfuResponse_3_bits_tag : 2'h0) | (responseDecodeVec_1_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_1_other ? _vfuResponse_otherDistributor_responseToSlot_bits_tag : 2'h0);
  assign selectResponse_1_bits_vxsat =
    (responseDecodeVec_1_adder ? vfuResponse_1_bits_vxsat : 4'h0) | (responseDecodeVec_1_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_1_multiplier ? vfuResponse_3_bits_vxsat : 4'h0)
    | (responseDecodeVec_1_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_1_other ? _vfuResponse_otherDistributor_responseToSlot_bits_vxsat : 4'h0);
  assign selectResponse_1_bits_adderMaskResp = responseDecodeVec_1_adder ? vfuResponse_1_bits_adderMaskResp : 4'h0;
  assign selectResponse_1_bits_ffoSuccess =
    responseDecodeVec_1_shift & _vfuResponse_shiftDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_1_divider & _vfuResponse_dividerDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_1_other
    & _vfuResponse_otherDistributor_responseToSlot_bits_ffoSuccess;
  assign selectResponse_1_bits_executeIndex = responseDecodeVec_1_adder ? vfuResponse_1_bits_executeIndex : 2'h0;
  assign selectResponse_1_bits_data =
    (responseDecodeVec_1_logic ? vfuResponse_0_bits_data : 32'h0) | (responseDecodeVec_1_adder ? vfuResponse_1_bits_data : 32'h0) | (responseDecodeVec_1_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_1_multiplier ? vfuResponse_3_bits_data : 32'h0) | (responseDecodeVec_1_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_1_other ? _vfuResponse_otherDistributor_responseToSlot_bits_data : 32'h0);
  wire          selectResponse_1_valid =
    responseDecodeVec_1_logic & vfuResponse_0_valid | responseDecodeVec_1_adder & vfuResponse_1_valid | responseDecodeVec_1_shift & _vfuResponse_shiftDistributor_responseToSlot_valid | responseDecodeVec_1_multiplier & vfuResponse_3_valid
    | responseDecodeVec_1_divider & _vfuResponse_dividerDistributor_responseToSlot_valid | responseDecodeVec_1_other & _vfuResponse_otherDistributor_responseToSlot_valid;
  assign responseVec_1_valid = selectResponse_1_valid & selectResponse_1_bits_tag == 2'h1;
  wire [31:0]   responseVec_2_bits_data = selectResponse_2_bits_data;
  wire [1:0]    responseVec_2_bits_executeIndex = selectResponse_2_bits_executeIndex;
  wire          responseVec_2_bits_ffoSuccess = selectResponse_2_bits_ffoSuccess;
  wire [3:0]    responseVec_2_bits_adderMaskResp = selectResponse_2_bits_adderMaskResp;
  assign responseVec_2_bits_vxsat = selectResponse_2_bits_vxsat;
  wire          responseDecodeVec_2_logic;
  wire [1:0]    responseVec_2_bits_tag = selectResponse_2_bits_tag;
  wire          responseDecodeVec_2_adder;
  wire          responseDecodeVec_2_shift;
  wire          responseDecodeVec_2_multiplier;
  wire          responseDecodeVec_2_divider;
  wire          responseDecodeVec_2_other;
  assign selectResponse_2_bits_tag =
    (responseDecodeVec_2_logic ? vfuResponse_0_bits_tag : 2'h0) | (responseDecodeVec_2_adder ? vfuResponse_1_bits_tag : 2'h0) | (responseDecodeVec_2_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_2_multiplier ? vfuResponse_3_bits_tag : 2'h0) | (responseDecodeVec_2_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_2_other ? _vfuResponse_otherDistributor_responseToSlot_bits_tag : 2'h0);
  assign selectResponse_2_bits_vxsat =
    (responseDecodeVec_2_adder ? vfuResponse_1_bits_vxsat : 4'h0) | (responseDecodeVec_2_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_2_multiplier ? vfuResponse_3_bits_vxsat : 4'h0)
    | (responseDecodeVec_2_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_2_other ? _vfuResponse_otherDistributor_responseToSlot_bits_vxsat : 4'h0);
  assign selectResponse_2_bits_adderMaskResp = responseDecodeVec_2_adder ? vfuResponse_1_bits_adderMaskResp : 4'h0;
  assign selectResponse_2_bits_ffoSuccess =
    responseDecodeVec_2_shift & _vfuResponse_shiftDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_2_divider & _vfuResponse_dividerDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_2_other
    & _vfuResponse_otherDistributor_responseToSlot_bits_ffoSuccess;
  assign selectResponse_2_bits_executeIndex = responseDecodeVec_2_adder ? vfuResponse_1_bits_executeIndex : 2'h0;
  assign selectResponse_2_bits_data =
    (responseDecodeVec_2_logic ? vfuResponse_0_bits_data : 32'h0) | (responseDecodeVec_2_adder ? vfuResponse_1_bits_data : 32'h0) | (responseDecodeVec_2_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_2_multiplier ? vfuResponse_3_bits_data : 32'h0) | (responseDecodeVec_2_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_2_other ? _vfuResponse_otherDistributor_responseToSlot_bits_data : 32'h0);
  wire          selectResponse_2_valid =
    responseDecodeVec_2_logic & vfuResponse_0_valid | responseDecodeVec_2_adder & vfuResponse_1_valid | responseDecodeVec_2_shift & _vfuResponse_shiftDistributor_responseToSlot_valid | responseDecodeVec_2_multiplier & vfuResponse_3_valid
    | responseDecodeVec_2_divider & _vfuResponse_dividerDistributor_responseToSlot_valid | responseDecodeVec_2_other & _vfuResponse_otherDistributor_responseToSlot_valid;
  assign responseVec_2_valid = selectResponse_2_valid & selectResponse_2_bits_tag == 2'h2;
  wire [31:0]   responseVec_3_bits_data = selectResponse_3_bits_data;
  wire [1:0]    responseVec_3_bits_executeIndex = selectResponse_3_bits_executeIndex;
  wire          responseVec_3_bits_ffoSuccess = selectResponse_3_bits_ffoSuccess;
  wire [3:0]    responseVec_3_bits_adderMaskResp = selectResponse_3_bits_adderMaskResp;
  assign responseVec_3_bits_vxsat = selectResponse_3_bits_vxsat;
  wire          responseDecodeVec_3_logic;
  wire [1:0]    responseVec_3_bits_tag = selectResponse_3_bits_tag;
  wire          responseDecodeVec_3_adder;
  wire          responseDecodeVec_3_shift;
  wire          responseDecodeVec_3_multiplier;
  wire          responseDecodeVec_3_divider;
  wire          responseDecodeVec_3_other;
  assign selectResponse_3_bits_tag =
    (responseDecodeVec_3_logic ? vfuResponse_0_bits_tag : 2'h0) | (responseDecodeVec_3_adder ? vfuResponse_1_bits_tag : 2'h0) | (responseDecodeVec_3_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_3_multiplier ? vfuResponse_3_bits_tag : 2'h0) | (responseDecodeVec_3_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_tag : 2'h0)
    | (responseDecodeVec_3_other ? _vfuResponse_otherDistributor_responseToSlot_bits_tag : 2'h0);
  assign selectResponse_3_bits_vxsat =
    (responseDecodeVec_3_adder ? vfuResponse_1_bits_vxsat : 4'h0) | (responseDecodeVec_3_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_3_multiplier ? vfuResponse_3_bits_vxsat : 4'h0)
    | (responseDecodeVec_3_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_vxsat : 4'h0) | (responseDecodeVec_3_other ? _vfuResponse_otherDistributor_responseToSlot_bits_vxsat : 4'h0);
  assign selectResponse_3_bits_adderMaskResp = responseDecodeVec_3_adder ? vfuResponse_1_bits_adderMaskResp : 4'h0;
  assign selectResponse_3_bits_ffoSuccess =
    responseDecodeVec_3_shift & _vfuResponse_shiftDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_3_divider & _vfuResponse_dividerDistributor_responseToSlot_bits_ffoSuccess | responseDecodeVec_3_other
    & _vfuResponse_otherDistributor_responseToSlot_bits_ffoSuccess;
  assign selectResponse_3_bits_executeIndex = responseDecodeVec_3_adder ? vfuResponse_1_bits_executeIndex : 2'h0;
  assign selectResponse_3_bits_data =
    (responseDecodeVec_3_logic ? vfuResponse_0_bits_data : 32'h0) | (responseDecodeVec_3_adder ? vfuResponse_1_bits_data : 32'h0) | (responseDecodeVec_3_shift ? _vfuResponse_shiftDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_3_multiplier ? vfuResponse_3_bits_data : 32'h0) | (responseDecodeVec_3_divider ? _vfuResponse_dividerDistributor_responseToSlot_bits_data : 32'h0)
    | (responseDecodeVec_3_other ? _vfuResponse_otherDistributor_responseToSlot_bits_data : 32'h0);
  wire          selectResponse_3_valid =
    responseDecodeVec_3_logic & vfuResponse_0_valid | responseDecodeVec_3_adder & vfuResponse_1_valid | responseDecodeVec_3_shift & _vfuResponse_shiftDistributor_responseToSlot_valid | responseDecodeVec_3_multiplier & vfuResponse_3_valid
    | responseDecodeVec_3_divider & _vfuResponse_dividerDistributor_responseToSlot_valid | responseDecodeVec_3_other & _vfuResponse_otherDistributor_responseToSlot_valid;
  assign responseVec_3_valid = selectResponse_3_valid & (&selectResponse_3_bits_tag);
  wire          queueBeforeMaskWrite_full;
  reg  [4:0]    queueBeforeMaskWrite_data_vd;
  wire [4:0]    queueBeforeMaskWrite_deq_bits_vd = queueBeforeMaskWrite_data_vd;
  reg  [5:0]    queueBeforeMaskWrite_data_offset;
  wire [5:0]    queueBeforeMaskWrite_deq_bits_offset = queueBeforeMaskWrite_data_offset;
  reg  [3:0]    queueBeforeMaskWrite_data_mask;
  wire [3:0]    queueBeforeMaskWrite_deq_bits_mask = queueBeforeMaskWrite_data_mask;
  reg  [31:0]   queueBeforeMaskWrite_data_data;
  wire [31:0]   queueBeforeMaskWrite_deq_bits_data = queueBeforeMaskWrite_data_data;
  reg           queueBeforeMaskWrite_data_last;
  wire          queueBeforeMaskWrite_deq_bits_last = queueBeforeMaskWrite_data_last;
  reg  [2:0]    queueBeforeMaskWrite_data_instructionIndex;
  wire [2:0]    queueBeforeMaskWrite_deq_bits_instructionIndex = queueBeforeMaskWrite_data_instructionIndex;
  reg           queueBeforeMaskWrite_empty;
  wire          queueBeforeMaskWrite_empty_0 = queueBeforeMaskWrite_empty;
  assign queueBeforeMaskWrite_full = ~queueBeforeMaskWrite_empty;
  wire          queueBeforeMaskWrite_enq_ready;
  wire          queueBeforeMaskWrite_enq_valid;
  wire          queueBeforeMaskWrite_deq_valid = queueBeforeMaskWrite_full;
  wire          queueBeforeMaskWrite_full_0 = queueBeforeMaskWrite_full;
  wire          queueBeforeMaskWrite_push = queueBeforeMaskWrite_enq_ready & queueBeforeMaskWrite_enq_valid;
  wire          queueBeforeMaskWrite_deq_ready;
  assign queueBeforeMaskWrite_enq_ready = queueBeforeMaskWrite_empty | queueBeforeMaskWrite_deq_ready;
  wire          queueBeforeMaskWrite_pop = queueBeforeMaskWrite_deq_ready & queueBeforeMaskWrite_full;
  wire [1:0]    writeCavitation_lo_hi = {allVrfWriteAfterCheck_2_mask == 4'h0, allVrfWriteAfterCheck_1_mask == 4'h0};
  wire [2:0]    writeCavitation_lo = {writeCavitation_lo_hi, allVrfWriteAfterCheck_0_mask == 4'h0};
  wire [1:0]    writeCavitation_hi_lo = {allVrfWriteAfterCheck_4_mask == 4'h0, allVrfWriteAfterCheck_3_mask == 4'h0};
  wire [1:0]    writeCavitation_hi_hi = {allVrfWriteAfterCheck_6_mask == 4'h0, allVrfWriteAfterCheck_5_mask == 4'h0};
  wire [3:0]    writeCavitation_hi = {writeCavitation_hi_hi, writeCavitation_hi_lo};
  wire [6:0]    writeCavitation = {writeCavitation_hi, writeCavitation_lo};
  wire          enqueueFire;
  wire          slot0EnqueueFire = slotEnqueueFire_0;
  wire          enqueueFire_1;
  wire          enqueueFire_2;
  wire          enqueueFire_3;
  assign enqReady = _vrf_writeAllow_0 & (~afterCheckValid_0 | afterCheckDequeueReady_0);
  wire          vrfWriteArbiter_0_ready = enqReady;
  wire          vrfWriteArbiter_0_valid;
  wire          enqFire = enqReady & vrfWriteArbiter_0_valid;
  assign enqReady_1 = _vrf_writeAllow_1 & (~afterCheckValid_1 | afterCheckDequeueReady_1);
  wire          vrfWriteArbiter_1_ready = enqReady_1;
  wire          vrfWriteArbiter_1_valid;
  wire          enqFire_1 = enqReady_1 & vrfWriteArbiter_1_valid;
  assign enqReady_2 = _vrf_writeAllow_2 & (~afterCheckValid_2 | afterCheckDequeueReady_2);
  wire          vrfWriteArbiter_2_ready = enqReady_2;
  wire          vrfWriteArbiter_2_valid;
  wire          enqFire_2 = enqReady_2 & vrfWriteArbiter_2_valid;
  assign enqReady_3 = _vrf_writeAllow_3 & (~afterCheckValid_3 | afterCheckDequeueReady_3);
  wire          vrfWriteArbiter_3_ready = enqReady_3;
  wire          vrfWriteArbiter_3_valid;
  wire          enqFire_3 = enqReady_3 & vrfWriteArbiter_3_valid;
  assign enqReady_4 = _vrf_writeAllow_4 & (~afterCheckValid_4 | afterCheckDequeueReady_4);
  assign vrfWriteArbiter_4_ready = enqReady_4;
  wire          enqFire_4 = enqReady_4 & vrfWriteArbiter_4_valid;
  assign enqReady_5 = _vrf_writeAllow_5 & (~afterCheckValid_5 | afterCheckDequeueReady_5);
  assign crossLaneWriteQueue_0_deq_ready = enqReady_5;
  wire          enqFire_5 = enqReady_5 & crossLaneWriteQueue_0_deq_valid;
  assign enqReady_6 = _vrf_writeAllow_6 & (~afterCheckValid_6 | afterCheckDequeueReady_6);
  assign crossLaneWriteQueue_1_deq_ready = enqReady_6;
  wire          enqFire_6 = enqReady_6 & crossLaneWriteQueue_1_deq_valid;
  wire [1:0]    writeSelect_lo_hi = {afterCheckValid_2, afterCheckValid_1};
  wire [2:0]    writeSelect_lo = {writeSelect_lo_hi, afterCheckValid_0};
  wire [1:0]    writeSelect_hi_lo = {afterCheckValid_4, afterCheckValid_3};
  wire [1:0]    writeSelect_hi_hi = {afterCheckValid_6, afterCheckValid_5};
  wire [3:0]    writeSelect_hi = {writeSelect_hi_hi, writeSelect_hi_lo};
  wire [6:0]    _writeSelect_T_2 = {writeSelect_hi, writeSelect_lo} & ~writeCavitation;
  wire [5:0]    _writeSelect_T_5 = _writeSelect_T_2[5:0] | {_writeSelect_T_2[4:0], 1'h0};
  wire [5:0]    _writeSelect_T_8 = _writeSelect_T_5 | {_writeSelect_T_5[3:0], 2'h0};
  wire [6:0]    writeSelect = {~(_writeSelect_T_8 | {_writeSelect_T_8[1:0], 4'h0}), 1'h1} & _writeSelect_T_2;
  assign afterCheckDequeueReady_0 = writeSelect[0] & queueBeforeMaskWrite_enq_ready | writeCavitation[0];
  assign afterCheckDequeueReady_1 = writeSelect[1] & queueBeforeMaskWrite_enq_ready | writeCavitation[1];
  assign afterCheckDequeueReady_2 = writeSelect[2] & queueBeforeMaskWrite_enq_ready | writeCavitation[2];
  assign afterCheckDequeueReady_3 = writeSelect[3] & queueBeforeMaskWrite_enq_ready | writeCavitation[3];
  assign afterCheckDequeueReady_4 = writeSelect[4] & queueBeforeMaskWrite_enq_ready | writeCavitation[4];
  assign afterCheckDequeueReady_5 = writeSelect[5] & queueBeforeMaskWrite_enq_ready | writeCavitation[5];
  assign afterCheckDequeueReady_6 = writeSelect[6] & queueBeforeMaskWrite_enq_ready | writeCavitation[6];
  assign queueBeforeMaskWrite_enq_valid = |writeSelect;
  wire [2:0]    queueBeforeMaskWrite_enq_bits_instructionIndex =
    (writeSelect[0] ? allVrfWriteAfterCheck_0_instructionIndex : 3'h0) | (writeSelect[1] ? allVrfWriteAfterCheck_1_instructionIndex : 3'h0) | (writeSelect[2] ? allVrfWriteAfterCheck_2_instructionIndex : 3'h0)
    | (writeSelect[3] ? allVrfWriteAfterCheck_3_instructionIndex : 3'h0) | (writeSelect[4] ? allVrfWriteAfterCheck_4_instructionIndex : 3'h0) | (writeSelect[5] ? allVrfWriteAfterCheck_5_instructionIndex : 3'h0)
    | (writeSelect[6] ? allVrfWriteAfterCheck_6_instructionIndex : 3'h0);
  wire          queueBeforeMaskWrite_enq_bits_last =
    writeSelect[0] & allVrfWriteAfterCheck_0_last | writeSelect[1] & allVrfWriteAfterCheck_1_last | writeSelect[2] & allVrfWriteAfterCheck_2_last | writeSelect[3] & allVrfWriteAfterCheck_3_last | writeSelect[4]
    & allVrfWriteAfterCheck_4_last | writeSelect[5] & allVrfWriteAfterCheck_5_last | writeSelect[6] & allVrfWriteAfterCheck_6_last;
  wire [31:0]   queueBeforeMaskWrite_enq_bits_data =
    (writeSelect[0] ? allVrfWriteAfterCheck_0_data : 32'h0) | (writeSelect[1] ? allVrfWriteAfterCheck_1_data : 32'h0) | (writeSelect[2] ? allVrfWriteAfterCheck_2_data : 32'h0) | (writeSelect[3] ? allVrfWriteAfterCheck_3_data : 32'h0)
    | (writeSelect[4] ? allVrfWriteAfterCheck_4_data : 32'h0) | (writeSelect[5] ? allVrfWriteAfterCheck_5_data : 32'h0) | (writeSelect[6] ? allVrfWriteAfterCheck_6_data : 32'h0);
  wire [3:0]    queueBeforeMaskWrite_enq_bits_mask =
    (writeSelect[0] ? allVrfWriteAfterCheck_0_mask : 4'h0) | (writeSelect[1] ? allVrfWriteAfterCheck_1_mask : 4'h0) | (writeSelect[2] ? allVrfWriteAfterCheck_2_mask : 4'h0) | (writeSelect[3] ? allVrfWriteAfterCheck_3_mask : 4'h0)
    | (writeSelect[4] ? allVrfWriteAfterCheck_4_mask : 4'h0) | (writeSelect[5] ? allVrfWriteAfterCheck_5_mask : 4'h0) | (writeSelect[6] ? allVrfWriteAfterCheck_6_mask : 4'h0);
  wire [5:0]    queueBeforeMaskWrite_enq_bits_offset =
    (writeSelect[0] ? allVrfWriteAfterCheck_0_offset : 6'h0) | (writeSelect[1] ? allVrfWriteAfterCheck_1_offset : 6'h0) | (writeSelect[2] ? allVrfWriteAfterCheck_2_offset : 6'h0) | (writeSelect[3] ? allVrfWriteAfterCheck_3_offset : 6'h0)
    | (writeSelect[4] ? allVrfWriteAfterCheck_4_offset : 6'h0) | (writeSelect[5] ? allVrfWriteAfterCheck_5_offset : 6'h0) | (writeSelect[6] ? allVrfWriteAfterCheck_6_offset : 6'h0);
  wire [4:0]    queueBeforeMaskWrite_enq_bits_vd =
    (writeSelect[0] ? allVrfWriteAfterCheck_0_vd : 5'h0) | (writeSelect[1] ? allVrfWriteAfterCheck_1_vd : 5'h0) | (writeSelect[2] ? allVrfWriteAfterCheck_2_vd : 5'h0) | (writeSelect[3] ? allVrfWriteAfterCheck_3_vd : 5'h0)
    | (writeSelect[4] ? allVrfWriteAfterCheck_4_vd : 5'h0) | (writeSelect[5] ? allVrfWriteAfterCheck_5_vd : 5'h0) | (writeSelect[6] ? allVrfWriteAfterCheck_6_vd : 5'h0);
  wire [1:0]    maskControlDataDeq_hitMaskControl_lo =
    {maskControlVec_1_index == slotControl_0_laneRequest_instructionIndex & maskControlVec_1_controlValid, maskControlVec_0_index == slotControl_0_laneRequest_instructionIndex & maskControlVec_0_controlValid};
  wire [1:0]    maskControlDataDeq_hitMaskControl_hi =
    {maskControlVec_3_index == slotControl_0_laneRequest_instructionIndex & maskControlVec_3_controlValid, maskControlVec_2_index == slotControl_0_laneRequest_instructionIndex & maskControlVec_2_controlValid};
  wire [3:0]    maskControlDataDeq_hitMaskControl = {maskControlDataDeq_hitMaskControl_hi, maskControlDataDeq_hitMaskControl_lo};
  wire          maskControlDataDeq_dataValid =
    maskControlDataDeq_hitMaskControl[0] & maskControlVec_0_dataValid | maskControlDataDeq_hitMaskControl[1] & maskControlVec_1_dataValid | maskControlDataDeq_hitMaskControl[2] & maskControlVec_2_dataValid
    | maskControlDataDeq_hitMaskControl[3] & maskControlVec_3_dataValid;
  assign maskControlDataDeq_data =
    (maskControlDataDeq_hitMaskControl[0] ? maskControlVec_0_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl[1] ? maskControlVec_1_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl[2] ? maskControlVec_2_maskData : 32'h0)
    | (maskControlDataDeq_hitMaskControl[3] ? maskControlVec_3_maskData : 32'h0);
  wire [31:0]   maskDataVec_0 = maskControlDataDeq_data;
  wire [7:0]    maskControlDataDeq_group =
    (maskControlDataDeq_hitMaskControl[0] ? maskControlVec_0_group : 8'h0) | (maskControlDataDeq_hitMaskControl[1] ? maskControlVec_1_group : 8'h0) | (maskControlDataDeq_hitMaskControl[2] ? maskControlVec_2_group : 8'h0)
    | (maskControlDataDeq_hitMaskControl[3] ? maskControlVec_3_group : 8'h0);
  wire [7:0]    slotMaskRequestVec_0_bits;
  wire          maskControlDataDeq_sameGroup = maskControlDataDeq_group == slotMaskRequestVec_0_bits;
  assign maskControlDataDeq_maskRequestFire = slotMaskRequestVec_0_valid & maskControlDataDeq_dataValid;
  assign maskRequestFireOH_0 = maskControlDataDeq_maskRequestFire;
  wire [1:0]    maskControlDataDeq_hitMaskControl_lo_1 =
    {maskControlVec_1_index == slotControl_1_laneRequest_instructionIndex & maskControlVec_1_controlValid, maskControlVec_0_index == slotControl_1_laneRequest_instructionIndex & maskControlVec_0_controlValid};
  wire [1:0]    maskControlDataDeq_hitMaskControl_hi_1 =
    {maskControlVec_3_index == slotControl_1_laneRequest_instructionIndex & maskControlVec_3_controlValid, maskControlVec_2_index == slotControl_1_laneRequest_instructionIndex & maskControlVec_2_controlValid};
  wire [3:0]    maskControlDataDeq_hitMaskControl_1 = {maskControlDataDeq_hitMaskControl_hi_1, maskControlDataDeq_hitMaskControl_lo_1};
  wire          maskControlDataDeq_dataValid_1 =
    maskControlDataDeq_hitMaskControl_1[0] & maskControlVec_0_dataValid | maskControlDataDeq_hitMaskControl_1[1] & maskControlVec_1_dataValid | maskControlDataDeq_hitMaskControl_1[2] & maskControlVec_2_dataValid
    | maskControlDataDeq_hitMaskControl_1[3] & maskControlVec_3_dataValid;
  assign maskControlDataDeq_data_1 =
    (maskControlDataDeq_hitMaskControl_1[0] ? maskControlVec_0_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl_1[1] ? maskControlVec_1_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl_1[2] ? maskControlVec_2_maskData : 32'h0)
    | (maskControlDataDeq_hitMaskControl_1[3] ? maskControlVec_3_maskData : 32'h0);
  wire [31:0]   maskDataVec_1 = maskControlDataDeq_data_1;
  wire [7:0]    maskControlDataDeq_group_1 =
    (maskControlDataDeq_hitMaskControl_1[0] ? maskControlVec_0_group : 8'h0) | (maskControlDataDeq_hitMaskControl_1[1] ? maskControlVec_1_group : 8'h0) | (maskControlDataDeq_hitMaskControl_1[2] ? maskControlVec_2_group : 8'h0)
    | (maskControlDataDeq_hitMaskControl_1[3] ? maskControlVec_3_group : 8'h0);
  wire [7:0]    slotMaskRequestVec_1_bits;
  wire          maskControlDataDeq_sameGroup_1 = maskControlDataDeq_group_1 == slotMaskRequestVec_1_bits;
  assign maskControlDataDeq_maskRequestFire_1 = slotMaskRequestVec_1_valid & maskControlDataDeq_dataValid_1 & ~slotEnqueueFire_0;
  assign maskRequestFireOH_1 = maskControlDataDeq_maskRequestFire_1;
  wire [1:0]    maskControlDataDeq_hitMaskControl_lo_2 =
    {maskControlVec_1_index == slotControl_2_laneRequest_instructionIndex & maskControlVec_1_controlValid, maskControlVec_0_index == slotControl_2_laneRequest_instructionIndex & maskControlVec_0_controlValid};
  wire [1:0]    maskControlDataDeq_hitMaskControl_hi_2 =
    {maskControlVec_3_index == slotControl_2_laneRequest_instructionIndex & maskControlVec_3_controlValid, maskControlVec_2_index == slotControl_2_laneRequest_instructionIndex & maskControlVec_2_controlValid};
  wire [3:0]    maskControlDataDeq_hitMaskControl_2 = {maskControlDataDeq_hitMaskControl_hi_2, maskControlDataDeq_hitMaskControl_lo_2};
  wire          maskControlDataDeq_dataValid_2 =
    maskControlDataDeq_hitMaskControl_2[0] & maskControlVec_0_dataValid | maskControlDataDeq_hitMaskControl_2[1] & maskControlVec_1_dataValid | maskControlDataDeq_hitMaskControl_2[2] & maskControlVec_2_dataValid
    | maskControlDataDeq_hitMaskControl_2[3] & maskControlVec_3_dataValid;
  assign maskControlDataDeq_data_2 =
    (maskControlDataDeq_hitMaskControl_2[0] ? maskControlVec_0_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl_2[1] ? maskControlVec_1_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl_2[2] ? maskControlVec_2_maskData : 32'h0)
    | (maskControlDataDeq_hitMaskControl_2[3] ? maskControlVec_3_maskData : 32'h0);
  wire [31:0]   maskDataVec_2 = maskControlDataDeq_data_2;
  wire [7:0]    maskControlDataDeq_group_2 =
    (maskControlDataDeq_hitMaskControl_2[0] ? maskControlVec_0_group : 8'h0) | (maskControlDataDeq_hitMaskControl_2[1] ? maskControlVec_1_group : 8'h0) | (maskControlDataDeq_hitMaskControl_2[2] ? maskControlVec_2_group : 8'h0)
    | (maskControlDataDeq_hitMaskControl_2[3] ? maskControlVec_3_group : 8'h0);
  wire [7:0]    slotMaskRequestVec_2_bits;
  wire          maskControlDataDeq_sameGroup_2 = maskControlDataDeq_group_2 == slotMaskRequestVec_2_bits;
  wire          slotEnqueueFire_1;
  assign maskControlDataDeq_maskRequestFire_2 = slotMaskRequestVec_2_valid & maskControlDataDeq_dataValid_2 & ~slotEnqueueFire_1;
  assign maskRequestFireOH_2 = maskControlDataDeq_maskRequestFire_2;
  wire [1:0]    maskControlDataDeq_hitMaskControl_lo_3 =
    {maskControlVec_1_index == slotControl_3_laneRequest_instructionIndex & maskControlVec_1_controlValid, maskControlVec_0_index == slotControl_3_laneRequest_instructionIndex & maskControlVec_0_controlValid};
  wire [1:0]    maskControlDataDeq_hitMaskControl_hi_3 =
    {maskControlVec_3_index == slotControl_3_laneRequest_instructionIndex & maskControlVec_3_controlValid, maskControlVec_2_index == slotControl_3_laneRequest_instructionIndex & maskControlVec_2_controlValid};
  wire [3:0]    maskControlDataDeq_hitMaskControl_3 = {maskControlDataDeq_hitMaskControl_hi_3, maskControlDataDeq_hitMaskControl_lo_3};
  wire          maskControlDataDeq_dataValid_3 =
    maskControlDataDeq_hitMaskControl_3[0] & maskControlVec_0_dataValid | maskControlDataDeq_hitMaskControl_3[1] & maskControlVec_1_dataValid | maskControlDataDeq_hitMaskControl_3[2] & maskControlVec_2_dataValid
    | maskControlDataDeq_hitMaskControl_3[3] & maskControlVec_3_dataValid;
  assign maskControlDataDeq_data_3 =
    (maskControlDataDeq_hitMaskControl_3[0] ? maskControlVec_0_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl_3[1] ? maskControlVec_1_maskData : 32'h0) | (maskControlDataDeq_hitMaskControl_3[2] ? maskControlVec_2_maskData : 32'h0)
    | (maskControlDataDeq_hitMaskControl_3[3] ? maskControlVec_3_maskData : 32'h0);
  wire [31:0]   maskDataVec_3 = maskControlDataDeq_data_3;
  wire [7:0]    maskControlDataDeq_group_3 =
    (maskControlDataDeq_hitMaskControl_3[0] ? maskControlVec_0_group : 8'h0) | (maskControlDataDeq_hitMaskControl_3[1] ? maskControlVec_1_group : 8'h0) | (maskControlDataDeq_hitMaskControl_3[2] ? maskControlVec_2_group : 8'h0)
    | (maskControlDataDeq_hitMaskControl_3[3] ? maskControlVec_3_group : 8'h0);
  wire [7:0]    slotMaskRequestVec_3_bits;
  wire          maskControlDataDeq_sameGroup_3 = maskControlDataDeq_group_3 == slotMaskRequestVec_3_bits;
  wire          slotEnqueueFire_2;
  assign maskControlDataDeq_maskRequestFire_3 = slotMaskRequestVec_3_valid & maskControlDataDeq_dataValid_3 & ~slotEnqueueFire_2;
  assign maskRequestFireOH_3 = maskControlDataDeq_maskRequestFire_3;
  wire [3:0]    maskControlDataDeq =
    (maskControlDataDeq_maskRequestFire ? maskControlDataDeq_hitMaskControl : 4'h0) | (maskControlDataDeq_maskRequestFire_1 ? maskControlDataDeq_hitMaskControl_1 : 4'h0)
    | (maskControlDataDeq_maskRequestFire_2 ? maskControlDataDeq_hitMaskControl_2 : 4'h0) | (maskControlDataDeq_maskRequestFire_3 ? maskControlDataDeq_hitMaskControl_3 : 4'h0);
  wire          maskLogicCompleted = laneRequest_bits_decodeResult_maskLogic_0 & {7'h0, laneIndex, 5'h0} >= laneRequest_bits_csrInterface_vl_0;
  wire [3:0]    _GEN_5 = {2'h0, laneRequest_bits_csrInterface_vSew_0};
  wire          _selectMask_T = laneRequest_bits_decodeResult_nr_0 | laneRequest_bits_lsWholeReg_0;
  wire          entranceControl_instructionFinished = ({10'h0, {laneIndex, 2'h0} >> _GEN_5} >= laneRequest_bits_csrInterface_vl_0 | maskLogicCompleted) & ~_selectMask_T;
  wire [12:0]   lastElementIndex = laneRequest_bits_csrInterface_vl_0[12:0] - {12'h0, |laneRequest_bits_csrInterface_vl_0};
  wire [3:0]    requestVSew1H = 4'h1 << _GEN_5;
  wire [10:0]   lastGroupForInstruction = {1'h0, {1'h0, requestVSew1H[0] ? lastElementIndex[12:4] : 9'h0} | (requestVSew1H[1] ? lastElementIndex[12:3] : 10'h0)} | (requestVSew1H[2] ? lastElementIndex[12:2] : 11'h0);
  wire [1:0]    lastLaneIndex = (requestVSew1H[0] ? lastElementIndex[3:2] : 2'h0) | (requestVSew1H[1] ? lastElementIndex[2:1] : 2'h0) | (requestVSew1H[2] ? lastElementIndex[1:0] : 2'h0);
  wire          lanePositionLargerThanEndLane = laneIndex > lastLaneIndex;
  wire          isEndLane = laneIndex == lastLaneIndex;
  wire [10:0]   lastGroupForLane = lastGroupForInstruction - {10'h0, lanePositionLargerThanEndLane};
  wire [4:0]    vlTail = laneRequest_bits_csrInterface_vl_0[4:0];
  wire [1:0]    vlBody = laneRequest_bits_csrInterface_vl_0[6:5];
  wire [6:0]    vlHead = laneRequest_bits_csrInterface_vl_0[13:7];
  wire [31:0]   _lastGroupMask_T = 32'h1 << vlTail;
  wire [29:0]   _GEN_6 = _lastGroupMask_T[30:1] | _lastGroupMask_T[31:2];
  wire [28:0]   _GEN_7 = _GEN_6[28:0] | {_lastGroupMask_T[31], _GEN_6[29:2]};
  wire [26:0]   _GEN_8 = _GEN_7[26:0] | {_lastGroupMask_T[31], _GEN_6[29], _GEN_7[28:4]};
  wire [22:0]   _GEN_9 = _GEN_8[22:0] | {_lastGroupMask_T[31], _GEN_6[29], _GEN_7[28:27], _GEN_8[26:8]};
  wire [30:0]   lastGroupMask = {_lastGroupMask_T[31], _GEN_6[29], _GEN_7[28:27], _GEN_8[26:23], _GEN_9[22:15], _GEN_9[14:0] | {_lastGroupMask_T[31], _GEN_6[29], _GEN_7[28:27], _GEN_8[26:23], _GEN_9[22:16]}};
  wire          dataPathMisaligned = |vlTail;
  wire [8:0]    maskeDataGroup = {vlHead, vlBody} - {8'h0, ~dataPathMisaligned};
  wire [1:0]    lastLaneIndexForMaskLogic = maskeDataGroup[1:0];
  wire          isLastLaneForMaskLogic = lastLaneIndexForMaskLogic == laneIndex;
  wire [6:0]    lastGroupCountForMaskLogic = maskeDataGroup[8:2] - {6'h0, ((|vlBody) | dataPathMisaligned) & laneIndex > lastLaneIndexForMaskLogic};
  wire          misalignedForOther = requestVSew1H[0] & (|(laneRequest_bits_csrInterface_vl_0[1:0])) | requestVSew1H[1] & laneRequest_bits_csrInterface_vl_0[0];
  wire [9:0]    entranceControl_lastGroupForInstruction = laneRequest_bits_decodeResult_maskLogic_0 ? {3'h0, lastGroupCountForMaskLogic} : lastGroupForLane[9:0];
  wire          entranceControl_isLastLaneForInstruction = laneRequest_bits_decodeResult_maskLogic_0 ? isLastLaneForMaskLogic & dataPathMisaligned : isEndLane & misalignedForOther;
  wire          entranceControl_additionalRW = (laneRequest_bits_decodeResult_crossRead_0 | laneRequest_bits_decodeResult_crossWrite_0) & lanePositionLargerThanEndLane & lastLaneIndex != 2'h3 & (|laneRequest_bits_csrInterface_vl_0);
  assign slotShiftValid_1 = ~slotOccupied_0 | ~slotOccupied_1;
  wire          _slotFree_T_3 = ~slotOccupied_0 | ~slotOccupied_1;
  assign slotShiftValid_2 = _slotFree_T_3 | ~slotOccupied_2;
  wire          _slotFree_T_5 = _slotFree_T_3 | ~slotOccupied_2;
  assign slotShiftValid_3 = _slotFree_T_5 | ~slotOccupied_3;
  assign slotFree = _slotFree_T_5 | ~slotOccupied_3;
  assign laneRequest_ready_0 = slotFree;
  assign enqueueFire = enqueueReady & enqueueValid;
  assign slotEnqueueFire_0 = enqueueFire;
  assign enqueueFire_1 = enqueueReady_1 & enqueueValid_1;
  assign slotEnqueueFire_1 = enqueueFire_1;
  assign enqueueFire_2 = enqueueReady_2 & enqueueValid_2;
  assign slotEnqueueFire_2 = enqueueFire_2;
  assign enqueueFire_3 = enqueueReady_3 & enqueueValid_3;
  wire          slotEnqueueFire_3 = enqueueFire_3;
  wire          slotDequeueFire_0 = slotCanShift_0 & slotOccupied_0;
  wire          instructionFinishAndNotReportByTop = entranceControl_instructionFinished & ~laneRequest_bits_decodeResult_readOnly_0 & writeCount == 10'h0;
  wire          needWaitCrossWrite = laneRequest_bits_decodeResult_crossWrite_0 & (|laneRequest_bits_csrInterface_vl_0);
  wire          _GEN_10 = laneRequest_bits_issueInst_0 & (~instructionFinishAndNotReportByTop | needWaitCrossWrite);
  wire          _GEN_11 = laneRequest_bits_loadStore_0 & ~laneRequest_bits_store_0;
  wire [127:0]  nrMask_lo_lo = {{64{laneRequest_bits_segment_0 == 3'h0}}, 64'h0};
  wire [127:0]  nrMask_lo_hi = {{64{laneRequest_bits_segment_0 < 3'h3}}, {64{laneRequest_bits_segment_0 < 3'h2}}};
  wire [255:0]  nrMask_lo = {nrMask_lo_hi, nrMask_lo_lo};
  wire [127:0]  nrMask_hi_lo = {{64{laneRequest_bits_segment_0 < 3'h5}}, {64{~(laneRequest_bits_segment_0[2])}}};
  wire [127:0]  nrMask_hi_hi = {{64{laneRequest_bits_segment_0 != 3'h7}}, {64{laneRequest_bits_segment_0[2:1] != 2'h3}}};
  wire [255:0]  nrMask_hi = {nrMask_hi_hi, nrMask_hi_lo};
  wire [511:0]  nrMask = {nrMask_hi, nrMask_lo};
  wire [1023:0] _lastWriteOH_T = 1024'h1 << writeCount;
  wire [511:0]  _lastWriteOH_T_4 = _lastWriteOH_T[511:0] | {_lastWriteOH_T[510:0], 1'h0};
  wire [511:0]  _lastWriteOH_T_7 = _lastWriteOH_T_4 | {_lastWriteOH_T_4[509:0], 2'h0};
  wire [511:0]  _lastWriteOH_T_10 = _lastWriteOH_T_7 | {_lastWriteOH_T_7[507:0], 4'h0};
  wire [511:0]  _lastWriteOH_T_13 = _lastWriteOH_T_10 | {_lastWriteOH_T_10[503:0], 8'h0};
  wire [511:0]  _lastWriteOH_T_16 = _lastWriteOH_T_13 | {_lastWriteOH_T_13[495:0], 16'h0};
  wire [511:0]  _lastWriteOH_T_19 = _lastWriteOH_T_16 | {_lastWriteOH_T_16[479:0], 32'h0};
  wire [511:0]  _lastWriteOH_T_22 = _lastWriteOH_T_19 | {_lastWriteOH_T_19[447:0], 64'h0};
  wire [511:0]  _lastWriteOH_T_25 = _lastWriteOH_T_22 | {_lastWriteOH_T_22[383:0], 128'h0};
  wire [511:0]  lastWriteOH = _lastWriteOH_T_25 | {_lastWriteOH_T_25[255:0], 256'h0};
  wire          segmentLS = laneRequest_bits_loadStore_0 & (|laneRequest_bits_segment_0) & ~laneRequest_bits_lsWholeReg_0;
  wire [1:0]    mul = laneRequest_bits_csrInterface_vlmul_0[2] ? 2'h0 : laneRequest_bits_csrInterface_vlmul_0[1:0];
  wire [3:0]    mul1H = 4'h1 << mul;
  wire [7:0]    seg1H = 8'h1 << laneRequest_bits_segment_0;
  wire [63:0]   segmentMask_writeOHGroup_0 = lastWriteOH[63:0];
  wire [63:0]   segmentMask_writeOHGroup_1 = lastWriteOH[127:64];
  wire [63:0]   segmentMask_writeOHGroup_2 = lastWriteOH[191:128];
  wire [63:0]   segmentMask_writeOHGroup_3 = lastWriteOH[255:192];
  wire [63:0]   segmentMask_writeOHGroup_4 = lastWriteOH[319:256];
  wire [63:0]   segmentMask_writeOHGroup_5 = lastWriteOH[383:320];
  wire [63:0]   segmentMask_writeOHGroup_6 = lastWriteOH[447:384];
  wire [63:0]   segmentMask_writeOHGroup_7 = lastWriteOH[511:448];
  wire [63:0]   segmentMask_segMask1 = (mul1H[2] | mul1H[1]) & seg1H[1] | mul1H[1] & (seg1H[2] | seg1H[3]) ? segmentMask_writeOHGroup_1 : segmentMask_writeOHGroup_0;
  wire [63:0]   segmentMask_segMask2 = mul1H[2] & seg1H[1] ? segmentMask_writeOHGroup_2 : mul1H[1] & seg1H[1] ? 64'hFFFFFFFFFFFFFFFF : segmentMask_writeOHGroup_0;
  wire          _GEN_12 = seg1H[6] | seg1H[5] | seg1H[4];
  wire [63:0]   segmentMask_segMask3 =
    mul1H[2] & seg1H[1] ? segmentMask_writeOHGroup_3 : mul1H[1] & (seg1H[1] | seg1H[2] | seg1H[3]) ? segmentMask_writeOHGroup_1 : mul1H[0] & seg1H[3] | seg1H[7] | _GEN_12 ? segmentMask_writeOHGroup_0 : 64'hFFFFFFFFFFFFFFFF;
  wire [63:0]   segmentMask_segMask4 = mul1H[2] & seg1H[1] | mul1H[1] & (seg1H[2] | seg1H[3]) | seg1H[7] | _GEN_12 ? segmentMask_writeOHGroup_0 : 64'hFFFFFFFFFFFFFFFF;
  wire [63:0]   segmentMask_segMask5 = mul1H[2] & seg1H[1] | mul1H[1] & (seg1H[2] | seg1H[3]) ? segmentMask_writeOHGroup_1 : mul1H[0] & (seg1H[7] | seg1H[6] | seg1H[5]) ? segmentMask_writeOHGroup_0 : 64'hFFFFFFFFFFFFFFFF;
  wire [63:0]   segmentMask_segMask6 = mul1H[2] & seg1H[1] ? segmentMask_writeOHGroup_2 : mul1H[1] & seg1H[3] | mul1H[0] & (seg1H[7] | seg1H[6]) ? segmentMask_writeOHGroup_0 : 64'hFFFFFFFFFFFFFFFF;
  wire [63:0]   segmentMask_segMask7 = mul1H[2] & seg1H[1] ? segmentMask_writeOHGroup_3 : mul1H[1] & seg1H[3] ? segmentMask_writeOHGroup_1 : mul1H[0] & seg1H[7] ? segmentMask_writeOHGroup_0 : 64'hFFFFFFFFFFFFFFFF;
  wire [511:0]  segmentMask = {segmentMask_segMask7, segmentMask_segMask6, segmentMask_segMask5, segmentMask_segMask4, segmentMask_segMask3, segmentMask_segMask2, segmentMask_segMask1, segmentMask_writeOHGroup_0};
  wire [511:0]  selectMask = segmentLS ? segmentMask : _selectMask_T ? nrMask : lastWriteOH;
  wire [7:0]    instructionValid;
  wire [7:0]    instructionFinishInSlot = ~instructionValid & instructionValidNext;
  reg           emptyInstValid;
  reg  [7:0]    emptyInstCount;
  wire [7:0]    emptyReport = emptyInstValid ? emptyInstCount : 8'h0;
  wire [7:0]    _instructionFinished_output = _vrf_vrfSlotRelease | emptyReport;
  wire          _GEN_13 = vrfWriteChannel_ready_0 & vrfWriteChannel_valid_0;
  wire [7:0]    instInSlot =
    (slotOccupied_0 ? 8'h1 << slotControl_0_laneRequest_instructionIndex : 8'h0) | (slotOccupied_1 ? 8'h1 << slotControl_1_laneRequest_instructionIndex : 8'h0) | (slotOccupied_2 ? 8'h1 << slotControl_2_laneRequest_instructionIndex : 8'h0)
    | (slotOccupied_3 ? 8'h1 << slotControl_3_laneRequest_instructionIndex : 8'h0);
  assign instructionValid = _tokenManager_instructionValid | instInSlot;
  wire [4:0]    vrfWriteArbiter_0_bits_vd;
  wire [5:0]    vrfWriteArbiter_0_bits_offset;
  wire [3:0]    vrfWriteArbiter_0_bits_mask;
  wire [31:0]   vrfWriteArbiter_0_bits_data;
  wire          vrfWriteArbiter_0_bits_last;
  wire [2:0]    vrfWriteArbiter_0_bits_instructionIndex;
  wire [4:0]    vrfWriteArbiter_1_bits_vd;
  wire [5:0]    vrfWriteArbiter_1_bits_offset;
  wire [3:0]    vrfWriteArbiter_1_bits_mask;
  wire [31:0]   vrfWriteArbiter_1_bits_data;
  wire          vrfWriteArbiter_1_bits_last;
  wire [2:0]    vrfWriteArbiter_1_bits_instructionIndex;
  wire [4:0]    vrfWriteArbiter_2_bits_vd;
  wire [5:0]    vrfWriteArbiter_2_bits_offset;
  wire [3:0]    vrfWriteArbiter_2_bits_mask;
  wire [31:0]   vrfWriteArbiter_2_bits_data;
  wire          vrfWriteArbiter_2_bits_last;
  wire [2:0]    vrfWriteArbiter_2_bits_instructionIndex;
  wire [4:0]    vrfWriteArbiter_3_bits_vd;
  wire [5:0]    vrfWriteArbiter_3_bits_offset;
  wire [3:0]    vrfWriteArbiter_3_bits_mask;
  wire [31:0]   vrfWriteArbiter_3_bits_data;
  wire          vrfWriteArbiter_3_bits_last;
  wire [2:0]    vrfWriteArbiter_3_bits_instructionIndex;
  always @(posedge clock) begin
    if (reset) begin
      slotOccupied_0 <= 1'h0;
      slotOccupied_1 <= 1'h0;
      slotOccupied_2 <= 1'h0;
      slotOccupied_3 <= 1'h0;
      maskGroupCountVec_0 <= 8'h0;
      maskGroupCountVec_1 <= 8'h0;
      maskGroupCountVec_2 <= 8'h0;
      maskGroupCountVec_3 <= 8'h0;
      maskIndexVec_0 <= 5'h0;
      maskIndexVec_1 <= 5'h0;
      maskIndexVec_2 <= 5'h0;
      maskIndexVec_3 <= 5'h0;
      allVrfWriteAfterCheck_0_vd <= 5'h0;
      allVrfWriteAfterCheck_0_offset <= 6'h0;
      allVrfWriteAfterCheck_0_mask <= 4'h0;
      allVrfWriteAfterCheck_0_data <= 32'h0;
      allVrfWriteAfterCheck_0_last <= 1'h0;
      allVrfWriteAfterCheck_0_instructionIndex <= 3'h0;
      allVrfWriteAfterCheck_1_vd <= 5'h0;
      allVrfWriteAfterCheck_1_offset <= 6'h0;
      allVrfWriteAfterCheck_1_mask <= 4'h0;
      allVrfWriteAfterCheck_1_data <= 32'h0;
      allVrfWriteAfterCheck_1_last <= 1'h0;
      allVrfWriteAfterCheck_1_instructionIndex <= 3'h0;
      allVrfWriteAfterCheck_2_vd <= 5'h0;
      allVrfWriteAfterCheck_2_offset <= 6'h0;
      allVrfWriteAfterCheck_2_mask <= 4'h0;
      allVrfWriteAfterCheck_2_data <= 32'h0;
      allVrfWriteAfterCheck_2_last <= 1'h0;
      allVrfWriteAfterCheck_2_instructionIndex <= 3'h0;
      allVrfWriteAfterCheck_3_vd <= 5'h0;
      allVrfWriteAfterCheck_3_offset <= 6'h0;
      allVrfWriteAfterCheck_3_mask <= 4'h0;
      allVrfWriteAfterCheck_3_data <= 32'h0;
      allVrfWriteAfterCheck_3_last <= 1'h0;
      allVrfWriteAfterCheck_3_instructionIndex <= 3'h0;
      allVrfWriteAfterCheck_4_vd <= 5'h0;
      allVrfWriteAfterCheck_4_offset <= 6'h0;
      allVrfWriteAfterCheck_4_mask <= 4'h0;
      allVrfWriteAfterCheck_4_data <= 32'h0;
      allVrfWriteAfterCheck_4_last <= 1'h0;
      allVrfWriteAfterCheck_4_instructionIndex <= 3'h0;
      allVrfWriteAfterCheck_5_vd <= 5'h0;
      allVrfWriteAfterCheck_5_offset <= 6'h0;
      allVrfWriteAfterCheck_5_mask <= 4'h0;
      allVrfWriteAfterCheck_5_data <= 32'h0;
      allVrfWriteAfterCheck_5_last <= 1'h0;
      allVrfWriteAfterCheck_5_instructionIndex <= 3'h0;
      allVrfWriteAfterCheck_6_vd <= 5'h0;
      allVrfWriteAfterCheck_6_offset <= 6'h0;
      allVrfWriteAfterCheck_6_mask <= 4'h0;
      allVrfWriteAfterCheck_6_data <= 32'h0;
      allVrfWriteAfterCheck_6_last <= 1'h0;
      allVrfWriteAfterCheck_6_instructionIndex <= 3'h0;
      afterCheckValid_0 <= 1'h0;
      afterCheckValid_1 <= 1'h0;
      afterCheckValid_2 <= 1'h0;
      afterCheckValid_3 <= 1'h0;
      afterCheckValid_4 <= 1'h0;
      afterCheckValid_5 <= 1'h0;
      afterCheckValid_6 <= 1'h0;
      maskControlVec_0_index <= 3'h0;
      maskControlVec_0_sew <= 2'h0;
      maskControlVec_0_maskData <= 32'h0;
      maskControlVec_0_group <= 8'h0;
      maskControlVec_0_dataValid <= 1'h0;
      maskControlVec_0_waiteResponse <= 1'h0;
      maskControlVec_0_controlValid <= 1'h0;
      maskControlVec_responseFire_pipe_v <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_v <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_v <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v <= 1'h0;
      maskControlVec_1_index <= 3'h0;
      maskControlVec_1_sew <= 2'h0;
      maskControlVec_1_maskData <= 32'h0;
      maskControlVec_1_group <= 8'h0;
      maskControlVec_1_dataValid <= 1'h0;
      maskControlVec_1_waiteResponse <= 1'h0;
      maskControlVec_1_controlValid <= 1'h0;
      maskControlVec_responseFire_pipe_v_1 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_v_1 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_v_1 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_1 <= 1'h0;
      maskControlVec_2_index <= 3'h0;
      maskControlVec_2_sew <= 2'h0;
      maskControlVec_2_maskData <= 32'h0;
      maskControlVec_2_group <= 8'h0;
      maskControlVec_2_dataValid <= 1'h0;
      maskControlVec_2_waiteResponse <= 1'h0;
      maskControlVec_2_controlValid <= 1'h0;
      maskControlVec_responseFire_pipe_v_2 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_v_2 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_v_2 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_2 <= 1'h0;
      maskControlVec_3_index <= 3'h0;
      maskControlVec_3_sew <= 2'h0;
      maskControlVec_3_maskData <= 32'h0;
      maskControlVec_3_group <= 8'h0;
      maskControlVec_3_dataValid <= 1'h0;
      maskControlVec_3_waiteResponse <= 1'h0;
      maskControlVec_3_controlValid <= 1'h0;
      maskControlVec_responseFire_pipe_v_3 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_v_3 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_v_3 <= 1'h0;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_3 <= 1'h0;
      slotControl_0_laneRequest_instructionIndex <= 3'h0;
      slotControl_0_laneRequest_decodeResult_specialSlot <= 1'h0;
      slotControl_0_laneRequest_decodeResult_topUop <= 5'h0;
      slotControl_0_laneRequest_decodeResult_popCount <= 1'h0;
      slotControl_0_laneRequest_decodeResult_ffo <= 1'h0;
      slotControl_0_laneRequest_decodeResult_average <= 1'h0;
      slotControl_0_laneRequest_decodeResult_reverse <= 1'h0;
      slotControl_0_laneRequest_decodeResult_dontNeedExecuteInLane <= 1'h0;
      slotControl_0_laneRequest_decodeResult_scheduler <= 1'h0;
      slotControl_0_laneRequest_decodeResult_sReadVD <= 1'h0;
      slotControl_0_laneRequest_decodeResult_vtype <= 1'h0;
      slotControl_0_laneRequest_decodeResult_sWrite <= 1'h0;
      slotControl_0_laneRequest_decodeResult_crossRead <= 1'h0;
      slotControl_0_laneRequest_decodeResult_crossWrite <= 1'h0;
      slotControl_0_laneRequest_decodeResult_maskUnit <= 1'h0;
      slotControl_0_laneRequest_decodeResult_special <= 1'h0;
      slotControl_0_laneRequest_decodeResult_saturate <= 1'h0;
      slotControl_0_laneRequest_decodeResult_vwmacc <= 1'h0;
      slotControl_0_laneRequest_decodeResult_readOnly <= 1'h0;
      slotControl_0_laneRequest_decodeResult_maskSource <= 1'h0;
      slotControl_0_laneRequest_decodeResult_maskDestination <= 1'h0;
      slotControl_0_laneRequest_decodeResult_maskLogic <= 1'h0;
      slotControl_0_laneRequest_decodeResult_uop <= 4'h0;
      slotControl_0_laneRequest_decodeResult_iota <= 1'h0;
      slotControl_0_laneRequest_decodeResult_mv <= 1'h0;
      slotControl_0_laneRequest_decodeResult_extend <= 1'h0;
      slotControl_0_laneRequest_decodeResult_unOrderWrite <= 1'h0;
      slotControl_0_laneRequest_decodeResult_compress <= 1'h0;
      slotControl_0_laneRequest_decodeResult_gather16 <= 1'h0;
      slotControl_0_laneRequest_decodeResult_gather <= 1'h0;
      slotControl_0_laneRequest_decodeResult_slid <= 1'h0;
      slotControl_0_laneRequest_decodeResult_targetRd <= 1'h0;
      slotControl_0_laneRequest_decodeResult_widenReduce <= 1'h0;
      slotControl_0_laneRequest_decodeResult_red <= 1'h0;
      slotControl_0_laneRequest_decodeResult_nr <= 1'h0;
      slotControl_0_laneRequest_decodeResult_itype <= 1'h0;
      slotControl_0_laneRequest_decodeResult_unsigned1 <= 1'h0;
      slotControl_0_laneRequest_decodeResult_unsigned0 <= 1'h0;
      slotControl_0_laneRequest_decodeResult_other <= 1'h0;
      slotControl_0_laneRequest_decodeResult_multiCycle <= 1'h0;
      slotControl_0_laneRequest_decodeResult_divider <= 1'h0;
      slotControl_0_laneRequest_decodeResult_multiplier <= 1'h0;
      slotControl_0_laneRequest_decodeResult_shift <= 1'h0;
      slotControl_0_laneRequest_decodeResult_adder <= 1'h0;
      slotControl_0_laneRequest_decodeResult_logic <= 1'h0;
      slotControl_0_laneRequest_loadStore <= 1'h0;
      slotControl_0_laneRequest_issueInst <= 1'h0;
      slotControl_0_laneRequest_store <= 1'h0;
      slotControl_0_laneRequest_special <= 1'h0;
      slotControl_0_laneRequest_lsWholeReg <= 1'h0;
      slotControl_0_laneRequest_vs1 <= 5'h0;
      slotControl_0_laneRequest_vs2 <= 5'h0;
      slotControl_0_laneRequest_vd <= 5'h0;
      slotControl_0_laneRequest_loadStoreEEW <= 2'h0;
      slotControl_0_laneRequest_mask <= 1'h0;
      slotControl_0_laneRequest_segment <= 3'h0;
      slotControl_0_laneRequest_readFromScalar <= 32'h0;
      slotControl_0_laneRequest_csrInterface_vl <= 14'h0;
      slotControl_0_laneRequest_csrInterface_vStart <= 14'h0;
      slotControl_0_laneRequest_csrInterface_vlmul <= 3'h0;
      slotControl_0_laneRequest_csrInterface_vSew <= 2'h0;
      slotControl_0_laneRequest_csrInterface_vxrm <= 2'h0;
      slotControl_0_laneRequest_csrInterface_vta <= 1'h0;
      slotControl_0_laneRequest_csrInterface_vma <= 1'h0;
      slotControl_0_lastGroupForInstruction <= 10'h0;
      slotControl_0_isLastLaneForInstruction <= 1'h0;
      slotControl_0_additionalRW <= 1'h0;
      slotControl_0_instructionFinished <= 1'h0;
      slotControl_0_mask_valid <= 1'h0;
      slotControl_0_mask_bits <= 32'h0;
      slotControl_1_laneRequest_instructionIndex <= 3'h0;
      slotControl_1_laneRequest_decodeResult_specialSlot <= 1'h0;
      slotControl_1_laneRequest_decodeResult_topUop <= 5'h0;
      slotControl_1_laneRequest_decodeResult_popCount <= 1'h0;
      slotControl_1_laneRequest_decodeResult_ffo <= 1'h0;
      slotControl_1_laneRequest_decodeResult_average <= 1'h0;
      slotControl_1_laneRequest_decodeResult_reverse <= 1'h0;
      slotControl_1_laneRequest_decodeResult_dontNeedExecuteInLane <= 1'h0;
      slotControl_1_laneRequest_decodeResult_scheduler <= 1'h0;
      slotControl_1_laneRequest_decodeResult_sReadVD <= 1'h0;
      slotControl_1_laneRequest_decodeResult_vtype <= 1'h0;
      slotControl_1_laneRequest_decodeResult_sWrite <= 1'h0;
      slotControl_1_laneRequest_decodeResult_crossRead <= 1'h0;
      slotControl_1_laneRequest_decodeResult_crossWrite <= 1'h0;
      slotControl_1_laneRequest_decodeResult_maskUnit <= 1'h0;
      slotControl_1_laneRequest_decodeResult_special <= 1'h0;
      slotControl_1_laneRequest_decodeResult_saturate <= 1'h0;
      slotControl_1_laneRequest_decodeResult_vwmacc <= 1'h0;
      slotControl_1_laneRequest_decodeResult_readOnly <= 1'h0;
      slotControl_1_laneRequest_decodeResult_maskSource <= 1'h0;
      slotControl_1_laneRequest_decodeResult_maskDestination <= 1'h0;
      slotControl_1_laneRequest_decodeResult_maskLogic <= 1'h0;
      slotControl_1_laneRequest_decodeResult_uop <= 4'h0;
      slotControl_1_laneRequest_decodeResult_iota <= 1'h0;
      slotControl_1_laneRequest_decodeResult_mv <= 1'h0;
      slotControl_1_laneRequest_decodeResult_extend <= 1'h0;
      slotControl_1_laneRequest_decodeResult_unOrderWrite <= 1'h0;
      slotControl_1_laneRequest_decodeResult_compress <= 1'h0;
      slotControl_1_laneRequest_decodeResult_gather16 <= 1'h0;
      slotControl_1_laneRequest_decodeResult_gather <= 1'h0;
      slotControl_1_laneRequest_decodeResult_slid <= 1'h0;
      slotControl_1_laneRequest_decodeResult_targetRd <= 1'h0;
      slotControl_1_laneRequest_decodeResult_widenReduce <= 1'h0;
      slotControl_1_laneRequest_decodeResult_red <= 1'h0;
      slotControl_1_laneRequest_decodeResult_nr <= 1'h0;
      slotControl_1_laneRequest_decodeResult_itype <= 1'h0;
      slotControl_1_laneRequest_decodeResult_unsigned1 <= 1'h0;
      slotControl_1_laneRequest_decodeResult_unsigned0 <= 1'h0;
      slotControl_1_laneRequest_decodeResult_other <= 1'h0;
      slotControl_1_laneRequest_decodeResult_multiCycle <= 1'h0;
      slotControl_1_laneRequest_decodeResult_divider <= 1'h0;
      slotControl_1_laneRequest_decodeResult_multiplier <= 1'h0;
      slotControl_1_laneRequest_decodeResult_shift <= 1'h0;
      slotControl_1_laneRequest_decodeResult_adder <= 1'h0;
      slotControl_1_laneRequest_decodeResult_logic <= 1'h0;
      slotControl_1_laneRequest_loadStore <= 1'h0;
      slotControl_1_laneRequest_issueInst <= 1'h0;
      slotControl_1_laneRequest_store <= 1'h0;
      slotControl_1_laneRequest_special <= 1'h0;
      slotControl_1_laneRequest_lsWholeReg <= 1'h0;
      slotControl_1_laneRequest_vs1 <= 5'h0;
      slotControl_1_laneRequest_vs2 <= 5'h0;
      slotControl_1_laneRequest_vd <= 5'h0;
      slotControl_1_laneRequest_loadStoreEEW <= 2'h0;
      slotControl_1_laneRequest_mask <= 1'h0;
      slotControl_1_laneRequest_segment <= 3'h0;
      slotControl_1_laneRequest_readFromScalar <= 32'h0;
      slotControl_1_laneRequest_csrInterface_vl <= 14'h0;
      slotControl_1_laneRequest_csrInterface_vStart <= 14'h0;
      slotControl_1_laneRequest_csrInterface_vlmul <= 3'h0;
      slotControl_1_laneRequest_csrInterface_vSew <= 2'h0;
      slotControl_1_laneRequest_csrInterface_vxrm <= 2'h0;
      slotControl_1_laneRequest_csrInterface_vta <= 1'h0;
      slotControl_1_laneRequest_csrInterface_vma <= 1'h0;
      slotControl_1_lastGroupForInstruction <= 10'h0;
      slotControl_1_isLastLaneForInstruction <= 1'h0;
      slotControl_1_additionalRW <= 1'h0;
      slotControl_1_instructionFinished <= 1'h0;
      slotControl_1_mask_valid <= 1'h0;
      slotControl_1_mask_bits <= 32'h0;
      slotControl_2_laneRequest_instructionIndex <= 3'h0;
      slotControl_2_laneRequest_decodeResult_specialSlot <= 1'h0;
      slotControl_2_laneRequest_decodeResult_topUop <= 5'h0;
      slotControl_2_laneRequest_decodeResult_popCount <= 1'h0;
      slotControl_2_laneRequest_decodeResult_ffo <= 1'h0;
      slotControl_2_laneRequest_decodeResult_average <= 1'h0;
      slotControl_2_laneRequest_decodeResult_reverse <= 1'h0;
      slotControl_2_laneRequest_decodeResult_dontNeedExecuteInLane <= 1'h0;
      slotControl_2_laneRequest_decodeResult_scheduler <= 1'h0;
      slotControl_2_laneRequest_decodeResult_sReadVD <= 1'h0;
      slotControl_2_laneRequest_decodeResult_vtype <= 1'h0;
      slotControl_2_laneRequest_decodeResult_sWrite <= 1'h0;
      slotControl_2_laneRequest_decodeResult_crossRead <= 1'h0;
      slotControl_2_laneRequest_decodeResult_crossWrite <= 1'h0;
      slotControl_2_laneRequest_decodeResult_maskUnit <= 1'h0;
      slotControl_2_laneRequest_decodeResult_special <= 1'h0;
      slotControl_2_laneRequest_decodeResult_saturate <= 1'h0;
      slotControl_2_laneRequest_decodeResult_vwmacc <= 1'h0;
      slotControl_2_laneRequest_decodeResult_readOnly <= 1'h0;
      slotControl_2_laneRequest_decodeResult_maskSource <= 1'h0;
      slotControl_2_laneRequest_decodeResult_maskDestination <= 1'h0;
      slotControl_2_laneRequest_decodeResult_maskLogic <= 1'h0;
      slotControl_2_laneRequest_decodeResult_uop <= 4'h0;
      slotControl_2_laneRequest_decodeResult_iota <= 1'h0;
      slotControl_2_laneRequest_decodeResult_mv <= 1'h0;
      slotControl_2_laneRequest_decodeResult_extend <= 1'h0;
      slotControl_2_laneRequest_decodeResult_unOrderWrite <= 1'h0;
      slotControl_2_laneRequest_decodeResult_compress <= 1'h0;
      slotControl_2_laneRequest_decodeResult_gather16 <= 1'h0;
      slotControl_2_laneRequest_decodeResult_gather <= 1'h0;
      slotControl_2_laneRequest_decodeResult_slid <= 1'h0;
      slotControl_2_laneRequest_decodeResult_targetRd <= 1'h0;
      slotControl_2_laneRequest_decodeResult_widenReduce <= 1'h0;
      slotControl_2_laneRequest_decodeResult_red <= 1'h0;
      slotControl_2_laneRequest_decodeResult_nr <= 1'h0;
      slotControl_2_laneRequest_decodeResult_itype <= 1'h0;
      slotControl_2_laneRequest_decodeResult_unsigned1 <= 1'h0;
      slotControl_2_laneRequest_decodeResult_unsigned0 <= 1'h0;
      slotControl_2_laneRequest_decodeResult_other <= 1'h0;
      slotControl_2_laneRequest_decodeResult_multiCycle <= 1'h0;
      slotControl_2_laneRequest_decodeResult_divider <= 1'h0;
      slotControl_2_laneRequest_decodeResult_multiplier <= 1'h0;
      slotControl_2_laneRequest_decodeResult_shift <= 1'h0;
      slotControl_2_laneRequest_decodeResult_adder <= 1'h0;
      slotControl_2_laneRequest_decodeResult_logic <= 1'h0;
      slotControl_2_laneRequest_loadStore <= 1'h0;
      slotControl_2_laneRequest_issueInst <= 1'h0;
      slotControl_2_laneRequest_store <= 1'h0;
      slotControl_2_laneRequest_special <= 1'h0;
      slotControl_2_laneRequest_lsWholeReg <= 1'h0;
      slotControl_2_laneRequest_vs1 <= 5'h0;
      slotControl_2_laneRequest_vs2 <= 5'h0;
      slotControl_2_laneRequest_vd <= 5'h0;
      slotControl_2_laneRequest_loadStoreEEW <= 2'h0;
      slotControl_2_laneRequest_mask <= 1'h0;
      slotControl_2_laneRequest_segment <= 3'h0;
      slotControl_2_laneRequest_readFromScalar <= 32'h0;
      slotControl_2_laneRequest_csrInterface_vl <= 14'h0;
      slotControl_2_laneRequest_csrInterface_vStart <= 14'h0;
      slotControl_2_laneRequest_csrInterface_vlmul <= 3'h0;
      slotControl_2_laneRequest_csrInterface_vSew <= 2'h0;
      slotControl_2_laneRequest_csrInterface_vxrm <= 2'h0;
      slotControl_2_laneRequest_csrInterface_vta <= 1'h0;
      slotControl_2_laneRequest_csrInterface_vma <= 1'h0;
      slotControl_2_lastGroupForInstruction <= 10'h0;
      slotControl_2_isLastLaneForInstruction <= 1'h0;
      slotControl_2_additionalRW <= 1'h0;
      slotControl_2_instructionFinished <= 1'h0;
      slotControl_2_mask_valid <= 1'h0;
      slotControl_2_mask_bits <= 32'h0;
      slotControl_3_laneRequest_instructionIndex <= 3'h0;
      slotControl_3_laneRequest_decodeResult_specialSlot <= 1'h0;
      slotControl_3_laneRequest_decodeResult_topUop <= 5'h0;
      slotControl_3_laneRequest_decodeResult_popCount <= 1'h0;
      slotControl_3_laneRequest_decodeResult_ffo <= 1'h0;
      slotControl_3_laneRequest_decodeResult_average <= 1'h0;
      slotControl_3_laneRequest_decodeResult_reverse <= 1'h0;
      slotControl_3_laneRequest_decodeResult_dontNeedExecuteInLane <= 1'h0;
      slotControl_3_laneRequest_decodeResult_scheduler <= 1'h0;
      slotControl_3_laneRequest_decodeResult_sReadVD <= 1'h0;
      slotControl_3_laneRequest_decodeResult_vtype <= 1'h0;
      slotControl_3_laneRequest_decodeResult_sWrite <= 1'h0;
      slotControl_3_laneRequest_decodeResult_crossRead <= 1'h0;
      slotControl_3_laneRequest_decodeResult_crossWrite <= 1'h0;
      slotControl_3_laneRequest_decodeResult_maskUnit <= 1'h0;
      slotControl_3_laneRequest_decodeResult_special <= 1'h0;
      slotControl_3_laneRequest_decodeResult_saturate <= 1'h0;
      slotControl_3_laneRequest_decodeResult_vwmacc <= 1'h0;
      slotControl_3_laneRequest_decodeResult_readOnly <= 1'h0;
      slotControl_3_laneRequest_decodeResult_maskSource <= 1'h0;
      slotControl_3_laneRequest_decodeResult_maskDestination <= 1'h0;
      slotControl_3_laneRequest_decodeResult_maskLogic <= 1'h0;
      slotControl_3_laneRequest_decodeResult_uop <= 4'h0;
      slotControl_3_laneRequest_decodeResult_iota <= 1'h0;
      slotControl_3_laneRequest_decodeResult_mv <= 1'h0;
      slotControl_3_laneRequest_decodeResult_extend <= 1'h0;
      slotControl_3_laneRequest_decodeResult_unOrderWrite <= 1'h0;
      slotControl_3_laneRequest_decodeResult_compress <= 1'h0;
      slotControl_3_laneRequest_decodeResult_gather16 <= 1'h0;
      slotControl_3_laneRequest_decodeResult_gather <= 1'h0;
      slotControl_3_laneRequest_decodeResult_slid <= 1'h0;
      slotControl_3_laneRequest_decodeResult_targetRd <= 1'h0;
      slotControl_3_laneRequest_decodeResult_widenReduce <= 1'h0;
      slotControl_3_laneRequest_decodeResult_red <= 1'h0;
      slotControl_3_laneRequest_decodeResult_nr <= 1'h0;
      slotControl_3_laneRequest_decodeResult_itype <= 1'h0;
      slotControl_3_laneRequest_decodeResult_unsigned1 <= 1'h0;
      slotControl_3_laneRequest_decodeResult_unsigned0 <= 1'h0;
      slotControl_3_laneRequest_decodeResult_other <= 1'h0;
      slotControl_3_laneRequest_decodeResult_multiCycle <= 1'h0;
      slotControl_3_laneRequest_decodeResult_divider <= 1'h0;
      slotControl_3_laneRequest_decodeResult_multiplier <= 1'h0;
      slotControl_3_laneRequest_decodeResult_shift <= 1'h0;
      slotControl_3_laneRequest_decodeResult_adder <= 1'h0;
      slotControl_3_laneRequest_decodeResult_logic <= 1'h0;
      slotControl_3_laneRequest_loadStore <= 1'h0;
      slotControl_3_laneRequest_issueInst <= 1'h0;
      slotControl_3_laneRequest_store <= 1'h0;
      slotControl_3_laneRequest_special <= 1'h0;
      slotControl_3_laneRequest_lsWholeReg <= 1'h0;
      slotControl_3_laneRequest_vs1 <= 5'h0;
      slotControl_3_laneRequest_vs2 <= 5'h0;
      slotControl_3_laneRequest_vd <= 5'h0;
      slotControl_3_laneRequest_loadStoreEEW <= 2'h0;
      slotControl_3_laneRequest_mask <= 1'h0;
      slotControl_3_laneRequest_segment <= 3'h0;
      slotControl_3_laneRequest_readFromScalar <= 32'h0;
      slotControl_3_laneRequest_csrInterface_vl <= 14'h0;
      slotControl_3_laneRequest_csrInterface_vStart <= 14'h0;
      slotControl_3_laneRequest_csrInterface_vlmul <= 3'h0;
      slotControl_3_laneRequest_csrInterface_vSew <= 2'h0;
      slotControl_3_laneRequest_csrInterface_vxrm <= 2'h0;
      slotControl_3_laneRequest_csrInterface_vta <= 1'h0;
      slotControl_3_laneRequest_csrInterface_vma <= 1'h0;
      slotControl_3_lastGroupForInstruction <= 10'h0;
      slotControl_3_isLastLaneForInstruction <= 1'h0;
      slotControl_3_additionalRW <= 1'h0;
      slotControl_3_instructionFinished <= 1'h0;
      slotControl_3_mask_valid <= 1'h0;
      slotControl_3_mask_bits <= 32'h0;
      instructionValidNext <= 8'h0;
      vxsatResult <= 8'h0;
      tokenReg <= 3'h0;
      tokenReg_1 <= 3'h0;
      tokenReg_2 <= 3'h0;
      tokenReg_3 <= 3'h0;
      queueBeforeMaskWrite_empty <= 1'h1;
      emptyInstValid <= 1'h0;
    end
    else begin
      slotOccupied_0 <= slotEnqueueFire_0 ^ slotDequeueFire_0 ? slotEnqueueFire_0 : ~(_maskFailure_T & _stage0_updateLaneState_outOfExecutionRange) & slotOccupied_0;
      slotOccupied_1 <= slotEnqueueFire_1 ^ slotEnqueueFire_0 ? slotEnqueueFire_1 : ~(_maskFailure_T_1 & _stage0_1_updateLaneState_outOfExecutionRange) & slotOccupied_1;
      slotOccupied_2 <= slotEnqueueFire_2 ^ slotEnqueueFire_1 ? slotEnqueueFire_2 : ~(_maskFailure_T_2 & _stage0_2_updateLaneState_outOfExecutionRange) & slotOccupied_2;
      slotOccupied_3 <= slotEnqueueFire_3 ^ slotEnqueueFire_2 ? slotEnqueueFire_3 : ~(_maskFailure_T_3 & _stage0_3_updateLaneState_outOfExecutionRange) & slotOccupied_3;
      if (enqueueFire) begin
        maskGroupCountVec_0 <= maskGroupCountVec_1;
        maskIndexVec_0 <= maskIndexVec_1;
        slotControl_0_laneRequest_instructionIndex <= slotControl_1_laneRequest_instructionIndex;
        slotControl_0_laneRequest_decodeResult_specialSlot <= slotControl_1_laneRequest_decodeResult_specialSlot;
        slotControl_0_laneRequest_decodeResult_topUop <= slotControl_1_laneRequest_decodeResult_topUop;
        slotControl_0_laneRequest_decodeResult_popCount <= slotControl_1_laneRequest_decodeResult_popCount;
        slotControl_0_laneRequest_decodeResult_ffo <= slotControl_1_laneRequest_decodeResult_ffo;
        slotControl_0_laneRequest_decodeResult_average <= slotControl_1_laneRequest_decodeResult_average;
        slotControl_0_laneRequest_decodeResult_reverse <= slotControl_1_laneRequest_decodeResult_reverse;
        slotControl_0_laneRequest_decodeResult_dontNeedExecuteInLane <= slotControl_1_laneRequest_decodeResult_dontNeedExecuteInLane;
        slotControl_0_laneRequest_decodeResult_scheduler <= slotControl_1_laneRequest_decodeResult_scheduler;
        slotControl_0_laneRequest_decodeResult_sReadVD <= slotControl_1_laneRequest_decodeResult_sReadVD;
        slotControl_0_laneRequest_decodeResult_vtype <= slotControl_1_laneRequest_decodeResult_vtype;
        slotControl_0_laneRequest_decodeResult_sWrite <= slotControl_1_laneRequest_decodeResult_sWrite;
        slotControl_0_laneRequest_decodeResult_crossRead <= slotControl_1_laneRequest_decodeResult_crossRead;
        slotControl_0_laneRequest_decodeResult_crossWrite <= slotControl_1_laneRequest_decodeResult_crossWrite;
        slotControl_0_laneRequest_decodeResult_maskUnit <= slotControl_1_laneRequest_decodeResult_maskUnit;
        slotControl_0_laneRequest_decodeResult_special <= slotControl_1_laneRequest_decodeResult_special;
        slotControl_0_laneRequest_decodeResult_saturate <= slotControl_1_laneRequest_decodeResult_saturate;
        slotControl_0_laneRequest_decodeResult_vwmacc <= slotControl_1_laneRequest_decodeResult_vwmacc;
        slotControl_0_laneRequest_decodeResult_readOnly <= slotControl_1_laneRequest_decodeResult_readOnly;
        slotControl_0_laneRequest_decodeResult_maskSource <= slotControl_1_laneRequest_decodeResult_maskSource;
        slotControl_0_laneRequest_decodeResult_maskDestination <= slotControl_1_laneRequest_decodeResult_maskDestination;
        slotControl_0_laneRequest_decodeResult_maskLogic <= slotControl_1_laneRequest_decodeResult_maskLogic;
        slotControl_0_laneRequest_decodeResult_uop <= slotControl_1_laneRequest_decodeResult_uop;
        slotControl_0_laneRequest_decodeResult_iota <= slotControl_1_laneRequest_decodeResult_iota;
        slotControl_0_laneRequest_decodeResult_mv <= slotControl_1_laneRequest_decodeResult_mv;
        slotControl_0_laneRequest_decodeResult_extend <= slotControl_1_laneRequest_decodeResult_extend;
        slotControl_0_laneRequest_decodeResult_unOrderWrite <= slotControl_1_laneRequest_decodeResult_unOrderWrite;
        slotControl_0_laneRequest_decodeResult_compress <= slotControl_1_laneRequest_decodeResult_compress;
        slotControl_0_laneRequest_decodeResult_gather16 <= slotControl_1_laneRequest_decodeResult_gather16;
        slotControl_0_laneRequest_decodeResult_gather <= slotControl_1_laneRequest_decodeResult_gather;
        slotControl_0_laneRequest_decodeResult_slid <= slotControl_1_laneRequest_decodeResult_slid;
        slotControl_0_laneRequest_decodeResult_targetRd <= slotControl_1_laneRequest_decodeResult_targetRd;
        slotControl_0_laneRequest_decodeResult_widenReduce <= slotControl_1_laneRequest_decodeResult_widenReduce;
        slotControl_0_laneRequest_decodeResult_red <= slotControl_1_laneRequest_decodeResult_red;
        slotControl_0_laneRequest_decodeResult_nr <= slotControl_1_laneRequest_decodeResult_nr;
        slotControl_0_laneRequest_decodeResult_itype <= slotControl_1_laneRequest_decodeResult_itype;
        slotControl_0_laneRequest_decodeResult_unsigned1 <= slotControl_1_laneRequest_decodeResult_unsigned1;
        slotControl_0_laneRequest_decodeResult_unsigned0 <= slotControl_1_laneRequest_decodeResult_unsigned0;
        slotControl_0_laneRequest_decodeResult_other <= slotControl_1_laneRequest_decodeResult_other;
        slotControl_0_laneRequest_decodeResult_multiCycle <= slotControl_1_laneRequest_decodeResult_multiCycle;
        slotControl_0_laneRequest_decodeResult_divider <= slotControl_1_laneRequest_decodeResult_divider;
        slotControl_0_laneRequest_decodeResult_multiplier <= slotControl_1_laneRequest_decodeResult_multiplier;
        slotControl_0_laneRequest_decodeResult_shift <= slotControl_1_laneRequest_decodeResult_shift;
        slotControl_0_laneRequest_decodeResult_adder <= slotControl_1_laneRequest_decodeResult_adder;
        slotControl_0_laneRequest_decodeResult_logic <= slotControl_1_laneRequest_decodeResult_logic;
        slotControl_0_laneRequest_loadStore <= slotControl_1_laneRequest_loadStore;
        slotControl_0_laneRequest_issueInst <= slotControl_1_laneRequest_issueInst;
        slotControl_0_laneRequest_store <= slotControl_1_laneRequest_store;
        slotControl_0_laneRequest_special <= slotControl_1_laneRequest_special;
        slotControl_0_laneRequest_lsWholeReg <= slotControl_1_laneRequest_lsWholeReg;
        slotControl_0_laneRequest_vs1 <= slotControl_1_laneRequest_vs1;
        slotControl_0_laneRequest_vs2 <= slotControl_1_laneRequest_vs2;
        slotControl_0_laneRequest_vd <= slotControl_1_laneRequest_vd;
        slotControl_0_laneRequest_loadStoreEEW <= slotControl_1_laneRequest_loadStoreEEW;
        slotControl_0_laneRequest_mask <= slotControl_1_laneRequest_mask;
        slotControl_0_laneRequest_segment <= slotControl_1_laneRequest_segment;
        slotControl_0_laneRequest_readFromScalar <= slotControl_1_laneRequest_readFromScalar;
        slotControl_0_laneRequest_csrInterface_vl <= slotControl_1_laneRequest_csrInterface_vl;
        slotControl_0_laneRequest_csrInterface_vStart <= slotControl_1_laneRequest_csrInterface_vStart;
        slotControl_0_laneRequest_csrInterface_vlmul <= slotControl_1_laneRequest_csrInterface_vlmul;
        slotControl_0_laneRequest_csrInterface_vSew <= slotControl_1_laneRequest_csrInterface_vSew;
        slotControl_0_laneRequest_csrInterface_vxrm <= slotControl_1_laneRequest_csrInterface_vxrm;
        slotControl_0_laneRequest_csrInterface_vta <= slotControl_1_laneRequest_csrInterface_vta;
        slotControl_0_laneRequest_csrInterface_vma <= slotControl_1_laneRequest_csrInterface_vma;
        slotControl_0_lastGroupForInstruction <= slotControl_1_lastGroupForInstruction;
        slotControl_0_isLastLaneForInstruction <= slotControl_1_isLastLaneForInstruction;
        slotControl_0_additionalRW <= slotControl_1_additionalRW;
        slotControl_0_instructionFinished <= slotControl_1_instructionFinished;
        slotControl_0_mask_valid <= slotControl_1_mask_valid;
        slotControl_0_mask_bits <= slotControl_1_mask_bits;
      end
      else begin
        if (_maskFailure_T) begin
          maskGroupCountVec_0 <= _stage0_updateLaneState_maskGroupCount;
          maskIndexVec_0 <= _stage0_updateLaneState_maskIndex;
        end
        if (maskUpdateFire ^ maskFailure)
          slotControl_0_mask_valid <= maskUpdateFire;
        if (maskUpdateFire)
          slotControl_0_mask_bits <= maskDataVec_0;
      end
      if (enqueueFire_1) begin
        maskGroupCountVec_1 <= maskGroupCountVec_2;
        maskIndexVec_1 <= maskIndexVec_2;
        slotControl_1_laneRequest_instructionIndex <= slotControl_2_laneRequest_instructionIndex;
        slotControl_1_laneRequest_decodeResult_specialSlot <= slotControl_2_laneRequest_decodeResult_specialSlot;
        slotControl_1_laneRequest_decodeResult_topUop <= slotControl_2_laneRequest_decodeResult_topUop;
        slotControl_1_laneRequest_decodeResult_popCount <= slotControl_2_laneRequest_decodeResult_popCount;
        slotControl_1_laneRequest_decodeResult_ffo <= slotControl_2_laneRequest_decodeResult_ffo;
        slotControl_1_laneRequest_decodeResult_average <= slotControl_2_laneRequest_decodeResult_average;
        slotControl_1_laneRequest_decodeResult_reverse <= slotControl_2_laneRequest_decodeResult_reverse;
        slotControl_1_laneRequest_decodeResult_dontNeedExecuteInLane <= slotControl_2_laneRequest_decodeResult_dontNeedExecuteInLane;
        slotControl_1_laneRequest_decodeResult_scheduler <= slotControl_2_laneRequest_decodeResult_scheduler;
        slotControl_1_laneRequest_decodeResult_sReadVD <= slotControl_2_laneRequest_decodeResult_sReadVD;
        slotControl_1_laneRequest_decodeResult_vtype <= slotControl_2_laneRequest_decodeResult_vtype;
        slotControl_1_laneRequest_decodeResult_sWrite <= slotControl_2_laneRequest_decodeResult_sWrite;
        slotControl_1_laneRequest_decodeResult_crossRead <= slotControl_2_laneRequest_decodeResult_crossRead;
        slotControl_1_laneRequest_decodeResult_crossWrite <= slotControl_2_laneRequest_decodeResult_crossWrite;
        slotControl_1_laneRequest_decodeResult_maskUnit <= slotControl_2_laneRequest_decodeResult_maskUnit;
        slotControl_1_laneRequest_decodeResult_special <= slotControl_2_laneRequest_decodeResult_special;
        slotControl_1_laneRequest_decodeResult_saturate <= slotControl_2_laneRequest_decodeResult_saturate;
        slotControl_1_laneRequest_decodeResult_vwmacc <= slotControl_2_laneRequest_decodeResult_vwmacc;
        slotControl_1_laneRequest_decodeResult_readOnly <= slotControl_2_laneRequest_decodeResult_readOnly;
        slotControl_1_laneRequest_decodeResult_maskSource <= slotControl_2_laneRequest_decodeResult_maskSource;
        slotControl_1_laneRequest_decodeResult_maskDestination <= slotControl_2_laneRequest_decodeResult_maskDestination;
        slotControl_1_laneRequest_decodeResult_maskLogic <= slotControl_2_laneRequest_decodeResult_maskLogic;
        slotControl_1_laneRequest_decodeResult_uop <= slotControl_2_laneRequest_decodeResult_uop;
        slotControl_1_laneRequest_decodeResult_iota <= slotControl_2_laneRequest_decodeResult_iota;
        slotControl_1_laneRequest_decodeResult_mv <= slotControl_2_laneRequest_decodeResult_mv;
        slotControl_1_laneRequest_decodeResult_extend <= slotControl_2_laneRequest_decodeResult_extend;
        slotControl_1_laneRequest_decodeResult_unOrderWrite <= slotControl_2_laneRequest_decodeResult_unOrderWrite;
        slotControl_1_laneRequest_decodeResult_compress <= slotControl_2_laneRequest_decodeResult_compress;
        slotControl_1_laneRequest_decodeResult_gather16 <= slotControl_2_laneRequest_decodeResult_gather16;
        slotControl_1_laneRequest_decodeResult_gather <= slotControl_2_laneRequest_decodeResult_gather;
        slotControl_1_laneRequest_decodeResult_slid <= slotControl_2_laneRequest_decodeResult_slid;
        slotControl_1_laneRequest_decodeResult_targetRd <= slotControl_2_laneRequest_decodeResult_targetRd;
        slotControl_1_laneRequest_decodeResult_widenReduce <= slotControl_2_laneRequest_decodeResult_widenReduce;
        slotControl_1_laneRequest_decodeResult_red <= slotControl_2_laneRequest_decodeResult_red;
        slotControl_1_laneRequest_decodeResult_nr <= slotControl_2_laneRequest_decodeResult_nr;
        slotControl_1_laneRequest_decodeResult_itype <= slotControl_2_laneRequest_decodeResult_itype;
        slotControl_1_laneRequest_decodeResult_unsigned1 <= slotControl_2_laneRequest_decodeResult_unsigned1;
        slotControl_1_laneRequest_decodeResult_unsigned0 <= slotControl_2_laneRequest_decodeResult_unsigned0;
        slotControl_1_laneRequest_decodeResult_other <= slotControl_2_laneRequest_decodeResult_other;
        slotControl_1_laneRequest_decodeResult_multiCycle <= slotControl_2_laneRequest_decodeResult_multiCycle;
        slotControl_1_laneRequest_decodeResult_divider <= slotControl_2_laneRequest_decodeResult_divider;
        slotControl_1_laneRequest_decodeResult_multiplier <= slotControl_2_laneRequest_decodeResult_multiplier;
        slotControl_1_laneRequest_decodeResult_shift <= slotControl_2_laneRequest_decodeResult_shift;
        slotControl_1_laneRequest_decodeResult_adder <= slotControl_2_laneRequest_decodeResult_adder;
        slotControl_1_laneRequest_decodeResult_logic <= slotControl_2_laneRequest_decodeResult_logic;
        slotControl_1_laneRequest_loadStore <= slotControl_2_laneRequest_loadStore;
        slotControl_1_laneRequest_issueInst <= slotControl_2_laneRequest_issueInst;
        slotControl_1_laneRequest_store <= slotControl_2_laneRequest_store;
        slotControl_1_laneRequest_special <= slotControl_2_laneRequest_special;
        slotControl_1_laneRequest_lsWholeReg <= slotControl_2_laneRequest_lsWholeReg;
        slotControl_1_laneRequest_vs1 <= slotControl_2_laneRequest_vs1;
        slotControl_1_laneRequest_vs2 <= slotControl_2_laneRequest_vs2;
        slotControl_1_laneRequest_vd <= slotControl_2_laneRequest_vd;
        slotControl_1_laneRequest_loadStoreEEW <= slotControl_2_laneRequest_loadStoreEEW;
        slotControl_1_laneRequest_mask <= slotControl_2_laneRequest_mask;
        slotControl_1_laneRequest_segment <= slotControl_2_laneRequest_segment;
        slotControl_1_laneRequest_readFromScalar <= slotControl_2_laneRequest_readFromScalar;
        slotControl_1_laneRequest_csrInterface_vl <= slotControl_2_laneRequest_csrInterface_vl;
        slotControl_1_laneRequest_csrInterface_vStart <= slotControl_2_laneRequest_csrInterface_vStart;
        slotControl_1_laneRequest_csrInterface_vlmul <= slotControl_2_laneRequest_csrInterface_vlmul;
        slotControl_1_laneRequest_csrInterface_vSew <= slotControl_2_laneRequest_csrInterface_vSew;
        slotControl_1_laneRequest_csrInterface_vxrm <= slotControl_2_laneRequest_csrInterface_vxrm;
        slotControl_1_laneRequest_csrInterface_vta <= slotControl_2_laneRequest_csrInterface_vta;
        slotControl_1_laneRequest_csrInterface_vma <= slotControl_2_laneRequest_csrInterface_vma;
        slotControl_1_lastGroupForInstruction <= slotControl_2_lastGroupForInstruction;
        slotControl_1_isLastLaneForInstruction <= slotControl_2_isLastLaneForInstruction;
        slotControl_1_additionalRW <= slotControl_2_additionalRW;
        slotControl_1_instructionFinished <= slotControl_2_instructionFinished;
        slotControl_1_mask_valid <= slotControl_2_mask_valid;
        slotControl_1_mask_bits <= slotControl_2_mask_bits;
      end
      else begin
        if (_maskFailure_T_1) begin
          maskGroupCountVec_1 <= _stage0_1_updateLaneState_maskGroupCount;
          maskIndexVec_1 <= _stage0_1_updateLaneState_maskIndex;
        end
        if (maskUpdateFire_1 ^ maskFailure_1)
          slotControl_1_mask_valid <= maskUpdateFire_1;
        if (maskUpdateFire_1)
          slotControl_1_mask_bits <= maskDataVec_1;
      end
      if (enqueueFire_2) begin
        maskGroupCountVec_2 <= maskGroupCountVec_3;
        maskIndexVec_2 <= maskIndexVec_3;
        slotControl_2_laneRequest_instructionIndex <= slotControl_3_laneRequest_instructionIndex;
        slotControl_2_laneRequest_decodeResult_specialSlot <= slotControl_3_laneRequest_decodeResult_specialSlot;
        slotControl_2_laneRequest_decodeResult_topUop <= slotControl_3_laneRequest_decodeResult_topUop;
        slotControl_2_laneRequest_decodeResult_popCount <= slotControl_3_laneRequest_decodeResult_popCount;
        slotControl_2_laneRequest_decodeResult_ffo <= slotControl_3_laneRequest_decodeResult_ffo;
        slotControl_2_laneRequest_decodeResult_average <= slotControl_3_laneRequest_decodeResult_average;
        slotControl_2_laneRequest_decodeResult_reverse <= slotControl_3_laneRequest_decodeResult_reverse;
        slotControl_2_laneRequest_decodeResult_dontNeedExecuteInLane <= slotControl_3_laneRequest_decodeResult_dontNeedExecuteInLane;
        slotControl_2_laneRequest_decodeResult_scheduler <= slotControl_3_laneRequest_decodeResult_scheduler;
        slotControl_2_laneRequest_decodeResult_sReadVD <= slotControl_3_laneRequest_decodeResult_sReadVD;
        slotControl_2_laneRequest_decodeResult_vtype <= slotControl_3_laneRequest_decodeResult_vtype;
        slotControl_2_laneRequest_decodeResult_sWrite <= slotControl_3_laneRequest_decodeResult_sWrite;
        slotControl_2_laneRequest_decodeResult_crossRead <= slotControl_3_laneRequest_decodeResult_crossRead;
        slotControl_2_laneRequest_decodeResult_crossWrite <= slotControl_3_laneRequest_decodeResult_crossWrite;
        slotControl_2_laneRequest_decodeResult_maskUnit <= slotControl_3_laneRequest_decodeResult_maskUnit;
        slotControl_2_laneRequest_decodeResult_special <= slotControl_3_laneRequest_decodeResult_special;
        slotControl_2_laneRequest_decodeResult_saturate <= slotControl_3_laneRequest_decodeResult_saturate;
        slotControl_2_laneRequest_decodeResult_vwmacc <= slotControl_3_laneRequest_decodeResult_vwmacc;
        slotControl_2_laneRequest_decodeResult_readOnly <= slotControl_3_laneRequest_decodeResult_readOnly;
        slotControl_2_laneRequest_decodeResult_maskSource <= slotControl_3_laneRequest_decodeResult_maskSource;
        slotControl_2_laneRequest_decodeResult_maskDestination <= slotControl_3_laneRequest_decodeResult_maskDestination;
        slotControl_2_laneRequest_decodeResult_maskLogic <= slotControl_3_laneRequest_decodeResult_maskLogic;
        slotControl_2_laneRequest_decodeResult_uop <= slotControl_3_laneRequest_decodeResult_uop;
        slotControl_2_laneRequest_decodeResult_iota <= slotControl_3_laneRequest_decodeResult_iota;
        slotControl_2_laneRequest_decodeResult_mv <= slotControl_3_laneRequest_decodeResult_mv;
        slotControl_2_laneRequest_decodeResult_extend <= slotControl_3_laneRequest_decodeResult_extend;
        slotControl_2_laneRequest_decodeResult_unOrderWrite <= slotControl_3_laneRequest_decodeResult_unOrderWrite;
        slotControl_2_laneRequest_decodeResult_compress <= slotControl_3_laneRequest_decodeResult_compress;
        slotControl_2_laneRequest_decodeResult_gather16 <= slotControl_3_laneRequest_decodeResult_gather16;
        slotControl_2_laneRequest_decodeResult_gather <= slotControl_3_laneRequest_decodeResult_gather;
        slotControl_2_laneRequest_decodeResult_slid <= slotControl_3_laneRequest_decodeResult_slid;
        slotControl_2_laneRequest_decodeResult_targetRd <= slotControl_3_laneRequest_decodeResult_targetRd;
        slotControl_2_laneRequest_decodeResult_widenReduce <= slotControl_3_laneRequest_decodeResult_widenReduce;
        slotControl_2_laneRequest_decodeResult_red <= slotControl_3_laneRequest_decodeResult_red;
        slotControl_2_laneRequest_decodeResult_nr <= slotControl_3_laneRequest_decodeResult_nr;
        slotControl_2_laneRequest_decodeResult_itype <= slotControl_3_laneRequest_decodeResult_itype;
        slotControl_2_laneRequest_decodeResult_unsigned1 <= slotControl_3_laneRequest_decodeResult_unsigned1;
        slotControl_2_laneRequest_decodeResult_unsigned0 <= slotControl_3_laneRequest_decodeResult_unsigned0;
        slotControl_2_laneRequest_decodeResult_other <= slotControl_3_laneRequest_decodeResult_other;
        slotControl_2_laneRequest_decodeResult_multiCycle <= slotControl_3_laneRequest_decodeResult_multiCycle;
        slotControl_2_laneRequest_decodeResult_divider <= slotControl_3_laneRequest_decodeResult_divider;
        slotControl_2_laneRequest_decodeResult_multiplier <= slotControl_3_laneRequest_decodeResult_multiplier;
        slotControl_2_laneRequest_decodeResult_shift <= slotControl_3_laneRequest_decodeResult_shift;
        slotControl_2_laneRequest_decodeResult_adder <= slotControl_3_laneRequest_decodeResult_adder;
        slotControl_2_laneRequest_decodeResult_logic <= slotControl_3_laneRequest_decodeResult_logic;
        slotControl_2_laneRequest_loadStore <= slotControl_3_laneRequest_loadStore;
        slotControl_2_laneRequest_issueInst <= slotControl_3_laneRequest_issueInst;
        slotControl_2_laneRequest_store <= slotControl_3_laneRequest_store;
        slotControl_2_laneRequest_special <= slotControl_3_laneRequest_special;
        slotControl_2_laneRequest_lsWholeReg <= slotControl_3_laneRequest_lsWholeReg;
        slotControl_2_laneRequest_vs1 <= slotControl_3_laneRequest_vs1;
        slotControl_2_laneRequest_vs2 <= slotControl_3_laneRequest_vs2;
        slotControl_2_laneRequest_vd <= slotControl_3_laneRequest_vd;
        slotControl_2_laneRequest_loadStoreEEW <= slotControl_3_laneRequest_loadStoreEEW;
        slotControl_2_laneRequest_mask <= slotControl_3_laneRequest_mask;
        slotControl_2_laneRequest_segment <= slotControl_3_laneRequest_segment;
        slotControl_2_laneRequest_readFromScalar <= slotControl_3_laneRequest_readFromScalar;
        slotControl_2_laneRequest_csrInterface_vl <= slotControl_3_laneRequest_csrInterface_vl;
        slotControl_2_laneRequest_csrInterface_vStart <= slotControl_3_laneRequest_csrInterface_vStart;
        slotControl_2_laneRequest_csrInterface_vlmul <= slotControl_3_laneRequest_csrInterface_vlmul;
        slotControl_2_laneRequest_csrInterface_vSew <= slotControl_3_laneRequest_csrInterface_vSew;
        slotControl_2_laneRequest_csrInterface_vxrm <= slotControl_3_laneRequest_csrInterface_vxrm;
        slotControl_2_laneRequest_csrInterface_vta <= slotControl_3_laneRequest_csrInterface_vta;
        slotControl_2_laneRequest_csrInterface_vma <= slotControl_3_laneRequest_csrInterface_vma;
        slotControl_2_lastGroupForInstruction <= slotControl_3_lastGroupForInstruction;
        slotControl_2_isLastLaneForInstruction <= slotControl_3_isLastLaneForInstruction;
        slotControl_2_additionalRW <= slotControl_3_additionalRW;
        slotControl_2_instructionFinished <= slotControl_3_instructionFinished;
        slotControl_2_mask_valid <= slotControl_3_mask_valid;
        slotControl_2_mask_bits <= slotControl_3_mask_bits;
      end
      else begin
        if (_maskFailure_T_2) begin
          maskGroupCountVec_2 <= _stage0_2_updateLaneState_maskGroupCount;
          maskIndexVec_2 <= _stage0_2_updateLaneState_maskIndex;
        end
        if (maskUpdateFire_2 ^ maskFailure_2)
          slotControl_2_mask_valid <= maskUpdateFire_2;
        if (maskUpdateFire_2)
          slotControl_2_mask_bits <= maskDataVec_2;
      end
      if (enqueueFire_3) begin
        maskGroupCountVec_3 <= 8'h0;
        maskIndexVec_3 <= 5'h0;
        slotControl_3_laneRequest_instructionIndex <= entranceControl_laneRequest_instructionIndex;
        slotControl_3_laneRequest_decodeResult_specialSlot <= entranceControl_laneRequest_decodeResult_specialSlot;
        slotControl_3_laneRequest_decodeResult_topUop <= entranceControl_laneRequest_decodeResult_topUop;
        slotControl_3_laneRequest_decodeResult_popCount <= entranceControl_laneRequest_decodeResult_popCount;
        slotControl_3_laneRequest_decodeResult_ffo <= entranceControl_laneRequest_decodeResult_ffo;
        slotControl_3_laneRequest_decodeResult_average <= entranceControl_laneRequest_decodeResult_average;
        slotControl_3_laneRequest_decodeResult_reverse <= entranceControl_laneRequest_decodeResult_reverse;
        slotControl_3_laneRequest_decodeResult_dontNeedExecuteInLane <= entranceControl_laneRequest_decodeResult_dontNeedExecuteInLane;
        slotControl_3_laneRequest_decodeResult_scheduler <= entranceControl_laneRequest_decodeResult_scheduler;
        slotControl_3_laneRequest_decodeResult_sReadVD <= entranceControl_laneRequest_decodeResult_sReadVD;
        slotControl_3_laneRequest_decodeResult_vtype <= entranceControl_laneRequest_decodeResult_vtype;
        slotControl_3_laneRequest_decodeResult_sWrite <= entranceControl_laneRequest_decodeResult_sWrite;
        slotControl_3_laneRequest_decodeResult_crossRead <= entranceControl_laneRequest_decodeResult_crossRead;
        slotControl_3_laneRequest_decodeResult_crossWrite <= entranceControl_laneRequest_decodeResult_crossWrite;
        slotControl_3_laneRequest_decodeResult_maskUnit <= entranceControl_laneRequest_decodeResult_maskUnit;
        slotControl_3_laneRequest_decodeResult_special <= entranceControl_laneRequest_decodeResult_special;
        slotControl_3_laneRequest_decodeResult_saturate <= entranceControl_laneRequest_decodeResult_saturate;
        slotControl_3_laneRequest_decodeResult_vwmacc <= entranceControl_laneRequest_decodeResult_vwmacc;
        slotControl_3_laneRequest_decodeResult_readOnly <= entranceControl_laneRequest_decodeResult_readOnly;
        slotControl_3_laneRequest_decodeResult_maskSource <= entranceControl_laneRequest_decodeResult_maskSource;
        slotControl_3_laneRequest_decodeResult_maskDestination <= entranceControl_laneRequest_decodeResult_maskDestination;
        slotControl_3_laneRequest_decodeResult_maskLogic <= entranceControl_laneRequest_decodeResult_maskLogic;
        slotControl_3_laneRequest_decodeResult_uop <= entranceControl_laneRequest_decodeResult_uop;
        slotControl_3_laneRequest_decodeResult_iota <= entranceControl_laneRequest_decodeResult_iota;
        slotControl_3_laneRequest_decodeResult_mv <= entranceControl_laneRequest_decodeResult_mv;
        slotControl_3_laneRequest_decodeResult_extend <= entranceControl_laneRequest_decodeResult_extend;
        slotControl_3_laneRequest_decodeResult_unOrderWrite <= entranceControl_laneRequest_decodeResult_unOrderWrite;
        slotControl_3_laneRequest_decodeResult_compress <= entranceControl_laneRequest_decodeResult_compress;
        slotControl_3_laneRequest_decodeResult_gather16 <= entranceControl_laneRequest_decodeResult_gather16;
        slotControl_3_laneRequest_decodeResult_gather <= entranceControl_laneRequest_decodeResult_gather;
        slotControl_3_laneRequest_decodeResult_slid <= entranceControl_laneRequest_decodeResult_slid;
        slotControl_3_laneRequest_decodeResult_targetRd <= entranceControl_laneRequest_decodeResult_targetRd;
        slotControl_3_laneRequest_decodeResult_widenReduce <= entranceControl_laneRequest_decodeResult_widenReduce;
        slotControl_3_laneRequest_decodeResult_red <= entranceControl_laneRequest_decodeResult_red;
        slotControl_3_laneRequest_decodeResult_nr <= entranceControl_laneRequest_decodeResult_nr;
        slotControl_3_laneRequest_decodeResult_itype <= entranceControl_laneRequest_decodeResult_itype;
        slotControl_3_laneRequest_decodeResult_unsigned1 <= entranceControl_laneRequest_decodeResult_unsigned1;
        slotControl_3_laneRequest_decodeResult_unsigned0 <= entranceControl_laneRequest_decodeResult_unsigned0;
        slotControl_3_laneRequest_decodeResult_other <= entranceControl_laneRequest_decodeResult_other;
        slotControl_3_laneRequest_decodeResult_multiCycle <= entranceControl_laneRequest_decodeResult_multiCycle;
        slotControl_3_laneRequest_decodeResult_divider <= entranceControl_laneRequest_decodeResult_divider;
        slotControl_3_laneRequest_decodeResult_multiplier <= entranceControl_laneRequest_decodeResult_multiplier;
        slotControl_3_laneRequest_decodeResult_shift <= entranceControl_laneRequest_decodeResult_shift;
        slotControl_3_laneRequest_decodeResult_adder <= entranceControl_laneRequest_decodeResult_adder;
        slotControl_3_laneRequest_decodeResult_logic <= entranceControl_laneRequest_decodeResult_logic;
        slotControl_3_laneRequest_loadStore <= entranceControl_laneRequest_loadStore;
        slotControl_3_laneRequest_issueInst <= entranceControl_laneRequest_issueInst;
        slotControl_3_laneRequest_store <= entranceControl_laneRequest_store;
        slotControl_3_laneRequest_special <= entranceControl_laneRequest_special;
        slotControl_3_laneRequest_lsWholeReg <= entranceControl_laneRequest_lsWholeReg;
        slotControl_3_laneRequest_vs1 <= entranceControl_laneRequest_vs1;
        slotControl_3_laneRequest_vs2 <= entranceControl_laneRequest_vs2;
        slotControl_3_laneRequest_vd <= entranceControl_laneRequest_vd;
        slotControl_3_laneRequest_loadStoreEEW <= entranceControl_laneRequest_loadStoreEEW;
        slotControl_3_laneRequest_mask <= entranceControl_laneRequest_mask;
        slotControl_3_laneRequest_segment <= entranceControl_laneRequest_segment;
        slotControl_3_laneRequest_readFromScalar <= entranceControl_laneRequest_readFromScalar;
        slotControl_3_laneRequest_csrInterface_vl <= entranceControl_laneRequest_csrInterface_vl;
        slotControl_3_laneRequest_csrInterface_vStart <= entranceControl_laneRequest_csrInterface_vStart;
        slotControl_3_laneRequest_csrInterface_vlmul <= entranceControl_laneRequest_csrInterface_vlmul;
        slotControl_3_laneRequest_csrInterface_vSew <= entranceControl_laneRequest_csrInterface_vSew;
        slotControl_3_laneRequest_csrInterface_vxrm <= entranceControl_laneRequest_csrInterface_vxrm;
        slotControl_3_laneRequest_csrInterface_vta <= entranceControl_laneRequest_csrInterface_vta;
        slotControl_3_laneRequest_csrInterface_vma <= entranceControl_laneRequest_csrInterface_vma;
        slotControl_3_lastGroupForInstruction <= entranceControl_lastGroupForInstruction;
        slotControl_3_isLastLaneForInstruction <= entranceControl_isLastLaneForInstruction;
        slotControl_3_additionalRW <= entranceControl_additionalRW;
        slotControl_3_instructionFinished <= entranceControl_instructionFinished;
        slotControl_3_mask_bits <= 32'h0;
      end
      else begin
        if (_maskFailure_T_3) begin
          maskGroupCountVec_3 <= _stage0_3_updateLaneState_maskGroupCount;
          maskIndexVec_3 <= _stage0_3_updateLaneState_maskIndex;
        end
        if (maskUpdateFire_3)
          slotControl_3_mask_bits <= maskDataVec_3;
      end
      if (enqFire) begin
        allVrfWriteAfterCheck_0_vd <= vrfWriteArbiter_0_bits_vd;
        allVrfWriteAfterCheck_0_offset <= vrfWriteArbiter_0_bits_offset;
        allVrfWriteAfterCheck_0_mask <= vrfWriteArbiter_0_bits_mask;
        allVrfWriteAfterCheck_0_data <= vrfWriteArbiter_0_bits_data;
        allVrfWriteAfterCheck_0_last <= vrfWriteArbiter_0_bits_last;
        allVrfWriteAfterCheck_0_instructionIndex <= vrfWriteArbiter_0_bits_instructionIndex;
      end
      if (enqFire_1) begin
        allVrfWriteAfterCheck_1_vd <= vrfWriteArbiter_1_bits_vd;
        allVrfWriteAfterCheck_1_offset <= vrfWriteArbiter_1_bits_offset;
        allVrfWriteAfterCheck_1_mask <= vrfWriteArbiter_1_bits_mask;
        allVrfWriteAfterCheck_1_data <= vrfWriteArbiter_1_bits_data;
        allVrfWriteAfterCheck_1_last <= vrfWriteArbiter_1_bits_last;
        allVrfWriteAfterCheck_1_instructionIndex <= vrfWriteArbiter_1_bits_instructionIndex;
      end
      if (enqFire_2) begin
        allVrfWriteAfterCheck_2_vd <= vrfWriteArbiter_2_bits_vd;
        allVrfWriteAfterCheck_2_offset <= vrfWriteArbiter_2_bits_offset;
        allVrfWriteAfterCheck_2_mask <= vrfWriteArbiter_2_bits_mask;
        allVrfWriteAfterCheck_2_data <= vrfWriteArbiter_2_bits_data;
        allVrfWriteAfterCheck_2_last <= vrfWriteArbiter_2_bits_last;
        allVrfWriteAfterCheck_2_instructionIndex <= vrfWriteArbiter_2_bits_instructionIndex;
      end
      if (enqFire_3) begin
        allVrfWriteAfterCheck_3_vd <= vrfWriteArbiter_3_bits_vd;
        allVrfWriteAfterCheck_3_offset <= vrfWriteArbiter_3_bits_offset;
        allVrfWriteAfterCheck_3_mask <= vrfWriteArbiter_3_bits_mask;
        allVrfWriteAfterCheck_3_data <= vrfWriteArbiter_3_bits_data;
        allVrfWriteAfterCheck_3_last <= vrfWriteArbiter_3_bits_last;
        allVrfWriteAfterCheck_3_instructionIndex <= vrfWriteArbiter_3_bits_instructionIndex;
      end
      if (enqFire_4) begin
        allVrfWriteAfterCheck_4_vd <= vrfWriteArbiter_4_bits_vd;
        allVrfWriteAfterCheck_4_offset <= vrfWriteArbiter_4_bits_offset;
        allVrfWriteAfterCheck_4_mask <= vrfWriteArbiter_4_bits_mask;
        allVrfWriteAfterCheck_4_data <= vrfWriteArbiter_4_bits_data;
        allVrfWriteAfterCheck_4_last <= vrfWriteArbiter_4_bits_last;
        allVrfWriteAfterCheck_4_instructionIndex <= vrfWriteArbiter_4_bits_instructionIndex;
      end
      if (enqFire_5) begin
        allVrfWriteAfterCheck_5_vd <= crossLaneWriteQueue_0_deq_bits_vd;
        allVrfWriteAfterCheck_5_offset <= crossLaneWriteQueue_0_deq_bits_offset;
        allVrfWriteAfterCheck_5_mask <= crossLaneWriteQueue_0_deq_bits_mask;
        allVrfWriteAfterCheck_5_data <= crossLaneWriteQueue_0_deq_bits_data;
        allVrfWriteAfterCheck_5_last <= crossLaneWriteQueue_0_deq_bits_last;
        allVrfWriteAfterCheck_5_instructionIndex <= crossLaneWriteQueue_0_deq_bits_instructionIndex;
      end
      if (enqFire_6) begin
        allVrfWriteAfterCheck_6_vd <= crossLaneWriteQueue_1_deq_bits_vd;
        allVrfWriteAfterCheck_6_offset <= crossLaneWriteQueue_1_deq_bits_offset;
        allVrfWriteAfterCheck_6_mask <= crossLaneWriteQueue_1_deq_bits_mask;
        allVrfWriteAfterCheck_6_data <= crossLaneWriteQueue_1_deq_bits_data;
        allVrfWriteAfterCheck_6_last <= crossLaneWriteQueue_1_deq_bits_last;
        allVrfWriteAfterCheck_6_instructionIndex <= crossLaneWriteQueue_1_deq_bits_instructionIndex;
      end
      if (afterCheckDequeueFire_0 ^ enqFire)
        afterCheckValid_0 <= enqFire;
      if (afterCheckDequeueFire_1 ^ enqFire_1)
        afterCheckValid_1 <= enqFire_1;
      if (afterCheckDequeueFire_2 ^ enqFire_2)
        afterCheckValid_2 <= enqFire_2;
      if (afterCheckDequeueFire_3 ^ enqFire_3)
        afterCheckValid_3 <= enqFire_3;
      if (afterCheckDequeueFire_4 ^ enqFire_4)
        afterCheckValid_4 <= enqFire_4;
      if (afterCheckDequeueFire_5 ^ enqFire_5)
        afterCheckValid_5 <= enqFire_5;
      if (afterCheckDequeueFire_6 ^ enqFire_6)
        afterCheckValid_6 <= enqFire_6;
      if (maskControlEnq[0]) begin
        maskControlVec_0_index <= laneRequest_bits_instructionIndex_0;
        maskControlVec_0_sew <= laneRequest_bits_csrInterface_vSew_0;
      end
      if (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_valid)
        maskControlVec_0_maskData <= maskInput;
      else if (maskControlEnq[0])
        maskControlVec_0_maskData <= 32'h0;
      if (maskControlReqSelect[0])
        maskControlVec_0_group <= maskControlVec_0_group + 8'h1;
      else if (maskControlEnq[0])
        maskControlVec_0_group <= 8'h0;
      maskControlVec_0_dataValid <= ~(maskControlDataDeq[0]) & (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_valid | ~(maskControlEnq[0]) & maskControlVec_0_dataValid);
      maskControlVec_0_waiteResponse <= ~maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_valid & (maskControlReqSelect[0] | ~(maskControlEnq[0]) & maskControlVec_0_waiteResponse);
      maskControlVec_0_controlValid <= ~(maskControlVec_0_controlValid & maskControlVec_releaseHit) & (maskControlEnq[0] | maskControlVec_0_controlValid);
      maskControlVec_responseFire_pipe_v <= maskControlReqSelect[0];
      maskControlVec_responseFire_pipe_pipe_v <= maskControlVec_responseFire_pipe_v;
      maskControlVec_responseFire_pipe_pipe_pipe_v <= maskControlVec_responseFire_pipe_pipe_v;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v <= maskControlVec_responseFire_pipe_pipe_pipe_v;
      if (maskControlEnq[1]) begin
        maskControlVec_1_index <= laneRequest_bits_instructionIndex_0;
        maskControlVec_1_sew <= laneRequest_bits_csrInterface_vSew_0;
      end
      if (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_1_valid)
        maskControlVec_1_maskData <= maskInput;
      else if (maskControlEnq[1])
        maskControlVec_1_maskData <= 32'h0;
      if (maskControlReqSelect[1])
        maskControlVec_1_group <= maskControlVec_1_group + 8'h1;
      else if (maskControlEnq[1])
        maskControlVec_1_group <= 8'h0;
      maskControlVec_1_dataValid <= ~(maskControlDataDeq[1]) & (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_1_valid | ~(maskControlEnq[1]) & maskControlVec_1_dataValid);
      maskControlVec_1_waiteResponse <= ~maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_1_valid & (maskControlReqSelect[1] | ~(maskControlEnq[1]) & maskControlVec_1_waiteResponse);
      maskControlVec_1_controlValid <= ~(maskControlVec_1_controlValid & maskControlVec_releaseHit_1) & (maskControlEnq[1] | maskControlVec_1_controlValid);
      maskControlVec_responseFire_pipe_v_1 <= maskControlReqSelect[1];
      maskControlVec_responseFire_pipe_pipe_v_1 <= maskControlVec_responseFire_pipe_v_1;
      maskControlVec_responseFire_pipe_pipe_pipe_v_1 <= maskControlVec_responseFire_pipe_pipe_v_1;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_1 <= maskControlVec_responseFire_pipe_pipe_pipe_v_1;
      if (maskControlEnq[2]) begin
        maskControlVec_2_index <= laneRequest_bits_instructionIndex_0;
        maskControlVec_2_sew <= laneRequest_bits_csrInterface_vSew_0;
      end
      if (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_2_valid)
        maskControlVec_2_maskData <= maskInput;
      else if (maskControlEnq[2])
        maskControlVec_2_maskData <= 32'h0;
      if (maskControlReqSelect[2])
        maskControlVec_2_group <= maskControlVec_2_group + 8'h1;
      else if (maskControlEnq[2])
        maskControlVec_2_group <= 8'h0;
      maskControlVec_2_dataValid <= ~(maskControlDataDeq[2]) & (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_2_valid | ~(maskControlEnq[2]) & maskControlVec_2_dataValid);
      maskControlVec_2_waiteResponse <= ~maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_2_valid & (maskControlReqSelect[2] | ~(maskControlEnq[2]) & maskControlVec_2_waiteResponse);
      maskControlVec_2_controlValid <= ~(maskControlVec_2_controlValid & maskControlVec_releaseHit_2) & (maskControlEnq[2] | maskControlVec_2_controlValid);
      maskControlVec_responseFire_pipe_v_2 <= maskControlReqSelect[2];
      maskControlVec_responseFire_pipe_pipe_v_2 <= maskControlVec_responseFire_pipe_v_2;
      maskControlVec_responseFire_pipe_pipe_pipe_v_2 <= maskControlVec_responseFire_pipe_pipe_v_2;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_2 <= maskControlVec_responseFire_pipe_pipe_pipe_v_2;
      if (maskControlEnq[3]) begin
        maskControlVec_3_index <= laneRequest_bits_instructionIndex_0;
        maskControlVec_3_sew <= laneRequest_bits_csrInterface_vSew_0;
      end
      if (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_3_valid)
        maskControlVec_3_maskData <= maskInput;
      else if (maskControlEnq[3])
        maskControlVec_3_maskData <= 32'h0;
      if (maskControlReqSelect[3])
        maskControlVec_3_group <= maskControlVec_3_group + 8'h1;
      else if (maskControlEnq[3])
        maskControlVec_3_group <= 8'h0;
      maskControlVec_3_dataValid <= ~(maskControlDataDeq[3]) & (maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_3_valid | ~(maskControlEnq[3]) & maskControlVec_3_dataValid);
      maskControlVec_3_waiteResponse <= ~maskControlVec_responseFire_pipe_pipe_pipe_pipe_out_3_valid & (maskControlReqSelect[3] | ~(maskControlEnq[3]) & maskControlVec_3_waiteResponse);
      maskControlVec_3_controlValid <= ~(maskControlVec_3_controlValid & maskControlVec_releaseHit_3) & (maskControlEnq[3] | maskControlVec_3_controlValid);
      maskControlVec_responseFire_pipe_v_3 <= maskControlReqSelect[3];
      maskControlVec_responseFire_pipe_pipe_v_3 <= maskControlVec_responseFire_pipe_v_3;
      maskControlVec_responseFire_pipe_pipe_pipe_v_3 <= maskControlVec_responseFire_pipe_pipe_v_3;
      maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_3 <= maskControlVec_responseFire_pipe_pipe_pipe_v_3;
      slotControl_3_mask_valid <= ~enqueueFire_3 & (maskUpdateFire_3 ^ maskFailure_3 ? maskUpdateFire_3 : slotControl_3_mask_valid);
      instructionValidNext <= instructionValid;
      vxsatResult <= (vxsatEnq_0 | vxsatEnq_1 | vxsatEnq_2 | vxsatEnq_3 | vxsatResult) & ~instructionFinishInSlot;
      if (readBusPort_0_deq_valid_0 ^ readBusPort_0_deqRelease_0)
        tokenReg <= tokenReg + tokenUpdate;
      if (readBusPort_1_deq_valid_0 ^ readBusPort_1_deqRelease_0)
        tokenReg_1 <= tokenReg_1 + tokenUpdate_1;
      if (writeBusPort_0_deq_valid_0 ^ writeBusPort_0_deqRelease_0)
        tokenReg_2 <= tokenReg_2 + tokenUpdate_2;
      if (writeBusPort_1_deq_valid_0 ^ writeBusPort_1_deqRelease_0)
        tokenReg_3 <= tokenReg_3 + tokenUpdate_3;
      if (~(queueBeforeMaskWrite_push == queueBeforeMaskWrite_pop))
        queueBeforeMaskWrite_empty <= queueBeforeMaskWrite_pop;
      emptyInstValid <= laneRequest_bits_issueInst_0 & ~_GEN_10;
    end
    if (queueBeforeMaskWrite_push) begin
      queueBeforeMaskWrite_data_vd <= queueBeforeMaskWrite_enq_bits_vd;
      queueBeforeMaskWrite_data_offset <= queueBeforeMaskWrite_enq_bits_offset;
      queueBeforeMaskWrite_data_mask <= queueBeforeMaskWrite_enq_bits_mask;
      queueBeforeMaskWrite_data_data <= queueBeforeMaskWrite_enq_bits_data;
      queueBeforeMaskWrite_data_last <= queueBeforeMaskWrite_enq_bits_last;
      queueBeforeMaskWrite_data_instructionIndex <= queueBeforeMaskWrite_enq_bits_instructionIndex;
    end
    emptyInstCount <= 8'h1 << laneRequest_bits_instructionIndex_0;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:48];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [5:0] i = 6'h0; i < 6'h31; i += 6'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        slotOccupied_0 = _RANDOM[6'h0][0];
        slotOccupied_1 = _RANDOM[6'h0][1];
        slotOccupied_2 = _RANDOM[6'h0][2];
        slotOccupied_3 = _RANDOM[6'h0][3];
        maskGroupCountVec_0 = _RANDOM[6'h0][11:4];
        maskGroupCountVec_1 = _RANDOM[6'h0][19:12];
        maskGroupCountVec_2 = _RANDOM[6'h0][27:20];
        maskGroupCountVec_3 = {_RANDOM[6'h0][31:28], _RANDOM[6'h1][3:0]};
        maskIndexVec_0 = _RANDOM[6'h1][8:4];
        maskIndexVec_1 = _RANDOM[6'h1][13:9];
        maskIndexVec_2 = _RANDOM[6'h1][18:14];
        maskIndexVec_3 = _RANDOM[6'h1][23:19];
        allVrfWriteAfterCheck_0_vd = _RANDOM[6'h2][28:24];
        allVrfWriteAfterCheck_0_offset = {_RANDOM[6'h2][31:29], _RANDOM[6'h3][2:0]};
        allVrfWriteAfterCheck_0_mask = _RANDOM[6'h3][6:3];
        allVrfWriteAfterCheck_0_data = {_RANDOM[6'h3][31:7], _RANDOM[6'h4][6:0]};
        allVrfWriteAfterCheck_0_last = _RANDOM[6'h4][7];
        allVrfWriteAfterCheck_0_instructionIndex = _RANDOM[6'h4][10:8];
        allVrfWriteAfterCheck_1_vd = _RANDOM[6'h4][15:11];
        allVrfWriteAfterCheck_1_offset = _RANDOM[6'h4][21:16];
        allVrfWriteAfterCheck_1_mask = _RANDOM[6'h4][25:22];
        allVrfWriteAfterCheck_1_data = {_RANDOM[6'h4][31:26], _RANDOM[6'h5][25:0]};
        allVrfWriteAfterCheck_1_last = _RANDOM[6'h5][26];
        allVrfWriteAfterCheck_1_instructionIndex = _RANDOM[6'h5][29:27];
        allVrfWriteAfterCheck_2_vd = {_RANDOM[6'h5][31:30], _RANDOM[6'h6][2:0]};
        allVrfWriteAfterCheck_2_offset = _RANDOM[6'h6][8:3];
        allVrfWriteAfterCheck_2_mask = _RANDOM[6'h6][12:9];
        allVrfWriteAfterCheck_2_data = {_RANDOM[6'h6][31:13], _RANDOM[6'h7][12:0]};
        allVrfWriteAfterCheck_2_last = _RANDOM[6'h7][13];
        allVrfWriteAfterCheck_2_instructionIndex = _RANDOM[6'h7][16:14];
        allVrfWriteAfterCheck_3_vd = _RANDOM[6'h7][21:17];
        allVrfWriteAfterCheck_3_offset = _RANDOM[6'h7][27:22];
        allVrfWriteAfterCheck_3_mask = _RANDOM[6'h7][31:28];
        allVrfWriteAfterCheck_3_data = _RANDOM[6'h8];
        allVrfWriteAfterCheck_3_last = _RANDOM[6'h9][0];
        allVrfWriteAfterCheck_3_instructionIndex = _RANDOM[6'h9][3:1];
        allVrfWriteAfterCheck_4_vd = _RANDOM[6'h9][8:4];
        allVrfWriteAfterCheck_4_offset = _RANDOM[6'h9][14:9];
        allVrfWriteAfterCheck_4_mask = _RANDOM[6'h9][18:15];
        allVrfWriteAfterCheck_4_data = {_RANDOM[6'h9][31:19], _RANDOM[6'hA][18:0]};
        allVrfWriteAfterCheck_4_last = _RANDOM[6'hA][19];
        allVrfWriteAfterCheck_4_instructionIndex = _RANDOM[6'hA][22:20];
        allVrfWriteAfterCheck_5_vd = _RANDOM[6'hA][27:23];
        allVrfWriteAfterCheck_5_offset = {_RANDOM[6'hA][31:28], _RANDOM[6'hB][1:0]};
        allVrfWriteAfterCheck_5_mask = _RANDOM[6'hB][5:2];
        allVrfWriteAfterCheck_5_data = {_RANDOM[6'hB][31:6], _RANDOM[6'hC][5:0]};
        allVrfWriteAfterCheck_5_last = _RANDOM[6'hC][6];
        allVrfWriteAfterCheck_5_instructionIndex = _RANDOM[6'hC][9:7];
        allVrfWriteAfterCheck_6_vd = _RANDOM[6'hC][14:10];
        allVrfWriteAfterCheck_6_offset = _RANDOM[6'hC][20:15];
        allVrfWriteAfterCheck_6_mask = _RANDOM[6'hC][24:21];
        allVrfWriteAfterCheck_6_data = {_RANDOM[6'hC][31:25], _RANDOM[6'hD][24:0]};
        allVrfWriteAfterCheck_6_last = _RANDOM[6'hD][25];
        allVrfWriteAfterCheck_6_instructionIndex = _RANDOM[6'hD][28:26];
        afterCheckValid_0 = _RANDOM[6'hD][29];
        afterCheckValid_1 = _RANDOM[6'hD][30];
        afterCheckValid_2 = _RANDOM[6'hD][31];
        afterCheckValid_3 = _RANDOM[6'hE][0];
        afterCheckValid_4 = _RANDOM[6'hE][1];
        afterCheckValid_5 = _RANDOM[6'hE][2];
        afterCheckValid_6 = _RANDOM[6'hE][3];
        maskControlVec_0_index = _RANDOM[6'hE][6:4];
        maskControlVec_0_sew = _RANDOM[6'hE][8:7];
        maskControlVec_0_maskData = {_RANDOM[6'hE][31:9], _RANDOM[6'hF][8:0]};
        maskControlVec_0_group = _RANDOM[6'hF][16:9];
        maskControlVec_0_dataValid = _RANDOM[6'hF][17];
        maskControlVec_0_waiteResponse = _RANDOM[6'hF][18];
        maskControlVec_0_controlValid = _RANDOM[6'hF][19];
        maskControlVec_responseFire_pipe_v = _RANDOM[6'hF][20];
        maskControlVec_responseFire_pipe_pipe_v = _RANDOM[6'hF][21];
        maskControlVec_responseFire_pipe_pipe_pipe_v = _RANDOM[6'hF][22];
        maskControlVec_responseFire_pipe_pipe_pipe_pipe_v = _RANDOM[6'hF][23];
        maskControlVec_1_index = _RANDOM[6'hF][26:24];
        maskControlVec_1_sew = _RANDOM[6'hF][28:27];
        maskControlVec_1_maskData = {_RANDOM[6'hF][31:29], _RANDOM[6'h10][28:0]};
        maskControlVec_1_group = {_RANDOM[6'h10][31:29], _RANDOM[6'h11][4:0]};
        maskControlVec_1_dataValid = _RANDOM[6'h11][5];
        maskControlVec_1_waiteResponse = _RANDOM[6'h11][6];
        maskControlVec_1_controlValid = _RANDOM[6'h11][7];
        maskControlVec_responseFire_pipe_v_1 = _RANDOM[6'h11][8];
        maskControlVec_responseFire_pipe_pipe_v_1 = _RANDOM[6'h11][9];
        maskControlVec_responseFire_pipe_pipe_pipe_v_1 = _RANDOM[6'h11][10];
        maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_1 = _RANDOM[6'h11][11];
        maskControlVec_2_index = _RANDOM[6'h11][14:12];
        maskControlVec_2_sew = _RANDOM[6'h11][16:15];
        maskControlVec_2_maskData = {_RANDOM[6'h11][31:17], _RANDOM[6'h12][16:0]};
        maskControlVec_2_group = _RANDOM[6'h12][24:17];
        maskControlVec_2_dataValid = _RANDOM[6'h12][25];
        maskControlVec_2_waiteResponse = _RANDOM[6'h12][26];
        maskControlVec_2_controlValid = _RANDOM[6'h12][27];
        maskControlVec_responseFire_pipe_v_2 = _RANDOM[6'h12][28];
        maskControlVec_responseFire_pipe_pipe_v_2 = _RANDOM[6'h12][29];
        maskControlVec_responseFire_pipe_pipe_pipe_v_2 = _RANDOM[6'h12][30];
        maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_2 = _RANDOM[6'h12][31];
        maskControlVec_3_index = _RANDOM[6'h13][2:0];
        maskControlVec_3_sew = _RANDOM[6'h13][4:3];
        maskControlVec_3_maskData = {_RANDOM[6'h13][31:5], _RANDOM[6'h14][4:0]};
        maskControlVec_3_group = _RANDOM[6'h14][12:5];
        maskControlVec_3_dataValid = _RANDOM[6'h14][13];
        maskControlVec_3_waiteResponse = _RANDOM[6'h14][14];
        maskControlVec_3_controlValid = _RANDOM[6'h14][15];
        maskControlVec_responseFire_pipe_v_3 = _RANDOM[6'h14][16];
        maskControlVec_responseFire_pipe_pipe_v_3 = _RANDOM[6'h14][17];
        maskControlVec_responseFire_pipe_pipe_pipe_v_3 = _RANDOM[6'h14][18];
        maskControlVec_responseFire_pipe_pipe_pipe_pipe_v_3 = _RANDOM[6'h14][19];
        slotControl_0_laneRequest_instructionIndex = _RANDOM[6'h14][22:20];
        slotControl_0_laneRequest_decodeResult_specialSlot = _RANDOM[6'h14][23];
        slotControl_0_laneRequest_decodeResult_topUop = _RANDOM[6'h14][28:24];
        slotControl_0_laneRequest_decodeResult_popCount = _RANDOM[6'h14][29];
        slotControl_0_laneRequest_decodeResult_ffo = _RANDOM[6'h14][30];
        slotControl_0_laneRequest_decodeResult_average = _RANDOM[6'h14][31];
        slotControl_0_laneRequest_decodeResult_reverse = _RANDOM[6'h15][0];
        slotControl_0_laneRequest_decodeResult_dontNeedExecuteInLane = _RANDOM[6'h15][1];
        slotControl_0_laneRequest_decodeResult_scheduler = _RANDOM[6'h15][2];
        slotControl_0_laneRequest_decodeResult_sReadVD = _RANDOM[6'h15][3];
        slotControl_0_laneRequest_decodeResult_vtype = _RANDOM[6'h15][4];
        slotControl_0_laneRequest_decodeResult_sWrite = _RANDOM[6'h15][5];
        slotControl_0_laneRequest_decodeResult_crossRead = _RANDOM[6'h15][6];
        slotControl_0_laneRequest_decodeResult_crossWrite = _RANDOM[6'h15][7];
        slotControl_0_laneRequest_decodeResult_maskUnit = _RANDOM[6'h15][8];
        slotControl_0_laneRequest_decodeResult_special = _RANDOM[6'h15][9];
        slotControl_0_laneRequest_decodeResult_saturate = _RANDOM[6'h15][10];
        slotControl_0_laneRequest_decodeResult_vwmacc = _RANDOM[6'h15][11];
        slotControl_0_laneRequest_decodeResult_readOnly = _RANDOM[6'h15][12];
        slotControl_0_laneRequest_decodeResult_maskSource = _RANDOM[6'h15][13];
        slotControl_0_laneRequest_decodeResult_maskDestination = _RANDOM[6'h15][14];
        slotControl_0_laneRequest_decodeResult_maskLogic = _RANDOM[6'h15][15];
        slotControl_0_laneRequest_decodeResult_uop = _RANDOM[6'h15][19:16];
        slotControl_0_laneRequest_decodeResult_iota = _RANDOM[6'h15][20];
        slotControl_0_laneRequest_decodeResult_mv = _RANDOM[6'h15][21];
        slotControl_0_laneRequest_decodeResult_extend = _RANDOM[6'h15][22];
        slotControl_0_laneRequest_decodeResult_unOrderWrite = _RANDOM[6'h15][23];
        slotControl_0_laneRequest_decodeResult_compress = _RANDOM[6'h15][24];
        slotControl_0_laneRequest_decodeResult_gather16 = _RANDOM[6'h15][25];
        slotControl_0_laneRequest_decodeResult_gather = _RANDOM[6'h15][26];
        slotControl_0_laneRequest_decodeResult_slid = _RANDOM[6'h15][27];
        slotControl_0_laneRequest_decodeResult_targetRd = _RANDOM[6'h15][28];
        slotControl_0_laneRequest_decodeResult_widenReduce = _RANDOM[6'h15][29];
        slotControl_0_laneRequest_decodeResult_red = _RANDOM[6'h15][30];
        slotControl_0_laneRequest_decodeResult_nr = _RANDOM[6'h15][31];
        slotControl_0_laneRequest_decodeResult_itype = _RANDOM[6'h16][0];
        slotControl_0_laneRequest_decodeResult_unsigned1 = _RANDOM[6'h16][1];
        slotControl_0_laneRequest_decodeResult_unsigned0 = _RANDOM[6'h16][2];
        slotControl_0_laneRequest_decodeResult_other = _RANDOM[6'h16][3];
        slotControl_0_laneRequest_decodeResult_multiCycle = _RANDOM[6'h16][4];
        slotControl_0_laneRequest_decodeResult_divider = _RANDOM[6'h16][5];
        slotControl_0_laneRequest_decodeResult_multiplier = _RANDOM[6'h16][6];
        slotControl_0_laneRequest_decodeResult_shift = _RANDOM[6'h16][7];
        slotControl_0_laneRequest_decodeResult_adder = _RANDOM[6'h16][8];
        slotControl_0_laneRequest_decodeResult_logic = _RANDOM[6'h16][9];
        slotControl_0_laneRequest_loadStore = _RANDOM[6'h16][10];
        slotControl_0_laneRequest_issueInst = _RANDOM[6'h16][11];
        slotControl_0_laneRequest_store = _RANDOM[6'h16][12];
        slotControl_0_laneRequest_special = _RANDOM[6'h16][13];
        slotControl_0_laneRequest_lsWholeReg = _RANDOM[6'h16][14];
        slotControl_0_laneRequest_vs1 = _RANDOM[6'h16][19:15];
        slotControl_0_laneRequest_vs2 = _RANDOM[6'h16][24:20];
        slotControl_0_laneRequest_vd = _RANDOM[6'h16][29:25];
        slotControl_0_laneRequest_loadStoreEEW = _RANDOM[6'h16][31:30];
        slotControl_0_laneRequest_mask = _RANDOM[6'h17][0];
        slotControl_0_laneRequest_segment = _RANDOM[6'h17][3:1];
        slotControl_0_laneRequest_readFromScalar = {_RANDOM[6'h17][31:4], _RANDOM[6'h18][3:0]};
        slotControl_0_laneRequest_csrInterface_vl = _RANDOM[6'h18][17:4];
        slotControl_0_laneRequest_csrInterface_vStart = _RANDOM[6'h18][31:18];
        slotControl_0_laneRequest_csrInterface_vlmul = _RANDOM[6'h19][2:0];
        slotControl_0_laneRequest_csrInterface_vSew = _RANDOM[6'h19][4:3];
        slotControl_0_laneRequest_csrInterface_vxrm = _RANDOM[6'h19][6:5];
        slotControl_0_laneRequest_csrInterface_vta = _RANDOM[6'h19][7];
        slotControl_0_laneRequest_csrInterface_vma = _RANDOM[6'h19][8];
        slotControl_0_lastGroupForInstruction = _RANDOM[6'h19][18:9];
        slotControl_0_isLastLaneForInstruction = _RANDOM[6'h19][19];
        slotControl_0_additionalRW = _RANDOM[6'h19][20];
        slotControl_0_instructionFinished = _RANDOM[6'h19][23];
        slotControl_0_mask_valid = _RANDOM[6'h19][24];
        slotControl_0_mask_bits = {_RANDOM[6'h19][31:25], _RANDOM[6'h1A][24:0]};
        slotControl_1_laneRequest_instructionIndex = _RANDOM[6'h1A][31:29];
        slotControl_1_laneRequest_decodeResult_specialSlot = _RANDOM[6'h1B][0];
        slotControl_1_laneRequest_decodeResult_topUop = _RANDOM[6'h1B][5:1];
        slotControl_1_laneRequest_decodeResult_popCount = _RANDOM[6'h1B][6];
        slotControl_1_laneRequest_decodeResult_ffo = _RANDOM[6'h1B][7];
        slotControl_1_laneRequest_decodeResult_average = _RANDOM[6'h1B][8];
        slotControl_1_laneRequest_decodeResult_reverse = _RANDOM[6'h1B][9];
        slotControl_1_laneRequest_decodeResult_dontNeedExecuteInLane = _RANDOM[6'h1B][10];
        slotControl_1_laneRequest_decodeResult_scheduler = _RANDOM[6'h1B][11];
        slotControl_1_laneRequest_decodeResult_sReadVD = _RANDOM[6'h1B][12];
        slotControl_1_laneRequest_decodeResult_vtype = _RANDOM[6'h1B][13];
        slotControl_1_laneRequest_decodeResult_sWrite = _RANDOM[6'h1B][14];
        slotControl_1_laneRequest_decodeResult_crossRead = _RANDOM[6'h1B][15];
        slotControl_1_laneRequest_decodeResult_crossWrite = _RANDOM[6'h1B][16];
        slotControl_1_laneRequest_decodeResult_maskUnit = _RANDOM[6'h1B][17];
        slotControl_1_laneRequest_decodeResult_special = _RANDOM[6'h1B][18];
        slotControl_1_laneRequest_decodeResult_saturate = _RANDOM[6'h1B][19];
        slotControl_1_laneRequest_decodeResult_vwmacc = _RANDOM[6'h1B][20];
        slotControl_1_laneRequest_decodeResult_readOnly = _RANDOM[6'h1B][21];
        slotControl_1_laneRequest_decodeResult_maskSource = _RANDOM[6'h1B][22];
        slotControl_1_laneRequest_decodeResult_maskDestination = _RANDOM[6'h1B][23];
        slotControl_1_laneRequest_decodeResult_maskLogic = _RANDOM[6'h1B][24];
        slotControl_1_laneRequest_decodeResult_uop = _RANDOM[6'h1B][28:25];
        slotControl_1_laneRequest_decodeResult_iota = _RANDOM[6'h1B][29];
        slotControl_1_laneRequest_decodeResult_mv = _RANDOM[6'h1B][30];
        slotControl_1_laneRequest_decodeResult_extend = _RANDOM[6'h1B][31];
        slotControl_1_laneRequest_decodeResult_unOrderWrite = _RANDOM[6'h1C][0];
        slotControl_1_laneRequest_decodeResult_compress = _RANDOM[6'h1C][1];
        slotControl_1_laneRequest_decodeResult_gather16 = _RANDOM[6'h1C][2];
        slotControl_1_laneRequest_decodeResult_gather = _RANDOM[6'h1C][3];
        slotControl_1_laneRequest_decodeResult_slid = _RANDOM[6'h1C][4];
        slotControl_1_laneRequest_decodeResult_targetRd = _RANDOM[6'h1C][5];
        slotControl_1_laneRequest_decodeResult_widenReduce = _RANDOM[6'h1C][6];
        slotControl_1_laneRequest_decodeResult_red = _RANDOM[6'h1C][7];
        slotControl_1_laneRequest_decodeResult_nr = _RANDOM[6'h1C][8];
        slotControl_1_laneRequest_decodeResult_itype = _RANDOM[6'h1C][9];
        slotControl_1_laneRequest_decodeResult_unsigned1 = _RANDOM[6'h1C][10];
        slotControl_1_laneRequest_decodeResult_unsigned0 = _RANDOM[6'h1C][11];
        slotControl_1_laneRequest_decodeResult_other = _RANDOM[6'h1C][12];
        slotControl_1_laneRequest_decodeResult_multiCycle = _RANDOM[6'h1C][13];
        slotControl_1_laneRequest_decodeResult_divider = _RANDOM[6'h1C][14];
        slotControl_1_laneRequest_decodeResult_multiplier = _RANDOM[6'h1C][15];
        slotControl_1_laneRequest_decodeResult_shift = _RANDOM[6'h1C][16];
        slotControl_1_laneRequest_decodeResult_adder = _RANDOM[6'h1C][17];
        slotControl_1_laneRequest_decodeResult_logic = _RANDOM[6'h1C][18];
        slotControl_1_laneRequest_loadStore = _RANDOM[6'h1C][19];
        slotControl_1_laneRequest_issueInst = _RANDOM[6'h1C][20];
        slotControl_1_laneRequest_store = _RANDOM[6'h1C][21];
        slotControl_1_laneRequest_special = _RANDOM[6'h1C][22];
        slotControl_1_laneRequest_lsWholeReg = _RANDOM[6'h1C][23];
        slotControl_1_laneRequest_vs1 = _RANDOM[6'h1C][28:24];
        slotControl_1_laneRequest_vs2 = {_RANDOM[6'h1C][31:29], _RANDOM[6'h1D][1:0]};
        slotControl_1_laneRequest_vd = _RANDOM[6'h1D][6:2];
        slotControl_1_laneRequest_loadStoreEEW = _RANDOM[6'h1D][8:7];
        slotControl_1_laneRequest_mask = _RANDOM[6'h1D][9];
        slotControl_1_laneRequest_segment = _RANDOM[6'h1D][12:10];
        slotControl_1_laneRequest_readFromScalar = {_RANDOM[6'h1D][31:13], _RANDOM[6'h1E][12:0]};
        slotControl_1_laneRequest_csrInterface_vl = _RANDOM[6'h1E][26:13];
        slotControl_1_laneRequest_csrInterface_vStart = {_RANDOM[6'h1E][31:27], _RANDOM[6'h1F][8:0]};
        slotControl_1_laneRequest_csrInterface_vlmul = _RANDOM[6'h1F][11:9];
        slotControl_1_laneRequest_csrInterface_vSew = _RANDOM[6'h1F][13:12];
        slotControl_1_laneRequest_csrInterface_vxrm = _RANDOM[6'h1F][15:14];
        slotControl_1_laneRequest_csrInterface_vta = _RANDOM[6'h1F][16];
        slotControl_1_laneRequest_csrInterface_vma = _RANDOM[6'h1F][17];
        slotControl_1_lastGroupForInstruction = _RANDOM[6'h1F][27:18];
        slotControl_1_isLastLaneForInstruction = _RANDOM[6'h1F][28];
        slotControl_1_additionalRW = _RANDOM[6'h1F][29];
        slotControl_1_instructionFinished = _RANDOM[6'h20][0];
        slotControl_1_mask_valid = _RANDOM[6'h20][1];
        slotControl_1_mask_bits = {_RANDOM[6'h20][31:2], _RANDOM[6'h21][1:0]};
        slotControl_2_laneRequest_instructionIndex = _RANDOM[6'h21][8:6];
        slotControl_2_laneRequest_decodeResult_specialSlot = _RANDOM[6'h21][9];
        slotControl_2_laneRequest_decodeResult_topUop = _RANDOM[6'h21][14:10];
        slotControl_2_laneRequest_decodeResult_popCount = _RANDOM[6'h21][15];
        slotControl_2_laneRequest_decodeResult_ffo = _RANDOM[6'h21][16];
        slotControl_2_laneRequest_decodeResult_average = _RANDOM[6'h21][17];
        slotControl_2_laneRequest_decodeResult_reverse = _RANDOM[6'h21][18];
        slotControl_2_laneRequest_decodeResult_dontNeedExecuteInLane = _RANDOM[6'h21][19];
        slotControl_2_laneRequest_decodeResult_scheduler = _RANDOM[6'h21][20];
        slotControl_2_laneRequest_decodeResult_sReadVD = _RANDOM[6'h21][21];
        slotControl_2_laneRequest_decodeResult_vtype = _RANDOM[6'h21][22];
        slotControl_2_laneRequest_decodeResult_sWrite = _RANDOM[6'h21][23];
        slotControl_2_laneRequest_decodeResult_crossRead = _RANDOM[6'h21][24];
        slotControl_2_laneRequest_decodeResult_crossWrite = _RANDOM[6'h21][25];
        slotControl_2_laneRequest_decodeResult_maskUnit = _RANDOM[6'h21][26];
        slotControl_2_laneRequest_decodeResult_special = _RANDOM[6'h21][27];
        slotControl_2_laneRequest_decodeResult_saturate = _RANDOM[6'h21][28];
        slotControl_2_laneRequest_decodeResult_vwmacc = _RANDOM[6'h21][29];
        slotControl_2_laneRequest_decodeResult_readOnly = _RANDOM[6'h21][30];
        slotControl_2_laneRequest_decodeResult_maskSource = _RANDOM[6'h21][31];
        slotControl_2_laneRequest_decodeResult_maskDestination = _RANDOM[6'h22][0];
        slotControl_2_laneRequest_decodeResult_maskLogic = _RANDOM[6'h22][1];
        slotControl_2_laneRequest_decodeResult_uop = _RANDOM[6'h22][5:2];
        slotControl_2_laneRequest_decodeResult_iota = _RANDOM[6'h22][6];
        slotControl_2_laneRequest_decodeResult_mv = _RANDOM[6'h22][7];
        slotControl_2_laneRequest_decodeResult_extend = _RANDOM[6'h22][8];
        slotControl_2_laneRequest_decodeResult_unOrderWrite = _RANDOM[6'h22][9];
        slotControl_2_laneRequest_decodeResult_compress = _RANDOM[6'h22][10];
        slotControl_2_laneRequest_decodeResult_gather16 = _RANDOM[6'h22][11];
        slotControl_2_laneRequest_decodeResult_gather = _RANDOM[6'h22][12];
        slotControl_2_laneRequest_decodeResult_slid = _RANDOM[6'h22][13];
        slotControl_2_laneRequest_decodeResult_targetRd = _RANDOM[6'h22][14];
        slotControl_2_laneRequest_decodeResult_widenReduce = _RANDOM[6'h22][15];
        slotControl_2_laneRequest_decodeResult_red = _RANDOM[6'h22][16];
        slotControl_2_laneRequest_decodeResult_nr = _RANDOM[6'h22][17];
        slotControl_2_laneRequest_decodeResult_itype = _RANDOM[6'h22][18];
        slotControl_2_laneRequest_decodeResult_unsigned1 = _RANDOM[6'h22][19];
        slotControl_2_laneRequest_decodeResult_unsigned0 = _RANDOM[6'h22][20];
        slotControl_2_laneRequest_decodeResult_other = _RANDOM[6'h22][21];
        slotControl_2_laneRequest_decodeResult_multiCycle = _RANDOM[6'h22][22];
        slotControl_2_laneRequest_decodeResult_divider = _RANDOM[6'h22][23];
        slotControl_2_laneRequest_decodeResult_multiplier = _RANDOM[6'h22][24];
        slotControl_2_laneRequest_decodeResult_shift = _RANDOM[6'h22][25];
        slotControl_2_laneRequest_decodeResult_adder = _RANDOM[6'h22][26];
        slotControl_2_laneRequest_decodeResult_logic = _RANDOM[6'h22][27];
        slotControl_2_laneRequest_loadStore = _RANDOM[6'h22][28];
        slotControl_2_laneRequest_issueInst = _RANDOM[6'h22][29];
        slotControl_2_laneRequest_store = _RANDOM[6'h22][30];
        slotControl_2_laneRequest_special = _RANDOM[6'h22][31];
        slotControl_2_laneRequest_lsWholeReg = _RANDOM[6'h23][0];
        slotControl_2_laneRequest_vs1 = _RANDOM[6'h23][5:1];
        slotControl_2_laneRequest_vs2 = _RANDOM[6'h23][10:6];
        slotControl_2_laneRequest_vd = _RANDOM[6'h23][15:11];
        slotControl_2_laneRequest_loadStoreEEW = _RANDOM[6'h23][17:16];
        slotControl_2_laneRequest_mask = _RANDOM[6'h23][18];
        slotControl_2_laneRequest_segment = _RANDOM[6'h23][21:19];
        slotControl_2_laneRequest_readFromScalar = {_RANDOM[6'h23][31:22], _RANDOM[6'h24][21:0]};
        slotControl_2_laneRequest_csrInterface_vl = {_RANDOM[6'h24][31:22], _RANDOM[6'h25][3:0]};
        slotControl_2_laneRequest_csrInterface_vStart = _RANDOM[6'h25][17:4];
        slotControl_2_laneRequest_csrInterface_vlmul = _RANDOM[6'h25][20:18];
        slotControl_2_laneRequest_csrInterface_vSew = _RANDOM[6'h25][22:21];
        slotControl_2_laneRequest_csrInterface_vxrm = _RANDOM[6'h25][24:23];
        slotControl_2_laneRequest_csrInterface_vta = _RANDOM[6'h25][25];
        slotControl_2_laneRequest_csrInterface_vma = _RANDOM[6'h25][26];
        slotControl_2_lastGroupForInstruction = {_RANDOM[6'h25][31:27], _RANDOM[6'h26][4:0]};
        slotControl_2_isLastLaneForInstruction = _RANDOM[6'h26][5];
        slotControl_2_additionalRW = _RANDOM[6'h26][6];
        slotControl_2_instructionFinished = _RANDOM[6'h26][9];
        slotControl_2_mask_valid = _RANDOM[6'h26][10];
        slotControl_2_mask_bits = {_RANDOM[6'h26][31:11], _RANDOM[6'h27][10:0]};
        slotControl_3_laneRequest_instructionIndex = _RANDOM[6'h27][17:15];
        slotControl_3_laneRequest_decodeResult_specialSlot = _RANDOM[6'h27][18];
        slotControl_3_laneRequest_decodeResult_topUop = _RANDOM[6'h27][23:19];
        slotControl_3_laneRequest_decodeResult_popCount = _RANDOM[6'h27][24];
        slotControl_3_laneRequest_decodeResult_ffo = _RANDOM[6'h27][25];
        slotControl_3_laneRequest_decodeResult_average = _RANDOM[6'h27][26];
        slotControl_3_laneRequest_decodeResult_reverse = _RANDOM[6'h27][27];
        slotControl_3_laneRequest_decodeResult_dontNeedExecuteInLane = _RANDOM[6'h27][28];
        slotControl_3_laneRequest_decodeResult_scheduler = _RANDOM[6'h27][29];
        slotControl_3_laneRequest_decodeResult_sReadVD = _RANDOM[6'h27][30];
        slotControl_3_laneRequest_decodeResult_vtype = _RANDOM[6'h27][31];
        slotControl_3_laneRequest_decodeResult_sWrite = _RANDOM[6'h28][0];
        slotControl_3_laneRequest_decodeResult_crossRead = _RANDOM[6'h28][1];
        slotControl_3_laneRequest_decodeResult_crossWrite = _RANDOM[6'h28][2];
        slotControl_3_laneRequest_decodeResult_maskUnit = _RANDOM[6'h28][3];
        slotControl_3_laneRequest_decodeResult_special = _RANDOM[6'h28][4];
        slotControl_3_laneRequest_decodeResult_saturate = _RANDOM[6'h28][5];
        slotControl_3_laneRequest_decodeResult_vwmacc = _RANDOM[6'h28][6];
        slotControl_3_laneRequest_decodeResult_readOnly = _RANDOM[6'h28][7];
        slotControl_3_laneRequest_decodeResult_maskSource = _RANDOM[6'h28][8];
        slotControl_3_laneRequest_decodeResult_maskDestination = _RANDOM[6'h28][9];
        slotControl_3_laneRequest_decodeResult_maskLogic = _RANDOM[6'h28][10];
        slotControl_3_laneRequest_decodeResult_uop = _RANDOM[6'h28][14:11];
        slotControl_3_laneRequest_decodeResult_iota = _RANDOM[6'h28][15];
        slotControl_3_laneRequest_decodeResult_mv = _RANDOM[6'h28][16];
        slotControl_3_laneRequest_decodeResult_extend = _RANDOM[6'h28][17];
        slotControl_3_laneRequest_decodeResult_unOrderWrite = _RANDOM[6'h28][18];
        slotControl_3_laneRequest_decodeResult_compress = _RANDOM[6'h28][19];
        slotControl_3_laneRequest_decodeResult_gather16 = _RANDOM[6'h28][20];
        slotControl_3_laneRequest_decodeResult_gather = _RANDOM[6'h28][21];
        slotControl_3_laneRequest_decodeResult_slid = _RANDOM[6'h28][22];
        slotControl_3_laneRequest_decodeResult_targetRd = _RANDOM[6'h28][23];
        slotControl_3_laneRequest_decodeResult_widenReduce = _RANDOM[6'h28][24];
        slotControl_3_laneRequest_decodeResult_red = _RANDOM[6'h28][25];
        slotControl_3_laneRequest_decodeResult_nr = _RANDOM[6'h28][26];
        slotControl_3_laneRequest_decodeResult_itype = _RANDOM[6'h28][27];
        slotControl_3_laneRequest_decodeResult_unsigned1 = _RANDOM[6'h28][28];
        slotControl_3_laneRequest_decodeResult_unsigned0 = _RANDOM[6'h28][29];
        slotControl_3_laneRequest_decodeResult_other = _RANDOM[6'h28][30];
        slotControl_3_laneRequest_decodeResult_multiCycle = _RANDOM[6'h28][31];
        slotControl_3_laneRequest_decodeResult_divider = _RANDOM[6'h29][0];
        slotControl_3_laneRequest_decodeResult_multiplier = _RANDOM[6'h29][1];
        slotControl_3_laneRequest_decodeResult_shift = _RANDOM[6'h29][2];
        slotControl_3_laneRequest_decodeResult_adder = _RANDOM[6'h29][3];
        slotControl_3_laneRequest_decodeResult_logic = _RANDOM[6'h29][4];
        slotControl_3_laneRequest_loadStore = _RANDOM[6'h29][5];
        slotControl_3_laneRequest_issueInst = _RANDOM[6'h29][6];
        slotControl_3_laneRequest_store = _RANDOM[6'h29][7];
        slotControl_3_laneRequest_special = _RANDOM[6'h29][8];
        slotControl_3_laneRequest_lsWholeReg = _RANDOM[6'h29][9];
        slotControl_3_laneRequest_vs1 = _RANDOM[6'h29][14:10];
        slotControl_3_laneRequest_vs2 = _RANDOM[6'h29][19:15];
        slotControl_3_laneRequest_vd = _RANDOM[6'h29][24:20];
        slotControl_3_laneRequest_loadStoreEEW = _RANDOM[6'h29][26:25];
        slotControl_3_laneRequest_mask = _RANDOM[6'h29][27];
        slotControl_3_laneRequest_segment = _RANDOM[6'h29][30:28];
        slotControl_3_laneRequest_readFromScalar = {_RANDOM[6'h29][31], _RANDOM[6'h2A][30:0]};
        slotControl_3_laneRequest_csrInterface_vl = {_RANDOM[6'h2A][31], _RANDOM[6'h2B][12:0]};
        slotControl_3_laneRequest_csrInterface_vStart = _RANDOM[6'h2B][26:13];
        slotControl_3_laneRequest_csrInterface_vlmul = _RANDOM[6'h2B][29:27];
        slotControl_3_laneRequest_csrInterface_vSew = _RANDOM[6'h2B][31:30];
        slotControl_3_laneRequest_csrInterface_vxrm = _RANDOM[6'h2C][1:0];
        slotControl_3_laneRequest_csrInterface_vta = _RANDOM[6'h2C][2];
        slotControl_3_laneRequest_csrInterface_vma = _RANDOM[6'h2C][3];
        slotControl_3_lastGroupForInstruction = _RANDOM[6'h2C][13:4];
        slotControl_3_isLastLaneForInstruction = _RANDOM[6'h2C][14];
        slotControl_3_additionalRW = _RANDOM[6'h2C][15];
        slotControl_3_instructionFinished = _RANDOM[6'h2C][18];
        slotControl_3_mask_valid = _RANDOM[6'h2C][19];
        slotControl_3_mask_bits = {_RANDOM[6'h2C][31:20], _RANDOM[6'h2D][19:0]};
        instructionValidNext = _RANDOM[6'h2D][31:24];
        vxsatResult = _RANDOM[6'h2E][7:0];
        tokenReg = _RANDOM[6'h2E][10:8];
        tokenReg_1 = _RANDOM[6'h2E][13:11];
        tokenReg_2 = _RANDOM[6'h2E][16:14];
        tokenReg_3 = _RANDOM[6'h2E][19:17];
        queueBeforeMaskWrite_data_vd = _RANDOM[6'h2E][24:20];
        queueBeforeMaskWrite_data_offset = _RANDOM[6'h2E][30:25];
        queueBeforeMaskWrite_data_mask = {_RANDOM[6'h2E][31], _RANDOM[6'h2F][2:0]};
        queueBeforeMaskWrite_data_data = {_RANDOM[6'h2F][31:3], _RANDOM[6'h30][2:0]};
        queueBeforeMaskWrite_data_last = _RANDOM[6'h30][3];
        queueBeforeMaskWrite_data_instructionIndex = _RANDOM[6'h30][6:4];
        queueBeforeMaskWrite_empty = _RANDOM[6'h30][7];
        emptyInstValid = _RANDOM[6'h30][8];
        emptyInstCount = _RANDOM[6'h30][16:9];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire [4:0]    readCheckRequestVec_0_vs;
  wire [5:0]    readCheckRequestVec_0_offset;
  wire [2:0]    readCheckRequestVec_0_instructionIndex;
  wire [4:0]    readCheckRequestVec_1_vs;
  wire [5:0]    readCheckRequestVec_1_offset;
  wire [2:0]    readCheckRequestVec_1_instructionIndex;
  wire [4:0]    readCheckRequestVec_2_vs;
  wire [5:0]    readCheckRequestVec_2_offset;
  wire [2:0]    readCheckRequestVec_2_instructionIndex;
  wire [4:0]    readCheckRequestVec_3_vs;
  wire [5:0]    readCheckRequestVec_3_offset;
  wire [2:0]    readCheckRequestVec_3_instructionIndex;
  wire [4:0]    readCheckRequestVec_4_vs;
  wire [5:0]    readCheckRequestVec_4_offset;
  wire [2:0]    readCheckRequestVec_4_instructionIndex;
  wire [4:0]    readCheckRequestVec_5_vs;
  wire [5:0]    readCheckRequestVec_5_offset;
  wire [2:0]    readCheckRequestVec_5_instructionIndex;
  wire [4:0]    readCheckRequestVec_6_vs;
  wire [5:0]    readCheckRequestVec_6_offset;
  wire [2:0]    readCheckRequestVec_6_instructionIndex;
  wire [4:0]    readCheckRequestVec_7_vs;
  wire [5:0]    readCheckRequestVec_7_offset;
  wire [2:0]    readCheckRequestVec_7_instructionIndex;
  wire [4:0]    readCheckRequestVec_8_vs;
  wire [5:0]    readCheckRequestVec_8_offset;
  wire [2:0]    readCheckRequestVec_8_instructionIndex;
  wire [4:0]    readCheckRequestVec_9_vs;
  wire [5:0]    readCheckRequestVec_9_offset;
  wire [2:0]    readCheckRequestVec_9_instructionIndex;
  wire [4:0]    readCheckRequestVec_10_vs;
  wire [5:0]    readCheckRequestVec_10_offset;
  wire [2:0]    readCheckRequestVec_10_instructionIndex;
  wire [4:0]    readCheckRequestVec_11_vs;
  wire [5:0]    readCheckRequestVec_11_offset;
  wire [2:0]    readCheckRequestVec_11_instructionIndex;
  wire [4:0]    readCheckRequestVec_12_vs;
  wire [5:0]    readCheckRequestVec_12_offset;
  wire [2:0]    readCheckRequestVec_12_instructionIndex;
  wire [4:0]    readCheckRequestVec_13_vs;
  wire [5:0]    readCheckRequestVec_13_offset;
  wire [2:0]    readCheckRequestVec_13_instructionIndex;
  wire          crossLaneWriteQueue_0_empty;
  assign crossLaneWriteQueue_0_empty = _crossLaneWriteQueue_fifo_empty;
  wire          crossLaneWriteQueue_0_full;
  assign crossLaneWriteQueue_0_full = _crossLaneWriteQueue_fifo_full;
  wire          crossLaneWriteQueue_1_empty;
  assign crossLaneWriteQueue_1_empty = _crossLaneWriteQueue_fifo_1_empty;
  wire          crossLaneWriteQueue_1_full;
  assign crossLaneWriteQueue_1_full = _crossLaneWriteQueue_fifo_1_full;
  wire          readBeforeMaskedWrite_ready;
  assign slotMaskRequestVec_0_bits = _stage0_updateLaneState_maskGroupCount;
  wire          vrfReadRequest_0_0_ready;
  wire          vrfReadRequest_0_1_ready;
  wire          vrfReadRequest_0_2_ready;
  assign executeEnqueueValid_0 = _executionUnit_vfuRequest_valid;
  wire          stage3EnqWire_valid;
  assign stage3EnqWire_valid = _executionUnit_dequeue_valid;
  assign vrfWriteArbiter_0_valid = _stage3_vrfWriteRequest_valid;
  assign vrfWriteArbiter_0_bits_mask = _stage3_vrfWriteRequest_bits_mask;
  assign vrfWriteArbiter_0_bits_instructionIndex = _stage3_vrfWriteRequest_bits_instructionIndex;
  wire          queue_empty;
  assign queue_empty = _queue_fifo_empty;
  wire          queue_full;
  assign queue_full = _queue_fifo_full;
  wire          queue_1_empty;
  assign queue_1_empty = _queue_fifo_1_empty;
  wire          queue_1_full;
  assign queue_1_full = _queue_fifo_1_full;
  assign slotMaskRequestVec_1_bits = _stage0_1_updateLaneState_maskGroupCount;
  wire          vrfReadRequest_1_0_ready;
  wire          vrfReadRequest_1_1_ready;
  wire          vrfReadRequest_1_2_ready;
  assign executeEnqueueValid_1 = _executionUnit_1_vfuRequest_valid;
  wire          stage3EnqWire_1_valid;
  assign stage3EnqWire_1_valid = _executionUnit_1_dequeue_valid;
  assign vrfWriteArbiter_1_valid = _stage3_1_vrfWriteRequest_valid;
  assign vrfWriteArbiter_1_bits_mask = _stage3_1_vrfWriteRequest_bits_mask;
  assign vrfWriteArbiter_1_bits_instructionIndex = _stage3_1_vrfWriteRequest_bits_instructionIndex;
  assign slotMaskRequestVec_2_bits = _stage0_2_updateLaneState_maskGroupCount;
  wire          vrfReadRequest_2_0_ready;
  wire          vrfReadRequest_2_1_ready;
  wire          vrfReadRequest_2_2_ready;
  assign executeEnqueueValid_2 = _executionUnit_2_vfuRequest_valid;
  wire          stage3EnqWire_2_valid;
  assign stage3EnqWire_2_valid = _executionUnit_2_dequeue_valid;
  assign vrfWriteArbiter_2_valid = _stage3_2_vrfWriteRequest_valid;
  assign vrfWriteArbiter_2_bits_mask = _stage3_2_vrfWriteRequest_bits_mask;
  assign vrfWriteArbiter_2_bits_instructionIndex = _stage3_2_vrfWriteRequest_bits_instructionIndex;
  assign slotMaskRequestVec_3_bits = _stage0_3_updateLaneState_maskGroupCount;
  wire          vrfReadRequest_3_0_ready;
  wire          vrfReadRequest_3_1_ready;
  wire          vrfReadRequest_3_2_ready;
  assign executeEnqueueValid_3 = _executionUnit_3_vfuRequest_valid;
  wire          stage3EnqWire_3_valid;
  assign stage3EnqWire_3_valid = _executionUnit_3_dequeue_valid;
  assign vrfWriteArbiter_3_valid = _stage3_3_vrfWriteRequest_valid;
  assign vrfWriteArbiter_3_bits_mask = _stage3_3_vrfWriteRequest_bits_mask;
  assign vrfWriteArbiter_3_bits_instructionIndex = _stage3_3_vrfWriteRequest_bits_instructionIndex;
  wire          executeOccupied_0;
  assign executeOccupied_0 = _vfuResponse_logicArbiter_io_out_valid;
  wire          executeOccupied_1;
  assign executeOccupied_1 = _vfuResponse_adderArbiter_io_out_valid;
  wire          executeOccupied_2;
  assign executeOccupied_2 = _vfuResponse_shiftDistributor_requestToVfu_valid;
  wire          executeOccupied_3;
  assign executeOccupied_3 = _vfuResponse_multiplierArbiter_io_out_valid;
  wire          executeOccupied_5;
  assign executeOccupied_5 = _vfuResponse_otherDistributor_requestToVfu_valid;
  VRF vrf (
    .clock                                              (clock),
    .reset                                              (reset),
    .readRequests_0_ready                               (_vrf_readRequests_0_ready),
    .readRequests_0_valid                               (_vrfReadArbiter_0_io_out_valid),
    .readRequests_0_bits_vs                             (_vrfReadArbiter_0_io_out_bits_vs),
    .readRequests_0_bits_readSource                     (_vrfReadArbiter_0_io_out_bits_readSource),
    .readRequests_0_bits_offset                         (_vrfReadArbiter_0_io_out_bits_offset),
    .readRequests_0_bits_instructionIndex               (_vrfReadArbiter_0_io_out_bits_instructionIndex),
    .readRequests_1_ready                               (_vrf_readRequests_1_ready),
    .readRequests_1_valid                               (_vrfReadArbiter_1_io_out_valid),
    .readRequests_1_bits_vs                             (_vrfReadArbiter_1_io_out_bits_vs),
    .readRequests_1_bits_readSource                     (_vrfReadArbiter_1_io_out_bits_readSource),
    .readRequests_1_bits_offset                         (_vrfReadArbiter_1_io_out_bits_offset),
    .readRequests_1_bits_instructionIndex               (_vrfReadArbiter_1_io_out_bits_instructionIndex),
    .readRequests_2_ready                               (_vrf_readRequests_2_ready),
    .readRequests_2_valid                               (_vrfReadArbiter_2_io_out_valid),
    .readRequests_2_bits_vs                             (_vrfReadArbiter_2_io_out_bits_vs),
    .readRequests_2_bits_readSource                     (_vrfReadArbiter_2_io_out_bits_readSource),
    .readRequests_2_bits_offset                         (_vrfReadArbiter_2_io_out_bits_offset),
    .readRequests_2_bits_instructionIndex               (_vrfReadArbiter_2_io_out_bits_instructionIndex),
    .readRequests_3_ready                               (_vrf_readRequests_3_ready),
    .readRequests_3_valid                               (_vrfReadArbiter_3_io_out_valid),
    .readRequests_3_bits_vs                             (_vrfReadArbiter_3_io_out_bits_vs),
    .readRequests_3_bits_readSource                     (_vrfReadArbiter_3_io_out_bits_readSource),
    .readRequests_3_bits_offset                         (_vrfReadArbiter_3_io_out_bits_offset),
    .readRequests_3_bits_instructionIndex               (_vrfReadArbiter_3_io_out_bits_instructionIndex),
    .readRequests_4_ready                               (_vrf_readRequests_4_ready),
    .readRequests_4_valid                               (_vrfReadArbiter_4_io_out_valid),
    .readRequests_4_bits_vs                             (_vrfReadArbiter_4_io_out_bits_vs),
    .readRequests_4_bits_readSource                     (_vrfReadArbiter_4_io_out_bits_readSource),
    .readRequests_4_bits_offset                         (_vrfReadArbiter_4_io_out_bits_offset),
    .readRequests_4_bits_instructionIndex               (_vrfReadArbiter_4_io_out_bits_instructionIndex),
    .readRequests_5_ready                               (_vrf_readRequests_5_ready),
    .readRequests_5_valid                               (_vrfReadArbiter_5_io_out_valid),
    .readRequests_5_bits_vs                             (_vrfReadArbiter_5_io_out_bits_vs),
    .readRequests_5_bits_readSource                     (_vrfReadArbiter_5_io_out_bits_readSource),
    .readRequests_5_bits_offset                         (_vrfReadArbiter_5_io_out_bits_offset),
    .readRequests_5_bits_instructionIndex               (_vrfReadArbiter_5_io_out_bits_instructionIndex),
    .readRequests_6_ready                               (_vrf_readRequests_6_ready),
    .readRequests_6_valid                               (_vrfReadArbiter_6_io_out_valid),
    .readRequests_6_bits_vs                             (_vrfReadArbiter_6_io_out_bits_vs),
    .readRequests_6_bits_readSource                     (_vrfReadArbiter_6_io_out_bits_readSource),
    .readRequests_6_bits_offset                         (_vrfReadArbiter_6_io_out_bits_offset),
    .readRequests_6_bits_instructionIndex               (_vrfReadArbiter_6_io_out_bits_instructionIndex),
    .readRequests_7_ready                               (_vrf_readRequests_7_ready),
    .readRequests_7_valid                               (_vrfReadArbiter_7_io_out_valid),
    .readRequests_7_bits_vs                             (_vrfReadArbiter_7_io_out_bits_vs),
    .readRequests_7_bits_readSource                     (_vrfReadArbiter_7_io_out_bits_readSource),
    .readRequests_7_bits_offset                         (_vrfReadArbiter_7_io_out_bits_offset),
    .readRequests_7_bits_instructionIndex               (_vrfReadArbiter_7_io_out_bits_instructionIndex),
    .readRequests_8_ready                               (_vrf_readRequests_8_ready),
    .readRequests_8_valid                               (_vrfReadArbiter_8_io_out_valid),
    .readRequests_8_bits_vs                             (_vrfReadArbiter_8_io_out_bits_vs),
    .readRequests_8_bits_readSource                     (_vrfReadArbiter_8_io_out_bits_readSource),
    .readRequests_8_bits_offset                         (_vrfReadArbiter_8_io_out_bits_offset),
    .readRequests_8_bits_instructionIndex               (_vrfReadArbiter_8_io_out_bits_instructionIndex),
    .readRequests_9_ready                               (_vrf_readRequests_9_ready),
    .readRequests_9_valid                               (_vrfReadArbiter_9_io_out_valid),
    .readRequests_9_bits_vs                             (_vrfReadArbiter_9_io_out_bits_vs),
    .readRequests_9_bits_readSource                     (_vrfReadArbiter_9_io_out_bits_readSource),
    .readRequests_9_bits_offset                         (_vrfReadArbiter_9_io_out_bits_offset),
    .readRequests_9_bits_instructionIndex               (_vrfReadArbiter_9_io_out_bits_instructionIndex),
    .readRequests_10_ready                              (_vrf_readRequests_10_ready),
    .readRequests_10_valid                              (_vrfReadArbiter_10_io_out_valid),
    .readRequests_10_bits_vs                            (_vrfReadArbiter_10_io_out_bits_vs),
    .readRequests_10_bits_readSource                    (_vrfReadArbiter_10_io_out_bits_readSource),
    .readRequests_10_bits_offset                        (_vrfReadArbiter_10_io_out_bits_offset),
    .readRequests_10_bits_instructionIndex              (_vrfReadArbiter_10_io_out_bits_instructionIndex),
    .readRequests_11_ready                              (_vrf_readRequests_11_ready),
    .readRequests_11_valid                              (_vrfReadArbiter_11_io_out_valid),
    .readRequests_11_bits_vs                            (_vrfReadArbiter_11_io_out_bits_vs),
    .readRequests_11_bits_readSource                    (_vrfReadArbiter_11_io_out_bits_readSource),
    .readRequests_11_bits_offset                        (_vrfReadArbiter_11_io_out_bits_offset),
    .readRequests_11_bits_instructionIndex              (_vrfReadArbiter_11_io_out_bits_instructionIndex),
    .readRequests_12_ready                              (_vrf_readRequests_12_ready),
    .readRequests_12_valid                              (_vrfReadArbiter_12_io_out_valid),
    .readRequests_12_bits_vs                            (_vrfReadArbiter_12_io_out_bits_vs),
    .readRequests_12_bits_readSource                    (_vrfReadArbiter_12_io_out_bits_readSource),
    .readRequests_12_bits_offset                        (_vrfReadArbiter_12_io_out_bits_offset),
    .readRequests_12_bits_instructionIndex              (_vrfReadArbiter_12_io_out_bits_instructionIndex),
    .readRequests_13_ready                              (_vrf_readRequests_13_ready),
    .readRequests_13_valid                              (_vrfReadArbiter_13_io_out_valid),
    .readRequests_13_bits_vs                            (_vrfReadArbiter_13_io_out_bits_vs),
    .readRequests_13_bits_readSource                    (_vrfReadArbiter_13_io_out_bits_readSource),
    .readRequests_13_bits_offset                        (_vrfReadArbiter_13_io_out_bits_offset),
    .readRequests_13_bits_instructionIndex              (_vrfReadArbiter_13_io_out_bits_instructionIndex),
    .readCheck_0_vs                                     (readCheckRequestVec_0_vs),
    .readCheck_0_offset                                 (readCheckRequestVec_0_offset),
    .readCheck_0_instructionIndex                       (readCheckRequestVec_0_instructionIndex),
    .readCheck_1_vs                                     (readCheckRequestVec_1_vs),
    .readCheck_1_offset                                 (readCheckRequestVec_1_offset),
    .readCheck_1_instructionIndex                       (readCheckRequestVec_1_instructionIndex),
    .readCheck_2_vs                                     (readCheckRequestVec_2_vs),
    .readCheck_2_offset                                 (readCheckRequestVec_2_offset),
    .readCheck_2_instructionIndex                       (readCheckRequestVec_2_instructionIndex),
    .readCheck_3_vs                                     (readCheckRequestVec_3_vs),
    .readCheck_3_offset                                 (readCheckRequestVec_3_offset),
    .readCheck_3_instructionIndex                       (readCheckRequestVec_3_instructionIndex),
    .readCheck_4_vs                                     (readCheckRequestVec_4_vs),
    .readCheck_4_offset                                 (readCheckRequestVec_4_offset),
    .readCheck_4_instructionIndex                       (readCheckRequestVec_4_instructionIndex),
    .readCheck_5_vs                                     (readCheckRequestVec_5_vs),
    .readCheck_5_offset                                 (readCheckRequestVec_5_offset),
    .readCheck_5_instructionIndex                       (readCheckRequestVec_5_instructionIndex),
    .readCheck_6_vs                                     (readCheckRequestVec_6_vs),
    .readCheck_6_offset                                 (readCheckRequestVec_6_offset),
    .readCheck_6_instructionIndex                       (readCheckRequestVec_6_instructionIndex),
    .readCheck_7_vs                                     (readCheckRequestVec_7_vs),
    .readCheck_7_offset                                 (readCheckRequestVec_7_offset),
    .readCheck_7_instructionIndex                       (readCheckRequestVec_7_instructionIndex),
    .readCheck_8_vs                                     (readCheckRequestVec_8_vs),
    .readCheck_8_offset                                 (readCheckRequestVec_8_offset),
    .readCheck_8_instructionIndex                       (readCheckRequestVec_8_instructionIndex),
    .readCheck_9_vs                                     (readCheckRequestVec_9_vs),
    .readCheck_9_offset                                 (readCheckRequestVec_9_offset),
    .readCheck_9_instructionIndex                       (readCheckRequestVec_9_instructionIndex),
    .readCheck_10_vs                                    (readCheckRequestVec_10_vs),
    .readCheck_10_offset                                (readCheckRequestVec_10_offset),
    .readCheck_10_instructionIndex                      (readCheckRequestVec_10_instructionIndex),
    .readCheck_11_vs                                    (readCheckRequestVec_11_vs),
    .readCheck_11_offset                                (readCheckRequestVec_11_offset),
    .readCheck_11_instructionIndex                      (readCheckRequestVec_11_instructionIndex),
    .readCheck_12_vs                                    (readCheckRequestVec_12_vs),
    .readCheck_12_offset                                (readCheckRequestVec_12_offset),
    .readCheck_12_instructionIndex                      (readCheckRequestVec_12_instructionIndex),
    .readCheck_13_vs                                    (readCheckRequestVec_13_vs),
    .readCheck_13_offset                                (readCheckRequestVec_13_offset),
    .readCheck_13_instructionIndex                      (readCheckRequestVec_13_instructionIndex),
    .readCheckResult_0                                  (readCheckResult_0),
    .readCheckResult_1                                  (readCheckResult_1),
    .readCheckResult_2                                  (readCheckResult_2),
    .readCheckResult_3                                  (readCheckResult_3),
    .readCheckResult_4                                  (readCheckResult_4),
    .readCheckResult_5                                  (readCheckResult_5),
    .readCheckResult_6                                  (readCheckResult_6),
    .readCheckResult_7                                  (readCheckResult_7),
    .readCheckResult_8                                  (readCheckResult_8),
    .readCheckResult_9                                  (readCheckResult_9),
    .readCheckResult_10                                 (readCheckResult_10),
    .readCheckResult_11                                 (readCheckResult_11),
    .readCheckResult_12                                 (readCheckResult_12),
    .readCheckResult_13                                 (readCheckResult_13),
    .readResults_0                                      (_vrf_readResults_0),
    .readResults_1                                      (vrfReadResult_0_0),
    .readResults_2                                      (vrfReadResult_0_1),
    .readResults_3                                      (vrfReadResult_0_2),
    .readResults_4                                      (vrfReadResult_1_0),
    .readResults_5                                      (vrfReadResult_1_1),
    .readResults_6                                      (vrfReadResult_1_2),
    .readResults_7                                      (vrfReadResult_2_0),
    .readResults_8                                      (vrfReadResult_2_1),
    .readResults_9                                      (vrfReadResult_2_2),
    .readResults_10                                     (vrfReadResult_3_0),
    .readResults_11                                     (vrfReadResult_3_1),
    .readResults_12                                     (vrfReadResult_3_2),
    .readResults_13                                     (vrfReadDataChannel),
    .write_ready                                        (_vrf_write_ready),
    .write_valid                                        (_maskedWriteUnit_dequeue_valid),
    .write_bits_vd                                      (_maskedWriteUnit_dequeue_bits_vd),
    .write_bits_offset                                  (_maskedWriteUnit_dequeue_bits_offset),
    .write_bits_mask                                    (_maskedWriteUnit_dequeue_bits_mask),
    .write_bits_data                                    (_maskedWriteUnit_dequeue_bits_data),
    .write_bits_last                                    (_maskedWriteUnit_dequeue_bits_last),
    .write_bits_instructionIndex                        (_maskedWriteUnit_dequeue_bits_instructionIndex),
    .writeCheck_0_vd                                    (vrfWriteArbiter_0_bits_vd),
    .writeCheck_0_offset                                (vrfWriteArbiter_0_bits_offset),
    .writeCheck_0_instructionIndex                      (vrfWriteArbiter_0_bits_instructionIndex),
    .writeCheck_1_vd                                    (vrfWriteArbiter_1_bits_vd),
    .writeCheck_1_offset                                (vrfWriteArbiter_1_bits_offset),
    .writeCheck_1_instructionIndex                      (vrfWriteArbiter_1_bits_instructionIndex),
    .writeCheck_2_vd                                    (vrfWriteArbiter_2_bits_vd),
    .writeCheck_2_offset                                (vrfWriteArbiter_2_bits_offset),
    .writeCheck_2_instructionIndex                      (vrfWriteArbiter_2_bits_instructionIndex),
    .writeCheck_3_vd                                    (vrfWriteArbiter_3_bits_vd),
    .writeCheck_3_offset                                (vrfWriteArbiter_3_bits_offset),
    .writeCheck_3_instructionIndex                      (vrfWriteArbiter_3_bits_instructionIndex),
    .writeCheck_4_vd                                    (vrfWriteArbiter_4_bits_vd),
    .writeCheck_4_offset                                (vrfWriteArbiter_4_bits_offset),
    .writeCheck_4_instructionIndex                      (vrfWriteArbiter_4_bits_instructionIndex),
    .writeCheck_5_vd                                    (crossLaneWriteQueue_0_deq_bits_vd),
    .writeCheck_5_offset                                (crossLaneWriteQueue_0_deq_bits_offset),
    .writeCheck_5_instructionIndex                      (crossLaneWriteQueue_0_deq_bits_instructionIndex),
    .writeCheck_6_vd                                    (crossLaneWriteQueue_1_deq_bits_vd),
    .writeCheck_6_offset                                (crossLaneWriteQueue_1_deq_bits_offset),
    .writeCheck_6_instructionIndex                      (crossLaneWriteQueue_1_deq_bits_instructionIndex),
    .writeAllow_0                                       (_vrf_writeAllow_0),
    .writeAllow_1                                       (_vrf_writeAllow_1),
    .writeAllow_2                                       (_vrf_writeAllow_2),
    .writeAllow_3                                       (_vrf_writeAllow_3),
    .writeAllow_4                                       (_vrf_writeAllow_4),
    .writeAllow_5                                       (_vrf_writeAllow_5),
    .writeAllow_6                                       (_vrf_writeAllow_6),
    .instructionWriteReport_valid                       (_GEN_10),
    .instructionWriteReport_bits_vd_valid               (~laneRequest_bits_decodeResult_targetRd_0 | _GEN_11),
    .instructionWriteReport_bits_vd_bits                (laneRequest_bits_vd_0),
    .instructionWriteReport_bits_vs1_valid              (laneRequest_bits_decodeResult_vtype_0),
    .instructionWriteReport_bits_vs1_bits               (laneRequest_bits_vs1_0),
    .instructionWriteReport_bits_vs2                    (laneRequest_bits_vs2_0),
    .instructionWriteReport_bits_instIndex              (laneRequest_bits_instructionIndex_0),
    .instructionWriteReport_bits_ls                     (laneRequest_bits_loadStore_0),
    .instructionWriteReport_bits_st                     (laneRequest_bits_store_0),
    .instructionWriteReport_bits_gather                 (laneRequest_bits_decodeResult_gather_0 & laneRequest_bits_decodeResult_vtype_0),
    .instructionWriteReport_bits_gather16               (laneRequest_bits_decodeResult_gather16_0),
    .instructionWriteReport_bits_crossWrite             (laneRequest_bits_decodeResult_crossWrite_0),
    .instructionWriteReport_bits_crossRead              (laneRequest_bits_decodeResult_crossRead_0),
    .instructionWriteReport_bits_indexType              (laneRequest_valid_0 & laneRequest_bits_loadStore_0),
    .instructionWriteReport_bits_ma                     (laneRequest_bits_decodeResult_multiplier_0 & ^(laneRequest_bits_decodeResult_uop_0[1:0]) & ~laneRequest_bits_decodeResult_vwmacc_0),
    .instructionWriteReport_bits_onlyRead               (laneRequest_bits_decodeResult_popCount_0),
    .instructionWriteReport_bits_slow                   (laneRequest_bits_decodeResult_special_0),
    .instructionWriteReport_bits_elementMask            (selectMask),
    .instructionWriteReport_bits_state_stFinish         (~laneRequest_bits_loadStore_0),
    .instructionWriteReport_bits_state_wWriteQueueClear (~_GEN_11),
    .instructionWriteReport_bits_state_wLaneLastReport  (~laneRequest_valid_0),
    .instructionWriteReport_bits_state_wTopLastReport   (~laneRequest_bits_decodeResult_maskUnit_0),
    .instructionLastReport                              (instructionFinishInSlot),
    .lsuLastReport                                      (lsuLastReport),
    .vrfSlotRelease                                     (_vrf_vrfSlotRelease),
    .dataInLane                                         (instructionValid),
    .loadDataInLSUWriteQueue                            (loadDataInLSUWriteQueue)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) crossLaneWriteQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(crossLaneWriteQueue_0_enq_ready & crossLaneWriteQueue_0_enq_valid)),
    .pop_req_n    (~(crossLaneWriteQueue_0_deq_ready & ~_crossLaneWriteQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (crossLaneWriteQueue_dataIn),
    .empty        (_crossLaneWriteQueue_fifo_empty),
    .almost_empty (crossLaneWriteQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (crossLaneWriteQueue_0_almostFull),
    .full         (_crossLaneWriteQueue_fifo_full),
    .error        (_crossLaneWriteQueue_fifo_error),
    .data_out     (_crossLaneWriteQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(51)
  ) crossLaneWriteQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(crossLaneWriteQueue_1_enq_ready & crossLaneWriteQueue_1_enq_valid)),
    .pop_req_n    (~(crossLaneWriteQueue_1_deq_ready & ~_crossLaneWriteQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (crossLaneWriteQueue_dataIn_1),
    .empty        (_crossLaneWriteQueue_fifo_1_empty),
    .almost_empty (crossLaneWriteQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (crossLaneWriteQueue_1_almostFull),
    .full         (_crossLaneWriteQueue_fifo_1_full),
    .error        (_crossLaneWriteQueue_fifo_1_error),
    .data_out     (_crossLaneWriteQueue_fifo_1_data_out)
  );
  MaskedWrite maskedWriteUnit (
    .clock                                (clock),
    .reset                                (reset),
    .enqueue_ready                        (queueBeforeMaskWrite_deq_ready),
    .enqueue_valid                        (queueBeforeMaskWrite_deq_valid),
    .enqueue_bits_vd                      (queueBeforeMaskWrite_deq_bits_vd),
    .enqueue_bits_offset                  (queueBeforeMaskWrite_deq_bits_offset),
    .enqueue_bits_mask                    (queueBeforeMaskWrite_deq_bits_mask),
    .enqueue_bits_data                    (queueBeforeMaskWrite_deq_bits_data),
    .enqueue_bits_last                    (queueBeforeMaskWrite_deq_bits_last),
    .enqueue_bits_instructionIndex        (queueBeforeMaskWrite_deq_bits_instructionIndex),
    .dequeue_ready                        (_vrf_write_ready),
    .dequeue_valid                        (_maskedWriteUnit_dequeue_valid),
    .dequeue_bits_vd                      (_maskedWriteUnit_dequeue_bits_vd),
    .dequeue_bits_offset                  (_maskedWriteUnit_dequeue_bits_offset),
    .dequeue_bits_mask                    (_maskedWriteUnit_dequeue_bits_mask),
    .dequeue_bits_data                    (_maskedWriteUnit_dequeue_bits_data),
    .dequeue_bits_last                    (_maskedWriteUnit_dequeue_bits_last),
    .dequeue_bits_instructionIndex        (_maskedWriteUnit_dequeue_bits_instructionIndex),
    .vrfReadRequest_ready                 (readBeforeMaskedWrite_ready),
    .vrfReadRequest_valid                 (readBeforeMaskedWrite_valid),
    .vrfReadRequest_bits_vs               (readBeforeMaskedWrite_bits_vs),
    .vrfReadRequest_bits_offset           (readBeforeMaskedWrite_bits_offset),
    .vrfReadRequest_bits_instructionIndex (readBeforeMaskedWrite_bits_instructionIndex),
    .vrfReadResult                        (_vrf_readResults_0)
  );
  SlotTokenManager tokenManager (
    .clock                                     (clock),
    .reset                                     (reset),
    .enqReports_0_valid                        (_stage0_tokenReport_valid),
    .enqReports_0_bits_decodeResult_sWrite     (_stage0_tokenReport_bits_decodeResult_sWrite),
    .enqReports_0_bits_decodeResult_crossWrite (_stage0_tokenReport_bits_decodeResult_crossWrite),
    .enqReports_0_bits_decodeResult_maskUnit   (_stage0_tokenReport_bits_decodeResult_maskUnit),
    .enqReports_0_bits_instructionIndex        (_stage0_tokenReport_bits_instructionIndex),
    .enqReports_0_bits_sSendResponse           (_stage0_tokenReport_bits_sSendResponse),
    .enqReports_1_valid                        (_stage0_1_tokenReport_valid),
    .enqReports_1_bits_decodeResult_sWrite     (_stage0_1_tokenReport_bits_decodeResult_sWrite),
    .enqReports_1_bits_decodeResult_maskUnit   (_stage0_1_tokenReport_bits_decodeResult_maskUnit),
    .enqReports_1_bits_instructionIndex        (_stage0_1_tokenReport_bits_instructionIndex),
    .enqReports_2_valid                        (_stage0_2_tokenReport_valid),
    .enqReports_2_bits_decodeResult_sWrite     (_stage0_2_tokenReport_bits_decodeResult_sWrite),
    .enqReports_2_bits_decodeResult_maskUnit   (_stage0_2_tokenReport_bits_decodeResult_maskUnit),
    .enqReports_2_bits_instructionIndex        (_stage0_2_tokenReport_bits_instructionIndex),
    .enqReports_3_valid                        (_stage0_3_tokenReport_valid),
    .enqReports_3_bits_decodeResult_sWrite     (_stage0_3_tokenReport_bits_decodeResult_sWrite),
    .enqReports_3_bits_decodeResult_maskUnit   (_stage0_3_tokenReport_bits_decodeResult_maskUnit),
    .enqReports_3_bits_instructionIndex        (_stage0_3_tokenReport_bits_instructionIndex),
    .crossWriteReports_0_valid                 (afterCheckDequeueFire_5),
    .crossWriteReports_0_bits                  (allVrfWriteAfterCheck_5_instructionIndex),
    .crossWriteReports_1_valid                 (afterCheckDequeueFire_6),
    .crossWriteReports_1_bits                  (allVrfWriteAfterCheck_6_instructionIndex),
    .responseReport_valid                      (_maskStage_maskReq_valid),
    .responseReport_bits                       (_maskStage_maskReq_bits_index),
    .responseFeedbackReport_valid              (_GEN_13 & writeFromMask),
    .responseFeedbackReport_bits               (vrfWriteChannel_bits_instructionIndex_0),
    .slotWriteReport_0_valid                   (afterCheckDequeueFire_0),
    .slotWriteReport_0_bits                    (allVrfWriteAfterCheck_0_instructionIndex),
    .slotWriteReport_1_valid                   (afterCheckDequeueFire_1),
    .slotWriteReport_1_bits                    (allVrfWriteAfterCheck_1_instructionIndex),
    .slotWriteReport_2_valid                   (afterCheckDequeueFire_2),
    .slotWriteReport_2_bits                    (allVrfWriteAfterCheck_2_instructionIndex),
    .slotWriteReport_3_valid                   (afterCheckDequeueFire_3),
    .slotWriteReport_3_bits                    (allVrfWriteAfterCheck_3_instructionIndex),
    .writePipeEnqReport_valid                  (queueBeforeMaskWrite_push),
    .writePipeEnqReport_bits                   (queueBeforeMaskWrite_enq_bits_instructionIndex),
    .writePipeDeqReport_valid                  (_vrf_write_ready & _maskedWriteUnit_dequeue_valid),
    .writePipeDeqReport_bits                   (_maskedWriteUnit_dequeue_bits_instructionIndex),
    .topWriteEnq_valid                         (_GEN_13),
    .topWriteEnq_bits                          (vrfWriteChannel_bits_instructionIndex_0),
    .topWriteDeq_valid                         (afterCheckDequeueFire_4),
    .topWriteDeq_bits                          (allVrfWriteAfterCheck_4_instructionIndex),
    .instructionValid                          (_tokenManager_instructionValid),
    .dataInWritePipe                           (writeQueueValid),
    .maskUnitLastReport                        (lsuLastReport)
  );
  LaneStage0 stage0 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage0_enqueue_ready),
    .enqueue_valid                                   (stage0_enqueue_valid),
    .enqueue_bits_maskIndex                          (maskIndexVec_0),
    .enqueue_bits_maskForMaskGroup                   (slotControl_0_mask_bits),
    .enqueue_bits_maskGroupCount                     (maskGroupCountVec_0),
    .enqueue_bits_readFromScalar                     (slotControl_0_laneRequest_readFromScalar),
    .enqueue_bits_vSew1H                             (laneState_vSew1H),
    .enqueue_bits_loadStore                          (laneState_loadStore),
    .enqueue_bits_laneIndex                          (laneState_laneIndex),
    .enqueue_bits_decodeResult_specialSlot           (laneState_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (laneState_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (laneState_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (laneState_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (laneState_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (laneState_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (laneState_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (laneState_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (laneState_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (laneState_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (laneState_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (laneState_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (laneState_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (laneState_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (laneState_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (laneState_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (laneState_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (laneState_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (laneState_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (laneState_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (laneState_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (laneState_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (laneState_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (laneState_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (laneState_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (laneState_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (laneState_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (laneState_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (laneState_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (laneState_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (laneState_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (laneState_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (laneState_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (laneState_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (laneState_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (laneState_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (laneState_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (laneState_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (laneState_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (laneState_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (laneState_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (laneState_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (laneState_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (laneState_decodeResult_logic),
    .enqueue_bits_lastGroupForInstruction            (laneState_lastGroupForInstruction),
    .enqueue_bits_isLastLaneForInstruction           (laneState_isLastLaneForInstruction),
    .enqueue_bits_instructionFinished                (laneState_instructionFinished),
    .enqueue_bits_csr_vl                             (laneState_csr_vl),
    .enqueue_bits_csr_vStart                         (laneState_csr_vStart),
    .enqueue_bits_csr_vlmul                          (laneState_csr_vlmul),
    .enqueue_bits_csr_vSew                           (laneState_csr_vSew),
    .enqueue_bits_csr_vxrm                           (laneState_csr_vxrm),
    .enqueue_bits_csr_vta                            (laneState_csr_vta),
    .enqueue_bits_csr_vma                            (laneState_csr_vma),
    .enqueue_bits_maskType                           (laneState_maskType),
    .enqueue_bits_maskNotMaskedElement               (laneState_maskNotMaskedElement),
    .enqueue_bits_vs1                                (laneState_vs1),
    .enqueue_bits_vs2                                (laneState_vs2),
    .enqueue_bits_vd                                 (laneState_vd),
    .enqueue_bits_instructionIndex                   (laneState_instructionIndex),
    .enqueue_bits_additionalRW                       (laneState_additionalRW),
    .enqueue_bits_skipRead                           (laneState_skipRead),
    .enqueue_bits_skipEnable                         (laneState_skipEnable),
    .dequeue_ready                                   (_stage1_enqueue_ready),
    .dequeue_valid                                   (_stage0_dequeue_valid),
    .dequeue_bits_maskForMaskInput                   (_stage0_dequeue_bits_maskForMaskInput),
    .dequeue_bits_boundaryMaskCorrection             (_stage0_dequeue_bits_boundaryMaskCorrection),
    .dequeue_bits_sSendResponse                      (_stage0_dequeue_bits_sSendResponse),
    .dequeue_bits_groupCounter                       (_stage0_dequeue_bits_groupCounter),
    .dequeue_bits_readFromScalar                     (_stage0_dequeue_bits_readFromScalar),
    .dequeue_bits_instructionIndex                   (_stage0_dequeue_bits_instructionIndex),
    .dequeue_bits_decodeResult_specialSlot           (_stage0_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage0_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage0_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage0_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage0_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage0_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage0_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage0_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage0_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage0_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage0_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage0_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage0_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage0_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage0_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage0_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage0_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage0_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage0_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage0_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage0_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage0_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage0_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage0_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage0_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage0_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage0_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage0_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage0_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage0_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage0_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage0_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage0_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage0_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage0_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage0_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage0_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage0_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage0_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage0_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage0_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage0_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage0_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage0_dequeue_bits_decodeResult_logic),
    .dequeue_bits_laneIndex                          (_stage0_dequeue_bits_laneIndex),
    .dequeue_bits_skipRead                           (_stage0_dequeue_bits_skipRead),
    .dequeue_bits_vs1                                (_stage0_dequeue_bits_vs1),
    .dequeue_bits_vs2                                (_stage0_dequeue_bits_vs2),
    .dequeue_bits_vd                                 (_stage0_dequeue_bits_vd),
    .dequeue_bits_vSew1H                             (_stage0_dequeue_bits_vSew1H),
    .dequeue_bits_maskNotMaskedElement               (_stage0_dequeue_bits_maskNotMaskedElement),
    .dequeue_bits_csr_vl                             (_stage0_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage0_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage0_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage0_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage0_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage0_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage0_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage0_dequeue_bits_maskType),
    .dequeue_bits_loadStore                          (_stage0_dequeue_bits_loadStore),
    .dequeue_bits_bordersForMaskLogic                (_stage0_dequeue_bits_bordersForMaskLogic),
    .updateLaneState_maskGroupCount                  (_stage0_updateLaneState_maskGroupCount),
    .updateLaneState_maskIndex                       (_stage0_updateLaneState_maskIndex),
    .updateLaneState_outOfExecutionRange             (_stage0_updateLaneState_outOfExecutionRange),
    .updateLaneState_maskExhausted                   (_stage0_updateLaneState_maskExhausted),
    .tokenReport_valid                               (_stage0_tokenReport_valid),
    .tokenReport_bits_decodeResult_sWrite            (_stage0_tokenReport_bits_decodeResult_sWrite),
    .tokenReport_bits_decodeResult_crossWrite        (_stage0_tokenReport_bits_decodeResult_crossWrite),
    .tokenReport_bits_decodeResult_maskUnit          (_stage0_tokenReport_bits_decodeResult_maskUnit),
    .tokenReport_bits_instructionIndex               (_stage0_tokenReport_bits_instructionIndex),
    .tokenReport_bits_sSendResponse                  (_stage0_tokenReport_bits_sSendResponse)
  );
  LaneStage1 stage1 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage1_enqueue_ready),
    .enqueue_valid                                   (_stage0_dequeue_valid),
    .enqueue_bits_groupCounter                       (_stage0_dequeue_bits_groupCounter),
    .enqueue_bits_maskForMaskInput                   (_stage0_dequeue_bits_maskForMaskInput),
    .enqueue_bits_boundaryMaskCorrection             (_stage0_dequeue_bits_boundaryMaskCorrection),
    .enqueue_bits_sSendResponse                      (_stage0_dequeue_bits_sSendResponse),
    .enqueue_bits_instructionIndex                   (_stage0_dequeue_bits_instructionIndex),
    .enqueue_bits_decodeResult_specialSlot           (_stage0_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage0_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage0_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage0_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage0_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage0_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage0_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage0_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage0_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage0_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage0_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage0_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage0_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage0_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage0_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage0_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage0_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage0_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage0_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage0_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage0_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage0_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage0_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage0_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage0_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage0_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage0_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage0_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage0_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage0_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage0_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage0_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage0_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage0_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage0_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage0_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage0_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage0_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage0_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage0_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage0_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage0_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage0_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage0_dequeue_bits_decodeResult_logic),
    .enqueue_bits_laneIndex                          (_stage0_dequeue_bits_laneIndex),
    .enqueue_bits_skipRead                           (_stage0_dequeue_bits_skipRead),
    .enqueue_bits_vs1                                (_stage0_dequeue_bits_vs1),
    .enqueue_bits_vs2                                (_stage0_dequeue_bits_vs2),
    .enqueue_bits_vd                                 (_stage0_dequeue_bits_vd),
    .enqueue_bits_vSew1H                             (_stage0_dequeue_bits_vSew1H),
    .enqueue_bits_maskNotMaskedElement               (_stage0_dequeue_bits_maskNotMaskedElement),
    .enqueue_bits_csr_vl                             (_stage0_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage0_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage0_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage0_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage0_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage0_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage0_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage0_dequeue_bits_maskType),
    .enqueue_bits_loadStore                          (_stage0_dequeue_bits_loadStore),
    .enqueue_bits_readFromScalar                     (_stage0_dequeue_bits_readFromScalar),
    .enqueue_bits_bordersForMaskLogic                (_stage0_dequeue_bits_bordersForMaskLogic),
    .dequeue_ready                                   (_stage2_enqueue_ready & _executionUnit_enqueue_ready),
    .dequeue_valid                                   (_stage1_dequeue_valid),
    .dequeue_bits_readBusDequeueGroup                (readBusDequeueGroup),
    .dequeue_bits_maskForFilter                      (_stage1_dequeue_bits_maskForFilter),
    .dequeue_bits_mask                               (_stage1_dequeue_bits_mask),
    .dequeue_bits_groupCounter                       (_stage1_dequeue_bits_groupCounter),
    .dequeue_bits_sSendResponse                      (_stage1_dequeue_bits_sSendResponse),
    .dequeue_bits_src_0                              (_stage1_dequeue_bits_src_0),
    .dequeue_bits_src_1                              (_stage1_dequeue_bits_src_1),
    .dequeue_bits_src_2                              (_stage1_dequeue_bits_src_2),
    .dequeue_bits_crossReadSource                    (_stage1_dequeue_bits_crossReadSource),
    .dequeue_bits_decodeResult_specialSlot           (_stage1_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage1_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage1_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage1_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage1_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage1_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage1_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage1_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage1_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage1_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage1_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage1_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage1_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage1_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage1_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage1_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage1_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage1_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage1_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage1_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage1_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage1_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage1_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage1_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage1_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage1_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage1_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage1_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage1_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage1_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage1_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage1_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage1_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage1_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage1_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage1_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage1_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage1_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage1_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage1_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage1_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage1_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage1_dequeue_bits_decodeResult_logic),
    .dequeue_bits_vSew1H                             (_stage1_dequeue_bits_vSew1H),
    .dequeue_bits_csr_vl                             (_stage1_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage1_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage1_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage1_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage1_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage1_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage1_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage1_dequeue_bits_maskType),
    .dequeue_bits_laneIndex                          (_stage1_dequeue_bits_laneIndex),
    .dequeue_bits_instructionIndex                   (_stage1_dequeue_bits_instructionIndex),
    .dequeue_bits_loadStore                          (_stage1_dequeue_bits_loadStore),
    .dequeue_bits_vd                                 (_stage1_dequeue_bits_vd),
    .dequeue_bits_bordersForMaskLogic                (_stage1_dequeue_bits_bordersForMaskLogic),
    .vrfReadRequest_0_ready                          (vrfReadRequest_0_0_ready),
    .vrfReadRequest_0_valid                          (vrfReadRequest_0_0_valid),
    .vrfReadRequest_0_bits_vs                        (vrfReadRequest_0_0_bits_vs),
    .vrfReadRequest_0_bits_readSource                (vrfReadRequest_0_0_bits_readSource),
    .vrfReadRequest_0_bits_offset                    (vrfReadRequest_0_0_bits_offset),
    .vrfReadRequest_0_bits_instructionIndex          (vrfReadRequest_0_0_bits_instructionIndex),
    .vrfReadRequest_1_ready                          (vrfReadRequest_0_1_ready),
    .vrfReadRequest_1_valid                          (vrfReadRequest_0_1_valid),
    .vrfReadRequest_1_bits_vs                        (vrfReadRequest_0_1_bits_vs),
    .vrfReadRequest_1_bits_readSource                (vrfReadRequest_0_1_bits_readSource),
    .vrfReadRequest_1_bits_offset                    (vrfReadRequest_0_1_bits_offset),
    .vrfReadRequest_1_bits_instructionIndex          (vrfReadRequest_0_1_bits_instructionIndex),
    .vrfReadRequest_2_ready                          (vrfReadRequest_0_2_ready),
    .vrfReadRequest_2_valid                          (vrfReadRequest_0_2_valid),
    .vrfReadRequest_2_bits_vs                        (vrfReadRequest_0_2_bits_vs),
    .vrfReadRequest_2_bits_readSource                (vrfReadRequest_0_2_bits_readSource),
    .vrfReadRequest_2_bits_offset                    (vrfReadRequest_0_2_bits_offset),
    .vrfReadRequest_2_bits_instructionIndex          (vrfReadRequest_0_2_bits_instructionIndex),
    .vrfCheckRequest_0_vs                            (readCheckRequestVec_9_vs),
    .vrfCheckRequest_0_readSource                    (readCheckRequestVec_9_readSource),
    .vrfCheckRequest_0_offset                        (readCheckRequestVec_9_offset),
    .vrfCheckRequest_0_instructionIndex              (readCheckRequestVec_9_instructionIndex),
    .vrfCheckRequest_1_vs                            (readCheckRequestVec_10_vs),
    .vrfCheckRequest_1_readSource                    (readCheckRequestVec_10_readSource),
    .vrfCheckRequest_1_offset                        (readCheckRequestVec_10_offset),
    .vrfCheckRequest_1_instructionIndex              (readCheckRequestVec_10_instructionIndex),
    .vrfCheckRequest_2_vs                            (readCheckRequestVec_11_vs),
    .vrfCheckRequest_2_readSource                    (readCheckRequestVec_11_readSource),
    .vrfCheckRequest_2_offset                        (readCheckRequestVec_11_offset),
    .vrfCheckRequest_2_instructionIndex              (readCheckRequestVec_11_instructionIndex),
    .vrfCheckRequest_3_vs                            (readCheckRequestVec_12_vs),
    .vrfCheckRequest_3_readSource                    (readCheckRequestVec_12_readSource),
    .vrfCheckRequest_3_offset                        (readCheckRequestVec_12_offset),
    .vrfCheckRequest_3_instructionIndex              (readCheckRequestVec_12_instructionIndex),
    .vrfCheckRequest_4_vs                            (readCheckRequestVec_13_vs),
    .vrfCheckRequest_4_readSource                    (readCheckRequestVec_13_readSource),
    .vrfCheckRequest_4_offset                        (readCheckRequestVec_13_offset),
    .vrfCheckRequest_4_instructionIndex              (readCheckRequestVec_13_instructionIndex),
    .checkResult_0                                   (readCheckResult_9),
    .checkResult_1                                   (readCheckResult_10),
    .checkResult_2                                   (readCheckResult_11),
    .checkResult_3                                   (readCheckResult_12),
    .checkResult_4                                   (readCheckResult_13),
    .vrfReadResult_0                                 (vrfReadResult_0_0),
    .vrfReadResult_1                                 (vrfReadResult_0_1),
    .vrfReadResult_2                                 (vrfReadResult_0_2),
    .readBusDequeue_0_ready                          (queue_deq_ready),
    .readBusDequeue_0_valid                          (queue_deq_valid),
    .readBusDequeue_0_bits_data                      (queue_deq_bits_data),
    .readBusDequeue_1_ready                          (queue_1_deq_ready),
    .readBusDequeue_1_valid                          (queue_1_deq_valid),
    .readBusDequeue_1_bits_data                      (queue_1_deq_bits_data),
    .readBusRequest_0_ready                          (tokenReady),
    .readBusRequest_0_valid                          (_stage1_readBusRequest_0_valid),
    .readBusRequest_0_bits_data                      (readBusPort_0_deq_bits_data_0),
    .readBusRequest_1_ready                          (tokenReady_1),
    .readBusRequest_1_valid                          (_stage1_readBusRequest_1_valid),
    .readBusRequest_1_bits_data                      (readBusPort_1_deq_bits_data_0)
  );
  LaneStage2 stage2 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage2_enqueue_ready),
    .enqueue_valid                                   (_stage1_dequeue_valid & _executionUnit_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_dequeue_bits_src_2),
    .enqueue_bits_groupCounter                       (_stage1_dequeue_bits_groupCounter),
    .enqueue_bits_maskForFilter                      (_stage1_dequeue_bits_maskForFilter),
    .enqueue_bits_mask                               (_stage1_dequeue_bits_mask),
    .enqueue_bits_sSendResponse                      (_stage1_dequeue_bits_sSendResponse),
    .enqueue_bits_bordersForMaskLogic                (_stage1_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_dequeue_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (_stage1_dequeue_bits_instructionIndex),
    .enqueue_bits_loadStore                          (_stage1_dequeue_bits_loadStore),
    .enqueue_bits_vd                                 (_stage1_dequeue_bits_vd),
    .enqueue_bits_csr_vl                             (_stage1_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_dequeue_bits_csr_vma),
    .enqueue_bits_vSew1H                             (_stage1_dequeue_bits_vSew1H),
    .enqueue_bits_maskType                           (_stage1_dequeue_bits_maskType),
    .dequeue_ready                                   (stage3EnqWire_ready & _executionUnit_dequeue_valid),
    .dequeue_valid                                   (_stage2_dequeue_valid),
    .dequeue_bits_groupCounter                       (stage3EnqWire_bits_groupCounter),
    .dequeue_bits_mask                               (stage3EnqWire_bits_mask),
    .dequeue_bits_sSendResponse                      (stage3EnqWire_bits_sSendResponse),
    .dequeue_bits_pipeData                           (stage3EnqWire_bits_pipeData),
    .dequeue_bits_decodeResult_specialSlot           (stage3EnqWire_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (stage3EnqWire_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (stage3EnqWire_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (stage3EnqWire_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (stage3EnqWire_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (stage3EnqWire_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (stage3EnqWire_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (stage3EnqWire_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (stage3EnqWire_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (stage3EnqWire_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (stage3EnqWire_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (stage3EnqWire_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (stage3EnqWire_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (stage3EnqWire_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (stage3EnqWire_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (stage3EnqWire_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (stage3EnqWire_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (stage3EnqWire_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (stage3EnqWire_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (stage3EnqWire_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (stage3EnqWire_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (stage3EnqWire_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (stage3EnqWire_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (stage3EnqWire_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (stage3EnqWire_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (stage3EnqWire_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (stage3EnqWire_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (stage3EnqWire_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (stage3EnqWire_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (stage3EnqWire_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (stage3EnqWire_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (stage3EnqWire_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (stage3EnqWire_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (stage3EnqWire_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (stage3EnqWire_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (stage3EnqWire_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (stage3EnqWire_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (stage3EnqWire_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (stage3EnqWire_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (stage3EnqWire_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (stage3EnqWire_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (stage3EnqWire_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (stage3EnqWire_bits_decodeResult_logic),
    .dequeue_bits_instructionIndex                   (stage3EnqWire_bits_instructionIndex),
    .dequeue_bits_loadStore                          (stage3EnqWire_bits_loadStore),
    .dequeue_bits_vd                                 (stage3EnqWire_bits_vd)
  );
  LaneExecutionBridge executionUnit (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_executionUnit_enqueue_ready),
    .enqueue_valid                                   (_stage1_dequeue_valid & _stage2_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_dequeue_bits_src_2),
    .enqueue_bits_crossReadSource                    (_stage1_dequeue_bits_crossReadSource),
    .enqueue_bits_bordersForMaskLogic                (_stage1_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_mask                               (_stage1_dequeue_bits_mask),
    .enqueue_bits_maskForFilter                      (_stage1_dequeue_bits_maskForFilter),
    .enqueue_bits_groupCounter                       (_stage1_dequeue_bits_groupCounter),
    .enqueue_bits_sSendResponse                      (_stage1_dequeue_bits_sSendResponse),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_dequeue_bits_decodeResult_logic),
    .enqueue_bits_vSew1H                             (_stage1_dequeue_bits_vSew1H),
    .enqueue_bits_csr_vl                             (_stage1_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage1_dequeue_bits_maskType),
    .enqueue_bits_laneIndex                          (_stage1_dequeue_bits_laneIndex),
    .enqueue_bits_instructionIndex                   (_stage1_dequeue_bits_instructionIndex),
    .dequeue_ready                                   (stage3EnqWire_ready),
    .dequeue_valid                                   (_executionUnit_dequeue_valid),
    .dequeue_bits_data                               (stage3EnqWire_bits_data),
    .dequeue_bits_ffoIndex                           (stage3EnqWire_bits_ffoIndex),
    .dequeue_bits_crossWriteData_0                   (stage3EnqWire_bits_crossWriteData_0),
    .dequeue_bits_crossWriteData_1                   (stage3EnqWire_bits_crossWriteData_1),
    .dequeue_bits_ffoSuccess                         (stage3EnqWire_bits_ffoSuccess),
    .vfuRequest_ready                                (executeEnqueueFire_0),
    .vfuRequest_valid                                (_executionUnit_vfuRequest_valid),
    .vfuRequest_bits_src_0                           (requestVec_0_src_0),
    .vfuRequest_bits_src_1                           (requestVec_0_src_1),
    .vfuRequest_bits_src_2                           (requestVec_0_src_2),
    .vfuRequest_bits_src_3                           (requestVec_0_src_3),
    .vfuRequest_bits_opcode                          (requestVec_0_opcode),
    .vfuRequest_bits_mask                            (requestVec_0_mask),
    .vfuRequest_bits_executeMask                     (requestVec_0_executeMask),
    .vfuRequest_bits_sign0                           (requestVec_0_sign0),
    .vfuRequest_bits_sign                            (requestVec_0_sign),
    .vfuRequest_bits_reverse                         (requestVec_0_reverse),
    .vfuRequest_bits_average                         (requestVec_0_average),
    .vfuRequest_bits_saturate                        (requestVec_0_saturate),
    .vfuRequest_bits_vxrm                            (requestVec_0_vxrm),
    .vfuRequest_bits_vSew                            (requestVec_0_vSew),
    .vfuRequest_bits_shifterSize                     (requestVec_0_shifterSize),
    .vfuRequest_bits_rem                             (requestVec_0_rem),
    .vfuRequest_bits_executeIndex                    (requestVec_0_executeIndex),
    .vfuRequest_bits_popInit                         (requestVec_0_popInit),
    .vfuRequest_bits_groupIndex                      (requestVec_0_groupIndex),
    .vfuRequest_bits_laneIndex                       (requestVec_0_laneIndex),
    .vfuRequest_bits_maskType                        (requestVec_0_maskType),
    .vfuRequest_bits_narrow                          (requestVec_0_narrow),
    .dataResponse_valid                              (responseVec_0_valid),
    .dataResponse_bits_data                          (responseVec_0_bits_data),
    .dataResponse_bits_executeIndex                  (responseVec_0_bits_executeIndex),
    .dataResponse_bits_ffoSuccess                    (responseVec_0_bits_ffoSuccess),
    .dataResponse_bits_adderMaskResp                 (responseVec_0_bits_adderMaskResp),
    .executeDecode_specialSlot                       (executeDecodeVec_0_specialSlot),
    .executeDecode_topUop                            (executeDecodeVec_0_topUop),
    .executeDecode_popCount                          (executeDecodeVec_0_popCount),
    .executeDecode_ffo                               (executeDecodeVec_0_ffo),
    .executeDecode_average                           (executeDecodeVec_0_average),
    .executeDecode_reverse                           (executeDecodeVec_0_reverse),
    .executeDecode_dontNeedExecuteInLane             (executeDecodeVec_0_dontNeedExecuteInLane),
    .executeDecode_scheduler                         (executeDecodeVec_0_scheduler),
    .executeDecode_sReadVD                           (executeDecodeVec_0_sReadVD),
    .executeDecode_vtype                             (executeDecodeVec_0_vtype),
    .executeDecode_sWrite                            (executeDecodeVec_0_sWrite),
    .executeDecode_crossRead                         (executeDecodeVec_0_crossRead),
    .executeDecode_crossWrite                        (executeDecodeVec_0_crossWrite),
    .executeDecode_maskUnit                          (executeDecodeVec_0_maskUnit),
    .executeDecode_special                           (executeDecodeVec_0_special),
    .executeDecode_saturate                          (executeDecodeVec_0_saturate),
    .executeDecode_vwmacc                            (executeDecodeVec_0_vwmacc),
    .executeDecode_readOnly                          (executeDecodeVec_0_readOnly),
    .executeDecode_maskSource                        (executeDecodeVec_0_maskSource),
    .executeDecode_maskDestination                   (executeDecodeVec_0_maskDestination),
    .executeDecode_maskLogic                         (executeDecodeVec_0_maskLogic),
    .executeDecode_uop                               (executeDecodeVec_0_uop),
    .executeDecode_iota                              (executeDecodeVec_0_iota),
    .executeDecode_mv                                (executeDecodeVec_0_mv),
    .executeDecode_extend                            (executeDecodeVec_0_extend),
    .executeDecode_unOrderWrite                      (executeDecodeVec_0_unOrderWrite),
    .executeDecode_compress                          (executeDecodeVec_0_compress),
    .executeDecode_gather16                          (executeDecodeVec_0_gather16),
    .executeDecode_gather                            (executeDecodeVec_0_gather),
    .executeDecode_slid                              (executeDecodeVec_0_slid),
    .executeDecode_targetRd                          (executeDecodeVec_0_targetRd),
    .executeDecode_widenReduce                       (executeDecodeVec_0_widenReduce),
    .executeDecode_red                               (executeDecodeVec_0_red),
    .executeDecode_nr                                (executeDecodeVec_0_nr),
    .executeDecode_itype                             (executeDecodeVec_0_itype),
    .executeDecode_unsigned1                         (executeDecodeVec_0_unsigned1),
    .executeDecode_unsigned0                         (executeDecodeVec_0_unsigned0),
    .executeDecode_other                             (executeDecodeVec_0_other),
    .executeDecode_multiCycle                        (executeDecodeVec_0_multiCycle),
    .executeDecode_divider                           (executeDecodeVec_0_divider),
    .executeDecode_multiplier                        (executeDecodeVec_0_multiplier),
    .executeDecode_shift                             (executeDecodeVec_0_shift),
    .executeDecode_adder                             (executeDecodeVec_0_adder),
    .executeDecode_logic                             (executeDecodeVec_0_logic),
    .responseDecode_specialSlot                      (responseDecodeVec_0_specialSlot),
    .responseDecode_topUop                           (responseDecodeVec_0_topUop),
    .responseDecode_popCount                         (responseDecodeVec_0_popCount),
    .responseDecode_ffo                              (responseDecodeVec_0_ffo),
    .responseDecode_average                          (responseDecodeVec_0_average),
    .responseDecode_reverse                          (responseDecodeVec_0_reverse),
    .responseDecode_dontNeedExecuteInLane            (responseDecodeVec_0_dontNeedExecuteInLane),
    .responseDecode_scheduler                        (responseDecodeVec_0_scheduler),
    .responseDecode_sReadVD                          (responseDecodeVec_0_sReadVD),
    .responseDecode_vtype                            (responseDecodeVec_0_vtype),
    .responseDecode_sWrite                           (responseDecodeVec_0_sWrite),
    .responseDecode_crossRead                        (responseDecodeVec_0_crossRead),
    .responseDecode_crossWrite                       (responseDecodeVec_0_crossWrite),
    .responseDecode_maskUnit                         (responseDecodeVec_0_maskUnit),
    .responseDecode_special                          (responseDecodeVec_0_special),
    .responseDecode_saturate                         (responseDecodeVec_0_saturate),
    .responseDecode_vwmacc                           (responseDecodeVec_0_vwmacc),
    .responseDecode_readOnly                         (responseDecodeVec_0_readOnly),
    .responseDecode_maskSource                       (responseDecodeVec_0_maskSource),
    .responseDecode_maskDestination                  (responseDecodeVec_0_maskDestination),
    .responseDecode_maskLogic                        (responseDecodeVec_0_maskLogic),
    .responseDecode_uop                              (responseDecodeVec_0_uop),
    .responseDecode_iota                             (responseDecodeVec_0_iota),
    .responseDecode_mv                               (responseDecodeVec_0_mv),
    .responseDecode_extend                           (responseDecodeVec_0_extend),
    .responseDecode_unOrderWrite                     (responseDecodeVec_0_unOrderWrite),
    .responseDecode_compress                         (responseDecodeVec_0_compress),
    .responseDecode_gather16                         (responseDecodeVec_0_gather16),
    .responseDecode_gather                           (responseDecodeVec_0_gather),
    .responseDecode_slid                             (responseDecodeVec_0_slid),
    .responseDecode_targetRd                         (responseDecodeVec_0_targetRd),
    .responseDecode_widenReduce                      (responseDecodeVec_0_widenReduce),
    .responseDecode_red                              (responseDecodeVec_0_red),
    .responseDecode_nr                               (responseDecodeVec_0_nr),
    .responseDecode_itype                            (responseDecodeVec_0_itype),
    .responseDecode_unsigned1                        (responseDecodeVec_0_unsigned1),
    .responseDecode_unsigned0                        (responseDecodeVec_0_unsigned0),
    .responseDecode_other                            (responseDecodeVec_0_other),
    .responseDecode_multiCycle                       (responseDecodeVec_0_multiCycle),
    .responseDecode_divider                          (responseDecodeVec_0_divider),
    .responseDecode_multiplier                       (responseDecodeVec_0_multiplier),
    .responseDecode_shift                            (responseDecodeVec_0_shift),
    .responseDecode_adder                            (responseDecodeVec_0_adder),
    .responseDecode_logic                            (responseDecodeVec_0_logic),
    .responseIndex                                   (_executionUnit_responseIndex)
  );
  MaskExchangeUnit maskStage (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (stage3EnqWire_ready),
    .enqueue_valid                                   (stage3EnqWire_valid),
    .enqueue_bits_groupCounter                       (stage3EnqWire_bits_groupCounter),
    .enqueue_bits_data                               (stage3EnqWire_bits_data),
    .enqueue_bits_pipeData                           (stage3EnqWire_bits_pipeData),
    .enqueue_bits_mask                               (stage3EnqWire_bits_mask),
    .enqueue_bits_ffoIndex                           (stage3EnqWire_bits_ffoIndex),
    .enqueue_bits_crossWriteData_0                   (stage3EnqWire_bits_crossWriteData_0),
    .enqueue_bits_crossWriteData_1                   (stage3EnqWire_bits_crossWriteData_1),
    .enqueue_bits_sSendResponse                      (stage3EnqWire_bits_sSendResponse),
    .enqueue_bits_ffoSuccess                         (stage3EnqWire_bits_ffoSuccess),
    .enqueue_bits_decodeResult_specialSlot           (stage3EnqWire_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (stage3EnqWire_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (stage3EnqWire_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (stage3EnqWire_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (stage3EnqWire_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (stage3EnqWire_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (stage3EnqWire_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (stage3EnqWire_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (stage3EnqWire_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (stage3EnqWire_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (stage3EnqWire_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (stage3EnqWire_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (stage3EnqWire_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (stage3EnqWire_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (stage3EnqWire_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (stage3EnqWire_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (stage3EnqWire_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (stage3EnqWire_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (stage3EnqWire_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (stage3EnqWire_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (stage3EnqWire_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (stage3EnqWire_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (stage3EnqWire_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (stage3EnqWire_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (stage3EnqWire_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (stage3EnqWire_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (stage3EnqWire_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (stage3EnqWire_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (stage3EnqWire_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (stage3EnqWire_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (stage3EnqWire_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (stage3EnqWire_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (stage3EnqWire_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (stage3EnqWire_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (stage3EnqWire_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (stage3EnqWire_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (stage3EnqWire_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (stage3EnqWire_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (stage3EnqWire_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (stage3EnqWire_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (stage3EnqWire_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (stage3EnqWire_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (stage3EnqWire_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (stage3EnqWire_bits_instructionIndex),
    .enqueue_bits_loadStore                          (stage3EnqWire_bits_loadStore),
    .enqueue_bits_vd                                 (stage3EnqWire_bits_vd),
    .dequeue_ready                                   (_stage3_enqueue_ready),
    .dequeue_valid                                   (_maskStage_dequeue_valid),
    .dequeue_bits_groupCounter                       (_maskStage_dequeue_bits_groupCounter),
    .dequeue_bits_data                               (_maskStage_dequeue_bits_data),
    .dequeue_bits_pipeData                           (_maskStage_dequeue_bits_pipeData),
    .dequeue_bits_mask                               (_maskStage_dequeue_bits_mask),
    .dequeue_bits_ffoIndex                           (_maskStage_dequeue_bits_ffoIndex),
    .dequeue_bits_crossWriteData_0                   (_maskStage_dequeue_bits_crossWriteData_0),
    .dequeue_bits_crossWriteData_1                   (_maskStage_dequeue_bits_crossWriteData_1),
    .dequeue_bits_sSendResponse                      (_maskStage_dequeue_bits_sSendResponse),
    .dequeue_bits_ffoSuccess                         (_maskStage_dequeue_bits_ffoSuccess),
    .dequeue_bits_decodeResult_specialSlot           (_maskStage_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_maskStage_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_maskStage_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_maskStage_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_maskStage_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_maskStage_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_maskStage_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_maskStage_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_maskStage_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_maskStage_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_maskStage_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_maskStage_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_maskStage_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_maskStage_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_maskStage_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_maskStage_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_maskStage_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_maskStage_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_maskStage_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_maskStage_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_maskStage_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_maskStage_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_maskStage_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_maskStage_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_maskStage_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_maskStage_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_maskStage_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_maskStage_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_maskStage_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_maskStage_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_maskStage_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_maskStage_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_maskStage_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_maskStage_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_maskStage_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_maskStage_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_maskStage_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_maskStage_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_maskStage_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_maskStage_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_maskStage_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_maskStage_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_maskStage_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_maskStage_dequeue_bits_decodeResult_logic),
    .dequeue_bits_instructionIndex                   (_maskStage_dequeue_bits_instructionIndex),
    .dequeue_bits_loadStore                          (_maskStage_dequeue_bits_loadStore),
    .dequeue_bits_vd                                 (_maskStage_dequeue_bits_vd),
    .maskReq_valid                                   (_maskStage_maskReq_valid),
    .maskReq_bits_source1                            (maskUnitRequest_bits_source1),
    .maskReq_bits_source2                            (maskUnitRequest_bits_source2),
    .maskReq_bits_index                              (_maskStage_maskReq_bits_index),
    .maskReq_bits_ffo                                (maskUnitRequest_bits_ffo),
    .maskRequestToLSU                                (maskRequestToLSU),
    .tokenIO_maskRequestRelease                      (tokenIO_maskRequestRelease_0)
  );
  LaneStage3 stage3 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage3_enqueue_ready),
    .enqueue_valid                                   (_maskStage_dequeue_valid),
    .enqueue_bits_groupCounter                       (_maskStage_dequeue_bits_groupCounter),
    .enqueue_bits_data                               (_maskStage_dequeue_bits_data),
    .enqueue_bits_pipeData                           (_maskStage_dequeue_bits_pipeData),
    .enqueue_bits_mask                               (_maskStage_dequeue_bits_mask),
    .enqueue_bits_ffoIndex                           (_maskStage_dequeue_bits_ffoIndex),
    .enqueue_bits_crossWriteData_0                   (_maskStage_dequeue_bits_crossWriteData_0),
    .enqueue_bits_crossWriteData_1                   (_maskStage_dequeue_bits_crossWriteData_1),
    .enqueue_bits_sSendResponse                      (_maskStage_dequeue_bits_sSendResponse),
    .enqueue_bits_ffoSuccess                         (_maskStage_dequeue_bits_ffoSuccess),
    .enqueue_bits_decodeResult_specialSlot           (_maskStage_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_maskStage_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_maskStage_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_maskStage_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_maskStage_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_maskStage_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_maskStage_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_maskStage_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_maskStage_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_maskStage_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_maskStage_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_maskStage_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_maskStage_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_maskStage_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_maskStage_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_maskStage_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_maskStage_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_maskStage_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_maskStage_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_maskStage_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_maskStage_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_maskStage_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_maskStage_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_maskStage_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_maskStage_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_maskStage_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_maskStage_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_maskStage_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_maskStage_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_maskStage_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_maskStage_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_maskStage_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_maskStage_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_maskStage_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_maskStage_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_maskStage_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_maskStage_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_maskStage_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_maskStage_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_maskStage_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_maskStage_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_maskStage_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_maskStage_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_maskStage_dequeue_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (_maskStage_dequeue_bits_instructionIndex),
    .enqueue_bits_loadStore                          (_maskStage_dequeue_bits_loadStore),
    .enqueue_bits_vd                                 (_maskStage_dequeue_bits_vd),
    .vrfWriteRequest_ready                           (vrfWriteArbiter_0_ready),
    .vrfWriteRequest_valid                           (_stage3_vrfWriteRequest_valid),
    .vrfWriteRequest_bits_vd                         (vrfWriteArbiter_0_bits_vd),
    .vrfWriteRequest_bits_offset                     (vrfWriteArbiter_0_bits_offset),
    .vrfWriteRequest_bits_mask                       (_stage3_vrfWriteRequest_bits_mask),
    .vrfWriteRequest_bits_data                       (vrfWriteArbiter_0_bits_data),
    .vrfWriteRequest_bits_last                       (vrfWriteArbiter_0_bits_last),
    .vrfWriteRequest_bits_instructionIndex           (_stage3_vrfWriteRequest_bits_instructionIndex),
    .crossWritePort_0_ready                          (tokenReady_2),
    .crossWritePort_0_valid                          (_stage3_crossWritePort_0_valid),
    .crossWritePort_0_bits_data                      (writeBusPort_0_deq_bits_data_0),
    .crossWritePort_0_bits_mask                      (writeBusPort_0_deq_bits_mask_0),
    .crossWritePort_0_bits_instructionIndex          (writeBusPort_0_deq_bits_instructionIndex_0),
    .crossWritePort_0_bits_counter                   (writeBusPort_0_deq_bits_counter_0),
    .crossWritePort_1_ready                          (tokenReady_3),
    .crossWritePort_1_valid                          (_stage3_crossWritePort_1_valid),
    .crossWritePort_1_bits_data                      (writeBusPort_1_deq_bits_data_0),
    .crossWritePort_1_bits_mask                      (writeBusPort_1_deq_bits_mask_0),
    .crossWritePort_1_bits_instructionIndex          (writeBusPort_1_deq_bits_instructionIndex_0),
    .crossWritePort_1_bits_counter                   (writeBusPort_1_deq_bits_counter_0)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_enq_ready & queue_enq_valid)),
    .pop_req_n    (~(queue_deq_ready & ~_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_enq_bits_data),
    .empty        (_queue_fifo_empty),
    .almost_empty (queue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_almostFull),
    .full         (_queue_fifo_full),
    .error        (_queue_fifo_error),
    .data_out     (queue_dataOut_data)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(queue_1_enq_ready & queue_1_enq_valid)),
    .pop_req_n    (~(queue_1_deq_ready & ~_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (queue_1_enq_bits_data),
    .empty        (_queue_fifo_1_empty),
    .almost_empty (queue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (queue_1_almostFull),
    .full         (_queue_fifo_1_full),
    .error        (_queue_fifo_1_error),
    .data_out     (queue_dataOut_1_data)
  );
  LaneStage0_1 stage0_1 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage0_1_enqueue_ready),
    .enqueue_valid                                   (stage0_1_enqueue_valid),
    .enqueue_bits_maskIndex                          (maskIndexVec_1),
    .enqueue_bits_maskForMaskGroup                   (slotControl_1_mask_bits),
    .enqueue_bits_maskGroupCount                     (maskGroupCountVec_1),
    .enqueue_bits_readFromScalar                     (slotControl_1_laneRequest_readFromScalar),
    .enqueue_bits_vSew1H                             (laneState_1_vSew1H),
    .enqueue_bits_loadStore                          (laneState_1_loadStore),
    .enqueue_bits_laneIndex                          (laneState_1_laneIndex),
    .enqueue_bits_decodeResult_specialSlot           (laneState_1_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (laneState_1_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (laneState_1_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (laneState_1_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (laneState_1_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (laneState_1_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (laneState_1_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (laneState_1_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (laneState_1_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (laneState_1_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (laneState_1_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (laneState_1_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (laneState_1_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (laneState_1_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (laneState_1_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (laneState_1_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (laneState_1_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (laneState_1_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (laneState_1_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (laneState_1_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (laneState_1_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (laneState_1_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (laneState_1_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (laneState_1_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (laneState_1_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (laneState_1_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (laneState_1_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (laneState_1_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (laneState_1_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (laneState_1_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (laneState_1_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (laneState_1_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (laneState_1_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (laneState_1_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (laneState_1_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (laneState_1_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (laneState_1_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (laneState_1_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (laneState_1_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (laneState_1_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (laneState_1_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (laneState_1_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (laneState_1_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (laneState_1_decodeResult_logic),
    .enqueue_bits_lastGroupForInstruction            (laneState_1_lastGroupForInstruction),
    .enqueue_bits_isLastLaneForInstruction           (laneState_1_isLastLaneForInstruction),
    .enqueue_bits_instructionFinished                (laneState_1_instructionFinished),
    .enqueue_bits_csr_vl                             (laneState_1_csr_vl),
    .enqueue_bits_csr_vStart                         (laneState_1_csr_vStart),
    .enqueue_bits_csr_vlmul                          (laneState_1_csr_vlmul),
    .enqueue_bits_csr_vSew                           (laneState_1_csr_vSew),
    .enqueue_bits_csr_vxrm                           (laneState_1_csr_vxrm),
    .enqueue_bits_csr_vta                            (laneState_1_csr_vta),
    .enqueue_bits_csr_vma                            (laneState_1_csr_vma),
    .enqueue_bits_maskType                           (laneState_1_maskType),
    .enqueue_bits_maskNotMaskedElement               (laneState_1_maskNotMaskedElement),
    .enqueue_bits_vs1                                (laneState_1_vs1),
    .enqueue_bits_vs2                                (laneState_1_vs2),
    .enqueue_bits_vd                                 (laneState_1_vd),
    .enqueue_bits_instructionIndex                   (laneState_1_instructionIndex),
    .enqueue_bits_additionalRW                       (laneState_1_additionalRW),
    .enqueue_bits_skipRead                           (laneState_1_skipRead),
    .enqueue_bits_skipEnable                         (laneState_1_skipEnable),
    .dequeue_ready                                   (_stage1_1_enqueue_ready),
    .dequeue_valid                                   (_stage0_1_dequeue_valid),
    .dequeue_bits_maskForMaskInput                   (_stage0_1_dequeue_bits_maskForMaskInput),
    .dequeue_bits_boundaryMaskCorrection             (_stage0_1_dequeue_bits_boundaryMaskCorrection),
    .dequeue_bits_groupCounter                       (_stage0_1_dequeue_bits_groupCounter),
    .dequeue_bits_readFromScalar                     (_stage0_1_dequeue_bits_readFromScalar),
    .dequeue_bits_instructionIndex                   (_stage0_1_dequeue_bits_instructionIndex),
    .dequeue_bits_decodeResult_specialSlot           (_stage0_1_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage0_1_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage0_1_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage0_1_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage0_1_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage0_1_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage0_1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage0_1_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage0_1_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage0_1_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage0_1_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage0_1_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage0_1_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage0_1_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage0_1_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage0_1_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage0_1_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage0_1_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage0_1_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage0_1_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage0_1_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage0_1_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage0_1_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage0_1_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage0_1_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage0_1_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage0_1_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage0_1_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage0_1_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage0_1_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage0_1_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage0_1_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage0_1_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage0_1_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage0_1_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage0_1_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage0_1_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage0_1_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage0_1_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage0_1_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage0_1_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage0_1_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage0_1_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage0_1_dequeue_bits_decodeResult_logic),
    .dequeue_bits_laneIndex                          (_stage0_1_dequeue_bits_laneIndex),
    .dequeue_bits_skipRead                           (_stage0_1_dequeue_bits_skipRead),
    .dequeue_bits_vs1                                (_stage0_1_dequeue_bits_vs1),
    .dequeue_bits_vs2                                (_stage0_1_dequeue_bits_vs2),
    .dequeue_bits_vd                                 (_stage0_1_dequeue_bits_vd),
    .dequeue_bits_vSew1H                             (_stage0_1_dequeue_bits_vSew1H),
    .dequeue_bits_maskNotMaskedElement               (_stage0_1_dequeue_bits_maskNotMaskedElement),
    .dequeue_bits_csr_vl                             (_stage0_1_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage0_1_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage0_1_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage0_1_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage0_1_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage0_1_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage0_1_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage0_1_dequeue_bits_maskType),
    .dequeue_bits_loadStore                          (_stage0_1_dequeue_bits_loadStore),
    .dequeue_bits_bordersForMaskLogic                (_stage0_1_dequeue_bits_bordersForMaskLogic),
    .updateLaneState_maskGroupCount                  (_stage0_1_updateLaneState_maskGroupCount),
    .updateLaneState_maskIndex                       (_stage0_1_updateLaneState_maskIndex),
    .updateLaneState_outOfExecutionRange             (_stage0_1_updateLaneState_outOfExecutionRange),
    .updateLaneState_maskExhausted                   (_stage0_1_updateLaneState_maskExhausted),
    .tokenReport_valid                               (_stage0_1_tokenReport_valid),
    .tokenReport_bits_decodeResult_sWrite            (_stage0_1_tokenReport_bits_decodeResult_sWrite),
    .tokenReport_bits_decodeResult_maskUnit          (_stage0_1_tokenReport_bits_decodeResult_maskUnit),
    .tokenReport_bits_instructionIndex               (_stage0_1_tokenReport_bits_instructionIndex)
  );
  LaneStage1_1 stage1_1 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage1_1_enqueue_ready),
    .enqueue_valid                                   (_stage0_1_dequeue_valid),
    .enqueue_bits_groupCounter                       (_stage0_1_dequeue_bits_groupCounter),
    .enqueue_bits_maskForMaskInput                   (_stage0_1_dequeue_bits_maskForMaskInput),
    .enqueue_bits_boundaryMaskCorrection             (_stage0_1_dequeue_bits_boundaryMaskCorrection),
    .enqueue_bits_instructionIndex                   (_stage0_1_dequeue_bits_instructionIndex),
    .enqueue_bits_decodeResult_specialSlot           (_stage0_1_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage0_1_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage0_1_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage0_1_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage0_1_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage0_1_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage0_1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage0_1_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage0_1_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage0_1_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage0_1_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage0_1_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage0_1_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage0_1_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage0_1_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage0_1_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage0_1_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage0_1_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage0_1_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage0_1_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage0_1_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage0_1_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage0_1_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage0_1_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage0_1_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage0_1_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage0_1_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage0_1_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage0_1_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage0_1_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage0_1_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage0_1_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage0_1_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage0_1_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage0_1_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage0_1_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage0_1_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage0_1_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage0_1_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage0_1_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage0_1_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage0_1_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage0_1_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage0_1_dequeue_bits_decodeResult_logic),
    .enqueue_bits_laneIndex                          (_stage0_1_dequeue_bits_laneIndex),
    .enqueue_bits_skipRead                           (_stage0_1_dequeue_bits_skipRead),
    .enqueue_bits_vs1                                (_stage0_1_dequeue_bits_vs1),
    .enqueue_bits_vs2                                (_stage0_1_dequeue_bits_vs2),
    .enqueue_bits_vd                                 (_stage0_1_dequeue_bits_vd),
    .enqueue_bits_vSew1H                             (_stage0_1_dequeue_bits_vSew1H),
    .enqueue_bits_maskNotMaskedElement               (_stage0_1_dequeue_bits_maskNotMaskedElement),
    .enqueue_bits_csr_vl                             (_stage0_1_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage0_1_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage0_1_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage0_1_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage0_1_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage0_1_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage0_1_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage0_1_dequeue_bits_maskType),
    .enqueue_bits_loadStore                          (_stage0_1_dequeue_bits_loadStore),
    .enqueue_bits_readFromScalar                     (_stage0_1_dequeue_bits_readFromScalar),
    .enqueue_bits_bordersForMaskLogic                (_stage0_1_dequeue_bits_bordersForMaskLogic),
    .dequeue_ready                                   (_stage2_1_enqueue_ready & _executionUnit_1_enqueue_ready),
    .dequeue_valid                                   (_stage1_1_dequeue_valid),
    .dequeue_bits_maskForFilter                      (_stage1_1_dequeue_bits_maskForFilter),
    .dequeue_bits_mask                               (_stage1_1_dequeue_bits_mask),
    .dequeue_bits_groupCounter                       (_stage1_1_dequeue_bits_groupCounter),
    .dequeue_bits_src_0                              (_stage1_1_dequeue_bits_src_0),
    .dequeue_bits_src_1                              (_stage1_1_dequeue_bits_src_1),
    .dequeue_bits_src_2                              (_stage1_1_dequeue_bits_src_2),
    .dequeue_bits_decodeResult_specialSlot           (_stage1_1_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage1_1_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage1_1_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage1_1_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage1_1_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage1_1_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage1_1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage1_1_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage1_1_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage1_1_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage1_1_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage1_1_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage1_1_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage1_1_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage1_1_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage1_1_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage1_1_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage1_1_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage1_1_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage1_1_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage1_1_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage1_1_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage1_1_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage1_1_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage1_1_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage1_1_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage1_1_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage1_1_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage1_1_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage1_1_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage1_1_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage1_1_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage1_1_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage1_1_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage1_1_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage1_1_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage1_1_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage1_1_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage1_1_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage1_1_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage1_1_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage1_1_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage1_1_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage1_1_dequeue_bits_decodeResult_logic),
    .dequeue_bits_vSew1H                             (_stage1_1_dequeue_bits_vSew1H),
    .dequeue_bits_csr_vl                             (_stage1_1_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage1_1_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage1_1_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage1_1_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage1_1_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage1_1_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage1_1_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage1_1_dequeue_bits_maskType),
    .dequeue_bits_laneIndex                          (_stage1_1_dequeue_bits_laneIndex),
    .dequeue_bits_instructionIndex                   (_stage1_1_dequeue_bits_instructionIndex),
    .dequeue_bits_loadStore                          (_stage1_1_dequeue_bits_loadStore),
    .dequeue_bits_vd                                 (_stage1_1_dequeue_bits_vd),
    .dequeue_bits_bordersForMaskLogic                (_stage1_1_dequeue_bits_bordersForMaskLogic),
    .vrfReadRequest_0_ready                          (vrfReadRequest_1_0_ready),
    .vrfReadRequest_0_valid                          (vrfReadRequest_1_0_valid),
    .vrfReadRequest_0_bits_vs                        (vrfReadRequest_1_0_bits_vs),
    .vrfReadRequest_0_bits_readSource                (vrfReadRequest_1_0_bits_readSource),
    .vrfReadRequest_0_bits_offset                    (vrfReadRequest_1_0_bits_offset),
    .vrfReadRequest_0_bits_instructionIndex          (vrfReadRequest_1_0_bits_instructionIndex),
    .vrfReadRequest_1_ready                          (vrfReadRequest_1_1_ready),
    .vrfReadRequest_1_valid                          (vrfReadRequest_1_1_valid),
    .vrfReadRequest_1_bits_vs                        (vrfReadRequest_1_1_bits_vs),
    .vrfReadRequest_1_bits_readSource                (vrfReadRequest_1_1_bits_readSource),
    .vrfReadRequest_1_bits_offset                    (vrfReadRequest_1_1_bits_offset),
    .vrfReadRequest_1_bits_instructionIndex          (vrfReadRequest_1_1_bits_instructionIndex),
    .vrfReadRequest_2_ready                          (vrfReadRequest_1_2_ready),
    .vrfReadRequest_2_valid                          (vrfReadRequest_1_2_valid),
    .vrfReadRequest_2_bits_vs                        (vrfReadRequest_1_2_bits_vs),
    .vrfReadRequest_2_bits_readSource                (vrfReadRequest_1_2_bits_readSource),
    .vrfReadRequest_2_bits_offset                    (vrfReadRequest_1_2_bits_offset),
    .vrfReadRequest_2_bits_instructionIndex          (vrfReadRequest_1_2_bits_instructionIndex),
    .vrfCheckRequest_0_vs                            (readCheckRequestVec_6_vs),
    .vrfCheckRequest_0_readSource                    (readCheckRequestVec_6_readSource),
    .vrfCheckRequest_0_offset                        (readCheckRequestVec_6_offset),
    .vrfCheckRequest_0_instructionIndex              (readCheckRequestVec_6_instructionIndex),
    .vrfCheckRequest_1_vs                            (readCheckRequestVec_7_vs),
    .vrfCheckRequest_1_readSource                    (readCheckRequestVec_7_readSource),
    .vrfCheckRequest_1_offset                        (readCheckRequestVec_7_offset),
    .vrfCheckRequest_1_instructionIndex              (readCheckRequestVec_7_instructionIndex),
    .vrfCheckRequest_2_vs                            (readCheckRequestVec_8_vs),
    .vrfCheckRequest_2_readSource                    (readCheckRequestVec_8_readSource),
    .vrfCheckRequest_2_offset                        (readCheckRequestVec_8_offset),
    .vrfCheckRequest_2_instructionIndex              (readCheckRequestVec_8_instructionIndex),
    .checkResult_0                                   (readCheckResult_6),
    .checkResult_1                                   (readCheckResult_7),
    .checkResult_2                                   (readCheckResult_8),
    .vrfReadResult_0                                 (vrfReadResult_1_0),
    .vrfReadResult_1                                 (vrfReadResult_1_1),
    .vrfReadResult_2                                 (vrfReadResult_1_2)
  );
  LaneStage2_1 stage2_1 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage2_1_enqueue_ready),
    .enqueue_valid                                   (_stage1_1_dequeue_valid & _executionUnit_1_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_1_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_1_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_1_dequeue_bits_src_2),
    .enqueue_bits_groupCounter                       (_stage1_1_dequeue_bits_groupCounter),
    .enqueue_bits_maskForFilter                      (_stage1_1_dequeue_bits_maskForFilter),
    .enqueue_bits_mask                               (_stage1_1_dequeue_bits_mask),
    .enqueue_bits_bordersForMaskLogic                (_stage1_1_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_1_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_1_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_1_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_1_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_1_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_1_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_1_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_1_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_1_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_1_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_1_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_1_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_1_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_1_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_1_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_1_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_1_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_1_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_1_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_1_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_1_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_1_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_1_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_1_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_1_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_1_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_1_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_1_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_1_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_1_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_1_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_1_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_1_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_1_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_1_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_1_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_1_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_1_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_1_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_1_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_1_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_1_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_1_dequeue_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (_stage1_1_dequeue_bits_instructionIndex),
    .enqueue_bits_loadStore                          (_stage1_1_dequeue_bits_loadStore),
    .enqueue_bits_vd                                 (_stage1_1_dequeue_bits_vd),
    .enqueue_bits_csr_vl                             (_stage1_1_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_1_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_1_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_1_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_1_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_1_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_1_dequeue_bits_csr_vma),
    .enqueue_bits_vSew1H                             (_stage1_1_dequeue_bits_vSew1H),
    .enqueue_bits_maskType                           (_stage1_1_dequeue_bits_maskType),
    .dequeue_ready                                   (stage3EnqWire_1_ready & _executionUnit_1_dequeue_valid),
    .dequeue_valid                                   (_stage2_1_dequeue_valid),
    .dequeue_bits_groupCounter                       (stage3EnqWire_1_bits_groupCounter),
    .dequeue_bits_mask                               (stage3EnqWire_1_bits_mask),
    .dequeue_bits_decodeResult_specialSlot           (stage3EnqWire_1_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (stage3EnqWire_1_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (stage3EnqWire_1_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (stage3EnqWire_1_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (stage3EnqWire_1_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (stage3EnqWire_1_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_1_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (stage3EnqWire_1_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (stage3EnqWire_1_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (stage3EnqWire_1_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (stage3EnqWire_1_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (stage3EnqWire_1_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (stage3EnqWire_1_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (stage3EnqWire_1_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (stage3EnqWire_1_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (stage3EnqWire_1_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (stage3EnqWire_1_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (stage3EnqWire_1_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (stage3EnqWire_1_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (stage3EnqWire_1_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (stage3EnqWire_1_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (stage3EnqWire_1_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (stage3EnqWire_1_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (stage3EnqWire_1_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (stage3EnqWire_1_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (stage3EnqWire_1_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (stage3EnqWire_1_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (stage3EnqWire_1_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (stage3EnqWire_1_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (stage3EnqWire_1_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (stage3EnqWire_1_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (stage3EnqWire_1_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (stage3EnqWire_1_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (stage3EnqWire_1_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (stage3EnqWire_1_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (stage3EnqWire_1_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (stage3EnqWire_1_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (stage3EnqWire_1_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (stage3EnqWire_1_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (stage3EnqWire_1_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (stage3EnqWire_1_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (stage3EnqWire_1_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (stage3EnqWire_1_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (stage3EnqWire_1_bits_decodeResult_logic),
    .dequeue_bits_instructionIndex                   (stage3EnqWire_1_bits_instructionIndex),
    .dequeue_bits_loadStore                          (stage3EnqWire_1_bits_loadStore),
    .dequeue_bits_vd                                 (stage3EnqWire_1_bits_vd)
  );
  LaneExecutionBridge_1 executionUnit_1 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_executionUnit_1_enqueue_ready),
    .enqueue_valid                                   (_stage1_1_dequeue_valid & _stage2_1_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_1_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_1_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_1_dequeue_bits_src_2),
    .enqueue_bits_bordersForMaskLogic                (_stage1_1_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_mask                               (_stage1_1_dequeue_bits_mask),
    .enqueue_bits_maskForFilter                      (_stage1_1_dequeue_bits_maskForFilter),
    .enqueue_bits_groupCounter                       (_stage1_1_dequeue_bits_groupCounter),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_1_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_1_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_1_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_1_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_1_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_1_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_1_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_1_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_1_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_1_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_1_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_1_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_1_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_1_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_1_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_1_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_1_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_1_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_1_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_1_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_1_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_1_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_1_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_1_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_1_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_1_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_1_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_1_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_1_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_1_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_1_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_1_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_1_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_1_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_1_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_1_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_1_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_1_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_1_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_1_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_1_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_1_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_1_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_1_dequeue_bits_decodeResult_logic),
    .enqueue_bits_vSew1H                             (_stage1_1_dequeue_bits_vSew1H),
    .enqueue_bits_csr_vl                             (_stage1_1_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_1_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_1_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_1_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_1_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_1_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_1_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage1_1_dequeue_bits_maskType),
    .enqueue_bits_laneIndex                          (_stage1_1_dequeue_bits_laneIndex),
    .enqueue_bits_instructionIndex                   (_stage1_1_dequeue_bits_instructionIndex),
    .dequeue_ready                                   (stage3EnqWire_1_ready),
    .dequeue_valid                                   (_executionUnit_1_dequeue_valid),
    .dequeue_bits_data                               (stage3EnqWire_1_bits_data),
    .dequeue_bits_ffoIndex                           (stage3EnqWire_1_bits_ffoIndex),
    .vfuRequest_ready                                (executeEnqueueFire_1),
    .vfuRequest_valid                                (_executionUnit_1_vfuRequest_valid),
    .vfuRequest_bits_src_0                           (requestVec_1_src_0),
    .vfuRequest_bits_src_1                           (requestVec_1_src_1),
    .vfuRequest_bits_src_2                           (requestVec_1_src_2),
    .vfuRequest_bits_src_3                           (requestVec_1_src_3),
    .vfuRequest_bits_opcode                          (requestVec_1_opcode),
    .vfuRequest_bits_mask                            (requestVec_1_mask),
    .vfuRequest_bits_executeMask                     (requestVec_1_executeMask),
    .vfuRequest_bits_sign0                           (requestVec_1_sign0),
    .vfuRequest_bits_sign                            (requestVec_1_sign),
    .vfuRequest_bits_reverse                         (requestVec_1_reverse),
    .vfuRequest_bits_average                         (requestVec_1_average),
    .vfuRequest_bits_saturate                        (requestVec_1_saturate),
    .vfuRequest_bits_vxrm                            (requestVec_1_vxrm),
    .vfuRequest_bits_vSew                            (requestVec_1_vSew),
    .vfuRequest_bits_shifterSize                     (requestVec_1_shifterSize),
    .vfuRequest_bits_rem                             (requestVec_1_rem),
    .vfuRequest_bits_groupIndex                      (requestVec_1_groupIndex),
    .vfuRequest_bits_laneIndex                       (requestVec_1_laneIndex),
    .vfuRequest_bits_maskType                        (requestVec_1_maskType),
    .vfuRequest_bits_narrow                          (requestVec_1_narrow),
    .dataResponse_valid                              (responseVec_1_valid),
    .dataResponse_bits_data                          (responseVec_1_bits_data),
    .executeDecode_specialSlot                       (executeDecodeVec_1_specialSlot),
    .executeDecode_topUop                            (executeDecodeVec_1_topUop),
    .executeDecode_popCount                          (executeDecodeVec_1_popCount),
    .executeDecode_ffo                               (executeDecodeVec_1_ffo),
    .executeDecode_average                           (executeDecodeVec_1_average),
    .executeDecode_reverse                           (executeDecodeVec_1_reverse),
    .executeDecode_dontNeedExecuteInLane             (executeDecodeVec_1_dontNeedExecuteInLane),
    .executeDecode_scheduler                         (executeDecodeVec_1_scheduler),
    .executeDecode_sReadVD                           (executeDecodeVec_1_sReadVD),
    .executeDecode_vtype                             (executeDecodeVec_1_vtype),
    .executeDecode_sWrite                            (executeDecodeVec_1_sWrite),
    .executeDecode_crossRead                         (executeDecodeVec_1_crossRead),
    .executeDecode_crossWrite                        (executeDecodeVec_1_crossWrite),
    .executeDecode_maskUnit                          (executeDecodeVec_1_maskUnit),
    .executeDecode_special                           (executeDecodeVec_1_special),
    .executeDecode_saturate                          (executeDecodeVec_1_saturate),
    .executeDecode_vwmacc                            (executeDecodeVec_1_vwmacc),
    .executeDecode_readOnly                          (executeDecodeVec_1_readOnly),
    .executeDecode_maskSource                        (executeDecodeVec_1_maskSource),
    .executeDecode_maskDestination                   (executeDecodeVec_1_maskDestination),
    .executeDecode_maskLogic                         (executeDecodeVec_1_maskLogic),
    .executeDecode_uop                               (executeDecodeVec_1_uop),
    .executeDecode_iota                              (executeDecodeVec_1_iota),
    .executeDecode_mv                                (executeDecodeVec_1_mv),
    .executeDecode_extend                            (executeDecodeVec_1_extend),
    .executeDecode_unOrderWrite                      (executeDecodeVec_1_unOrderWrite),
    .executeDecode_compress                          (executeDecodeVec_1_compress),
    .executeDecode_gather16                          (executeDecodeVec_1_gather16),
    .executeDecode_gather                            (executeDecodeVec_1_gather),
    .executeDecode_slid                              (executeDecodeVec_1_slid),
    .executeDecode_targetRd                          (executeDecodeVec_1_targetRd),
    .executeDecode_widenReduce                       (executeDecodeVec_1_widenReduce),
    .executeDecode_red                               (executeDecodeVec_1_red),
    .executeDecode_nr                                (executeDecodeVec_1_nr),
    .executeDecode_itype                             (executeDecodeVec_1_itype),
    .executeDecode_unsigned1                         (executeDecodeVec_1_unsigned1),
    .executeDecode_unsigned0                         (executeDecodeVec_1_unsigned0),
    .executeDecode_other                             (executeDecodeVec_1_other),
    .executeDecode_multiCycle                        (executeDecodeVec_1_multiCycle),
    .executeDecode_divider                           (executeDecodeVec_1_divider),
    .executeDecode_multiplier                        (executeDecodeVec_1_multiplier),
    .executeDecode_shift                             (executeDecodeVec_1_shift),
    .executeDecode_adder                             (executeDecodeVec_1_adder),
    .executeDecode_logic                             (executeDecodeVec_1_logic),
    .responseDecode_specialSlot                      (responseDecodeVec_1_specialSlot),
    .responseDecode_topUop                           (responseDecodeVec_1_topUop),
    .responseDecode_popCount                         (responseDecodeVec_1_popCount),
    .responseDecode_ffo                              (responseDecodeVec_1_ffo),
    .responseDecode_average                          (responseDecodeVec_1_average),
    .responseDecode_reverse                          (responseDecodeVec_1_reverse),
    .responseDecode_dontNeedExecuteInLane            (responseDecodeVec_1_dontNeedExecuteInLane),
    .responseDecode_scheduler                        (responseDecodeVec_1_scheduler),
    .responseDecode_sReadVD                          (responseDecodeVec_1_sReadVD),
    .responseDecode_vtype                            (responseDecodeVec_1_vtype),
    .responseDecode_sWrite                           (responseDecodeVec_1_sWrite),
    .responseDecode_crossRead                        (responseDecodeVec_1_crossRead),
    .responseDecode_crossWrite                       (responseDecodeVec_1_crossWrite),
    .responseDecode_maskUnit                         (responseDecodeVec_1_maskUnit),
    .responseDecode_special                          (responseDecodeVec_1_special),
    .responseDecode_saturate                         (responseDecodeVec_1_saturate),
    .responseDecode_vwmacc                           (responseDecodeVec_1_vwmacc),
    .responseDecode_readOnly                         (responseDecodeVec_1_readOnly),
    .responseDecode_maskSource                       (responseDecodeVec_1_maskSource),
    .responseDecode_maskDestination                  (responseDecodeVec_1_maskDestination),
    .responseDecode_maskLogic                        (responseDecodeVec_1_maskLogic),
    .responseDecode_uop                              (responseDecodeVec_1_uop),
    .responseDecode_iota                             (responseDecodeVec_1_iota),
    .responseDecode_mv                               (responseDecodeVec_1_mv),
    .responseDecode_extend                           (responseDecodeVec_1_extend),
    .responseDecode_unOrderWrite                     (responseDecodeVec_1_unOrderWrite),
    .responseDecode_compress                         (responseDecodeVec_1_compress),
    .responseDecode_gather16                         (responseDecodeVec_1_gather16),
    .responseDecode_gather                           (responseDecodeVec_1_gather),
    .responseDecode_slid                             (responseDecodeVec_1_slid),
    .responseDecode_targetRd                         (responseDecodeVec_1_targetRd),
    .responseDecode_widenReduce                      (responseDecodeVec_1_widenReduce),
    .responseDecode_red                              (responseDecodeVec_1_red),
    .responseDecode_nr                               (responseDecodeVec_1_nr),
    .responseDecode_itype                            (responseDecodeVec_1_itype),
    .responseDecode_unsigned1                        (responseDecodeVec_1_unsigned1),
    .responseDecode_unsigned0                        (responseDecodeVec_1_unsigned0),
    .responseDecode_other                            (responseDecodeVec_1_other),
    .responseDecode_multiCycle                       (responseDecodeVec_1_multiCycle),
    .responseDecode_divider                          (responseDecodeVec_1_divider),
    .responseDecode_multiplier                       (responseDecodeVec_1_multiplier),
    .responseDecode_shift                            (responseDecodeVec_1_shift),
    .responseDecode_adder                            (responseDecodeVec_1_adder),
    .responseDecode_logic                            (responseDecodeVec_1_logic),
    .responseIndex                                   (_executionUnit_1_responseIndex)
  );
  LaneStage3_1 stage3_1 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (stage3EnqWire_1_ready),
    .enqueue_valid                                   (stage3EnqWire_1_valid),
    .enqueue_bits_groupCounter                       (stage3EnqWire_1_bits_groupCounter),
    .enqueue_bits_data                               (stage3EnqWire_1_bits_data),
    .enqueue_bits_mask                               (stage3EnqWire_1_bits_mask),
    .enqueue_bits_ffoIndex                           (stage3EnqWire_1_bits_ffoIndex),
    .enqueue_bits_decodeResult_specialSlot           (stage3EnqWire_1_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (stage3EnqWire_1_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (stage3EnqWire_1_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (stage3EnqWire_1_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (stage3EnqWire_1_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (stage3EnqWire_1_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_1_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (stage3EnqWire_1_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (stage3EnqWire_1_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (stage3EnqWire_1_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (stage3EnqWire_1_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (stage3EnqWire_1_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (stage3EnqWire_1_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (stage3EnqWire_1_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (stage3EnqWire_1_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (stage3EnqWire_1_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (stage3EnqWire_1_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (stage3EnqWire_1_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (stage3EnqWire_1_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (stage3EnqWire_1_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (stage3EnqWire_1_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (stage3EnqWire_1_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (stage3EnqWire_1_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (stage3EnqWire_1_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (stage3EnqWire_1_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (stage3EnqWire_1_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (stage3EnqWire_1_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (stage3EnqWire_1_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (stage3EnqWire_1_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (stage3EnqWire_1_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (stage3EnqWire_1_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (stage3EnqWire_1_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (stage3EnqWire_1_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (stage3EnqWire_1_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (stage3EnqWire_1_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (stage3EnqWire_1_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (stage3EnqWire_1_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (stage3EnqWire_1_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (stage3EnqWire_1_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (stage3EnqWire_1_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (stage3EnqWire_1_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (stage3EnqWire_1_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (stage3EnqWire_1_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (stage3EnqWire_1_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (stage3EnqWire_1_bits_instructionIndex),
    .enqueue_bits_loadStore                          (stage3EnqWire_1_bits_loadStore),
    .enqueue_bits_vd                                 (stage3EnqWire_1_bits_vd),
    .vrfWriteRequest_ready                           (vrfWriteArbiter_1_ready),
    .vrfWriteRequest_valid                           (_stage3_1_vrfWriteRequest_valid),
    .vrfWriteRequest_bits_vd                         (vrfWriteArbiter_1_bits_vd),
    .vrfWriteRequest_bits_offset                     (vrfWriteArbiter_1_bits_offset),
    .vrfWriteRequest_bits_mask                       (_stage3_1_vrfWriteRequest_bits_mask),
    .vrfWriteRequest_bits_data                       (vrfWriteArbiter_1_bits_data),
    .vrfWriteRequest_bits_last                       (vrfWriteArbiter_1_bits_last),
    .vrfWriteRequest_bits_instructionIndex           (_stage3_1_vrfWriteRequest_bits_instructionIndex)
  );
  LaneStage0_1 stage0_2 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage0_2_enqueue_ready),
    .enqueue_valid                                   (stage0_2_enqueue_valid),
    .enqueue_bits_maskIndex                          (maskIndexVec_2),
    .enqueue_bits_maskForMaskGroup                   (slotControl_2_mask_bits),
    .enqueue_bits_maskGroupCount                     (maskGroupCountVec_2),
    .enqueue_bits_readFromScalar                     (slotControl_2_laneRequest_readFromScalar),
    .enqueue_bits_vSew1H                             (laneState_2_vSew1H),
    .enqueue_bits_loadStore                          (laneState_2_loadStore),
    .enqueue_bits_laneIndex                          (laneState_2_laneIndex),
    .enqueue_bits_decodeResult_specialSlot           (laneState_2_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (laneState_2_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (laneState_2_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (laneState_2_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (laneState_2_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (laneState_2_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (laneState_2_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (laneState_2_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (laneState_2_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (laneState_2_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (laneState_2_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (laneState_2_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (laneState_2_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (laneState_2_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (laneState_2_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (laneState_2_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (laneState_2_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (laneState_2_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (laneState_2_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (laneState_2_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (laneState_2_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (laneState_2_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (laneState_2_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (laneState_2_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (laneState_2_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (laneState_2_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (laneState_2_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (laneState_2_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (laneState_2_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (laneState_2_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (laneState_2_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (laneState_2_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (laneState_2_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (laneState_2_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (laneState_2_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (laneState_2_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (laneState_2_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (laneState_2_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (laneState_2_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (laneState_2_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (laneState_2_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (laneState_2_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (laneState_2_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (laneState_2_decodeResult_logic),
    .enqueue_bits_lastGroupForInstruction            (laneState_2_lastGroupForInstruction),
    .enqueue_bits_isLastLaneForInstruction           (laneState_2_isLastLaneForInstruction),
    .enqueue_bits_instructionFinished                (laneState_2_instructionFinished),
    .enqueue_bits_csr_vl                             (laneState_2_csr_vl),
    .enqueue_bits_csr_vStart                         (laneState_2_csr_vStart),
    .enqueue_bits_csr_vlmul                          (laneState_2_csr_vlmul),
    .enqueue_bits_csr_vSew                           (laneState_2_csr_vSew),
    .enqueue_bits_csr_vxrm                           (laneState_2_csr_vxrm),
    .enqueue_bits_csr_vta                            (laneState_2_csr_vta),
    .enqueue_bits_csr_vma                            (laneState_2_csr_vma),
    .enqueue_bits_maskType                           (laneState_2_maskType),
    .enqueue_bits_maskNotMaskedElement               (laneState_2_maskNotMaskedElement),
    .enqueue_bits_vs1                                (laneState_2_vs1),
    .enqueue_bits_vs2                                (laneState_2_vs2),
    .enqueue_bits_vd                                 (laneState_2_vd),
    .enqueue_bits_instructionIndex                   (laneState_2_instructionIndex),
    .enqueue_bits_additionalRW                       (laneState_2_additionalRW),
    .enqueue_bits_skipRead                           (laneState_2_skipRead),
    .enqueue_bits_skipEnable                         (laneState_2_skipEnable),
    .dequeue_ready                                   (_stage1_2_enqueue_ready),
    .dequeue_valid                                   (_stage0_2_dequeue_valid),
    .dequeue_bits_maskForMaskInput                   (_stage0_2_dequeue_bits_maskForMaskInput),
    .dequeue_bits_boundaryMaskCorrection             (_stage0_2_dequeue_bits_boundaryMaskCorrection),
    .dequeue_bits_groupCounter                       (_stage0_2_dequeue_bits_groupCounter),
    .dequeue_bits_readFromScalar                     (_stage0_2_dequeue_bits_readFromScalar),
    .dequeue_bits_instructionIndex                   (_stage0_2_dequeue_bits_instructionIndex),
    .dequeue_bits_decodeResult_specialSlot           (_stage0_2_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage0_2_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage0_2_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage0_2_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage0_2_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage0_2_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage0_2_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage0_2_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage0_2_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage0_2_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage0_2_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage0_2_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage0_2_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage0_2_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage0_2_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage0_2_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage0_2_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage0_2_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage0_2_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage0_2_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage0_2_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage0_2_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage0_2_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage0_2_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage0_2_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage0_2_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage0_2_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage0_2_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage0_2_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage0_2_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage0_2_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage0_2_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage0_2_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage0_2_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage0_2_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage0_2_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage0_2_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage0_2_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage0_2_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage0_2_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage0_2_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage0_2_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage0_2_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage0_2_dequeue_bits_decodeResult_logic),
    .dequeue_bits_laneIndex                          (_stage0_2_dequeue_bits_laneIndex),
    .dequeue_bits_skipRead                           (_stage0_2_dequeue_bits_skipRead),
    .dequeue_bits_vs1                                (_stage0_2_dequeue_bits_vs1),
    .dequeue_bits_vs2                                (_stage0_2_dequeue_bits_vs2),
    .dequeue_bits_vd                                 (_stage0_2_dequeue_bits_vd),
    .dequeue_bits_vSew1H                             (_stage0_2_dequeue_bits_vSew1H),
    .dequeue_bits_maskNotMaskedElement               (_stage0_2_dequeue_bits_maskNotMaskedElement),
    .dequeue_bits_csr_vl                             (_stage0_2_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage0_2_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage0_2_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage0_2_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage0_2_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage0_2_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage0_2_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage0_2_dequeue_bits_maskType),
    .dequeue_bits_loadStore                          (_stage0_2_dequeue_bits_loadStore),
    .dequeue_bits_bordersForMaskLogic                (_stage0_2_dequeue_bits_bordersForMaskLogic),
    .updateLaneState_maskGroupCount                  (_stage0_2_updateLaneState_maskGroupCount),
    .updateLaneState_maskIndex                       (_stage0_2_updateLaneState_maskIndex),
    .updateLaneState_outOfExecutionRange             (_stage0_2_updateLaneState_outOfExecutionRange),
    .updateLaneState_maskExhausted                   (_stage0_2_updateLaneState_maskExhausted),
    .tokenReport_valid                               (_stage0_2_tokenReport_valid),
    .tokenReport_bits_decodeResult_sWrite            (_stage0_2_tokenReport_bits_decodeResult_sWrite),
    .tokenReport_bits_decodeResult_maskUnit          (_stage0_2_tokenReport_bits_decodeResult_maskUnit),
    .tokenReport_bits_instructionIndex               (_stage0_2_tokenReport_bits_instructionIndex)
  );
  LaneStage1_1 stage1_2 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage1_2_enqueue_ready),
    .enqueue_valid                                   (_stage0_2_dequeue_valid),
    .enqueue_bits_groupCounter                       (_stage0_2_dequeue_bits_groupCounter),
    .enqueue_bits_maskForMaskInput                   (_stage0_2_dequeue_bits_maskForMaskInput),
    .enqueue_bits_boundaryMaskCorrection             (_stage0_2_dequeue_bits_boundaryMaskCorrection),
    .enqueue_bits_instructionIndex                   (_stage0_2_dequeue_bits_instructionIndex),
    .enqueue_bits_decodeResult_specialSlot           (_stage0_2_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage0_2_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage0_2_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage0_2_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage0_2_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage0_2_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage0_2_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage0_2_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage0_2_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage0_2_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage0_2_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage0_2_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage0_2_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage0_2_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage0_2_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage0_2_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage0_2_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage0_2_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage0_2_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage0_2_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage0_2_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage0_2_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage0_2_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage0_2_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage0_2_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage0_2_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage0_2_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage0_2_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage0_2_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage0_2_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage0_2_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage0_2_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage0_2_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage0_2_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage0_2_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage0_2_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage0_2_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage0_2_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage0_2_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage0_2_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage0_2_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage0_2_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage0_2_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage0_2_dequeue_bits_decodeResult_logic),
    .enqueue_bits_laneIndex                          (_stage0_2_dequeue_bits_laneIndex),
    .enqueue_bits_skipRead                           (_stage0_2_dequeue_bits_skipRead),
    .enqueue_bits_vs1                                (_stage0_2_dequeue_bits_vs1),
    .enqueue_bits_vs2                                (_stage0_2_dequeue_bits_vs2),
    .enqueue_bits_vd                                 (_stage0_2_dequeue_bits_vd),
    .enqueue_bits_vSew1H                             (_stage0_2_dequeue_bits_vSew1H),
    .enqueue_bits_maskNotMaskedElement               (_stage0_2_dequeue_bits_maskNotMaskedElement),
    .enqueue_bits_csr_vl                             (_stage0_2_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage0_2_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage0_2_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage0_2_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage0_2_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage0_2_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage0_2_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage0_2_dequeue_bits_maskType),
    .enqueue_bits_loadStore                          (_stage0_2_dequeue_bits_loadStore),
    .enqueue_bits_readFromScalar                     (_stage0_2_dequeue_bits_readFromScalar),
    .enqueue_bits_bordersForMaskLogic                (_stage0_2_dequeue_bits_bordersForMaskLogic),
    .dequeue_ready                                   (_stage2_2_enqueue_ready & _executionUnit_2_enqueue_ready),
    .dequeue_valid                                   (_stage1_2_dequeue_valid),
    .dequeue_bits_maskForFilter                      (_stage1_2_dequeue_bits_maskForFilter),
    .dequeue_bits_mask                               (_stage1_2_dequeue_bits_mask),
    .dequeue_bits_groupCounter                       (_stage1_2_dequeue_bits_groupCounter),
    .dequeue_bits_src_0                              (_stage1_2_dequeue_bits_src_0),
    .dequeue_bits_src_1                              (_stage1_2_dequeue_bits_src_1),
    .dequeue_bits_src_2                              (_stage1_2_dequeue_bits_src_2),
    .dequeue_bits_decodeResult_specialSlot           (_stage1_2_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage1_2_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage1_2_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage1_2_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage1_2_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage1_2_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage1_2_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage1_2_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage1_2_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage1_2_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage1_2_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage1_2_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage1_2_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage1_2_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage1_2_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage1_2_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage1_2_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage1_2_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage1_2_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage1_2_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage1_2_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage1_2_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage1_2_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage1_2_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage1_2_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage1_2_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage1_2_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage1_2_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage1_2_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage1_2_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage1_2_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage1_2_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage1_2_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage1_2_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage1_2_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage1_2_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage1_2_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage1_2_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage1_2_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage1_2_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage1_2_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage1_2_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage1_2_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage1_2_dequeue_bits_decodeResult_logic),
    .dequeue_bits_vSew1H                             (_stage1_2_dequeue_bits_vSew1H),
    .dequeue_bits_csr_vl                             (_stage1_2_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage1_2_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage1_2_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage1_2_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage1_2_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage1_2_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage1_2_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage1_2_dequeue_bits_maskType),
    .dequeue_bits_laneIndex                          (_stage1_2_dequeue_bits_laneIndex),
    .dequeue_bits_instructionIndex                   (_stage1_2_dequeue_bits_instructionIndex),
    .dequeue_bits_loadStore                          (_stage1_2_dequeue_bits_loadStore),
    .dequeue_bits_vd                                 (_stage1_2_dequeue_bits_vd),
    .dequeue_bits_bordersForMaskLogic                (_stage1_2_dequeue_bits_bordersForMaskLogic),
    .vrfReadRequest_0_ready                          (vrfReadRequest_2_0_ready),
    .vrfReadRequest_0_valid                          (vrfReadRequest_2_0_valid),
    .vrfReadRequest_0_bits_vs                        (vrfReadRequest_2_0_bits_vs),
    .vrfReadRequest_0_bits_readSource                (vrfReadRequest_2_0_bits_readSource),
    .vrfReadRequest_0_bits_offset                    (vrfReadRequest_2_0_bits_offset),
    .vrfReadRequest_0_bits_instructionIndex          (vrfReadRequest_2_0_bits_instructionIndex),
    .vrfReadRequest_1_ready                          (vrfReadRequest_2_1_ready),
    .vrfReadRequest_1_valid                          (vrfReadRequest_2_1_valid),
    .vrfReadRequest_1_bits_vs                        (vrfReadRequest_2_1_bits_vs),
    .vrfReadRequest_1_bits_readSource                (vrfReadRequest_2_1_bits_readSource),
    .vrfReadRequest_1_bits_offset                    (vrfReadRequest_2_1_bits_offset),
    .vrfReadRequest_1_bits_instructionIndex          (vrfReadRequest_2_1_bits_instructionIndex),
    .vrfReadRequest_2_ready                          (vrfReadRequest_2_2_ready),
    .vrfReadRequest_2_valid                          (vrfReadRequest_2_2_valid),
    .vrfReadRequest_2_bits_vs                        (vrfReadRequest_2_2_bits_vs),
    .vrfReadRequest_2_bits_readSource                (vrfReadRequest_2_2_bits_readSource),
    .vrfReadRequest_2_bits_offset                    (vrfReadRequest_2_2_bits_offset),
    .vrfReadRequest_2_bits_instructionIndex          (vrfReadRequest_2_2_bits_instructionIndex),
    .vrfCheckRequest_0_vs                            (readCheckRequestVec_3_vs),
    .vrfCheckRequest_0_readSource                    (readCheckRequestVec_3_readSource),
    .vrfCheckRequest_0_offset                        (readCheckRequestVec_3_offset),
    .vrfCheckRequest_0_instructionIndex              (readCheckRequestVec_3_instructionIndex),
    .vrfCheckRequest_1_vs                            (readCheckRequestVec_4_vs),
    .vrfCheckRequest_1_readSource                    (readCheckRequestVec_4_readSource),
    .vrfCheckRequest_1_offset                        (readCheckRequestVec_4_offset),
    .vrfCheckRequest_1_instructionIndex              (readCheckRequestVec_4_instructionIndex),
    .vrfCheckRequest_2_vs                            (readCheckRequestVec_5_vs),
    .vrfCheckRequest_2_readSource                    (readCheckRequestVec_5_readSource),
    .vrfCheckRequest_2_offset                        (readCheckRequestVec_5_offset),
    .vrfCheckRequest_2_instructionIndex              (readCheckRequestVec_5_instructionIndex),
    .checkResult_0                                   (readCheckResult_3),
    .checkResult_1                                   (readCheckResult_4),
    .checkResult_2                                   (readCheckResult_5),
    .vrfReadResult_0                                 (vrfReadResult_2_0),
    .vrfReadResult_1                                 (vrfReadResult_2_1),
    .vrfReadResult_2                                 (vrfReadResult_2_2)
  );
  LaneStage2_1 stage2_2 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage2_2_enqueue_ready),
    .enqueue_valid                                   (_stage1_2_dequeue_valid & _executionUnit_2_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_2_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_2_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_2_dequeue_bits_src_2),
    .enqueue_bits_groupCounter                       (_stage1_2_dequeue_bits_groupCounter),
    .enqueue_bits_maskForFilter                      (_stage1_2_dequeue_bits_maskForFilter),
    .enqueue_bits_mask                               (_stage1_2_dequeue_bits_mask),
    .enqueue_bits_bordersForMaskLogic                (_stage1_2_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_2_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_2_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_2_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_2_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_2_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_2_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_2_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_2_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_2_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_2_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_2_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_2_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_2_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_2_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_2_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_2_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_2_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_2_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_2_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_2_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_2_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_2_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_2_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_2_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_2_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_2_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_2_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_2_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_2_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_2_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_2_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_2_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_2_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_2_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_2_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_2_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_2_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_2_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_2_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_2_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_2_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_2_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_2_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_2_dequeue_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (_stage1_2_dequeue_bits_instructionIndex),
    .enqueue_bits_loadStore                          (_stage1_2_dequeue_bits_loadStore),
    .enqueue_bits_vd                                 (_stage1_2_dequeue_bits_vd),
    .enqueue_bits_csr_vl                             (_stage1_2_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_2_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_2_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_2_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_2_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_2_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_2_dequeue_bits_csr_vma),
    .enqueue_bits_vSew1H                             (_stage1_2_dequeue_bits_vSew1H),
    .enqueue_bits_maskType                           (_stage1_2_dequeue_bits_maskType),
    .dequeue_ready                                   (stage3EnqWire_2_ready & _executionUnit_2_dequeue_valid),
    .dequeue_valid                                   (_stage2_2_dequeue_valid),
    .dequeue_bits_groupCounter                       (stage3EnqWire_2_bits_groupCounter),
    .dequeue_bits_mask                               (stage3EnqWire_2_bits_mask),
    .dequeue_bits_decodeResult_specialSlot           (stage3EnqWire_2_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (stage3EnqWire_2_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (stage3EnqWire_2_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (stage3EnqWire_2_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (stage3EnqWire_2_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (stage3EnqWire_2_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_2_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (stage3EnqWire_2_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (stage3EnqWire_2_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (stage3EnqWire_2_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (stage3EnqWire_2_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (stage3EnqWire_2_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (stage3EnqWire_2_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (stage3EnqWire_2_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (stage3EnqWire_2_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (stage3EnqWire_2_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (stage3EnqWire_2_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (stage3EnqWire_2_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (stage3EnqWire_2_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (stage3EnqWire_2_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (stage3EnqWire_2_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (stage3EnqWire_2_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (stage3EnqWire_2_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (stage3EnqWire_2_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (stage3EnqWire_2_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (stage3EnqWire_2_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (stage3EnqWire_2_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (stage3EnqWire_2_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (stage3EnqWire_2_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (stage3EnqWire_2_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (stage3EnqWire_2_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (stage3EnqWire_2_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (stage3EnqWire_2_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (stage3EnqWire_2_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (stage3EnqWire_2_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (stage3EnqWire_2_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (stage3EnqWire_2_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (stage3EnqWire_2_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (stage3EnqWire_2_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (stage3EnqWire_2_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (stage3EnqWire_2_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (stage3EnqWire_2_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (stage3EnqWire_2_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (stage3EnqWire_2_bits_decodeResult_logic),
    .dequeue_bits_instructionIndex                   (stage3EnqWire_2_bits_instructionIndex),
    .dequeue_bits_loadStore                          (stage3EnqWire_2_bits_loadStore),
    .dequeue_bits_vd                                 (stage3EnqWire_2_bits_vd)
  );
  LaneExecutionBridge_2 executionUnit_2 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_executionUnit_2_enqueue_ready),
    .enqueue_valid                                   (_stage1_2_dequeue_valid & _stage2_2_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_2_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_2_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_2_dequeue_bits_src_2),
    .enqueue_bits_bordersForMaskLogic                (_stage1_2_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_mask                               (_stage1_2_dequeue_bits_mask),
    .enqueue_bits_maskForFilter                      (_stage1_2_dequeue_bits_maskForFilter),
    .enqueue_bits_groupCounter                       (_stage1_2_dequeue_bits_groupCounter),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_2_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_2_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_2_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_2_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_2_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_2_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_2_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_2_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_2_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_2_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_2_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_2_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_2_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_2_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_2_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_2_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_2_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_2_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_2_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_2_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_2_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_2_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_2_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_2_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_2_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_2_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_2_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_2_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_2_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_2_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_2_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_2_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_2_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_2_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_2_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_2_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_2_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_2_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_2_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_2_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_2_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_2_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_2_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_2_dequeue_bits_decodeResult_logic),
    .enqueue_bits_vSew1H                             (_stage1_2_dequeue_bits_vSew1H),
    .enqueue_bits_csr_vl                             (_stage1_2_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_2_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_2_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_2_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_2_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_2_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_2_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage1_2_dequeue_bits_maskType),
    .enqueue_bits_laneIndex                          (_stage1_2_dequeue_bits_laneIndex),
    .enqueue_bits_instructionIndex                   (_stage1_2_dequeue_bits_instructionIndex),
    .dequeue_ready                                   (stage3EnqWire_2_ready),
    .dequeue_valid                                   (_executionUnit_2_dequeue_valid),
    .dequeue_bits_data                               (stage3EnqWire_2_bits_data),
    .dequeue_bits_ffoIndex                           (stage3EnqWire_2_bits_ffoIndex),
    .vfuRequest_ready                                (executeEnqueueFire_2),
    .vfuRequest_valid                                (_executionUnit_2_vfuRequest_valid),
    .vfuRequest_bits_src_0                           (requestVec_2_src_0),
    .vfuRequest_bits_src_1                           (requestVec_2_src_1),
    .vfuRequest_bits_src_2                           (requestVec_2_src_2),
    .vfuRequest_bits_src_3                           (requestVec_2_src_3),
    .vfuRequest_bits_opcode                          (requestVec_2_opcode),
    .vfuRequest_bits_mask                            (requestVec_2_mask),
    .vfuRequest_bits_executeMask                     (requestVec_2_executeMask),
    .vfuRequest_bits_sign0                           (requestVec_2_sign0),
    .vfuRequest_bits_sign                            (requestVec_2_sign),
    .vfuRequest_bits_reverse                         (requestVec_2_reverse),
    .vfuRequest_bits_average                         (requestVec_2_average),
    .vfuRequest_bits_saturate                        (requestVec_2_saturate),
    .vfuRequest_bits_vxrm                            (requestVec_2_vxrm),
    .vfuRequest_bits_vSew                            (requestVec_2_vSew),
    .vfuRequest_bits_shifterSize                     (requestVec_2_shifterSize),
    .vfuRequest_bits_rem                             (requestVec_2_rem),
    .vfuRequest_bits_groupIndex                      (requestVec_2_groupIndex),
    .vfuRequest_bits_laneIndex                       (requestVec_2_laneIndex),
    .vfuRequest_bits_maskType                        (requestVec_2_maskType),
    .vfuRequest_bits_narrow                          (requestVec_2_narrow),
    .dataResponse_valid                              (responseVec_2_valid),
    .dataResponse_bits_data                          (responseVec_2_bits_data),
    .executeDecode_specialSlot                       (executeDecodeVec_2_specialSlot),
    .executeDecode_topUop                            (executeDecodeVec_2_topUop),
    .executeDecode_popCount                          (executeDecodeVec_2_popCount),
    .executeDecode_ffo                               (executeDecodeVec_2_ffo),
    .executeDecode_average                           (executeDecodeVec_2_average),
    .executeDecode_reverse                           (executeDecodeVec_2_reverse),
    .executeDecode_dontNeedExecuteInLane             (executeDecodeVec_2_dontNeedExecuteInLane),
    .executeDecode_scheduler                         (executeDecodeVec_2_scheduler),
    .executeDecode_sReadVD                           (executeDecodeVec_2_sReadVD),
    .executeDecode_vtype                             (executeDecodeVec_2_vtype),
    .executeDecode_sWrite                            (executeDecodeVec_2_sWrite),
    .executeDecode_crossRead                         (executeDecodeVec_2_crossRead),
    .executeDecode_crossWrite                        (executeDecodeVec_2_crossWrite),
    .executeDecode_maskUnit                          (executeDecodeVec_2_maskUnit),
    .executeDecode_special                           (executeDecodeVec_2_special),
    .executeDecode_saturate                          (executeDecodeVec_2_saturate),
    .executeDecode_vwmacc                            (executeDecodeVec_2_vwmacc),
    .executeDecode_readOnly                          (executeDecodeVec_2_readOnly),
    .executeDecode_maskSource                        (executeDecodeVec_2_maskSource),
    .executeDecode_maskDestination                   (executeDecodeVec_2_maskDestination),
    .executeDecode_maskLogic                         (executeDecodeVec_2_maskLogic),
    .executeDecode_uop                               (executeDecodeVec_2_uop),
    .executeDecode_iota                              (executeDecodeVec_2_iota),
    .executeDecode_mv                                (executeDecodeVec_2_mv),
    .executeDecode_extend                            (executeDecodeVec_2_extend),
    .executeDecode_unOrderWrite                      (executeDecodeVec_2_unOrderWrite),
    .executeDecode_compress                          (executeDecodeVec_2_compress),
    .executeDecode_gather16                          (executeDecodeVec_2_gather16),
    .executeDecode_gather                            (executeDecodeVec_2_gather),
    .executeDecode_slid                              (executeDecodeVec_2_slid),
    .executeDecode_targetRd                          (executeDecodeVec_2_targetRd),
    .executeDecode_widenReduce                       (executeDecodeVec_2_widenReduce),
    .executeDecode_red                               (executeDecodeVec_2_red),
    .executeDecode_nr                                (executeDecodeVec_2_nr),
    .executeDecode_itype                             (executeDecodeVec_2_itype),
    .executeDecode_unsigned1                         (executeDecodeVec_2_unsigned1),
    .executeDecode_unsigned0                         (executeDecodeVec_2_unsigned0),
    .executeDecode_other                             (executeDecodeVec_2_other),
    .executeDecode_multiCycle                        (executeDecodeVec_2_multiCycle),
    .executeDecode_divider                           (executeDecodeVec_2_divider),
    .executeDecode_multiplier                        (executeDecodeVec_2_multiplier),
    .executeDecode_shift                             (executeDecodeVec_2_shift),
    .executeDecode_adder                             (executeDecodeVec_2_adder),
    .executeDecode_logic                             (executeDecodeVec_2_logic),
    .responseDecode_specialSlot                      (responseDecodeVec_2_specialSlot),
    .responseDecode_topUop                           (responseDecodeVec_2_topUop),
    .responseDecode_popCount                         (responseDecodeVec_2_popCount),
    .responseDecode_ffo                              (responseDecodeVec_2_ffo),
    .responseDecode_average                          (responseDecodeVec_2_average),
    .responseDecode_reverse                          (responseDecodeVec_2_reverse),
    .responseDecode_dontNeedExecuteInLane            (responseDecodeVec_2_dontNeedExecuteInLane),
    .responseDecode_scheduler                        (responseDecodeVec_2_scheduler),
    .responseDecode_sReadVD                          (responseDecodeVec_2_sReadVD),
    .responseDecode_vtype                            (responseDecodeVec_2_vtype),
    .responseDecode_sWrite                           (responseDecodeVec_2_sWrite),
    .responseDecode_crossRead                        (responseDecodeVec_2_crossRead),
    .responseDecode_crossWrite                       (responseDecodeVec_2_crossWrite),
    .responseDecode_maskUnit                         (responseDecodeVec_2_maskUnit),
    .responseDecode_special                          (responseDecodeVec_2_special),
    .responseDecode_saturate                         (responseDecodeVec_2_saturate),
    .responseDecode_vwmacc                           (responseDecodeVec_2_vwmacc),
    .responseDecode_readOnly                         (responseDecodeVec_2_readOnly),
    .responseDecode_maskSource                       (responseDecodeVec_2_maskSource),
    .responseDecode_maskDestination                  (responseDecodeVec_2_maskDestination),
    .responseDecode_maskLogic                        (responseDecodeVec_2_maskLogic),
    .responseDecode_uop                              (responseDecodeVec_2_uop),
    .responseDecode_iota                             (responseDecodeVec_2_iota),
    .responseDecode_mv                               (responseDecodeVec_2_mv),
    .responseDecode_extend                           (responseDecodeVec_2_extend),
    .responseDecode_unOrderWrite                     (responseDecodeVec_2_unOrderWrite),
    .responseDecode_compress                         (responseDecodeVec_2_compress),
    .responseDecode_gather16                         (responseDecodeVec_2_gather16),
    .responseDecode_gather                           (responseDecodeVec_2_gather),
    .responseDecode_slid                             (responseDecodeVec_2_slid),
    .responseDecode_targetRd                         (responseDecodeVec_2_targetRd),
    .responseDecode_widenReduce                      (responseDecodeVec_2_widenReduce),
    .responseDecode_red                              (responseDecodeVec_2_red),
    .responseDecode_nr                               (responseDecodeVec_2_nr),
    .responseDecode_itype                            (responseDecodeVec_2_itype),
    .responseDecode_unsigned1                        (responseDecodeVec_2_unsigned1),
    .responseDecode_unsigned0                        (responseDecodeVec_2_unsigned0),
    .responseDecode_other                            (responseDecodeVec_2_other),
    .responseDecode_multiCycle                       (responseDecodeVec_2_multiCycle),
    .responseDecode_divider                          (responseDecodeVec_2_divider),
    .responseDecode_multiplier                       (responseDecodeVec_2_multiplier),
    .responseDecode_shift                            (responseDecodeVec_2_shift),
    .responseDecode_adder                            (responseDecodeVec_2_adder),
    .responseDecode_logic                            (responseDecodeVec_2_logic),
    .responseIndex                                   (_executionUnit_2_responseIndex)
  );
  LaneStage3_1 stage3_2 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (stage3EnqWire_2_ready),
    .enqueue_valid                                   (stage3EnqWire_2_valid),
    .enqueue_bits_groupCounter                       (stage3EnqWire_2_bits_groupCounter),
    .enqueue_bits_data                               (stage3EnqWire_2_bits_data),
    .enqueue_bits_mask                               (stage3EnqWire_2_bits_mask),
    .enqueue_bits_ffoIndex                           (stage3EnqWire_2_bits_ffoIndex),
    .enqueue_bits_decodeResult_specialSlot           (stage3EnqWire_2_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (stage3EnqWire_2_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (stage3EnqWire_2_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (stage3EnqWire_2_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (stage3EnqWire_2_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (stage3EnqWire_2_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_2_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (stage3EnqWire_2_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (stage3EnqWire_2_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (stage3EnqWire_2_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (stage3EnqWire_2_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (stage3EnqWire_2_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (stage3EnqWire_2_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (stage3EnqWire_2_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (stage3EnqWire_2_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (stage3EnqWire_2_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (stage3EnqWire_2_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (stage3EnqWire_2_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (stage3EnqWire_2_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (stage3EnqWire_2_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (stage3EnqWire_2_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (stage3EnqWire_2_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (stage3EnqWire_2_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (stage3EnqWire_2_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (stage3EnqWire_2_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (stage3EnqWire_2_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (stage3EnqWire_2_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (stage3EnqWire_2_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (stage3EnqWire_2_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (stage3EnqWire_2_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (stage3EnqWire_2_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (stage3EnqWire_2_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (stage3EnqWire_2_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (stage3EnqWire_2_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (stage3EnqWire_2_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (stage3EnqWire_2_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (stage3EnqWire_2_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (stage3EnqWire_2_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (stage3EnqWire_2_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (stage3EnqWire_2_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (stage3EnqWire_2_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (stage3EnqWire_2_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (stage3EnqWire_2_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (stage3EnqWire_2_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (stage3EnqWire_2_bits_instructionIndex),
    .enqueue_bits_loadStore                          (stage3EnqWire_2_bits_loadStore),
    .enqueue_bits_vd                                 (stage3EnqWire_2_bits_vd),
    .vrfWriteRequest_ready                           (vrfWriteArbiter_2_ready),
    .vrfWriteRequest_valid                           (_stage3_2_vrfWriteRequest_valid),
    .vrfWriteRequest_bits_vd                         (vrfWriteArbiter_2_bits_vd),
    .vrfWriteRequest_bits_offset                     (vrfWriteArbiter_2_bits_offset),
    .vrfWriteRequest_bits_mask                       (_stage3_2_vrfWriteRequest_bits_mask),
    .vrfWriteRequest_bits_data                       (vrfWriteArbiter_2_bits_data),
    .vrfWriteRequest_bits_last                       (vrfWriteArbiter_2_bits_last),
    .vrfWriteRequest_bits_instructionIndex           (_stage3_2_vrfWriteRequest_bits_instructionIndex)
  );
  LaneStage0_1 stage0_3 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage0_3_enqueue_ready),
    .enqueue_valid                                   (stage0_3_enqueue_valid),
    .enqueue_bits_maskIndex                          (maskIndexVec_3),
    .enqueue_bits_maskForMaskGroup                   (slotControl_3_mask_bits),
    .enqueue_bits_maskGroupCount                     (maskGroupCountVec_3),
    .enqueue_bits_readFromScalar                     (slotControl_3_laneRequest_readFromScalar),
    .enqueue_bits_vSew1H                             (laneState_3_vSew1H),
    .enqueue_bits_loadStore                          (laneState_3_loadStore),
    .enqueue_bits_laneIndex                          (laneState_3_laneIndex),
    .enqueue_bits_decodeResult_specialSlot           (laneState_3_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (laneState_3_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (laneState_3_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (laneState_3_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (laneState_3_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (laneState_3_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (laneState_3_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (laneState_3_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (laneState_3_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (laneState_3_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (laneState_3_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (laneState_3_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (laneState_3_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (laneState_3_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (laneState_3_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (laneState_3_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (laneState_3_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (laneState_3_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (laneState_3_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (laneState_3_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (laneState_3_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (laneState_3_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (laneState_3_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (laneState_3_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (laneState_3_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (laneState_3_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (laneState_3_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (laneState_3_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (laneState_3_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (laneState_3_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (laneState_3_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (laneState_3_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (laneState_3_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (laneState_3_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (laneState_3_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (laneState_3_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (laneState_3_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (laneState_3_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (laneState_3_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (laneState_3_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (laneState_3_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (laneState_3_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (laneState_3_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (laneState_3_decodeResult_logic),
    .enqueue_bits_lastGroupForInstruction            (laneState_3_lastGroupForInstruction),
    .enqueue_bits_isLastLaneForInstruction           (laneState_3_isLastLaneForInstruction),
    .enqueue_bits_instructionFinished                (laneState_3_instructionFinished),
    .enqueue_bits_csr_vl                             (laneState_3_csr_vl),
    .enqueue_bits_csr_vStart                         (laneState_3_csr_vStart),
    .enqueue_bits_csr_vlmul                          (laneState_3_csr_vlmul),
    .enqueue_bits_csr_vSew                           (laneState_3_csr_vSew),
    .enqueue_bits_csr_vxrm                           (laneState_3_csr_vxrm),
    .enqueue_bits_csr_vta                            (laneState_3_csr_vta),
    .enqueue_bits_csr_vma                            (laneState_3_csr_vma),
    .enqueue_bits_maskType                           (laneState_3_maskType),
    .enqueue_bits_maskNotMaskedElement               (laneState_3_maskNotMaskedElement),
    .enqueue_bits_vs1                                (laneState_3_vs1),
    .enqueue_bits_vs2                                (laneState_3_vs2),
    .enqueue_bits_vd                                 (laneState_3_vd),
    .enqueue_bits_instructionIndex                   (laneState_3_instructionIndex),
    .enqueue_bits_additionalRW                       (laneState_3_additionalRW),
    .enqueue_bits_skipRead                           (laneState_3_skipRead),
    .enqueue_bits_skipEnable                         (laneState_3_skipEnable),
    .dequeue_ready                                   (_stage1_3_enqueue_ready),
    .dequeue_valid                                   (_stage0_3_dequeue_valid),
    .dequeue_bits_maskForMaskInput                   (_stage0_3_dequeue_bits_maskForMaskInput),
    .dequeue_bits_boundaryMaskCorrection             (_stage0_3_dequeue_bits_boundaryMaskCorrection),
    .dequeue_bits_groupCounter                       (_stage0_3_dequeue_bits_groupCounter),
    .dequeue_bits_readFromScalar                     (_stage0_3_dequeue_bits_readFromScalar),
    .dequeue_bits_instructionIndex                   (_stage0_3_dequeue_bits_instructionIndex),
    .dequeue_bits_decodeResult_specialSlot           (_stage0_3_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage0_3_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage0_3_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage0_3_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage0_3_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage0_3_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage0_3_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage0_3_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage0_3_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage0_3_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage0_3_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage0_3_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage0_3_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage0_3_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage0_3_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage0_3_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage0_3_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage0_3_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage0_3_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage0_3_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage0_3_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage0_3_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage0_3_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage0_3_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage0_3_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage0_3_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage0_3_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage0_3_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage0_3_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage0_3_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage0_3_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage0_3_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage0_3_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage0_3_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage0_3_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage0_3_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage0_3_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage0_3_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage0_3_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage0_3_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage0_3_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage0_3_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage0_3_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage0_3_dequeue_bits_decodeResult_logic),
    .dequeue_bits_laneIndex                          (_stage0_3_dequeue_bits_laneIndex),
    .dequeue_bits_skipRead                           (_stage0_3_dequeue_bits_skipRead),
    .dequeue_bits_vs1                                (_stage0_3_dequeue_bits_vs1),
    .dequeue_bits_vs2                                (_stage0_3_dequeue_bits_vs2),
    .dequeue_bits_vd                                 (_stage0_3_dequeue_bits_vd),
    .dequeue_bits_vSew1H                             (_stage0_3_dequeue_bits_vSew1H),
    .dequeue_bits_maskNotMaskedElement               (_stage0_3_dequeue_bits_maskNotMaskedElement),
    .dequeue_bits_csr_vl                             (_stage0_3_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage0_3_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage0_3_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage0_3_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage0_3_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage0_3_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage0_3_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage0_3_dequeue_bits_maskType),
    .dequeue_bits_loadStore                          (_stage0_3_dequeue_bits_loadStore),
    .dequeue_bits_bordersForMaskLogic                (_stage0_3_dequeue_bits_bordersForMaskLogic),
    .updateLaneState_maskGroupCount                  (_stage0_3_updateLaneState_maskGroupCount),
    .updateLaneState_maskIndex                       (_stage0_3_updateLaneState_maskIndex),
    .updateLaneState_outOfExecutionRange             (_stage0_3_updateLaneState_outOfExecutionRange),
    .updateLaneState_maskExhausted                   (_stage0_3_updateLaneState_maskExhausted),
    .tokenReport_valid                               (_stage0_3_tokenReport_valid),
    .tokenReport_bits_decodeResult_sWrite            (_stage0_3_tokenReport_bits_decodeResult_sWrite),
    .tokenReport_bits_decodeResult_maskUnit          (_stage0_3_tokenReport_bits_decodeResult_maskUnit),
    .tokenReport_bits_instructionIndex               (_stage0_3_tokenReport_bits_instructionIndex)
  );
  LaneStage1_1 stage1_3 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage1_3_enqueue_ready),
    .enqueue_valid                                   (_stage0_3_dequeue_valid),
    .enqueue_bits_groupCounter                       (_stage0_3_dequeue_bits_groupCounter),
    .enqueue_bits_maskForMaskInput                   (_stage0_3_dequeue_bits_maskForMaskInput),
    .enqueue_bits_boundaryMaskCorrection             (_stage0_3_dequeue_bits_boundaryMaskCorrection),
    .enqueue_bits_instructionIndex                   (_stage0_3_dequeue_bits_instructionIndex),
    .enqueue_bits_decodeResult_specialSlot           (_stage0_3_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage0_3_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage0_3_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage0_3_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage0_3_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage0_3_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage0_3_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage0_3_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage0_3_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage0_3_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage0_3_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage0_3_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage0_3_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage0_3_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage0_3_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage0_3_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage0_3_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage0_3_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage0_3_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage0_3_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage0_3_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage0_3_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage0_3_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage0_3_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage0_3_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage0_3_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage0_3_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage0_3_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage0_3_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage0_3_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage0_3_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage0_3_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage0_3_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage0_3_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage0_3_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage0_3_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage0_3_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage0_3_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage0_3_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage0_3_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage0_3_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage0_3_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage0_3_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage0_3_dequeue_bits_decodeResult_logic),
    .enqueue_bits_laneIndex                          (_stage0_3_dequeue_bits_laneIndex),
    .enqueue_bits_skipRead                           (_stage0_3_dequeue_bits_skipRead),
    .enqueue_bits_vs1                                (_stage0_3_dequeue_bits_vs1),
    .enqueue_bits_vs2                                (_stage0_3_dequeue_bits_vs2),
    .enqueue_bits_vd                                 (_stage0_3_dequeue_bits_vd),
    .enqueue_bits_vSew1H                             (_stage0_3_dequeue_bits_vSew1H),
    .enqueue_bits_maskNotMaskedElement               (_stage0_3_dequeue_bits_maskNotMaskedElement),
    .enqueue_bits_csr_vl                             (_stage0_3_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage0_3_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage0_3_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage0_3_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage0_3_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage0_3_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage0_3_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage0_3_dequeue_bits_maskType),
    .enqueue_bits_loadStore                          (_stage0_3_dequeue_bits_loadStore),
    .enqueue_bits_readFromScalar                     (_stage0_3_dequeue_bits_readFromScalar),
    .enqueue_bits_bordersForMaskLogic                (_stage0_3_dequeue_bits_bordersForMaskLogic),
    .dequeue_ready                                   (_stage2_3_enqueue_ready & _executionUnit_3_enqueue_ready),
    .dequeue_valid                                   (_stage1_3_dequeue_valid),
    .dequeue_bits_maskForFilter                      (_stage1_3_dequeue_bits_maskForFilter),
    .dequeue_bits_mask                               (_stage1_3_dequeue_bits_mask),
    .dequeue_bits_groupCounter                       (_stage1_3_dequeue_bits_groupCounter),
    .dequeue_bits_src_0                              (_stage1_3_dequeue_bits_src_0),
    .dequeue_bits_src_1                              (_stage1_3_dequeue_bits_src_1),
    .dequeue_bits_src_2                              (_stage1_3_dequeue_bits_src_2),
    .dequeue_bits_decodeResult_specialSlot           (_stage1_3_dequeue_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (_stage1_3_dequeue_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (_stage1_3_dequeue_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (_stage1_3_dequeue_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (_stage1_3_dequeue_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (_stage1_3_dequeue_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (_stage1_3_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (_stage1_3_dequeue_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (_stage1_3_dequeue_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (_stage1_3_dequeue_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (_stage1_3_dequeue_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (_stage1_3_dequeue_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (_stage1_3_dequeue_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (_stage1_3_dequeue_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (_stage1_3_dequeue_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (_stage1_3_dequeue_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (_stage1_3_dequeue_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (_stage1_3_dequeue_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (_stage1_3_dequeue_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (_stage1_3_dequeue_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (_stage1_3_dequeue_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (_stage1_3_dequeue_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (_stage1_3_dequeue_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (_stage1_3_dequeue_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (_stage1_3_dequeue_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (_stage1_3_dequeue_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (_stage1_3_dequeue_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (_stage1_3_dequeue_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (_stage1_3_dequeue_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (_stage1_3_dequeue_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (_stage1_3_dequeue_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (_stage1_3_dequeue_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (_stage1_3_dequeue_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (_stage1_3_dequeue_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (_stage1_3_dequeue_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (_stage1_3_dequeue_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (_stage1_3_dequeue_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (_stage1_3_dequeue_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (_stage1_3_dequeue_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (_stage1_3_dequeue_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (_stage1_3_dequeue_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (_stage1_3_dequeue_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (_stage1_3_dequeue_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (_stage1_3_dequeue_bits_decodeResult_logic),
    .dequeue_bits_vSew1H                             (_stage1_3_dequeue_bits_vSew1H),
    .dequeue_bits_csr_vl                             (_stage1_3_dequeue_bits_csr_vl),
    .dequeue_bits_csr_vStart                         (_stage1_3_dequeue_bits_csr_vStart),
    .dequeue_bits_csr_vlmul                          (_stage1_3_dequeue_bits_csr_vlmul),
    .dequeue_bits_csr_vSew                           (_stage1_3_dequeue_bits_csr_vSew),
    .dequeue_bits_csr_vxrm                           (_stage1_3_dequeue_bits_csr_vxrm),
    .dequeue_bits_csr_vta                            (_stage1_3_dequeue_bits_csr_vta),
    .dequeue_bits_csr_vma                            (_stage1_3_dequeue_bits_csr_vma),
    .dequeue_bits_maskType                           (_stage1_3_dequeue_bits_maskType),
    .dequeue_bits_laneIndex                          (_stage1_3_dequeue_bits_laneIndex),
    .dequeue_bits_instructionIndex                   (_stage1_3_dequeue_bits_instructionIndex),
    .dequeue_bits_loadStore                          (_stage1_3_dequeue_bits_loadStore),
    .dequeue_bits_vd                                 (_stage1_3_dequeue_bits_vd),
    .dequeue_bits_bordersForMaskLogic                (_stage1_3_dequeue_bits_bordersForMaskLogic),
    .vrfReadRequest_0_ready                          (vrfReadRequest_3_0_ready),
    .vrfReadRequest_0_valid                          (vrfReadRequest_3_0_valid),
    .vrfReadRequest_0_bits_vs                        (vrfReadRequest_3_0_bits_vs),
    .vrfReadRequest_0_bits_readSource                (vrfReadRequest_3_0_bits_readSource),
    .vrfReadRequest_0_bits_offset                    (vrfReadRequest_3_0_bits_offset),
    .vrfReadRequest_0_bits_instructionIndex          (vrfReadRequest_3_0_bits_instructionIndex),
    .vrfReadRequest_1_ready                          (vrfReadRequest_3_1_ready),
    .vrfReadRequest_1_valid                          (vrfReadRequest_3_1_valid),
    .vrfReadRequest_1_bits_vs                        (vrfReadRequest_3_1_bits_vs),
    .vrfReadRequest_1_bits_readSource                (vrfReadRequest_3_1_bits_readSource),
    .vrfReadRequest_1_bits_offset                    (vrfReadRequest_3_1_bits_offset),
    .vrfReadRequest_1_bits_instructionIndex          (vrfReadRequest_3_1_bits_instructionIndex),
    .vrfReadRequest_2_ready                          (vrfReadRequest_3_2_ready),
    .vrfReadRequest_2_valid                          (vrfReadRequest_3_2_valid),
    .vrfReadRequest_2_bits_vs                        (vrfReadRequest_3_2_bits_vs),
    .vrfReadRequest_2_bits_readSource                (vrfReadRequest_3_2_bits_readSource),
    .vrfReadRequest_2_bits_offset                    (vrfReadRequest_3_2_bits_offset),
    .vrfReadRequest_2_bits_instructionIndex          (vrfReadRequest_3_2_bits_instructionIndex),
    .vrfCheckRequest_0_vs                            (readCheckRequestVec_0_vs),
    .vrfCheckRequest_0_readSource                    (readCheckRequestVec_0_readSource),
    .vrfCheckRequest_0_offset                        (readCheckRequestVec_0_offset),
    .vrfCheckRequest_0_instructionIndex              (readCheckRequestVec_0_instructionIndex),
    .vrfCheckRequest_1_vs                            (readCheckRequestVec_1_vs),
    .vrfCheckRequest_1_readSource                    (readCheckRequestVec_1_readSource),
    .vrfCheckRequest_1_offset                        (readCheckRequestVec_1_offset),
    .vrfCheckRequest_1_instructionIndex              (readCheckRequestVec_1_instructionIndex),
    .vrfCheckRequest_2_vs                            (readCheckRequestVec_2_vs),
    .vrfCheckRequest_2_readSource                    (readCheckRequestVec_2_readSource),
    .vrfCheckRequest_2_offset                        (readCheckRequestVec_2_offset),
    .vrfCheckRequest_2_instructionIndex              (readCheckRequestVec_2_instructionIndex),
    .checkResult_0                                   (readCheckResult_0),
    .checkResult_1                                   (readCheckResult_1),
    .checkResult_2                                   (readCheckResult_2),
    .vrfReadResult_0                                 (vrfReadResult_3_0),
    .vrfReadResult_1                                 (vrfReadResult_3_1),
    .vrfReadResult_2                                 (vrfReadResult_3_2)
  );
  LaneStage2_1 stage2_3 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_stage2_3_enqueue_ready),
    .enqueue_valid                                   (_stage1_3_dequeue_valid & _executionUnit_3_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_3_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_3_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_3_dequeue_bits_src_2),
    .enqueue_bits_groupCounter                       (_stage1_3_dequeue_bits_groupCounter),
    .enqueue_bits_maskForFilter                      (_stage1_3_dequeue_bits_maskForFilter),
    .enqueue_bits_mask                               (_stage1_3_dequeue_bits_mask),
    .enqueue_bits_bordersForMaskLogic                (_stage1_3_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_3_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_3_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_3_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_3_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_3_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_3_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_3_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_3_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_3_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_3_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_3_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_3_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_3_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_3_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_3_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_3_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_3_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_3_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_3_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_3_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_3_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_3_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_3_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_3_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_3_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_3_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_3_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_3_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_3_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_3_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_3_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_3_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_3_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_3_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_3_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_3_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_3_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_3_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_3_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_3_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_3_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_3_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_3_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_3_dequeue_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (_stage1_3_dequeue_bits_instructionIndex),
    .enqueue_bits_loadStore                          (_stage1_3_dequeue_bits_loadStore),
    .enqueue_bits_vd                                 (_stage1_3_dequeue_bits_vd),
    .enqueue_bits_csr_vl                             (_stage1_3_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_3_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_3_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_3_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_3_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_3_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_3_dequeue_bits_csr_vma),
    .enqueue_bits_vSew1H                             (_stage1_3_dequeue_bits_vSew1H),
    .enqueue_bits_maskType                           (_stage1_3_dequeue_bits_maskType),
    .dequeue_ready                                   (stage3EnqWire_3_ready & _executionUnit_3_dequeue_valid),
    .dequeue_valid                                   (_stage2_3_dequeue_valid),
    .dequeue_bits_groupCounter                       (stage3EnqWire_3_bits_groupCounter),
    .dequeue_bits_mask                               (stage3EnqWire_3_bits_mask),
    .dequeue_bits_decodeResult_specialSlot           (stage3EnqWire_3_bits_decodeResult_specialSlot),
    .dequeue_bits_decodeResult_topUop                (stage3EnqWire_3_bits_decodeResult_topUop),
    .dequeue_bits_decodeResult_popCount              (stage3EnqWire_3_bits_decodeResult_popCount),
    .dequeue_bits_decodeResult_ffo                   (stage3EnqWire_3_bits_decodeResult_ffo),
    .dequeue_bits_decodeResult_average               (stage3EnqWire_3_bits_decodeResult_average),
    .dequeue_bits_decodeResult_reverse               (stage3EnqWire_3_bits_decodeResult_reverse),
    .dequeue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_3_bits_decodeResult_dontNeedExecuteInLane),
    .dequeue_bits_decodeResult_scheduler             (stage3EnqWire_3_bits_decodeResult_scheduler),
    .dequeue_bits_decodeResult_sReadVD               (stage3EnqWire_3_bits_decodeResult_sReadVD),
    .dequeue_bits_decodeResult_vtype                 (stage3EnqWire_3_bits_decodeResult_vtype),
    .dequeue_bits_decodeResult_sWrite                (stage3EnqWire_3_bits_decodeResult_sWrite),
    .dequeue_bits_decodeResult_crossRead             (stage3EnqWire_3_bits_decodeResult_crossRead),
    .dequeue_bits_decodeResult_crossWrite            (stage3EnqWire_3_bits_decodeResult_crossWrite),
    .dequeue_bits_decodeResult_maskUnit              (stage3EnqWire_3_bits_decodeResult_maskUnit),
    .dequeue_bits_decodeResult_special               (stage3EnqWire_3_bits_decodeResult_special),
    .dequeue_bits_decodeResult_saturate              (stage3EnqWire_3_bits_decodeResult_saturate),
    .dequeue_bits_decodeResult_vwmacc                (stage3EnqWire_3_bits_decodeResult_vwmacc),
    .dequeue_bits_decodeResult_readOnly              (stage3EnqWire_3_bits_decodeResult_readOnly),
    .dequeue_bits_decodeResult_maskSource            (stage3EnqWire_3_bits_decodeResult_maskSource),
    .dequeue_bits_decodeResult_maskDestination       (stage3EnqWire_3_bits_decodeResult_maskDestination),
    .dequeue_bits_decodeResult_maskLogic             (stage3EnqWire_3_bits_decodeResult_maskLogic),
    .dequeue_bits_decodeResult_uop                   (stage3EnqWire_3_bits_decodeResult_uop),
    .dequeue_bits_decodeResult_iota                  (stage3EnqWire_3_bits_decodeResult_iota),
    .dequeue_bits_decodeResult_mv                    (stage3EnqWire_3_bits_decodeResult_mv),
    .dequeue_bits_decodeResult_extend                (stage3EnqWire_3_bits_decodeResult_extend),
    .dequeue_bits_decodeResult_unOrderWrite          (stage3EnqWire_3_bits_decodeResult_unOrderWrite),
    .dequeue_bits_decodeResult_compress              (stage3EnqWire_3_bits_decodeResult_compress),
    .dequeue_bits_decodeResult_gather16              (stage3EnqWire_3_bits_decodeResult_gather16),
    .dequeue_bits_decodeResult_gather                (stage3EnqWire_3_bits_decodeResult_gather),
    .dequeue_bits_decodeResult_slid                  (stage3EnqWire_3_bits_decodeResult_slid),
    .dequeue_bits_decodeResult_targetRd              (stage3EnqWire_3_bits_decodeResult_targetRd),
    .dequeue_bits_decodeResult_widenReduce           (stage3EnqWire_3_bits_decodeResult_widenReduce),
    .dequeue_bits_decodeResult_red                   (stage3EnqWire_3_bits_decodeResult_red),
    .dequeue_bits_decodeResult_nr                    (stage3EnqWire_3_bits_decodeResult_nr),
    .dequeue_bits_decodeResult_itype                 (stage3EnqWire_3_bits_decodeResult_itype),
    .dequeue_bits_decodeResult_unsigned1             (stage3EnqWire_3_bits_decodeResult_unsigned1),
    .dequeue_bits_decodeResult_unsigned0             (stage3EnqWire_3_bits_decodeResult_unsigned0),
    .dequeue_bits_decodeResult_other                 (stage3EnqWire_3_bits_decodeResult_other),
    .dequeue_bits_decodeResult_multiCycle            (stage3EnqWire_3_bits_decodeResult_multiCycle),
    .dequeue_bits_decodeResult_divider               (stage3EnqWire_3_bits_decodeResult_divider),
    .dequeue_bits_decodeResult_multiplier            (stage3EnqWire_3_bits_decodeResult_multiplier),
    .dequeue_bits_decodeResult_shift                 (stage3EnqWire_3_bits_decodeResult_shift),
    .dequeue_bits_decodeResult_adder                 (stage3EnqWire_3_bits_decodeResult_adder),
    .dequeue_bits_decodeResult_logic                 (stage3EnqWire_3_bits_decodeResult_logic),
    .dequeue_bits_instructionIndex                   (stage3EnqWire_3_bits_instructionIndex),
    .dequeue_bits_loadStore                          (stage3EnqWire_3_bits_loadStore),
    .dequeue_bits_vd                                 (stage3EnqWire_3_bits_vd)
  );
  LaneExecutionBridge_3 executionUnit_3 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (_executionUnit_3_enqueue_ready),
    .enqueue_valid                                   (_stage1_3_dequeue_valid & _stage2_3_enqueue_ready),
    .enqueue_bits_src_0                              (_stage1_3_dequeue_bits_src_0),
    .enqueue_bits_src_1                              (_stage1_3_dequeue_bits_src_1),
    .enqueue_bits_src_2                              (_stage1_3_dequeue_bits_src_2),
    .enqueue_bits_bordersForMaskLogic                (_stage1_3_dequeue_bits_bordersForMaskLogic),
    .enqueue_bits_mask                               (_stage1_3_dequeue_bits_mask),
    .enqueue_bits_maskForFilter                      (_stage1_3_dequeue_bits_maskForFilter),
    .enqueue_bits_groupCounter                       (_stage1_3_dequeue_bits_groupCounter),
    .enqueue_bits_decodeResult_specialSlot           (_stage1_3_dequeue_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (_stage1_3_dequeue_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (_stage1_3_dequeue_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (_stage1_3_dequeue_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (_stage1_3_dequeue_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (_stage1_3_dequeue_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (_stage1_3_dequeue_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (_stage1_3_dequeue_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (_stage1_3_dequeue_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (_stage1_3_dequeue_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (_stage1_3_dequeue_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (_stage1_3_dequeue_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (_stage1_3_dequeue_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (_stage1_3_dequeue_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (_stage1_3_dequeue_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (_stage1_3_dequeue_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (_stage1_3_dequeue_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (_stage1_3_dequeue_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (_stage1_3_dequeue_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (_stage1_3_dequeue_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (_stage1_3_dequeue_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (_stage1_3_dequeue_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (_stage1_3_dequeue_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (_stage1_3_dequeue_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (_stage1_3_dequeue_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (_stage1_3_dequeue_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (_stage1_3_dequeue_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (_stage1_3_dequeue_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (_stage1_3_dequeue_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (_stage1_3_dequeue_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (_stage1_3_dequeue_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (_stage1_3_dequeue_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (_stage1_3_dequeue_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (_stage1_3_dequeue_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (_stage1_3_dequeue_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (_stage1_3_dequeue_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (_stage1_3_dequeue_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (_stage1_3_dequeue_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (_stage1_3_dequeue_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (_stage1_3_dequeue_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (_stage1_3_dequeue_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (_stage1_3_dequeue_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (_stage1_3_dequeue_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (_stage1_3_dequeue_bits_decodeResult_logic),
    .enqueue_bits_vSew1H                             (_stage1_3_dequeue_bits_vSew1H),
    .enqueue_bits_csr_vl                             (_stage1_3_dequeue_bits_csr_vl),
    .enqueue_bits_csr_vStart                         (_stage1_3_dequeue_bits_csr_vStart),
    .enqueue_bits_csr_vlmul                          (_stage1_3_dequeue_bits_csr_vlmul),
    .enqueue_bits_csr_vSew                           (_stage1_3_dequeue_bits_csr_vSew),
    .enqueue_bits_csr_vxrm                           (_stage1_3_dequeue_bits_csr_vxrm),
    .enqueue_bits_csr_vta                            (_stage1_3_dequeue_bits_csr_vta),
    .enqueue_bits_csr_vma                            (_stage1_3_dequeue_bits_csr_vma),
    .enqueue_bits_maskType                           (_stage1_3_dequeue_bits_maskType),
    .enqueue_bits_laneIndex                          (_stage1_3_dequeue_bits_laneIndex),
    .enqueue_bits_instructionIndex                   (_stage1_3_dequeue_bits_instructionIndex),
    .dequeue_ready                                   (stage3EnqWire_3_ready),
    .dequeue_valid                                   (_executionUnit_3_dequeue_valid),
    .dequeue_bits_data                               (stage3EnqWire_3_bits_data),
    .dequeue_bits_ffoIndex                           (stage3EnqWire_3_bits_ffoIndex),
    .vfuRequest_ready                                (executeEnqueueFire_3),
    .vfuRequest_valid                                (_executionUnit_3_vfuRequest_valid),
    .vfuRequest_bits_src_0                           (requestVec_3_src_0),
    .vfuRequest_bits_src_1                           (requestVec_3_src_1),
    .vfuRequest_bits_src_2                           (requestVec_3_src_2),
    .vfuRequest_bits_src_3                           (requestVec_3_src_3),
    .vfuRequest_bits_opcode                          (requestVec_3_opcode),
    .vfuRequest_bits_mask                            (requestVec_3_mask),
    .vfuRequest_bits_executeMask                     (requestVec_3_executeMask),
    .vfuRequest_bits_sign0                           (requestVec_3_sign0),
    .vfuRequest_bits_sign                            (requestVec_3_sign),
    .vfuRequest_bits_reverse                         (requestVec_3_reverse),
    .vfuRequest_bits_average                         (requestVec_3_average),
    .vfuRequest_bits_saturate                        (requestVec_3_saturate),
    .vfuRequest_bits_vxrm                            (requestVec_3_vxrm),
    .vfuRequest_bits_vSew                            (requestVec_3_vSew),
    .vfuRequest_bits_shifterSize                     (requestVec_3_shifterSize),
    .vfuRequest_bits_rem                             (requestVec_3_rem),
    .vfuRequest_bits_groupIndex                      (requestVec_3_groupIndex),
    .vfuRequest_bits_laneIndex                       (requestVec_3_laneIndex),
    .vfuRequest_bits_maskType                        (requestVec_3_maskType),
    .vfuRequest_bits_narrow                          (requestVec_3_narrow),
    .dataResponse_valid                              (responseVec_3_valid),
    .dataResponse_bits_data                          (responseVec_3_bits_data),
    .executeDecode_specialSlot                       (executeDecodeVec_3_specialSlot),
    .executeDecode_topUop                            (executeDecodeVec_3_topUop),
    .executeDecode_popCount                          (executeDecodeVec_3_popCount),
    .executeDecode_ffo                               (executeDecodeVec_3_ffo),
    .executeDecode_average                           (executeDecodeVec_3_average),
    .executeDecode_reverse                           (executeDecodeVec_3_reverse),
    .executeDecode_dontNeedExecuteInLane             (executeDecodeVec_3_dontNeedExecuteInLane),
    .executeDecode_scheduler                         (executeDecodeVec_3_scheduler),
    .executeDecode_sReadVD                           (executeDecodeVec_3_sReadVD),
    .executeDecode_vtype                             (executeDecodeVec_3_vtype),
    .executeDecode_sWrite                            (executeDecodeVec_3_sWrite),
    .executeDecode_crossRead                         (executeDecodeVec_3_crossRead),
    .executeDecode_crossWrite                        (executeDecodeVec_3_crossWrite),
    .executeDecode_maskUnit                          (executeDecodeVec_3_maskUnit),
    .executeDecode_special                           (executeDecodeVec_3_special),
    .executeDecode_saturate                          (executeDecodeVec_3_saturate),
    .executeDecode_vwmacc                            (executeDecodeVec_3_vwmacc),
    .executeDecode_readOnly                          (executeDecodeVec_3_readOnly),
    .executeDecode_maskSource                        (executeDecodeVec_3_maskSource),
    .executeDecode_maskDestination                   (executeDecodeVec_3_maskDestination),
    .executeDecode_maskLogic                         (executeDecodeVec_3_maskLogic),
    .executeDecode_uop                               (executeDecodeVec_3_uop),
    .executeDecode_iota                              (executeDecodeVec_3_iota),
    .executeDecode_mv                                (executeDecodeVec_3_mv),
    .executeDecode_extend                            (executeDecodeVec_3_extend),
    .executeDecode_unOrderWrite                      (executeDecodeVec_3_unOrderWrite),
    .executeDecode_compress                          (executeDecodeVec_3_compress),
    .executeDecode_gather16                          (executeDecodeVec_3_gather16),
    .executeDecode_gather                            (executeDecodeVec_3_gather),
    .executeDecode_slid                              (executeDecodeVec_3_slid),
    .executeDecode_targetRd                          (executeDecodeVec_3_targetRd),
    .executeDecode_widenReduce                       (executeDecodeVec_3_widenReduce),
    .executeDecode_red                               (executeDecodeVec_3_red),
    .executeDecode_nr                                (executeDecodeVec_3_nr),
    .executeDecode_itype                             (executeDecodeVec_3_itype),
    .executeDecode_unsigned1                         (executeDecodeVec_3_unsigned1),
    .executeDecode_unsigned0                         (executeDecodeVec_3_unsigned0),
    .executeDecode_other                             (executeDecodeVec_3_other),
    .executeDecode_multiCycle                        (executeDecodeVec_3_multiCycle),
    .executeDecode_divider                           (executeDecodeVec_3_divider),
    .executeDecode_multiplier                        (executeDecodeVec_3_multiplier),
    .executeDecode_shift                             (executeDecodeVec_3_shift),
    .executeDecode_adder                             (executeDecodeVec_3_adder),
    .executeDecode_logic                             (executeDecodeVec_3_logic),
    .responseDecode_specialSlot                      (responseDecodeVec_3_specialSlot),
    .responseDecode_topUop                           (responseDecodeVec_3_topUop),
    .responseDecode_popCount                         (responseDecodeVec_3_popCount),
    .responseDecode_ffo                              (responseDecodeVec_3_ffo),
    .responseDecode_average                          (responseDecodeVec_3_average),
    .responseDecode_reverse                          (responseDecodeVec_3_reverse),
    .responseDecode_dontNeedExecuteInLane            (responseDecodeVec_3_dontNeedExecuteInLane),
    .responseDecode_scheduler                        (responseDecodeVec_3_scheduler),
    .responseDecode_sReadVD                          (responseDecodeVec_3_sReadVD),
    .responseDecode_vtype                            (responseDecodeVec_3_vtype),
    .responseDecode_sWrite                           (responseDecodeVec_3_sWrite),
    .responseDecode_crossRead                        (responseDecodeVec_3_crossRead),
    .responseDecode_crossWrite                       (responseDecodeVec_3_crossWrite),
    .responseDecode_maskUnit                         (responseDecodeVec_3_maskUnit),
    .responseDecode_special                          (responseDecodeVec_3_special),
    .responseDecode_saturate                         (responseDecodeVec_3_saturate),
    .responseDecode_vwmacc                           (responseDecodeVec_3_vwmacc),
    .responseDecode_readOnly                         (responseDecodeVec_3_readOnly),
    .responseDecode_maskSource                       (responseDecodeVec_3_maskSource),
    .responseDecode_maskDestination                  (responseDecodeVec_3_maskDestination),
    .responseDecode_maskLogic                        (responseDecodeVec_3_maskLogic),
    .responseDecode_uop                              (responseDecodeVec_3_uop),
    .responseDecode_iota                             (responseDecodeVec_3_iota),
    .responseDecode_mv                               (responseDecodeVec_3_mv),
    .responseDecode_extend                           (responseDecodeVec_3_extend),
    .responseDecode_unOrderWrite                     (responseDecodeVec_3_unOrderWrite),
    .responseDecode_compress                         (responseDecodeVec_3_compress),
    .responseDecode_gather16                         (responseDecodeVec_3_gather16),
    .responseDecode_gather                           (responseDecodeVec_3_gather),
    .responseDecode_slid                             (responseDecodeVec_3_slid),
    .responseDecode_targetRd                         (responseDecodeVec_3_targetRd),
    .responseDecode_widenReduce                      (responseDecodeVec_3_widenReduce),
    .responseDecode_red                              (responseDecodeVec_3_red),
    .responseDecode_nr                               (responseDecodeVec_3_nr),
    .responseDecode_itype                            (responseDecodeVec_3_itype),
    .responseDecode_unsigned1                        (responseDecodeVec_3_unsigned1),
    .responseDecode_unsigned0                        (responseDecodeVec_3_unsigned0),
    .responseDecode_other                            (responseDecodeVec_3_other),
    .responseDecode_multiCycle                       (responseDecodeVec_3_multiCycle),
    .responseDecode_divider                          (responseDecodeVec_3_divider),
    .responseDecode_multiplier                       (responseDecodeVec_3_multiplier),
    .responseDecode_shift                            (responseDecodeVec_3_shift),
    .responseDecode_adder                            (responseDecodeVec_3_adder),
    .responseDecode_logic                            (responseDecodeVec_3_logic),
    .responseIndex                                   (_executionUnit_3_responseIndex)
  );
  LaneStage3_1 stage3_3 (
    .clock                                           (clock),
    .reset                                           (reset),
    .enqueue_ready                                   (stage3EnqWire_3_ready),
    .enqueue_valid                                   (stage3EnqWire_3_valid),
    .enqueue_bits_groupCounter                       (stage3EnqWire_3_bits_groupCounter),
    .enqueue_bits_data                               (stage3EnqWire_3_bits_data),
    .enqueue_bits_mask                               (stage3EnqWire_3_bits_mask),
    .enqueue_bits_ffoIndex                           (stage3EnqWire_3_bits_ffoIndex),
    .enqueue_bits_decodeResult_specialSlot           (stage3EnqWire_3_bits_decodeResult_specialSlot),
    .enqueue_bits_decodeResult_topUop                (stage3EnqWire_3_bits_decodeResult_topUop),
    .enqueue_bits_decodeResult_popCount              (stage3EnqWire_3_bits_decodeResult_popCount),
    .enqueue_bits_decodeResult_ffo                   (stage3EnqWire_3_bits_decodeResult_ffo),
    .enqueue_bits_decodeResult_average               (stage3EnqWire_3_bits_decodeResult_average),
    .enqueue_bits_decodeResult_reverse               (stage3EnqWire_3_bits_decodeResult_reverse),
    .enqueue_bits_decodeResult_dontNeedExecuteInLane (stage3EnqWire_3_bits_decodeResult_dontNeedExecuteInLane),
    .enqueue_bits_decodeResult_scheduler             (stage3EnqWire_3_bits_decodeResult_scheduler),
    .enqueue_bits_decodeResult_sReadVD               (stage3EnqWire_3_bits_decodeResult_sReadVD),
    .enqueue_bits_decodeResult_vtype                 (stage3EnqWire_3_bits_decodeResult_vtype),
    .enqueue_bits_decodeResult_sWrite                (stage3EnqWire_3_bits_decodeResult_sWrite),
    .enqueue_bits_decodeResult_crossRead             (stage3EnqWire_3_bits_decodeResult_crossRead),
    .enqueue_bits_decodeResult_crossWrite            (stage3EnqWire_3_bits_decodeResult_crossWrite),
    .enqueue_bits_decodeResult_maskUnit              (stage3EnqWire_3_bits_decodeResult_maskUnit),
    .enqueue_bits_decodeResult_special               (stage3EnqWire_3_bits_decodeResult_special),
    .enqueue_bits_decodeResult_saturate              (stage3EnqWire_3_bits_decodeResult_saturate),
    .enqueue_bits_decodeResult_vwmacc                (stage3EnqWire_3_bits_decodeResult_vwmacc),
    .enqueue_bits_decodeResult_readOnly              (stage3EnqWire_3_bits_decodeResult_readOnly),
    .enqueue_bits_decodeResult_maskSource            (stage3EnqWire_3_bits_decodeResult_maskSource),
    .enqueue_bits_decodeResult_maskDestination       (stage3EnqWire_3_bits_decodeResult_maskDestination),
    .enqueue_bits_decodeResult_maskLogic             (stage3EnqWire_3_bits_decodeResult_maskLogic),
    .enqueue_bits_decodeResult_uop                   (stage3EnqWire_3_bits_decodeResult_uop),
    .enqueue_bits_decodeResult_iota                  (stage3EnqWire_3_bits_decodeResult_iota),
    .enqueue_bits_decodeResult_mv                    (stage3EnqWire_3_bits_decodeResult_mv),
    .enqueue_bits_decodeResult_extend                (stage3EnqWire_3_bits_decodeResult_extend),
    .enqueue_bits_decodeResult_unOrderWrite          (stage3EnqWire_3_bits_decodeResult_unOrderWrite),
    .enqueue_bits_decodeResult_compress              (stage3EnqWire_3_bits_decodeResult_compress),
    .enqueue_bits_decodeResult_gather16              (stage3EnqWire_3_bits_decodeResult_gather16),
    .enqueue_bits_decodeResult_gather                (stage3EnqWire_3_bits_decodeResult_gather),
    .enqueue_bits_decodeResult_slid                  (stage3EnqWire_3_bits_decodeResult_slid),
    .enqueue_bits_decodeResult_targetRd              (stage3EnqWire_3_bits_decodeResult_targetRd),
    .enqueue_bits_decodeResult_widenReduce           (stage3EnqWire_3_bits_decodeResult_widenReduce),
    .enqueue_bits_decodeResult_red                   (stage3EnqWire_3_bits_decodeResult_red),
    .enqueue_bits_decodeResult_nr                    (stage3EnqWire_3_bits_decodeResult_nr),
    .enqueue_bits_decodeResult_itype                 (stage3EnqWire_3_bits_decodeResult_itype),
    .enqueue_bits_decodeResult_unsigned1             (stage3EnqWire_3_bits_decodeResult_unsigned1),
    .enqueue_bits_decodeResult_unsigned0             (stage3EnqWire_3_bits_decodeResult_unsigned0),
    .enqueue_bits_decodeResult_other                 (stage3EnqWire_3_bits_decodeResult_other),
    .enqueue_bits_decodeResult_multiCycle            (stage3EnqWire_3_bits_decodeResult_multiCycle),
    .enqueue_bits_decodeResult_divider               (stage3EnqWire_3_bits_decodeResult_divider),
    .enqueue_bits_decodeResult_multiplier            (stage3EnqWire_3_bits_decodeResult_multiplier),
    .enqueue_bits_decodeResult_shift                 (stage3EnqWire_3_bits_decodeResult_shift),
    .enqueue_bits_decodeResult_adder                 (stage3EnqWire_3_bits_decodeResult_adder),
    .enqueue_bits_decodeResult_logic                 (stage3EnqWire_3_bits_decodeResult_logic),
    .enqueue_bits_instructionIndex                   (stage3EnqWire_3_bits_instructionIndex),
    .enqueue_bits_loadStore                          (stage3EnqWire_3_bits_loadStore),
    .enqueue_bits_vd                                 (stage3EnqWire_3_bits_vd),
    .vrfWriteRequest_ready                           (vrfWriteArbiter_3_ready),
    .vrfWriteRequest_valid                           (_stage3_3_vrfWriteRequest_valid),
    .vrfWriteRequest_bits_vd                         (vrfWriteArbiter_3_bits_vd),
    .vrfWriteRequest_bits_offset                     (vrfWriteArbiter_3_bits_offset),
    .vrfWriteRequest_bits_mask                       (_stage3_3_vrfWriteRequest_bits_mask),
    .vrfWriteRequest_bits_data                       (vrfWriteArbiter_3_bits_data),
    .vrfWriteRequest_bits_last                       (vrfWriteArbiter_3_bits_last),
    .vrfWriteRequest_bits_instructionIndex           (_stage3_3_vrfWriteRequest_bits_instructionIndex)
  );
  MaskedLogic logic_0 (
    .clock                 (clock),
    .reset                 (reset),
    .requestIO_valid       (_vfuResponse_logicArbiter_io_out_valid),
    .requestIO_bits_tag    (_vfuResponse_logicArbiter_io_out_bits_tag),
    .requestIO_bits_src_0  (_vfuResponse_logicArbiter_io_out_bits_src_0[31:0]),
    .requestIO_bits_src_1  (_vfuResponse_logicArbiter_io_out_bits_src_1[31:0]),
    .requestIO_bits_src_2  (_vfuResponse_logicArbiter_io_out_bits_src_2[31:0]),
    .requestIO_bits_src_3  (_vfuResponse_logicArbiter_io_out_bits_src_3[31:0]),
    .requestIO_bits_opcode (_vfuResponse_logicArbiter_io_out_bits_opcode),
    .responseIO_valid      (vfuResponse_0_valid),
    .responseIO_bits_tag   (vfuResponse_0_bits_tag),
    .responseIO_bits_data  (vfuResponse_0_bits_data)
  );
  LaneAdder adder (
    .clock                         (clock),
    .reset                         (reset),
    .requestIO_valid               (_vfuResponse_adderArbiter_io_out_valid),
    .requestIO_bits_tag            (_vfuResponse_adderArbiter_io_out_bits_tag),
    .requestIO_bits_src_0          (_vfuResponse_adderArbiter_io_out_bits_src_0[31:0]),
    .requestIO_bits_src_1          (_vfuResponse_adderArbiter_io_out_bits_src_1[31:0]),
    .requestIO_bits_mask           (_vfuResponse_adderArbiter_io_out_bits_mask),
    .requestIO_bits_opcode         (_vfuResponse_adderArbiter_io_out_bits_opcode),
    .requestIO_bits_sign           (_vfuResponse_adderArbiter_io_out_bits_sign),
    .requestIO_bits_reverse        (_vfuResponse_adderArbiter_io_out_bits_reverse),
    .requestIO_bits_average        (_vfuResponse_adderArbiter_io_out_bits_average),
    .requestIO_bits_saturate       (_vfuResponse_adderArbiter_io_out_bits_saturate),
    .requestIO_bits_vxrm           (_vfuResponse_adderArbiter_io_out_bits_vxrm),
    .requestIO_bits_vSew           (_vfuResponse_adderArbiter_io_out_bits_vSew),
    .requestIO_bits_executeIndex   (_vfuResponse_adderArbiter_io_out_bits_executeIndex),
    .responseIO_valid              (vfuResponse_1_valid),
    .responseIO_bits_tag           (vfuResponse_1_bits_tag),
    .responseIO_bits_data          (vfuResponse_1_bits_data),
    .responseIO_bits_adderMaskResp (vfuResponse_1_bits_adderMaskResp),
    .responseIO_bits_vxsat         (vfuResponse_1_bits_vxsat),
    .responseIO_bits_executeIndex  (vfuResponse_1_bits_executeIndex)
  );
  LaneShifter shift (
    .clock                      (clock),
    .reset                      (reset),
    .requestIO_valid            (_vfuResponse_shiftDistributor_requestToVfu_valid),
    .requestIO_bits_tag         (_vfuResponse_shiftDistributor_requestToVfu_bits_tag),
    .requestIO_bits_src_0       (_vfuResponse_shiftDistributor_requestToVfu_bits_src_0[31:0]),
    .requestIO_bits_src_1       (_vfuResponse_shiftDistributor_requestToVfu_bits_src_1[31:0]),
    .requestIO_bits_shifterSize (_vfuResponse_shiftDistributor_requestToVfu_bits_shifterSize[4:0]),
    .requestIO_bits_opcode      (_vfuResponse_shiftDistributor_requestToVfu_bits_opcode[2:0]),
    .requestIO_bits_vxrm        (_vfuResponse_shiftDistributor_requestToVfu_bits_vxrm),
    .responseIO_valid           (vfuResponse_responseBundle_valid),
    .responseIO_bits_tag        (vfuResponse_responseBundle_bits_tag),
    .responseIO_bits_data       (vfuResponse_responseBundle_bits_data)
  );
  LaneMul multiplier (
    .clock                   (clock),
    .reset                   (reset),
    .requestIO_valid         (_vfuResponse_multiplierArbiter_io_out_valid),
    .requestIO_bits_tag      (_vfuResponse_multiplierArbiter_io_out_bits_tag),
    .requestIO_bits_src_0    (_vfuResponse_multiplierArbiter_io_out_bits_src_0[31:0]),
    .requestIO_bits_src_1    (_vfuResponse_multiplierArbiter_io_out_bits_src_1[31:0]),
    .requestIO_bits_src_2    (_vfuResponse_multiplierArbiter_io_out_bits_src_2[31:0]),
    .requestIO_bits_opcode   (_vfuResponse_multiplierArbiter_io_out_bits_opcode),
    .requestIO_bits_saturate (_vfuResponse_multiplierArbiter_io_out_bits_saturate),
    .requestIO_bits_vSew     (_vfuResponse_multiplierArbiter_io_out_bits_vSew),
    .requestIO_bits_sign0    (_vfuResponse_multiplierArbiter_io_out_bits_sign0),
    .requestIO_bits_sign     (_vfuResponse_multiplierArbiter_io_out_bits_sign),
    .requestIO_bits_vxrm     (_vfuResponse_multiplierArbiter_io_out_bits_vxrm),
    .responseIO_valid        (vfuResponse_3_valid),
    .responseIO_bits_tag     (vfuResponse_3_bits_tag),
    .responseIO_bits_data    (vfuResponse_3_bits_data),
    .responseIO_bits_vxsat   (_multiplier_responseIO_bits_vxsat)
  );
  LaneDiv divider (
    .clock                        (clock),
    .reset                        (reset),
    .requestIO_ready              (_divider_requestIO_ready),
    .requestIO_valid              (_vfuResponse_dividerDistributor_requestToVfu_valid),
    .requestIO_bits_tag           (_vfuResponse_dividerDistributor_requestToVfu_bits_tag),
    .requestIO_bits_src_0         (_vfuResponse_dividerDistributor_requestToVfu_bits_src_0[31:0]),
    .requestIO_bits_src_1         (_vfuResponse_dividerDistributor_requestToVfu_bits_src_1[31:0]),
    .requestIO_bits_opcode        (_vfuResponse_dividerDistributor_requestToVfu_bits_opcode),
    .requestIO_bits_sign          (_vfuResponse_dividerDistributor_requestToVfu_bits_sign),
    .requestIO_bits_executeIndex  (_vfuResponse_dividerDistributor_requestToVfu_bits_executeIndex),
    .responseIO_valid             (vfuResponse_responseBundle_1_valid),
    .responseIO_bits_tag          (vfuResponse_responseBundle_1_bits_tag),
    .responseIO_bits_data         (vfuResponse_responseBundle_1_bits_data),
    .responseIO_bits_executeIndex (vfuResponse_responseBundle_1_bits_executeIndex),
    .responseIO_bits_busy         (vrfIsBusy_4)
  );
  OtherUnit other (
    .clock                       (clock),
    .reset                       (reset),
    .requestIO_valid             (_vfuResponse_otherDistributor_requestToVfu_valid),
    .requestIO_bits_tag          (_vfuResponse_otherDistributor_requestToVfu_bits_tag),
    .requestIO_bits_src_0        (_vfuResponse_otherDistributor_requestToVfu_bits_src_0[31:0]),
    .requestIO_bits_src_1        (_vfuResponse_otherDistributor_requestToVfu_bits_src_1[31:0]),
    .requestIO_bits_src_2        (_vfuResponse_otherDistributor_requestToVfu_bits_src_2[31:0]),
    .requestIO_bits_src_3        (_vfuResponse_otherDistributor_requestToVfu_bits_src_3[31:0]),
    .requestIO_bits_popInit      (_vfuResponse_otherDistributor_requestToVfu_bits_popInit),
    .requestIO_bits_opcode       (_vfuResponse_otherDistributor_requestToVfu_bits_opcode),
    .requestIO_bits_groupIndex   (_vfuResponse_otherDistributor_requestToVfu_bits_groupIndex[8:0]),
    .requestIO_bits_laneIndex    (_vfuResponse_otherDistributor_requestToVfu_bits_laneIndex),
    .requestIO_bits_executeIndex (_vfuResponse_otherDistributor_requestToVfu_bits_executeIndex),
    .requestIO_bits_sign         (_vfuResponse_otherDistributor_requestToVfu_bits_sign),
    .requestIO_bits_mask         (_vfuResponse_otherDistributor_requestToVfu_bits_mask[0]),
    .requestIO_bits_maskType     (_vfuResponse_otherDistributor_requestToVfu_bits_maskType),
    .requestIO_bits_vSew         (_vfuResponse_otherDistributor_requestToVfu_bits_vSew),
    .requestIO_bits_vxrm         (_vfuResponse_otherDistributor_requestToVfu_bits_vxrm),
    .requestIO_bits_narrow       (_vfuResponse_otherDistributor_requestToVfu_bits_narrow),
    .responseIO_valid            (vfuResponse_responseBundle_2_valid),
    .responseIO_bits_tag         (vfuResponse_responseBundle_2_bits_tag),
    .responseIO_bits_data        (vfuResponse_responseBundle_2_bits_data),
    .responseIO_bits_clipFail    (vfuResponse_responseBundle_2_bits_clipFail),
    .responseIO_bits_ffoSuccess  (vfuResponse_responseBundle_2_bits_ffoSuccess)
  );
  Arbiter4_SlotRequestToVFU vfuResponse_logicArbiter (
    .io_in_0_ready             (requestVecFromSlot_0_logic_ready),
    .io_in_0_valid             (requestVecFromSlot_0_logic_valid),
    .io_in_0_bits_src_0        (requestVecFromSlot_0_logic_bits_src_0),
    .io_in_0_bits_src_1        (requestVecFromSlot_0_logic_bits_src_1),
    .io_in_0_bits_src_2        (requestVecFromSlot_0_logic_bits_src_2),
    .io_in_0_bits_src_3        (requestVecFromSlot_0_logic_bits_src_3),
    .io_in_0_bits_opcode       (requestVecFromSlot_0_logic_bits_opcode),
    .io_in_0_bits_mask         (requestVecFromSlot_0_logic_bits_mask),
    .io_in_0_bits_executeMask  (requestVecFromSlot_0_logic_bits_executeMask),
    .io_in_0_bits_sign0        (requestVecFromSlot_0_logic_bits_sign0),
    .io_in_0_bits_sign         (requestVecFromSlot_0_logic_bits_sign),
    .io_in_0_bits_reverse      (requestVecFromSlot_0_logic_bits_reverse),
    .io_in_0_bits_average      (requestVecFromSlot_0_logic_bits_average),
    .io_in_0_bits_saturate     (requestVecFromSlot_0_logic_bits_saturate),
    .io_in_0_bits_vxrm         (requestVecFromSlot_0_logic_bits_vxrm),
    .io_in_0_bits_vSew         (requestVecFromSlot_0_logic_bits_vSew),
    .io_in_0_bits_shifterSize  (requestVecFromSlot_0_logic_bits_shifterSize),
    .io_in_0_bits_rem          (requestVecFromSlot_0_logic_bits_rem),
    .io_in_0_bits_executeIndex (requestVecFromSlot_0_logic_bits_executeIndex),
    .io_in_0_bits_popInit      (requestVecFromSlot_0_logic_bits_popInit),
    .io_in_0_bits_groupIndex   (requestVecFromSlot_0_logic_bits_groupIndex),
    .io_in_0_bits_laneIndex    (requestVecFromSlot_0_logic_bits_laneIndex),
    .io_in_0_bits_maskType     (requestVecFromSlot_0_logic_bits_maskType),
    .io_in_0_bits_narrow       (requestVecFromSlot_0_logic_bits_narrow),
    .io_in_1_ready             (requestVecFromSlot_1_logic_ready),
    .io_in_1_valid             (requestVecFromSlot_1_logic_valid),
    .io_in_1_bits_src_0        (requestVecFromSlot_1_logic_bits_src_0),
    .io_in_1_bits_src_1        (requestVecFromSlot_1_logic_bits_src_1),
    .io_in_1_bits_src_2        (requestVecFromSlot_1_logic_bits_src_2),
    .io_in_1_bits_src_3        (requestVecFromSlot_1_logic_bits_src_3),
    .io_in_1_bits_opcode       (requestVecFromSlot_1_logic_bits_opcode),
    .io_in_1_bits_mask         (requestVecFromSlot_1_logic_bits_mask),
    .io_in_1_bits_executeMask  (requestVecFromSlot_1_logic_bits_executeMask),
    .io_in_1_bits_sign0        (requestVecFromSlot_1_logic_bits_sign0),
    .io_in_1_bits_sign         (requestVecFromSlot_1_logic_bits_sign),
    .io_in_1_bits_reverse      (requestVecFromSlot_1_logic_bits_reverse),
    .io_in_1_bits_average      (requestVecFromSlot_1_logic_bits_average),
    .io_in_1_bits_saturate     (requestVecFromSlot_1_logic_bits_saturate),
    .io_in_1_bits_vxrm         (requestVecFromSlot_1_logic_bits_vxrm),
    .io_in_1_bits_vSew         (requestVecFromSlot_1_logic_bits_vSew),
    .io_in_1_bits_shifterSize  (requestVecFromSlot_1_logic_bits_shifterSize),
    .io_in_1_bits_rem          (requestVecFromSlot_1_logic_bits_rem),
    .io_in_1_bits_groupIndex   (requestVecFromSlot_1_logic_bits_groupIndex),
    .io_in_1_bits_laneIndex    (requestVecFromSlot_1_logic_bits_laneIndex),
    .io_in_1_bits_maskType     (requestVecFromSlot_1_logic_bits_maskType),
    .io_in_1_bits_narrow       (requestVecFromSlot_1_logic_bits_narrow),
    .io_in_2_ready             (requestVecFromSlot_2_logic_ready),
    .io_in_2_valid             (requestVecFromSlot_2_logic_valid),
    .io_in_2_bits_src_0        (requestVecFromSlot_2_logic_bits_src_0),
    .io_in_2_bits_src_1        (requestVecFromSlot_2_logic_bits_src_1),
    .io_in_2_bits_src_2        (requestVecFromSlot_2_logic_bits_src_2),
    .io_in_2_bits_src_3        (requestVecFromSlot_2_logic_bits_src_3),
    .io_in_2_bits_opcode       (requestVecFromSlot_2_logic_bits_opcode),
    .io_in_2_bits_mask         (requestVecFromSlot_2_logic_bits_mask),
    .io_in_2_bits_executeMask  (requestVecFromSlot_2_logic_bits_executeMask),
    .io_in_2_bits_sign0        (requestVecFromSlot_2_logic_bits_sign0),
    .io_in_2_bits_sign         (requestVecFromSlot_2_logic_bits_sign),
    .io_in_2_bits_reverse      (requestVecFromSlot_2_logic_bits_reverse),
    .io_in_2_bits_average      (requestVecFromSlot_2_logic_bits_average),
    .io_in_2_bits_saturate     (requestVecFromSlot_2_logic_bits_saturate),
    .io_in_2_bits_vxrm         (requestVecFromSlot_2_logic_bits_vxrm),
    .io_in_2_bits_vSew         (requestVecFromSlot_2_logic_bits_vSew),
    .io_in_2_bits_shifterSize  (requestVecFromSlot_2_logic_bits_shifterSize),
    .io_in_2_bits_rem          (requestVecFromSlot_2_logic_bits_rem),
    .io_in_2_bits_groupIndex   (requestVecFromSlot_2_logic_bits_groupIndex),
    .io_in_2_bits_laneIndex    (requestVecFromSlot_2_logic_bits_laneIndex),
    .io_in_2_bits_maskType     (requestVecFromSlot_2_logic_bits_maskType),
    .io_in_2_bits_narrow       (requestVecFromSlot_2_logic_bits_narrow),
    .io_in_3_ready             (requestVecFromSlot_3_logic_ready),
    .io_in_3_valid             (requestVecFromSlot_3_logic_valid),
    .io_in_3_bits_src_0        (requestVecFromSlot_3_logic_bits_src_0),
    .io_in_3_bits_src_1        (requestVecFromSlot_3_logic_bits_src_1),
    .io_in_3_bits_src_2        (requestVecFromSlot_3_logic_bits_src_2),
    .io_in_3_bits_src_3        (requestVecFromSlot_3_logic_bits_src_3),
    .io_in_3_bits_opcode       (requestVecFromSlot_3_logic_bits_opcode),
    .io_in_3_bits_mask         (requestVecFromSlot_3_logic_bits_mask),
    .io_in_3_bits_executeMask  (requestVecFromSlot_3_logic_bits_executeMask),
    .io_in_3_bits_sign0        (requestVecFromSlot_3_logic_bits_sign0),
    .io_in_3_bits_sign         (requestVecFromSlot_3_logic_bits_sign),
    .io_in_3_bits_reverse      (requestVecFromSlot_3_logic_bits_reverse),
    .io_in_3_bits_average      (requestVecFromSlot_3_logic_bits_average),
    .io_in_3_bits_saturate     (requestVecFromSlot_3_logic_bits_saturate),
    .io_in_3_bits_vxrm         (requestVecFromSlot_3_logic_bits_vxrm),
    .io_in_3_bits_vSew         (requestVecFromSlot_3_logic_bits_vSew),
    .io_in_3_bits_shifterSize  (requestVecFromSlot_3_logic_bits_shifterSize),
    .io_in_3_bits_rem          (requestVecFromSlot_3_logic_bits_rem),
    .io_in_3_bits_groupIndex   (requestVecFromSlot_3_logic_bits_groupIndex),
    .io_in_3_bits_laneIndex    (requestVecFromSlot_3_logic_bits_laneIndex),
    .io_in_3_bits_maskType     (requestVecFromSlot_3_logic_bits_maskType),
    .io_in_3_bits_narrow       (requestVecFromSlot_3_logic_bits_narrow),
    .io_out_ready              (1'h1),
    .io_out_valid              (_vfuResponse_logicArbiter_io_out_valid),
    .io_out_bits_src_0         (_vfuResponse_logicArbiter_io_out_bits_src_0),
    .io_out_bits_src_1         (_vfuResponse_logicArbiter_io_out_bits_src_1),
    .io_out_bits_src_2         (_vfuResponse_logicArbiter_io_out_bits_src_2),
    .io_out_bits_src_3         (_vfuResponse_logicArbiter_io_out_bits_src_3),
    .io_out_bits_opcode        (_vfuResponse_logicArbiter_io_out_bits_opcode),
    .io_out_bits_mask          (/* unused */),
    .io_out_bits_executeMask   (/* unused */),
    .io_out_bits_sign0         (/* unused */),
    .io_out_bits_sign          (/* unused */),
    .io_out_bits_reverse       (/* unused */),
    .io_out_bits_average       (/* unused */),
    .io_out_bits_saturate      (/* unused */),
    .io_out_bits_vxrm          (/* unused */),
    .io_out_bits_vSew          (/* unused */),
    .io_out_bits_shifterSize   (/* unused */),
    .io_out_bits_rem           (/* unused */),
    .io_out_bits_executeIndex  (/* unused */),
    .io_out_bits_popInit       (/* unused */),
    .io_out_bits_groupIndex    (/* unused */),
    .io_out_bits_laneIndex     (/* unused */),
    .io_out_bits_maskType      (/* unused */),
    .io_out_bits_narrow        (/* unused */),
    .io_out_bits_tag           (_vfuResponse_logicArbiter_io_out_bits_tag)
  );
  Arbiter4_SlotRequestToVFU vfuResponse_adderArbiter (
    .io_in_0_ready             (requestVecFromSlot_0_adder_ready),
    .io_in_0_valid             (requestVecFromSlot_0_adder_valid),
    .io_in_0_bits_src_0        (requestVecFromSlot_0_adder_bits_src_0),
    .io_in_0_bits_src_1        (requestVecFromSlot_0_adder_bits_src_1),
    .io_in_0_bits_src_2        (requestVecFromSlot_0_adder_bits_src_2),
    .io_in_0_bits_src_3        (requestVecFromSlot_0_adder_bits_src_3),
    .io_in_0_bits_opcode       (requestVecFromSlot_0_adder_bits_opcode),
    .io_in_0_bits_mask         (requestVecFromSlot_0_adder_bits_mask),
    .io_in_0_bits_executeMask  (requestVecFromSlot_0_adder_bits_executeMask),
    .io_in_0_bits_sign0        (requestVecFromSlot_0_adder_bits_sign0),
    .io_in_0_bits_sign         (requestVecFromSlot_0_adder_bits_sign),
    .io_in_0_bits_reverse      (requestVecFromSlot_0_adder_bits_reverse),
    .io_in_0_bits_average      (requestVecFromSlot_0_adder_bits_average),
    .io_in_0_bits_saturate     (requestVecFromSlot_0_adder_bits_saturate),
    .io_in_0_bits_vxrm         (requestVecFromSlot_0_adder_bits_vxrm),
    .io_in_0_bits_vSew         (requestVecFromSlot_0_adder_bits_vSew),
    .io_in_0_bits_shifterSize  (requestVecFromSlot_0_adder_bits_shifterSize),
    .io_in_0_bits_rem          (requestVecFromSlot_0_adder_bits_rem),
    .io_in_0_bits_executeIndex (requestVecFromSlot_0_adder_bits_executeIndex),
    .io_in_0_bits_popInit      (requestVecFromSlot_0_adder_bits_popInit),
    .io_in_0_bits_groupIndex   (requestVecFromSlot_0_adder_bits_groupIndex),
    .io_in_0_bits_laneIndex    (requestVecFromSlot_0_adder_bits_laneIndex),
    .io_in_0_bits_maskType     (requestVecFromSlot_0_adder_bits_maskType),
    .io_in_0_bits_narrow       (requestVecFromSlot_0_adder_bits_narrow),
    .io_in_1_ready             (requestVecFromSlot_1_adder_ready),
    .io_in_1_valid             (requestVecFromSlot_1_adder_valid),
    .io_in_1_bits_src_0        (requestVecFromSlot_1_adder_bits_src_0),
    .io_in_1_bits_src_1        (requestVecFromSlot_1_adder_bits_src_1),
    .io_in_1_bits_src_2        (requestVecFromSlot_1_adder_bits_src_2),
    .io_in_1_bits_src_3        (requestVecFromSlot_1_adder_bits_src_3),
    .io_in_1_bits_opcode       (requestVecFromSlot_1_adder_bits_opcode),
    .io_in_1_bits_mask         (requestVecFromSlot_1_adder_bits_mask),
    .io_in_1_bits_executeMask  (requestVecFromSlot_1_adder_bits_executeMask),
    .io_in_1_bits_sign0        (requestVecFromSlot_1_adder_bits_sign0),
    .io_in_1_bits_sign         (requestVecFromSlot_1_adder_bits_sign),
    .io_in_1_bits_reverse      (requestVecFromSlot_1_adder_bits_reverse),
    .io_in_1_bits_average      (requestVecFromSlot_1_adder_bits_average),
    .io_in_1_bits_saturate     (requestVecFromSlot_1_adder_bits_saturate),
    .io_in_1_bits_vxrm         (requestVecFromSlot_1_adder_bits_vxrm),
    .io_in_1_bits_vSew         (requestVecFromSlot_1_adder_bits_vSew),
    .io_in_1_bits_shifterSize  (requestVecFromSlot_1_adder_bits_shifterSize),
    .io_in_1_bits_rem          (requestVecFromSlot_1_adder_bits_rem),
    .io_in_1_bits_groupIndex   (requestVecFromSlot_1_adder_bits_groupIndex),
    .io_in_1_bits_laneIndex    (requestVecFromSlot_1_adder_bits_laneIndex),
    .io_in_1_bits_maskType     (requestVecFromSlot_1_adder_bits_maskType),
    .io_in_1_bits_narrow       (requestVecFromSlot_1_adder_bits_narrow),
    .io_in_2_ready             (requestVecFromSlot_2_adder_ready),
    .io_in_2_valid             (requestVecFromSlot_2_adder_valid),
    .io_in_2_bits_src_0        (requestVecFromSlot_2_adder_bits_src_0),
    .io_in_2_bits_src_1        (requestVecFromSlot_2_adder_bits_src_1),
    .io_in_2_bits_src_2        (requestVecFromSlot_2_adder_bits_src_2),
    .io_in_2_bits_src_3        (requestVecFromSlot_2_adder_bits_src_3),
    .io_in_2_bits_opcode       (requestVecFromSlot_2_adder_bits_opcode),
    .io_in_2_bits_mask         (requestVecFromSlot_2_adder_bits_mask),
    .io_in_2_bits_executeMask  (requestVecFromSlot_2_adder_bits_executeMask),
    .io_in_2_bits_sign0        (requestVecFromSlot_2_adder_bits_sign0),
    .io_in_2_bits_sign         (requestVecFromSlot_2_adder_bits_sign),
    .io_in_2_bits_reverse      (requestVecFromSlot_2_adder_bits_reverse),
    .io_in_2_bits_average      (requestVecFromSlot_2_adder_bits_average),
    .io_in_2_bits_saturate     (requestVecFromSlot_2_adder_bits_saturate),
    .io_in_2_bits_vxrm         (requestVecFromSlot_2_adder_bits_vxrm),
    .io_in_2_bits_vSew         (requestVecFromSlot_2_adder_bits_vSew),
    .io_in_2_bits_shifterSize  (requestVecFromSlot_2_adder_bits_shifterSize),
    .io_in_2_bits_rem          (requestVecFromSlot_2_adder_bits_rem),
    .io_in_2_bits_groupIndex   (requestVecFromSlot_2_adder_bits_groupIndex),
    .io_in_2_bits_laneIndex    (requestVecFromSlot_2_adder_bits_laneIndex),
    .io_in_2_bits_maskType     (requestVecFromSlot_2_adder_bits_maskType),
    .io_in_2_bits_narrow       (requestVecFromSlot_2_adder_bits_narrow),
    .io_in_3_ready             (requestVecFromSlot_3_adder_ready),
    .io_in_3_valid             (requestVecFromSlot_3_adder_valid),
    .io_in_3_bits_src_0        (requestVecFromSlot_3_adder_bits_src_0),
    .io_in_3_bits_src_1        (requestVecFromSlot_3_adder_bits_src_1),
    .io_in_3_bits_src_2        (requestVecFromSlot_3_adder_bits_src_2),
    .io_in_3_bits_src_3        (requestVecFromSlot_3_adder_bits_src_3),
    .io_in_3_bits_opcode       (requestVecFromSlot_3_adder_bits_opcode),
    .io_in_3_bits_mask         (requestVecFromSlot_3_adder_bits_mask),
    .io_in_3_bits_executeMask  (requestVecFromSlot_3_adder_bits_executeMask),
    .io_in_3_bits_sign0        (requestVecFromSlot_3_adder_bits_sign0),
    .io_in_3_bits_sign         (requestVecFromSlot_3_adder_bits_sign),
    .io_in_3_bits_reverse      (requestVecFromSlot_3_adder_bits_reverse),
    .io_in_3_bits_average      (requestVecFromSlot_3_adder_bits_average),
    .io_in_3_bits_saturate     (requestVecFromSlot_3_adder_bits_saturate),
    .io_in_3_bits_vxrm         (requestVecFromSlot_3_adder_bits_vxrm),
    .io_in_3_bits_vSew         (requestVecFromSlot_3_adder_bits_vSew),
    .io_in_3_bits_shifterSize  (requestVecFromSlot_3_adder_bits_shifterSize),
    .io_in_3_bits_rem          (requestVecFromSlot_3_adder_bits_rem),
    .io_in_3_bits_groupIndex   (requestVecFromSlot_3_adder_bits_groupIndex),
    .io_in_3_bits_laneIndex    (requestVecFromSlot_3_adder_bits_laneIndex),
    .io_in_3_bits_maskType     (requestVecFromSlot_3_adder_bits_maskType),
    .io_in_3_bits_narrow       (requestVecFromSlot_3_adder_bits_narrow),
    .io_out_ready              (1'h1),
    .io_out_valid              (_vfuResponse_adderArbiter_io_out_valid),
    .io_out_bits_src_0         (_vfuResponse_adderArbiter_io_out_bits_src_0),
    .io_out_bits_src_1         (_vfuResponse_adderArbiter_io_out_bits_src_1),
    .io_out_bits_src_2         (/* unused */),
    .io_out_bits_src_3         (/* unused */),
    .io_out_bits_opcode        (_vfuResponse_adderArbiter_io_out_bits_opcode),
    .io_out_bits_mask          (_vfuResponse_adderArbiter_io_out_bits_mask),
    .io_out_bits_executeMask   (/* unused */),
    .io_out_bits_sign0         (/* unused */),
    .io_out_bits_sign          (_vfuResponse_adderArbiter_io_out_bits_sign),
    .io_out_bits_reverse       (_vfuResponse_adderArbiter_io_out_bits_reverse),
    .io_out_bits_average       (_vfuResponse_adderArbiter_io_out_bits_average),
    .io_out_bits_saturate      (_vfuResponse_adderArbiter_io_out_bits_saturate),
    .io_out_bits_vxrm          (_vfuResponse_adderArbiter_io_out_bits_vxrm),
    .io_out_bits_vSew          (_vfuResponse_adderArbiter_io_out_bits_vSew),
    .io_out_bits_shifterSize   (/* unused */),
    .io_out_bits_rem           (/* unused */),
    .io_out_bits_executeIndex  (_vfuResponse_adderArbiter_io_out_bits_executeIndex),
    .io_out_bits_popInit       (/* unused */),
    .io_out_bits_groupIndex    (/* unused */),
    .io_out_bits_laneIndex     (/* unused */),
    .io_out_bits_maskType      (/* unused */),
    .io_out_bits_narrow        (/* unused */),
    .io_out_bits_tag           (_vfuResponse_adderArbiter_io_out_bits_tag)
  );
  Distributor vfuResponse_shiftDistributor (
    .clock                             (clock),
    .reset                             (reset),
    .requestToVfu_ready                (1'h1),
    .requestToVfu_valid                (_vfuResponse_shiftDistributor_requestToVfu_valid),
    .requestToVfu_bits_src_0           (_vfuResponse_shiftDistributor_requestToVfu_bits_src_0),
    .requestToVfu_bits_src_1           (_vfuResponse_shiftDistributor_requestToVfu_bits_src_1),
    .requestToVfu_bits_src_2           (/* unused */),
    .requestToVfu_bits_src_3           (/* unused */),
    .requestToVfu_bits_opcode          (_vfuResponse_shiftDistributor_requestToVfu_bits_opcode),
    .requestToVfu_bits_mask            (/* unused */),
    .requestToVfu_bits_sign            (/* unused */),
    .requestToVfu_bits_vxrm            (_vfuResponse_shiftDistributor_requestToVfu_bits_vxrm),
    .requestToVfu_bits_vSew            (/* unused */),
    .requestToVfu_bits_shifterSize     (_vfuResponse_shiftDistributor_requestToVfu_bits_shifterSize),
    .requestToVfu_bits_executeIndex    (/* unused */),
    .requestToVfu_bits_popInit         (/* unused */),
    .requestToVfu_bits_groupIndex      (/* unused */),
    .requestToVfu_bits_laneIndex       (/* unused */),
    .requestToVfu_bits_maskType        (/* unused */),
    .requestToVfu_bits_narrow          (/* unused */),
    .requestToVfu_bits_tag             (_vfuResponse_shiftDistributor_requestToVfu_bits_tag),
    .responseFromVfu_valid             (vfuResponse_responseBundle_valid),
    .responseFromVfu_bits_data         (vfuResponse_responseBundle_bits_data),
    .responseFromVfu_bits_clipFail     (1'h0),
    .responseFromVfu_bits_ffoSuccess   (1'h0),
    .requestFromSlot_ready             (_vfuResponse_shiftDistributor_requestFromSlot_ready),
    .requestFromSlot_valid             (_vfuResponse_shiftArbiter_io_out_valid),
    .requestFromSlot_bits_src_0        (_vfuResponse_shiftArbiter_io_out_bits_src_0),
    .requestFromSlot_bits_src_1        (_vfuResponse_shiftArbiter_io_out_bits_src_1),
    .requestFromSlot_bits_src_2        (_vfuResponse_shiftArbiter_io_out_bits_src_2),
    .requestFromSlot_bits_src_3        (_vfuResponse_shiftArbiter_io_out_bits_src_3),
    .requestFromSlot_bits_opcode       (_vfuResponse_shiftArbiter_io_out_bits_opcode),
    .requestFromSlot_bits_mask         (_vfuResponse_shiftArbiter_io_out_bits_mask),
    .requestFromSlot_bits_executeMask  (_vfuResponse_shiftArbiter_io_out_bits_executeMask),
    .requestFromSlot_bits_sign0        (_vfuResponse_shiftArbiter_io_out_bits_sign0),
    .requestFromSlot_bits_sign         (_vfuResponse_shiftArbiter_io_out_bits_sign),
    .requestFromSlot_bits_reverse      (_vfuResponse_shiftArbiter_io_out_bits_reverse),
    .requestFromSlot_bits_average      (_vfuResponse_shiftArbiter_io_out_bits_average),
    .requestFromSlot_bits_saturate     (_vfuResponse_shiftArbiter_io_out_bits_saturate),
    .requestFromSlot_bits_vxrm         (_vfuResponse_shiftArbiter_io_out_bits_vxrm),
    .requestFromSlot_bits_vSew         (_vfuResponse_shiftArbiter_io_out_bits_vSew),
    .requestFromSlot_bits_shifterSize  (_vfuResponse_shiftArbiter_io_out_bits_shifterSize),
    .requestFromSlot_bits_rem          (_vfuResponse_shiftArbiter_io_out_bits_rem),
    .requestFromSlot_bits_executeIndex (_vfuResponse_shiftArbiter_io_out_bits_executeIndex),
    .requestFromSlot_bits_popInit      (_vfuResponse_shiftArbiter_io_out_bits_popInit),
    .requestFromSlot_bits_groupIndex   (_vfuResponse_shiftArbiter_io_out_bits_groupIndex),
    .requestFromSlot_bits_laneIndex    (_vfuResponse_shiftArbiter_io_out_bits_laneIndex),
    .requestFromSlot_bits_maskType     (_vfuResponse_shiftArbiter_io_out_bits_maskType),
    .requestFromSlot_bits_narrow       (_vfuResponse_shiftArbiter_io_out_bits_narrow),
    .requestFromSlot_bits_tag          (_vfuResponse_shiftArbiter_io_out_bits_tag),
    .responseToSlot_valid              (_vfuResponse_shiftDistributor_responseToSlot_valid),
    .responseToSlot_bits_data          (_vfuResponse_shiftDistributor_responseToSlot_bits_data),
    .responseToSlot_bits_ffoSuccess    (_vfuResponse_shiftDistributor_responseToSlot_bits_ffoSuccess),
    .responseToSlot_bits_vxsat         (_vfuResponse_shiftDistributor_responseToSlot_bits_vxsat),
    .responseToSlot_bits_tag           (_vfuResponse_shiftDistributor_responseToSlot_bits_tag)
  );
  Arbiter4_SlotRequestToVFU vfuResponse_shiftArbiter (
    .io_in_0_ready             (requestVecFromSlot_0_shift_ready),
    .io_in_0_valid             (requestVecFromSlot_0_shift_valid),
    .io_in_0_bits_src_0        (requestVecFromSlot_0_shift_bits_src_0),
    .io_in_0_bits_src_1        (requestVecFromSlot_0_shift_bits_src_1),
    .io_in_0_bits_src_2        (requestVecFromSlot_0_shift_bits_src_2),
    .io_in_0_bits_src_3        (requestVecFromSlot_0_shift_bits_src_3),
    .io_in_0_bits_opcode       (requestVecFromSlot_0_shift_bits_opcode),
    .io_in_0_bits_mask         (requestVecFromSlot_0_shift_bits_mask),
    .io_in_0_bits_executeMask  (requestVecFromSlot_0_shift_bits_executeMask),
    .io_in_0_bits_sign0        (requestVecFromSlot_0_shift_bits_sign0),
    .io_in_0_bits_sign         (requestVecFromSlot_0_shift_bits_sign),
    .io_in_0_bits_reverse      (requestVecFromSlot_0_shift_bits_reverse),
    .io_in_0_bits_average      (requestVecFromSlot_0_shift_bits_average),
    .io_in_0_bits_saturate     (requestVecFromSlot_0_shift_bits_saturate),
    .io_in_0_bits_vxrm         (requestVecFromSlot_0_shift_bits_vxrm),
    .io_in_0_bits_vSew         (requestVecFromSlot_0_shift_bits_vSew),
    .io_in_0_bits_shifterSize  (requestVecFromSlot_0_shift_bits_shifterSize),
    .io_in_0_bits_rem          (requestVecFromSlot_0_shift_bits_rem),
    .io_in_0_bits_executeIndex (requestVecFromSlot_0_shift_bits_executeIndex),
    .io_in_0_bits_popInit      (requestVecFromSlot_0_shift_bits_popInit),
    .io_in_0_bits_groupIndex   (requestVecFromSlot_0_shift_bits_groupIndex),
    .io_in_0_bits_laneIndex    (requestVecFromSlot_0_shift_bits_laneIndex),
    .io_in_0_bits_maskType     (requestVecFromSlot_0_shift_bits_maskType),
    .io_in_0_bits_narrow       (requestVecFromSlot_0_shift_bits_narrow),
    .io_in_1_ready             (requestVecFromSlot_1_shift_ready),
    .io_in_1_valid             (requestVecFromSlot_1_shift_valid),
    .io_in_1_bits_src_0        (requestVecFromSlot_1_shift_bits_src_0),
    .io_in_1_bits_src_1        (requestVecFromSlot_1_shift_bits_src_1),
    .io_in_1_bits_src_2        (requestVecFromSlot_1_shift_bits_src_2),
    .io_in_1_bits_src_3        (requestVecFromSlot_1_shift_bits_src_3),
    .io_in_1_bits_opcode       (requestVecFromSlot_1_shift_bits_opcode),
    .io_in_1_bits_mask         (requestVecFromSlot_1_shift_bits_mask),
    .io_in_1_bits_executeMask  (requestVecFromSlot_1_shift_bits_executeMask),
    .io_in_1_bits_sign0        (requestVecFromSlot_1_shift_bits_sign0),
    .io_in_1_bits_sign         (requestVecFromSlot_1_shift_bits_sign),
    .io_in_1_bits_reverse      (requestVecFromSlot_1_shift_bits_reverse),
    .io_in_1_bits_average      (requestVecFromSlot_1_shift_bits_average),
    .io_in_1_bits_saturate     (requestVecFromSlot_1_shift_bits_saturate),
    .io_in_1_bits_vxrm         (requestVecFromSlot_1_shift_bits_vxrm),
    .io_in_1_bits_vSew         (requestVecFromSlot_1_shift_bits_vSew),
    .io_in_1_bits_shifterSize  (requestVecFromSlot_1_shift_bits_shifterSize),
    .io_in_1_bits_rem          (requestVecFromSlot_1_shift_bits_rem),
    .io_in_1_bits_groupIndex   (requestVecFromSlot_1_shift_bits_groupIndex),
    .io_in_1_bits_laneIndex    (requestVecFromSlot_1_shift_bits_laneIndex),
    .io_in_1_bits_maskType     (requestVecFromSlot_1_shift_bits_maskType),
    .io_in_1_bits_narrow       (requestVecFromSlot_1_shift_bits_narrow),
    .io_in_2_ready             (requestVecFromSlot_2_shift_ready),
    .io_in_2_valid             (requestVecFromSlot_2_shift_valid),
    .io_in_2_bits_src_0        (requestVecFromSlot_2_shift_bits_src_0),
    .io_in_2_bits_src_1        (requestVecFromSlot_2_shift_bits_src_1),
    .io_in_2_bits_src_2        (requestVecFromSlot_2_shift_bits_src_2),
    .io_in_2_bits_src_3        (requestVecFromSlot_2_shift_bits_src_3),
    .io_in_2_bits_opcode       (requestVecFromSlot_2_shift_bits_opcode),
    .io_in_2_bits_mask         (requestVecFromSlot_2_shift_bits_mask),
    .io_in_2_bits_executeMask  (requestVecFromSlot_2_shift_bits_executeMask),
    .io_in_2_bits_sign0        (requestVecFromSlot_2_shift_bits_sign0),
    .io_in_2_bits_sign         (requestVecFromSlot_2_shift_bits_sign),
    .io_in_2_bits_reverse      (requestVecFromSlot_2_shift_bits_reverse),
    .io_in_2_bits_average      (requestVecFromSlot_2_shift_bits_average),
    .io_in_2_bits_saturate     (requestVecFromSlot_2_shift_bits_saturate),
    .io_in_2_bits_vxrm         (requestVecFromSlot_2_shift_bits_vxrm),
    .io_in_2_bits_vSew         (requestVecFromSlot_2_shift_bits_vSew),
    .io_in_2_bits_shifterSize  (requestVecFromSlot_2_shift_bits_shifterSize),
    .io_in_2_bits_rem          (requestVecFromSlot_2_shift_bits_rem),
    .io_in_2_bits_groupIndex   (requestVecFromSlot_2_shift_bits_groupIndex),
    .io_in_2_bits_laneIndex    (requestVecFromSlot_2_shift_bits_laneIndex),
    .io_in_2_bits_maskType     (requestVecFromSlot_2_shift_bits_maskType),
    .io_in_2_bits_narrow       (requestVecFromSlot_2_shift_bits_narrow),
    .io_in_3_ready             (requestVecFromSlot_3_shift_ready),
    .io_in_3_valid             (requestVecFromSlot_3_shift_valid),
    .io_in_3_bits_src_0        (requestVecFromSlot_3_shift_bits_src_0),
    .io_in_3_bits_src_1        (requestVecFromSlot_3_shift_bits_src_1),
    .io_in_3_bits_src_2        (requestVecFromSlot_3_shift_bits_src_2),
    .io_in_3_bits_src_3        (requestVecFromSlot_3_shift_bits_src_3),
    .io_in_3_bits_opcode       (requestVecFromSlot_3_shift_bits_opcode),
    .io_in_3_bits_mask         (requestVecFromSlot_3_shift_bits_mask),
    .io_in_3_bits_executeMask  (requestVecFromSlot_3_shift_bits_executeMask),
    .io_in_3_bits_sign0        (requestVecFromSlot_3_shift_bits_sign0),
    .io_in_3_bits_sign         (requestVecFromSlot_3_shift_bits_sign),
    .io_in_3_bits_reverse      (requestVecFromSlot_3_shift_bits_reverse),
    .io_in_3_bits_average      (requestVecFromSlot_3_shift_bits_average),
    .io_in_3_bits_saturate     (requestVecFromSlot_3_shift_bits_saturate),
    .io_in_3_bits_vxrm         (requestVecFromSlot_3_shift_bits_vxrm),
    .io_in_3_bits_vSew         (requestVecFromSlot_3_shift_bits_vSew),
    .io_in_3_bits_shifterSize  (requestVecFromSlot_3_shift_bits_shifterSize),
    .io_in_3_bits_rem          (requestVecFromSlot_3_shift_bits_rem),
    .io_in_3_bits_groupIndex   (requestVecFromSlot_3_shift_bits_groupIndex),
    .io_in_3_bits_laneIndex    (requestVecFromSlot_3_shift_bits_laneIndex),
    .io_in_3_bits_maskType     (requestVecFromSlot_3_shift_bits_maskType),
    .io_in_3_bits_narrow       (requestVecFromSlot_3_shift_bits_narrow),
    .io_out_ready              (_vfuResponse_shiftDistributor_requestFromSlot_ready),
    .io_out_valid              (_vfuResponse_shiftArbiter_io_out_valid),
    .io_out_bits_src_0         (_vfuResponse_shiftArbiter_io_out_bits_src_0),
    .io_out_bits_src_1         (_vfuResponse_shiftArbiter_io_out_bits_src_1),
    .io_out_bits_src_2         (_vfuResponse_shiftArbiter_io_out_bits_src_2),
    .io_out_bits_src_3         (_vfuResponse_shiftArbiter_io_out_bits_src_3),
    .io_out_bits_opcode        (_vfuResponse_shiftArbiter_io_out_bits_opcode),
    .io_out_bits_mask          (_vfuResponse_shiftArbiter_io_out_bits_mask),
    .io_out_bits_executeMask   (_vfuResponse_shiftArbiter_io_out_bits_executeMask),
    .io_out_bits_sign0         (_vfuResponse_shiftArbiter_io_out_bits_sign0),
    .io_out_bits_sign          (_vfuResponse_shiftArbiter_io_out_bits_sign),
    .io_out_bits_reverse       (_vfuResponse_shiftArbiter_io_out_bits_reverse),
    .io_out_bits_average       (_vfuResponse_shiftArbiter_io_out_bits_average),
    .io_out_bits_saturate      (_vfuResponse_shiftArbiter_io_out_bits_saturate),
    .io_out_bits_vxrm          (_vfuResponse_shiftArbiter_io_out_bits_vxrm),
    .io_out_bits_vSew          (_vfuResponse_shiftArbiter_io_out_bits_vSew),
    .io_out_bits_shifterSize   (_vfuResponse_shiftArbiter_io_out_bits_shifterSize),
    .io_out_bits_rem           (_vfuResponse_shiftArbiter_io_out_bits_rem),
    .io_out_bits_executeIndex  (_vfuResponse_shiftArbiter_io_out_bits_executeIndex),
    .io_out_bits_popInit       (_vfuResponse_shiftArbiter_io_out_bits_popInit),
    .io_out_bits_groupIndex    (_vfuResponse_shiftArbiter_io_out_bits_groupIndex),
    .io_out_bits_laneIndex     (_vfuResponse_shiftArbiter_io_out_bits_laneIndex),
    .io_out_bits_maskType      (_vfuResponse_shiftArbiter_io_out_bits_maskType),
    .io_out_bits_narrow        (_vfuResponse_shiftArbiter_io_out_bits_narrow),
    .io_out_bits_tag           (_vfuResponse_shiftArbiter_io_out_bits_tag)
  );
  Arbiter4_SlotRequestToVFU vfuResponse_multiplierArbiter (
    .io_in_0_ready             (requestVecFromSlot_0_multiplier_ready),
    .io_in_0_valid             (requestVecFromSlot_0_multiplier_valid),
    .io_in_0_bits_src_0        (requestVecFromSlot_0_multiplier_bits_src_0),
    .io_in_0_bits_src_1        (requestVecFromSlot_0_multiplier_bits_src_1),
    .io_in_0_bits_src_2        (requestVecFromSlot_0_multiplier_bits_src_2),
    .io_in_0_bits_src_3        (requestVecFromSlot_0_multiplier_bits_src_3),
    .io_in_0_bits_opcode       (requestVecFromSlot_0_multiplier_bits_opcode),
    .io_in_0_bits_mask         (requestVecFromSlot_0_multiplier_bits_mask),
    .io_in_0_bits_executeMask  (requestVecFromSlot_0_multiplier_bits_executeMask),
    .io_in_0_bits_sign0        (requestVecFromSlot_0_multiplier_bits_sign0),
    .io_in_0_bits_sign         (requestVecFromSlot_0_multiplier_bits_sign),
    .io_in_0_bits_reverse      (requestVecFromSlot_0_multiplier_bits_reverse),
    .io_in_0_bits_average      (requestVecFromSlot_0_multiplier_bits_average),
    .io_in_0_bits_saturate     (requestVecFromSlot_0_multiplier_bits_saturate),
    .io_in_0_bits_vxrm         (requestVecFromSlot_0_multiplier_bits_vxrm),
    .io_in_0_bits_vSew         (requestVecFromSlot_0_multiplier_bits_vSew),
    .io_in_0_bits_shifterSize  (requestVecFromSlot_0_multiplier_bits_shifterSize),
    .io_in_0_bits_rem          (requestVecFromSlot_0_multiplier_bits_rem),
    .io_in_0_bits_executeIndex (requestVecFromSlot_0_multiplier_bits_executeIndex),
    .io_in_0_bits_popInit      (requestVecFromSlot_0_multiplier_bits_popInit),
    .io_in_0_bits_groupIndex   (requestVecFromSlot_0_multiplier_bits_groupIndex),
    .io_in_0_bits_laneIndex    (requestVecFromSlot_0_multiplier_bits_laneIndex),
    .io_in_0_bits_maskType     (requestVecFromSlot_0_multiplier_bits_maskType),
    .io_in_0_bits_narrow       (requestVecFromSlot_0_multiplier_bits_narrow),
    .io_in_1_ready             (requestVecFromSlot_1_multiplier_ready),
    .io_in_1_valid             (requestVecFromSlot_1_multiplier_valid),
    .io_in_1_bits_src_0        (requestVecFromSlot_1_multiplier_bits_src_0),
    .io_in_1_bits_src_1        (requestVecFromSlot_1_multiplier_bits_src_1),
    .io_in_1_bits_src_2        (requestVecFromSlot_1_multiplier_bits_src_2),
    .io_in_1_bits_src_3        (requestVecFromSlot_1_multiplier_bits_src_3),
    .io_in_1_bits_opcode       (requestVecFromSlot_1_multiplier_bits_opcode),
    .io_in_1_bits_mask         (requestVecFromSlot_1_multiplier_bits_mask),
    .io_in_1_bits_executeMask  (requestVecFromSlot_1_multiplier_bits_executeMask),
    .io_in_1_bits_sign0        (requestVecFromSlot_1_multiplier_bits_sign0),
    .io_in_1_bits_sign         (requestVecFromSlot_1_multiplier_bits_sign),
    .io_in_1_bits_reverse      (requestVecFromSlot_1_multiplier_bits_reverse),
    .io_in_1_bits_average      (requestVecFromSlot_1_multiplier_bits_average),
    .io_in_1_bits_saturate     (requestVecFromSlot_1_multiplier_bits_saturate),
    .io_in_1_bits_vxrm         (requestVecFromSlot_1_multiplier_bits_vxrm),
    .io_in_1_bits_vSew         (requestVecFromSlot_1_multiplier_bits_vSew),
    .io_in_1_bits_shifterSize  (requestVecFromSlot_1_multiplier_bits_shifterSize),
    .io_in_1_bits_rem          (requestVecFromSlot_1_multiplier_bits_rem),
    .io_in_1_bits_groupIndex   (requestVecFromSlot_1_multiplier_bits_groupIndex),
    .io_in_1_bits_laneIndex    (requestVecFromSlot_1_multiplier_bits_laneIndex),
    .io_in_1_bits_maskType     (requestVecFromSlot_1_multiplier_bits_maskType),
    .io_in_1_bits_narrow       (requestVecFromSlot_1_multiplier_bits_narrow),
    .io_in_2_ready             (requestVecFromSlot_2_multiplier_ready),
    .io_in_2_valid             (requestVecFromSlot_2_multiplier_valid),
    .io_in_2_bits_src_0        (requestVecFromSlot_2_multiplier_bits_src_0),
    .io_in_2_bits_src_1        (requestVecFromSlot_2_multiplier_bits_src_1),
    .io_in_2_bits_src_2        (requestVecFromSlot_2_multiplier_bits_src_2),
    .io_in_2_bits_src_3        (requestVecFromSlot_2_multiplier_bits_src_3),
    .io_in_2_bits_opcode       (requestVecFromSlot_2_multiplier_bits_opcode),
    .io_in_2_bits_mask         (requestVecFromSlot_2_multiplier_bits_mask),
    .io_in_2_bits_executeMask  (requestVecFromSlot_2_multiplier_bits_executeMask),
    .io_in_2_bits_sign0        (requestVecFromSlot_2_multiplier_bits_sign0),
    .io_in_2_bits_sign         (requestVecFromSlot_2_multiplier_bits_sign),
    .io_in_2_bits_reverse      (requestVecFromSlot_2_multiplier_bits_reverse),
    .io_in_2_bits_average      (requestVecFromSlot_2_multiplier_bits_average),
    .io_in_2_bits_saturate     (requestVecFromSlot_2_multiplier_bits_saturate),
    .io_in_2_bits_vxrm         (requestVecFromSlot_2_multiplier_bits_vxrm),
    .io_in_2_bits_vSew         (requestVecFromSlot_2_multiplier_bits_vSew),
    .io_in_2_bits_shifterSize  (requestVecFromSlot_2_multiplier_bits_shifterSize),
    .io_in_2_bits_rem          (requestVecFromSlot_2_multiplier_bits_rem),
    .io_in_2_bits_groupIndex   (requestVecFromSlot_2_multiplier_bits_groupIndex),
    .io_in_2_bits_laneIndex    (requestVecFromSlot_2_multiplier_bits_laneIndex),
    .io_in_2_bits_maskType     (requestVecFromSlot_2_multiplier_bits_maskType),
    .io_in_2_bits_narrow       (requestVecFromSlot_2_multiplier_bits_narrow),
    .io_in_3_ready             (requestVecFromSlot_3_multiplier_ready),
    .io_in_3_valid             (requestVecFromSlot_3_multiplier_valid),
    .io_in_3_bits_src_0        (requestVecFromSlot_3_multiplier_bits_src_0),
    .io_in_3_bits_src_1        (requestVecFromSlot_3_multiplier_bits_src_1),
    .io_in_3_bits_src_2        (requestVecFromSlot_3_multiplier_bits_src_2),
    .io_in_3_bits_src_3        (requestVecFromSlot_3_multiplier_bits_src_3),
    .io_in_3_bits_opcode       (requestVecFromSlot_3_multiplier_bits_opcode),
    .io_in_3_bits_mask         (requestVecFromSlot_3_multiplier_bits_mask),
    .io_in_3_bits_executeMask  (requestVecFromSlot_3_multiplier_bits_executeMask),
    .io_in_3_bits_sign0        (requestVecFromSlot_3_multiplier_bits_sign0),
    .io_in_3_bits_sign         (requestVecFromSlot_3_multiplier_bits_sign),
    .io_in_3_bits_reverse      (requestVecFromSlot_3_multiplier_bits_reverse),
    .io_in_3_bits_average      (requestVecFromSlot_3_multiplier_bits_average),
    .io_in_3_bits_saturate     (requestVecFromSlot_3_multiplier_bits_saturate),
    .io_in_3_bits_vxrm         (requestVecFromSlot_3_multiplier_bits_vxrm),
    .io_in_3_bits_vSew         (requestVecFromSlot_3_multiplier_bits_vSew),
    .io_in_3_bits_shifterSize  (requestVecFromSlot_3_multiplier_bits_shifterSize),
    .io_in_3_bits_rem          (requestVecFromSlot_3_multiplier_bits_rem),
    .io_in_3_bits_groupIndex   (requestVecFromSlot_3_multiplier_bits_groupIndex),
    .io_in_3_bits_laneIndex    (requestVecFromSlot_3_multiplier_bits_laneIndex),
    .io_in_3_bits_maskType     (requestVecFromSlot_3_multiplier_bits_maskType),
    .io_in_3_bits_narrow       (requestVecFromSlot_3_multiplier_bits_narrow),
    .io_out_ready              (1'h1),
    .io_out_valid              (_vfuResponse_multiplierArbiter_io_out_valid),
    .io_out_bits_src_0         (_vfuResponse_multiplierArbiter_io_out_bits_src_0),
    .io_out_bits_src_1         (_vfuResponse_multiplierArbiter_io_out_bits_src_1),
    .io_out_bits_src_2         (_vfuResponse_multiplierArbiter_io_out_bits_src_2),
    .io_out_bits_src_3         (/* unused */),
    .io_out_bits_opcode        (_vfuResponse_multiplierArbiter_io_out_bits_opcode),
    .io_out_bits_mask          (/* unused */),
    .io_out_bits_executeMask   (/* unused */),
    .io_out_bits_sign0         (_vfuResponse_multiplierArbiter_io_out_bits_sign0),
    .io_out_bits_sign          (_vfuResponse_multiplierArbiter_io_out_bits_sign),
    .io_out_bits_reverse       (/* unused */),
    .io_out_bits_average       (/* unused */),
    .io_out_bits_saturate      (_vfuResponse_multiplierArbiter_io_out_bits_saturate),
    .io_out_bits_vxrm          (_vfuResponse_multiplierArbiter_io_out_bits_vxrm),
    .io_out_bits_vSew          (_vfuResponse_multiplierArbiter_io_out_bits_vSew),
    .io_out_bits_shifterSize   (/* unused */),
    .io_out_bits_rem           (/* unused */),
    .io_out_bits_executeIndex  (/* unused */),
    .io_out_bits_popInit       (/* unused */),
    .io_out_bits_groupIndex    (/* unused */),
    .io_out_bits_laneIndex     (/* unused */),
    .io_out_bits_maskType      (/* unused */),
    .io_out_bits_narrow        (/* unused */),
    .io_out_bits_tag           (_vfuResponse_multiplierArbiter_io_out_bits_tag)
  );
  Distributor vfuResponse_dividerDistributor (
    .clock                             (clock),
    .reset                             (reset),
    .requestToVfu_ready                (_divider_requestIO_ready),
    .requestToVfu_valid                (_vfuResponse_dividerDistributor_requestToVfu_valid),
    .requestToVfu_bits_src_0           (_vfuResponse_dividerDistributor_requestToVfu_bits_src_0),
    .requestToVfu_bits_src_1           (_vfuResponse_dividerDistributor_requestToVfu_bits_src_1),
    .requestToVfu_bits_src_2           (/* unused */),
    .requestToVfu_bits_src_3           (/* unused */),
    .requestToVfu_bits_opcode          (_vfuResponse_dividerDistributor_requestToVfu_bits_opcode),
    .requestToVfu_bits_mask            (/* unused */),
    .requestToVfu_bits_sign            (_vfuResponse_dividerDistributor_requestToVfu_bits_sign),
    .requestToVfu_bits_vxrm            (/* unused */),
    .requestToVfu_bits_vSew            (/* unused */),
    .requestToVfu_bits_shifterSize     (/* unused */),
    .requestToVfu_bits_executeIndex    (_vfuResponse_dividerDistributor_requestToVfu_bits_executeIndex),
    .requestToVfu_bits_popInit         (/* unused */),
    .requestToVfu_bits_groupIndex      (/* unused */),
    .requestToVfu_bits_laneIndex       (/* unused */),
    .requestToVfu_bits_maskType        (/* unused */),
    .requestToVfu_bits_narrow          (/* unused */),
    .requestToVfu_bits_tag             (_vfuResponse_dividerDistributor_requestToVfu_bits_tag),
    .responseFromVfu_valid             (vfuResponse_responseBundle_1_valid),
    .responseFromVfu_bits_data         (vfuResponse_responseBundle_1_bits_data),
    .responseFromVfu_bits_clipFail     (1'h0),
    .responseFromVfu_bits_ffoSuccess   (1'h0),
    .requestFromSlot_ready             (_vfuResponse_dividerDistributor_requestFromSlot_ready),
    .requestFromSlot_valid             (_vfuResponse_dividerArbiter_io_out_valid),
    .requestFromSlot_bits_src_0        (_vfuResponse_dividerArbiter_io_out_bits_src_0),
    .requestFromSlot_bits_src_1        (_vfuResponse_dividerArbiter_io_out_bits_src_1),
    .requestFromSlot_bits_src_2        (_vfuResponse_dividerArbiter_io_out_bits_src_2),
    .requestFromSlot_bits_src_3        (_vfuResponse_dividerArbiter_io_out_bits_src_3),
    .requestFromSlot_bits_opcode       (_vfuResponse_dividerArbiter_io_out_bits_opcode),
    .requestFromSlot_bits_mask         (_vfuResponse_dividerArbiter_io_out_bits_mask),
    .requestFromSlot_bits_executeMask  (_vfuResponse_dividerArbiter_io_out_bits_executeMask),
    .requestFromSlot_bits_sign0        (_vfuResponse_dividerArbiter_io_out_bits_sign0),
    .requestFromSlot_bits_sign         (_vfuResponse_dividerArbiter_io_out_bits_sign),
    .requestFromSlot_bits_reverse      (_vfuResponse_dividerArbiter_io_out_bits_reverse),
    .requestFromSlot_bits_average      (_vfuResponse_dividerArbiter_io_out_bits_average),
    .requestFromSlot_bits_saturate     (_vfuResponse_dividerArbiter_io_out_bits_saturate),
    .requestFromSlot_bits_vxrm         (_vfuResponse_dividerArbiter_io_out_bits_vxrm),
    .requestFromSlot_bits_vSew         (_vfuResponse_dividerArbiter_io_out_bits_vSew),
    .requestFromSlot_bits_shifterSize  (_vfuResponse_dividerArbiter_io_out_bits_shifterSize),
    .requestFromSlot_bits_rem          (_vfuResponse_dividerArbiter_io_out_bits_rem),
    .requestFromSlot_bits_executeIndex (_vfuResponse_dividerArbiter_io_out_bits_executeIndex),
    .requestFromSlot_bits_popInit      (_vfuResponse_dividerArbiter_io_out_bits_popInit),
    .requestFromSlot_bits_groupIndex   (_vfuResponse_dividerArbiter_io_out_bits_groupIndex),
    .requestFromSlot_bits_laneIndex    (_vfuResponse_dividerArbiter_io_out_bits_laneIndex),
    .requestFromSlot_bits_maskType     (_vfuResponse_dividerArbiter_io_out_bits_maskType),
    .requestFromSlot_bits_narrow       (_vfuResponse_dividerArbiter_io_out_bits_narrow),
    .requestFromSlot_bits_tag          (_vfuResponse_dividerArbiter_io_out_bits_tag),
    .responseToSlot_valid              (_vfuResponse_dividerDistributor_responseToSlot_valid),
    .responseToSlot_bits_data          (_vfuResponse_dividerDistributor_responseToSlot_bits_data),
    .responseToSlot_bits_ffoSuccess    (_vfuResponse_dividerDistributor_responseToSlot_bits_ffoSuccess),
    .responseToSlot_bits_vxsat         (_vfuResponse_dividerDistributor_responseToSlot_bits_vxsat),
    .responseToSlot_bits_tag           (_vfuResponse_dividerDistributor_responseToSlot_bits_tag)
  );
  Arbiter4_SlotRequestToVFU vfuResponse_dividerArbiter (
    .io_in_0_ready             (requestVecFromSlot_0_divider_ready),
    .io_in_0_valid             (requestVecFromSlot_0_divider_valid),
    .io_in_0_bits_src_0        (requestVecFromSlot_0_divider_bits_src_0),
    .io_in_0_bits_src_1        (requestVecFromSlot_0_divider_bits_src_1),
    .io_in_0_bits_src_2        (requestVecFromSlot_0_divider_bits_src_2),
    .io_in_0_bits_src_3        (requestVecFromSlot_0_divider_bits_src_3),
    .io_in_0_bits_opcode       (requestVecFromSlot_0_divider_bits_opcode),
    .io_in_0_bits_mask         (requestVecFromSlot_0_divider_bits_mask),
    .io_in_0_bits_executeMask  (requestVecFromSlot_0_divider_bits_executeMask),
    .io_in_0_bits_sign0        (requestVecFromSlot_0_divider_bits_sign0),
    .io_in_0_bits_sign         (requestVecFromSlot_0_divider_bits_sign),
    .io_in_0_bits_reverse      (requestVecFromSlot_0_divider_bits_reverse),
    .io_in_0_bits_average      (requestVecFromSlot_0_divider_bits_average),
    .io_in_0_bits_saturate     (requestVecFromSlot_0_divider_bits_saturate),
    .io_in_0_bits_vxrm         (requestVecFromSlot_0_divider_bits_vxrm),
    .io_in_0_bits_vSew         (requestVecFromSlot_0_divider_bits_vSew),
    .io_in_0_bits_shifterSize  (requestVecFromSlot_0_divider_bits_shifterSize),
    .io_in_0_bits_rem          (requestVecFromSlot_0_divider_bits_rem),
    .io_in_0_bits_executeIndex (requestVecFromSlot_0_divider_bits_executeIndex),
    .io_in_0_bits_popInit      (requestVecFromSlot_0_divider_bits_popInit),
    .io_in_0_bits_groupIndex   (requestVecFromSlot_0_divider_bits_groupIndex),
    .io_in_0_bits_laneIndex    (requestVecFromSlot_0_divider_bits_laneIndex),
    .io_in_0_bits_maskType     (requestVecFromSlot_0_divider_bits_maskType),
    .io_in_0_bits_narrow       (requestVecFromSlot_0_divider_bits_narrow),
    .io_in_1_ready             (requestVecFromSlot_1_divider_ready),
    .io_in_1_valid             (requestVecFromSlot_1_divider_valid),
    .io_in_1_bits_src_0        (requestVecFromSlot_1_divider_bits_src_0),
    .io_in_1_bits_src_1        (requestVecFromSlot_1_divider_bits_src_1),
    .io_in_1_bits_src_2        (requestVecFromSlot_1_divider_bits_src_2),
    .io_in_1_bits_src_3        (requestVecFromSlot_1_divider_bits_src_3),
    .io_in_1_bits_opcode       (requestVecFromSlot_1_divider_bits_opcode),
    .io_in_1_bits_mask         (requestVecFromSlot_1_divider_bits_mask),
    .io_in_1_bits_executeMask  (requestVecFromSlot_1_divider_bits_executeMask),
    .io_in_1_bits_sign0        (requestVecFromSlot_1_divider_bits_sign0),
    .io_in_1_bits_sign         (requestVecFromSlot_1_divider_bits_sign),
    .io_in_1_bits_reverse      (requestVecFromSlot_1_divider_bits_reverse),
    .io_in_1_bits_average      (requestVecFromSlot_1_divider_bits_average),
    .io_in_1_bits_saturate     (requestVecFromSlot_1_divider_bits_saturate),
    .io_in_1_bits_vxrm         (requestVecFromSlot_1_divider_bits_vxrm),
    .io_in_1_bits_vSew         (requestVecFromSlot_1_divider_bits_vSew),
    .io_in_1_bits_shifterSize  (requestVecFromSlot_1_divider_bits_shifterSize),
    .io_in_1_bits_rem          (requestVecFromSlot_1_divider_bits_rem),
    .io_in_1_bits_groupIndex   (requestVecFromSlot_1_divider_bits_groupIndex),
    .io_in_1_bits_laneIndex    (requestVecFromSlot_1_divider_bits_laneIndex),
    .io_in_1_bits_maskType     (requestVecFromSlot_1_divider_bits_maskType),
    .io_in_1_bits_narrow       (requestVecFromSlot_1_divider_bits_narrow),
    .io_in_2_ready             (requestVecFromSlot_2_divider_ready),
    .io_in_2_valid             (requestVecFromSlot_2_divider_valid),
    .io_in_2_bits_src_0        (requestVecFromSlot_2_divider_bits_src_0),
    .io_in_2_bits_src_1        (requestVecFromSlot_2_divider_bits_src_1),
    .io_in_2_bits_src_2        (requestVecFromSlot_2_divider_bits_src_2),
    .io_in_2_bits_src_3        (requestVecFromSlot_2_divider_bits_src_3),
    .io_in_2_bits_opcode       (requestVecFromSlot_2_divider_bits_opcode),
    .io_in_2_bits_mask         (requestVecFromSlot_2_divider_bits_mask),
    .io_in_2_bits_executeMask  (requestVecFromSlot_2_divider_bits_executeMask),
    .io_in_2_bits_sign0        (requestVecFromSlot_2_divider_bits_sign0),
    .io_in_2_bits_sign         (requestVecFromSlot_2_divider_bits_sign),
    .io_in_2_bits_reverse      (requestVecFromSlot_2_divider_bits_reverse),
    .io_in_2_bits_average      (requestVecFromSlot_2_divider_bits_average),
    .io_in_2_bits_saturate     (requestVecFromSlot_2_divider_bits_saturate),
    .io_in_2_bits_vxrm         (requestVecFromSlot_2_divider_bits_vxrm),
    .io_in_2_bits_vSew         (requestVecFromSlot_2_divider_bits_vSew),
    .io_in_2_bits_shifterSize  (requestVecFromSlot_2_divider_bits_shifterSize),
    .io_in_2_bits_rem          (requestVecFromSlot_2_divider_bits_rem),
    .io_in_2_bits_groupIndex   (requestVecFromSlot_2_divider_bits_groupIndex),
    .io_in_2_bits_laneIndex    (requestVecFromSlot_2_divider_bits_laneIndex),
    .io_in_2_bits_maskType     (requestVecFromSlot_2_divider_bits_maskType),
    .io_in_2_bits_narrow       (requestVecFromSlot_2_divider_bits_narrow),
    .io_in_3_ready             (requestVecFromSlot_3_divider_ready),
    .io_in_3_valid             (requestVecFromSlot_3_divider_valid),
    .io_in_3_bits_src_0        (requestVecFromSlot_3_divider_bits_src_0),
    .io_in_3_bits_src_1        (requestVecFromSlot_3_divider_bits_src_1),
    .io_in_3_bits_src_2        (requestVecFromSlot_3_divider_bits_src_2),
    .io_in_3_bits_src_3        (requestVecFromSlot_3_divider_bits_src_3),
    .io_in_3_bits_opcode       (requestVecFromSlot_3_divider_bits_opcode),
    .io_in_3_bits_mask         (requestVecFromSlot_3_divider_bits_mask),
    .io_in_3_bits_executeMask  (requestVecFromSlot_3_divider_bits_executeMask),
    .io_in_3_bits_sign0        (requestVecFromSlot_3_divider_bits_sign0),
    .io_in_3_bits_sign         (requestVecFromSlot_3_divider_bits_sign),
    .io_in_3_bits_reverse      (requestVecFromSlot_3_divider_bits_reverse),
    .io_in_3_bits_average      (requestVecFromSlot_3_divider_bits_average),
    .io_in_3_bits_saturate     (requestVecFromSlot_3_divider_bits_saturate),
    .io_in_3_bits_vxrm         (requestVecFromSlot_3_divider_bits_vxrm),
    .io_in_3_bits_vSew         (requestVecFromSlot_3_divider_bits_vSew),
    .io_in_3_bits_shifterSize  (requestVecFromSlot_3_divider_bits_shifterSize),
    .io_in_3_bits_rem          (requestVecFromSlot_3_divider_bits_rem),
    .io_in_3_bits_groupIndex   (requestVecFromSlot_3_divider_bits_groupIndex),
    .io_in_3_bits_laneIndex    (requestVecFromSlot_3_divider_bits_laneIndex),
    .io_in_3_bits_maskType     (requestVecFromSlot_3_divider_bits_maskType),
    .io_in_3_bits_narrow       (requestVecFromSlot_3_divider_bits_narrow),
    .io_out_ready              (_vfuResponse_dividerDistributor_requestFromSlot_ready),
    .io_out_valid              (_vfuResponse_dividerArbiter_io_out_valid),
    .io_out_bits_src_0         (_vfuResponse_dividerArbiter_io_out_bits_src_0),
    .io_out_bits_src_1         (_vfuResponse_dividerArbiter_io_out_bits_src_1),
    .io_out_bits_src_2         (_vfuResponse_dividerArbiter_io_out_bits_src_2),
    .io_out_bits_src_3         (_vfuResponse_dividerArbiter_io_out_bits_src_3),
    .io_out_bits_opcode        (_vfuResponse_dividerArbiter_io_out_bits_opcode),
    .io_out_bits_mask          (_vfuResponse_dividerArbiter_io_out_bits_mask),
    .io_out_bits_executeMask   (_vfuResponse_dividerArbiter_io_out_bits_executeMask),
    .io_out_bits_sign0         (_vfuResponse_dividerArbiter_io_out_bits_sign0),
    .io_out_bits_sign          (_vfuResponse_dividerArbiter_io_out_bits_sign),
    .io_out_bits_reverse       (_vfuResponse_dividerArbiter_io_out_bits_reverse),
    .io_out_bits_average       (_vfuResponse_dividerArbiter_io_out_bits_average),
    .io_out_bits_saturate      (_vfuResponse_dividerArbiter_io_out_bits_saturate),
    .io_out_bits_vxrm          (_vfuResponse_dividerArbiter_io_out_bits_vxrm),
    .io_out_bits_vSew          (_vfuResponse_dividerArbiter_io_out_bits_vSew),
    .io_out_bits_shifterSize   (_vfuResponse_dividerArbiter_io_out_bits_shifterSize),
    .io_out_bits_rem           (_vfuResponse_dividerArbiter_io_out_bits_rem),
    .io_out_bits_executeIndex  (_vfuResponse_dividerArbiter_io_out_bits_executeIndex),
    .io_out_bits_popInit       (_vfuResponse_dividerArbiter_io_out_bits_popInit),
    .io_out_bits_groupIndex    (_vfuResponse_dividerArbiter_io_out_bits_groupIndex),
    .io_out_bits_laneIndex     (_vfuResponse_dividerArbiter_io_out_bits_laneIndex),
    .io_out_bits_maskType      (_vfuResponse_dividerArbiter_io_out_bits_maskType),
    .io_out_bits_narrow        (_vfuResponse_dividerArbiter_io_out_bits_narrow),
    .io_out_bits_tag           (_vfuResponse_dividerArbiter_io_out_bits_tag)
  );
  Distributor vfuResponse_otherDistributor (
    .clock                             (clock),
    .reset                             (reset),
    .requestToVfu_ready                (1'h1),
    .requestToVfu_valid                (_vfuResponse_otherDistributor_requestToVfu_valid),
    .requestToVfu_bits_src_0           (_vfuResponse_otherDistributor_requestToVfu_bits_src_0),
    .requestToVfu_bits_src_1           (_vfuResponse_otherDistributor_requestToVfu_bits_src_1),
    .requestToVfu_bits_src_2           (_vfuResponse_otherDistributor_requestToVfu_bits_src_2),
    .requestToVfu_bits_src_3           (_vfuResponse_otherDistributor_requestToVfu_bits_src_3),
    .requestToVfu_bits_opcode          (_vfuResponse_otherDistributor_requestToVfu_bits_opcode),
    .requestToVfu_bits_mask            (_vfuResponse_otherDistributor_requestToVfu_bits_mask),
    .requestToVfu_bits_sign            (_vfuResponse_otherDistributor_requestToVfu_bits_sign),
    .requestToVfu_bits_vxrm            (_vfuResponse_otherDistributor_requestToVfu_bits_vxrm),
    .requestToVfu_bits_vSew            (_vfuResponse_otherDistributor_requestToVfu_bits_vSew),
    .requestToVfu_bits_shifterSize     (/* unused */),
    .requestToVfu_bits_executeIndex    (_vfuResponse_otherDistributor_requestToVfu_bits_executeIndex),
    .requestToVfu_bits_popInit         (_vfuResponse_otherDistributor_requestToVfu_bits_popInit),
    .requestToVfu_bits_groupIndex      (_vfuResponse_otherDistributor_requestToVfu_bits_groupIndex),
    .requestToVfu_bits_laneIndex       (_vfuResponse_otherDistributor_requestToVfu_bits_laneIndex),
    .requestToVfu_bits_maskType        (_vfuResponse_otherDistributor_requestToVfu_bits_maskType),
    .requestToVfu_bits_narrow          (_vfuResponse_otherDistributor_requestToVfu_bits_narrow),
    .requestToVfu_bits_tag             (_vfuResponse_otherDistributor_requestToVfu_bits_tag),
    .responseFromVfu_valid             (vfuResponse_responseBundle_2_valid),
    .responseFromVfu_bits_data         (vfuResponse_responseBundle_2_bits_data),
    .responseFromVfu_bits_clipFail     (vfuResponse_responseBundle_2_bits_clipFail),
    .responseFromVfu_bits_ffoSuccess   (vfuResponse_responseBundle_2_bits_ffoSuccess),
    .requestFromSlot_ready             (_vfuResponse_otherDistributor_requestFromSlot_ready),
    .requestFromSlot_valid             (_vfuResponse_otherArbiter_io_out_valid),
    .requestFromSlot_bits_src_0        (_vfuResponse_otherArbiter_io_out_bits_src_0),
    .requestFromSlot_bits_src_1        (_vfuResponse_otherArbiter_io_out_bits_src_1),
    .requestFromSlot_bits_src_2        (_vfuResponse_otherArbiter_io_out_bits_src_2),
    .requestFromSlot_bits_src_3        (_vfuResponse_otherArbiter_io_out_bits_src_3),
    .requestFromSlot_bits_opcode       (_vfuResponse_otherArbiter_io_out_bits_opcode),
    .requestFromSlot_bits_mask         (_vfuResponse_otherArbiter_io_out_bits_mask),
    .requestFromSlot_bits_executeMask  (_vfuResponse_otherArbiter_io_out_bits_executeMask),
    .requestFromSlot_bits_sign0        (_vfuResponse_otherArbiter_io_out_bits_sign0),
    .requestFromSlot_bits_sign         (_vfuResponse_otherArbiter_io_out_bits_sign),
    .requestFromSlot_bits_reverse      (_vfuResponse_otherArbiter_io_out_bits_reverse),
    .requestFromSlot_bits_average      (_vfuResponse_otherArbiter_io_out_bits_average),
    .requestFromSlot_bits_saturate     (_vfuResponse_otherArbiter_io_out_bits_saturate),
    .requestFromSlot_bits_vxrm         (_vfuResponse_otherArbiter_io_out_bits_vxrm),
    .requestFromSlot_bits_vSew         (_vfuResponse_otherArbiter_io_out_bits_vSew),
    .requestFromSlot_bits_shifterSize  (_vfuResponse_otherArbiter_io_out_bits_shifterSize),
    .requestFromSlot_bits_rem          (_vfuResponse_otherArbiter_io_out_bits_rem),
    .requestFromSlot_bits_executeIndex (_vfuResponse_otherArbiter_io_out_bits_executeIndex),
    .requestFromSlot_bits_popInit      (_vfuResponse_otherArbiter_io_out_bits_popInit),
    .requestFromSlot_bits_groupIndex   (_vfuResponse_otherArbiter_io_out_bits_groupIndex),
    .requestFromSlot_bits_laneIndex    (_vfuResponse_otherArbiter_io_out_bits_laneIndex),
    .requestFromSlot_bits_maskType     (_vfuResponse_otherArbiter_io_out_bits_maskType),
    .requestFromSlot_bits_narrow       (_vfuResponse_otherArbiter_io_out_bits_narrow),
    .requestFromSlot_bits_tag          (_vfuResponse_otherArbiter_io_out_bits_tag),
    .responseToSlot_valid              (_vfuResponse_otherDistributor_responseToSlot_valid),
    .responseToSlot_bits_data          (_vfuResponse_otherDistributor_responseToSlot_bits_data),
    .responseToSlot_bits_ffoSuccess    (_vfuResponse_otherDistributor_responseToSlot_bits_ffoSuccess),
    .responseToSlot_bits_vxsat         (_vfuResponse_otherDistributor_responseToSlot_bits_vxsat),
    .responseToSlot_bits_tag           (_vfuResponse_otherDistributor_responseToSlot_bits_tag)
  );
  Arbiter4_SlotRequestToVFU vfuResponse_otherArbiter (
    .io_in_0_ready             (requestVecFromSlot_0_other_ready),
    .io_in_0_valid             (requestVecFromSlot_0_other_valid),
    .io_in_0_bits_src_0        (requestVecFromSlot_0_other_bits_src_0),
    .io_in_0_bits_src_1        (requestVecFromSlot_0_other_bits_src_1),
    .io_in_0_bits_src_2        (requestVecFromSlot_0_other_bits_src_2),
    .io_in_0_bits_src_3        (requestVecFromSlot_0_other_bits_src_3),
    .io_in_0_bits_opcode       (requestVecFromSlot_0_other_bits_opcode),
    .io_in_0_bits_mask         (requestVecFromSlot_0_other_bits_mask),
    .io_in_0_bits_executeMask  (requestVecFromSlot_0_other_bits_executeMask),
    .io_in_0_bits_sign0        (requestVecFromSlot_0_other_bits_sign0),
    .io_in_0_bits_sign         (requestVecFromSlot_0_other_bits_sign),
    .io_in_0_bits_reverse      (requestVecFromSlot_0_other_bits_reverse),
    .io_in_0_bits_average      (requestVecFromSlot_0_other_bits_average),
    .io_in_0_bits_saturate     (requestVecFromSlot_0_other_bits_saturate),
    .io_in_0_bits_vxrm         (requestVecFromSlot_0_other_bits_vxrm),
    .io_in_0_bits_vSew         (requestVecFromSlot_0_other_bits_vSew),
    .io_in_0_bits_shifterSize  (requestVecFromSlot_0_other_bits_shifterSize),
    .io_in_0_bits_rem          (requestVecFromSlot_0_other_bits_rem),
    .io_in_0_bits_executeIndex (requestVecFromSlot_0_other_bits_executeIndex),
    .io_in_0_bits_popInit      (requestVecFromSlot_0_other_bits_popInit),
    .io_in_0_bits_groupIndex   (requestVecFromSlot_0_other_bits_groupIndex),
    .io_in_0_bits_laneIndex    (requestVecFromSlot_0_other_bits_laneIndex),
    .io_in_0_bits_maskType     (requestVecFromSlot_0_other_bits_maskType),
    .io_in_0_bits_narrow       (requestVecFromSlot_0_other_bits_narrow),
    .io_in_1_ready             (requestVecFromSlot_1_other_ready),
    .io_in_1_valid             (requestVecFromSlot_1_other_valid),
    .io_in_1_bits_src_0        (requestVecFromSlot_1_other_bits_src_0),
    .io_in_1_bits_src_1        (requestVecFromSlot_1_other_bits_src_1),
    .io_in_1_bits_src_2        (requestVecFromSlot_1_other_bits_src_2),
    .io_in_1_bits_src_3        (requestVecFromSlot_1_other_bits_src_3),
    .io_in_1_bits_opcode       (requestVecFromSlot_1_other_bits_opcode),
    .io_in_1_bits_mask         (requestVecFromSlot_1_other_bits_mask),
    .io_in_1_bits_executeMask  (requestVecFromSlot_1_other_bits_executeMask),
    .io_in_1_bits_sign0        (requestVecFromSlot_1_other_bits_sign0),
    .io_in_1_bits_sign         (requestVecFromSlot_1_other_bits_sign),
    .io_in_1_bits_reverse      (requestVecFromSlot_1_other_bits_reverse),
    .io_in_1_bits_average      (requestVecFromSlot_1_other_bits_average),
    .io_in_1_bits_saturate     (requestVecFromSlot_1_other_bits_saturate),
    .io_in_1_bits_vxrm         (requestVecFromSlot_1_other_bits_vxrm),
    .io_in_1_bits_vSew         (requestVecFromSlot_1_other_bits_vSew),
    .io_in_1_bits_shifterSize  (requestVecFromSlot_1_other_bits_shifterSize),
    .io_in_1_bits_rem          (requestVecFromSlot_1_other_bits_rem),
    .io_in_1_bits_groupIndex   (requestVecFromSlot_1_other_bits_groupIndex),
    .io_in_1_bits_laneIndex    (requestVecFromSlot_1_other_bits_laneIndex),
    .io_in_1_bits_maskType     (requestVecFromSlot_1_other_bits_maskType),
    .io_in_1_bits_narrow       (requestVecFromSlot_1_other_bits_narrow),
    .io_in_2_ready             (requestVecFromSlot_2_other_ready),
    .io_in_2_valid             (requestVecFromSlot_2_other_valid),
    .io_in_2_bits_src_0        (requestVecFromSlot_2_other_bits_src_0),
    .io_in_2_bits_src_1        (requestVecFromSlot_2_other_bits_src_1),
    .io_in_2_bits_src_2        (requestVecFromSlot_2_other_bits_src_2),
    .io_in_2_bits_src_3        (requestVecFromSlot_2_other_bits_src_3),
    .io_in_2_bits_opcode       (requestVecFromSlot_2_other_bits_opcode),
    .io_in_2_bits_mask         (requestVecFromSlot_2_other_bits_mask),
    .io_in_2_bits_executeMask  (requestVecFromSlot_2_other_bits_executeMask),
    .io_in_2_bits_sign0        (requestVecFromSlot_2_other_bits_sign0),
    .io_in_2_bits_sign         (requestVecFromSlot_2_other_bits_sign),
    .io_in_2_bits_reverse      (requestVecFromSlot_2_other_bits_reverse),
    .io_in_2_bits_average      (requestVecFromSlot_2_other_bits_average),
    .io_in_2_bits_saturate     (requestVecFromSlot_2_other_bits_saturate),
    .io_in_2_bits_vxrm         (requestVecFromSlot_2_other_bits_vxrm),
    .io_in_2_bits_vSew         (requestVecFromSlot_2_other_bits_vSew),
    .io_in_2_bits_shifterSize  (requestVecFromSlot_2_other_bits_shifterSize),
    .io_in_2_bits_rem          (requestVecFromSlot_2_other_bits_rem),
    .io_in_2_bits_groupIndex   (requestVecFromSlot_2_other_bits_groupIndex),
    .io_in_2_bits_laneIndex    (requestVecFromSlot_2_other_bits_laneIndex),
    .io_in_2_bits_maskType     (requestVecFromSlot_2_other_bits_maskType),
    .io_in_2_bits_narrow       (requestVecFromSlot_2_other_bits_narrow),
    .io_in_3_ready             (requestVecFromSlot_3_other_ready),
    .io_in_3_valid             (requestVecFromSlot_3_other_valid),
    .io_in_3_bits_src_0        (requestVecFromSlot_3_other_bits_src_0),
    .io_in_3_bits_src_1        (requestVecFromSlot_3_other_bits_src_1),
    .io_in_3_bits_src_2        (requestVecFromSlot_3_other_bits_src_2),
    .io_in_3_bits_src_3        (requestVecFromSlot_3_other_bits_src_3),
    .io_in_3_bits_opcode       (requestVecFromSlot_3_other_bits_opcode),
    .io_in_3_bits_mask         (requestVecFromSlot_3_other_bits_mask),
    .io_in_3_bits_executeMask  (requestVecFromSlot_3_other_bits_executeMask),
    .io_in_3_bits_sign0        (requestVecFromSlot_3_other_bits_sign0),
    .io_in_3_bits_sign         (requestVecFromSlot_3_other_bits_sign),
    .io_in_3_bits_reverse      (requestVecFromSlot_3_other_bits_reverse),
    .io_in_3_bits_average      (requestVecFromSlot_3_other_bits_average),
    .io_in_3_bits_saturate     (requestVecFromSlot_3_other_bits_saturate),
    .io_in_3_bits_vxrm         (requestVecFromSlot_3_other_bits_vxrm),
    .io_in_3_bits_vSew         (requestVecFromSlot_3_other_bits_vSew),
    .io_in_3_bits_shifterSize  (requestVecFromSlot_3_other_bits_shifterSize),
    .io_in_3_bits_rem          (requestVecFromSlot_3_other_bits_rem),
    .io_in_3_bits_groupIndex   (requestVecFromSlot_3_other_bits_groupIndex),
    .io_in_3_bits_laneIndex    (requestVecFromSlot_3_other_bits_laneIndex),
    .io_in_3_bits_maskType     (requestVecFromSlot_3_other_bits_maskType),
    .io_in_3_bits_narrow       (requestVecFromSlot_3_other_bits_narrow),
    .io_out_ready              (_vfuResponse_otherDistributor_requestFromSlot_ready),
    .io_out_valid              (_vfuResponse_otherArbiter_io_out_valid),
    .io_out_bits_src_0         (_vfuResponse_otherArbiter_io_out_bits_src_0),
    .io_out_bits_src_1         (_vfuResponse_otherArbiter_io_out_bits_src_1),
    .io_out_bits_src_2         (_vfuResponse_otherArbiter_io_out_bits_src_2),
    .io_out_bits_src_3         (_vfuResponse_otherArbiter_io_out_bits_src_3),
    .io_out_bits_opcode        (_vfuResponse_otherArbiter_io_out_bits_opcode),
    .io_out_bits_mask          (_vfuResponse_otherArbiter_io_out_bits_mask),
    .io_out_bits_executeMask   (_vfuResponse_otherArbiter_io_out_bits_executeMask),
    .io_out_bits_sign0         (_vfuResponse_otherArbiter_io_out_bits_sign0),
    .io_out_bits_sign          (_vfuResponse_otherArbiter_io_out_bits_sign),
    .io_out_bits_reverse       (_vfuResponse_otherArbiter_io_out_bits_reverse),
    .io_out_bits_average       (_vfuResponse_otherArbiter_io_out_bits_average),
    .io_out_bits_saturate      (_vfuResponse_otherArbiter_io_out_bits_saturate),
    .io_out_bits_vxrm          (_vfuResponse_otherArbiter_io_out_bits_vxrm),
    .io_out_bits_vSew          (_vfuResponse_otherArbiter_io_out_bits_vSew),
    .io_out_bits_shifterSize   (_vfuResponse_otherArbiter_io_out_bits_shifterSize),
    .io_out_bits_rem           (_vfuResponse_otherArbiter_io_out_bits_rem),
    .io_out_bits_executeIndex  (_vfuResponse_otherArbiter_io_out_bits_executeIndex),
    .io_out_bits_popInit       (_vfuResponse_otherArbiter_io_out_bits_popInit),
    .io_out_bits_groupIndex    (_vfuResponse_otherArbiter_io_out_bits_groupIndex),
    .io_out_bits_laneIndex     (_vfuResponse_otherArbiter_io_out_bits_laneIndex),
    .io_out_bits_maskType      (_vfuResponse_otherArbiter_io_out_bits_maskType),
    .io_out_bits_narrow        (_vfuResponse_otherArbiter_io_out_bits_narrow),
    .io_out_bits_tag           (_vfuResponse_otherArbiter_io_out_bits_tag)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_0 (
    .io_in_0_ready                 (readBeforeMaskedWrite_ready),
    .io_in_0_valid                 (readBeforeMaskedWrite_valid),
    .io_in_0_bits_vs               (readBeforeMaskedWrite_bits_vs),
    .io_in_0_bits_readSource       (2'h2),
    .io_in_0_bits_offset           (readBeforeMaskedWrite_bits_offset),
    .io_in_0_bits_instructionIndex (readBeforeMaskedWrite_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_0_ready),
    .io_out_valid                  (_vrfReadArbiter_0_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_0_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_0_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_0_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_0_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_1 (
    .io_in_0_ready                 (vrfReadRequest_0_0_ready),
    .io_in_0_valid                 (vrfReadRequest_0_0_valid),
    .io_in_0_bits_vs               (vrfReadRequest_0_0_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_0_0_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_0_0_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_0_0_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_1_ready),
    .io_out_valid                  (_vrfReadArbiter_1_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_1_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_1_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_1_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_1_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_2 (
    .io_in_0_ready                 (vrfReadRequest_0_1_ready),
    .io_in_0_valid                 (vrfReadRequest_0_1_valid),
    .io_in_0_bits_vs               (vrfReadRequest_0_1_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_0_1_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_0_1_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_0_1_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_2_ready),
    .io_out_valid                  (_vrfReadArbiter_2_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_2_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_2_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_2_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_2_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_3 (
    .io_in_0_ready                 (vrfReadRequest_0_2_ready),
    .io_in_0_valid                 (vrfReadRequest_0_2_valid),
    .io_in_0_bits_vs               (vrfReadRequest_0_2_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_0_2_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_0_2_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_0_2_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_3_ready),
    .io_out_valid                  (_vrfReadArbiter_3_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_3_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_3_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_3_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_3_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_4 (
    .io_in_0_ready                 (vrfReadRequest_1_0_ready),
    .io_in_0_valid                 (vrfReadRequest_1_0_valid),
    .io_in_0_bits_vs               (vrfReadRequest_1_0_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_1_0_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_1_0_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_1_0_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_4_ready),
    .io_out_valid                  (_vrfReadArbiter_4_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_4_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_4_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_4_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_4_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_5 (
    .io_in_0_ready                 (vrfReadRequest_1_1_ready),
    .io_in_0_valid                 (vrfReadRequest_1_1_valid),
    .io_in_0_bits_vs               (vrfReadRequest_1_1_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_1_1_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_1_1_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_1_1_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_5_ready),
    .io_out_valid                  (_vrfReadArbiter_5_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_5_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_5_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_5_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_5_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_6 (
    .io_in_0_ready                 (vrfReadRequest_1_2_ready),
    .io_in_0_valid                 (vrfReadRequest_1_2_valid),
    .io_in_0_bits_vs               (vrfReadRequest_1_2_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_1_2_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_1_2_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_1_2_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_6_ready),
    .io_out_valid                  (_vrfReadArbiter_6_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_6_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_6_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_6_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_6_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_7 (
    .io_in_0_ready                 (vrfReadRequest_2_0_ready),
    .io_in_0_valid                 (vrfReadRequest_2_0_valid),
    .io_in_0_bits_vs               (vrfReadRequest_2_0_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_2_0_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_2_0_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_2_0_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_7_ready),
    .io_out_valid                  (_vrfReadArbiter_7_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_7_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_7_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_7_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_7_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_8 (
    .io_in_0_ready                 (vrfReadRequest_2_1_ready),
    .io_in_0_valid                 (vrfReadRequest_2_1_valid),
    .io_in_0_bits_vs               (vrfReadRequest_2_1_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_2_1_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_2_1_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_2_1_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_8_ready),
    .io_out_valid                  (_vrfReadArbiter_8_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_8_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_8_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_8_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_8_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_9 (
    .io_in_0_ready                 (vrfReadRequest_2_2_ready),
    .io_in_0_valid                 (vrfReadRequest_2_2_valid),
    .io_in_0_bits_vs               (vrfReadRequest_2_2_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_2_2_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_2_2_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_2_2_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_9_ready),
    .io_out_valid                  (_vrfReadArbiter_9_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_9_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_9_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_9_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_9_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_10 (
    .io_in_0_ready                 (vrfReadRequest_3_0_ready),
    .io_in_0_valid                 (vrfReadRequest_3_0_valid),
    .io_in_0_bits_vs               (vrfReadRequest_3_0_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_3_0_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_3_0_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_3_0_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_10_ready),
    .io_out_valid                  (_vrfReadArbiter_10_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_10_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_10_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_10_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_10_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_11 (
    .io_in_0_ready                 (vrfReadRequest_3_1_ready),
    .io_in_0_valid                 (vrfReadRequest_3_1_valid),
    .io_in_0_bits_vs               (vrfReadRequest_3_1_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_3_1_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_3_1_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_3_1_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_11_ready),
    .io_out_valid                  (_vrfReadArbiter_11_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_11_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_11_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_11_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_11_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_12 (
    .io_in_0_ready                 (vrfReadRequest_3_2_ready),
    .io_in_0_valid                 (vrfReadRequest_3_2_valid),
    .io_in_0_bits_vs               (vrfReadRequest_3_2_bits_vs),
    .io_in_0_bits_readSource       (vrfReadRequest_3_2_bits_readSource),
    .io_in_0_bits_offset           (vrfReadRequest_3_2_bits_offset),
    .io_in_0_bits_instructionIndex (vrfReadRequest_3_2_bits_instructionIndex),
    .io_out_ready                  (_vrf_readRequests_12_ready),
    .io_out_valid                  (_vrfReadArbiter_12_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_12_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_12_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_12_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_12_io_out_bits_instructionIndex)
  );
  Arbiter1_VRFReadRequest vrfReadArbiter_13 (
    .io_in_0_ready                 (vrfReadAddressChannel_ready_0),
    .io_in_0_valid                 (vrfReadAddressChannel_valid_0),
    .io_in_0_bits_vs               (vrfReadAddressChannel_bits_vs_0),
    .io_in_0_bits_readSource       (vrfReadAddressChannel_bits_readSource_0),
    .io_in_0_bits_offset           (vrfReadAddressChannel_bits_offset_0),
    .io_in_0_bits_instructionIndex (vrfReadAddressChannel_bits_instructionIndex_0),
    .io_out_ready                  (_vrf_readRequests_13_ready),
    .io_out_valid                  (_vrfReadArbiter_13_io_out_valid),
    .io_out_bits_vs                (_vrfReadArbiter_13_io_out_bits_vs),
    .io_out_bits_readSource        (_vrfReadArbiter_13_io_out_bits_readSource),
    .io_out_bits_offset            (_vrfReadArbiter_13_io_out_bits_offset),
    .io_out_bits_instructionIndex  (_vrfReadArbiter_13_io_out_bits_instructionIndex)
  );
  assign readBusPort_0_enqRelease = readBusPort_0_enqRelease_0;
  assign readBusPort_0_deq_valid = readBusPort_0_deq_valid_0;
  assign readBusPort_0_deq_bits_data = readBusPort_0_deq_bits_data_0;
  assign readBusPort_1_enqRelease = readBusPort_1_enqRelease_0;
  assign readBusPort_1_deq_valid = readBusPort_1_deq_valid_0;
  assign readBusPort_1_deq_bits_data = readBusPort_1_deq_bits_data_0;
  assign writeBusPort_0_enqRelease = writeBusPort_0_enqRelease_0;
  assign writeBusPort_0_deq_valid = writeBusPort_0_deq_valid_0;
  assign writeBusPort_0_deq_bits_data = writeBusPort_0_deq_bits_data_0;
  assign writeBusPort_0_deq_bits_mask = writeBusPort_0_deq_bits_mask_0;
  assign writeBusPort_0_deq_bits_instructionIndex = writeBusPort_0_deq_bits_instructionIndex_0;
  assign writeBusPort_0_deq_bits_counter = writeBusPort_0_deq_bits_counter_0;
  assign writeBusPort_1_enqRelease = writeBusPort_1_enqRelease_0;
  assign writeBusPort_1_deq_valid = writeBusPort_1_deq_valid_0;
  assign writeBusPort_1_deq_bits_data = writeBusPort_1_deq_bits_data_0;
  assign writeBusPort_1_deq_bits_mask = writeBusPort_1_deq_bits_mask_0;
  assign writeBusPort_1_deq_bits_instructionIndex = writeBusPort_1_deq_bits_instructionIndex_0;
  assign writeBusPort_1_deq_bits_counter = writeBusPort_1_deq_bits_counter_0;
  assign laneRequest_ready = laneRequest_ready_0;
  assign maskUnitRequest_valid = _maskStage_maskReq_valid;
  assign maskUnitRequest_bits_index = _maskStage_maskReq_bits_index;
  assign vrfReadAddressChannel_ready = vrfReadAddressChannel_ready_0;
  assign vrfWriteChannel_ready = vrfWriteChannel_ready_0;
  assign instructionFinished = _instructionFinished_output;
  assign vxsatReport = vxsatResult;
  assign v0Update_valid = _maskedWriteUnit_dequeue_valid & _maskedWriteUnit_dequeue_bits_vd == 5'h0;
  assign v0Update_bits_data = _maskedWriteUnit_dequeue_bits_data;
  assign v0Update_bits_offset = _maskedWriteUnit_dequeue_bits_offset;
  assign v0Update_bits_mask = _maskedWriteUnit_dequeue_bits_mask;
  assign maskSelect =
    (maskControlReqSelect[0] ? maskControlVec_0_group : 8'h0) | (maskControlReqSelect[1] ? maskControlVec_1_group : 8'h0) | (maskControlReqSelect[2] ? maskControlVec_2_group : 8'h0)
    | (maskControlReqSelect[3] ? maskControlVec_3_group : 8'h0);
  assign maskSelectSew =
    (maskControlReqSelect[0] ? maskControlVec_0_sew : 2'h0) | (maskControlReqSelect[1] ? maskControlVec_1_sew : 2'h0) | (maskControlReqSelect[2] ? maskControlVec_2_sew : 2'h0) | (maskControlReqSelect[3] ? maskControlVec_3_sew : 2'h0);
endmodule

