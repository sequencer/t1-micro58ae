
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module StoreUnit(
  input          clock,
                 reset,
                 lsuRequest_valid,
  input  [2:0]   lsuRequest_bits_instructionInformation_nf,
  input          lsuRequest_bits_instructionInformation_mew,
  input  [1:0]   lsuRequest_bits_instructionInformation_mop,
  input  [4:0]   lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]   lsuRequest_bits_instructionInformation_eew,
  input  [4:0]   lsuRequest_bits_instructionInformation_vs3,
  input          lsuRequest_bits_instructionInformation_isStore,
                 lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]  lsuRequest_bits_rs1Data,
                 lsuRequest_bits_rs2Data,
  input  [2:0]   lsuRequest_bits_instructionIndex,
  input  [11:0]  csrInterface_vl,
                 csrInterface_vStart,
  input  [2:0]   csrInterface_vlmul,
  input  [1:0]   csrInterface_vSew,
                 csrInterface_vxrm,
  input          csrInterface_vta,
                 csrInterface_vma,
  input  [31:0]  maskInput,
  output         maskSelect_valid,
  output [5:0]   maskSelect_bits,
  input          memRequest_ready,
  output         memRequest_valid,
  output [255:0] memRequest_bits_data,
  output [31:0]  memRequest_bits_mask,
  output [6:0]   memRequest_bits_index,
  output [31:0]  memRequest_bits_address,
  output         status_idle,
                 status_last,
  output [2:0]   status_instructionIndex,
  output         status_changeMaskGroup,
  output [31:0]  status_startAddress,
                 status_endAddress,
  input          vrfReadDataPorts_0_ready,
  output         vrfReadDataPorts_0_valid,
  output [4:0]   vrfReadDataPorts_0_bits_vs,
  output [2:0]   vrfReadDataPorts_0_bits_offset,
                 vrfReadDataPorts_0_bits_instructionIndex,
  input          vrfReadDataPorts_1_ready,
  output         vrfReadDataPorts_1_valid,
  output [4:0]   vrfReadDataPorts_1_bits_vs,
  output [2:0]   vrfReadDataPorts_1_bits_offset,
                 vrfReadDataPorts_1_bits_instructionIndex,
  input          vrfReadDataPorts_2_ready,
  output         vrfReadDataPorts_2_valid,
  output [4:0]   vrfReadDataPorts_2_bits_vs,
  output [2:0]   vrfReadDataPorts_2_bits_offset,
                 vrfReadDataPorts_2_bits_instructionIndex,
  input          vrfReadDataPorts_3_ready,
  output         vrfReadDataPorts_3_valid,
  output [4:0]   vrfReadDataPorts_3_bits_vs,
  output [2:0]   vrfReadDataPorts_3_bits_offset,
                 vrfReadDataPorts_3_bits_instructionIndex,
  input          vrfReadDataPorts_4_ready,
  output         vrfReadDataPorts_4_valid,
  output [4:0]   vrfReadDataPorts_4_bits_vs,
  output [2:0]   vrfReadDataPorts_4_bits_offset,
                 vrfReadDataPorts_4_bits_instructionIndex,
  input          vrfReadDataPorts_5_ready,
  output         vrfReadDataPorts_5_valid,
  output [4:0]   vrfReadDataPorts_5_bits_vs,
  output [2:0]   vrfReadDataPorts_5_bits_offset,
                 vrfReadDataPorts_5_bits_instructionIndex,
  input          vrfReadDataPorts_6_ready,
  output         vrfReadDataPorts_6_valid,
  output [4:0]   vrfReadDataPorts_6_bits_vs,
  output [2:0]   vrfReadDataPorts_6_bits_offset,
                 vrfReadDataPorts_6_bits_instructionIndex,
  input          vrfReadDataPorts_7_ready,
  output         vrfReadDataPorts_7_valid,
  output [4:0]   vrfReadDataPorts_7_bits_vs,
  output [2:0]   vrfReadDataPorts_7_bits_offset,
                 vrfReadDataPorts_7_bits_instructionIndex,
  input          vrfReadResults_0_valid,
  input  [31:0]  vrfReadResults_0_bits,
  input          vrfReadResults_1_valid,
  input  [31:0]  vrfReadResults_1_bits,
  input          vrfReadResults_2_valid,
  input  [31:0]  vrfReadResults_2_bits,
  input          vrfReadResults_3_valid,
  input  [31:0]  vrfReadResults_3_bits,
  input          vrfReadResults_4_valid,
  input  [31:0]  vrfReadResults_4_bits,
  input          vrfReadResults_5_valid,
  input  [31:0]  vrfReadResults_5_bits,
  input          vrfReadResults_6_valid,
  input  [31:0]  vrfReadResults_6_bits,
  input          vrfReadResults_7_valid,
  input  [31:0]  vrfReadResults_7_bits,
  input          storeResponse
);

  wire             _addressQueue_fifo_empty;
  wire             _addressQueue_fifo_full;
  wire             _addressQueue_fifo_error;
  wire             _vrfReadQueueVec_fifo_7_empty;
  wire             _vrfReadQueueVec_fifo_7_full;
  wire             _vrfReadQueueVec_fifo_7_error;
  wire [31:0]      _vrfReadQueueVec_fifo_7_data_out;
  wire             _vrfReadQueueVec_fifo_6_empty;
  wire             _vrfReadQueueVec_fifo_6_full;
  wire             _vrfReadQueueVec_fifo_6_error;
  wire [31:0]      _vrfReadQueueVec_fifo_6_data_out;
  wire             _vrfReadQueueVec_fifo_5_empty;
  wire             _vrfReadQueueVec_fifo_5_full;
  wire             _vrfReadQueueVec_fifo_5_error;
  wire [31:0]      _vrfReadQueueVec_fifo_5_data_out;
  wire             _vrfReadQueueVec_fifo_4_empty;
  wire             _vrfReadQueueVec_fifo_4_full;
  wire             _vrfReadQueueVec_fifo_4_error;
  wire [31:0]      _vrfReadQueueVec_fifo_4_data_out;
  wire             _vrfReadQueueVec_fifo_3_empty;
  wire             _vrfReadQueueVec_fifo_3_full;
  wire             _vrfReadQueueVec_fifo_3_error;
  wire [31:0]      _vrfReadQueueVec_fifo_3_data_out;
  wire             _vrfReadQueueVec_fifo_2_empty;
  wire             _vrfReadQueueVec_fifo_2_full;
  wire             _vrfReadQueueVec_fifo_2_error;
  wire [31:0]      _vrfReadQueueVec_fifo_2_data_out;
  wire             _vrfReadQueueVec_fifo_1_empty;
  wire             _vrfReadQueueVec_fifo_1_full;
  wire             _vrfReadQueueVec_fifo_1_error;
  wire [31:0]      _vrfReadQueueVec_fifo_1_data_out;
  wire             _vrfReadQueueVec_fifo_empty;
  wire             _vrfReadQueueVec_fifo_full;
  wire             _vrfReadQueueVec_fifo_error;
  wire [31:0]      _vrfReadQueueVec_fifo_data_out;
  wire             addressQueue_almostFull;
  wire             addressQueue_almostEmpty;
  wire             vrfReadQueueVec_7_almostFull;
  wire             vrfReadQueueVec_7_almostEmpty;
  wire             vrfReadQueueVec_6_almostFull;
  wire             vrfReadQueueVec_6_almostEmpty;
  wire             vrfReadQueueVec_5_almostFull;
  wire             vrfReadQueueVec_5_almostEmpty;
  wire             vrfReadQueueVec_4_almostFull;
  wire             vrfReadQueueVec_4_almostEmpty;
  wire             vrfReadQueueVec_3_almostFull;
  wire             vrfReadQueueVec_3_almostEmpty;
  wire             vrfReadQueueVec_2_almostFull;
  wire             vrfReadQueueVec_2_almostEmpty;
  wire             vrfReadQueueVec_1_almostFull;
  wire             vrfReadQueueVec_1_almostEmpty;
  wire             vrfReadQueueVec_0_almostFull;
  wire             vrfReadQueueVec_0_almostEmpty;
  wire             memRequest_ready_0 = memRequest_ready;
  wire             vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire             vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire             vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire             vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire             vrfReadDataPorts_4_ready_0 = vrfReadDataPorts_4_ready;
  wire             vrfReadDataPorts_5_ready_0 = vrfReadDataPorts_5_ready;
  wire             vrfReadDataPorts_6_ready_0 = vrfReadDataPorts_6_ready;
  wire             vrfReadDataPorts_7_ready_0 = vrfReadDataPorts_7_ready;
  wire             vrfReadQueueVec_0_enq_valid = vrfReadResults_0_valid;
  wire [31:0]      vrfReadQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire             vrfReadQueueVec_1_enq_valid = vrfReadResults_1_valid;
  wire [31:0]      vrfReadQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire             vrfReadQueueVec_2_enq_valid = vrfReadResults_2_valid;
  wire [31:0]      vrfReadQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire             vrfReadQueueVec_3_enq_valid = vrfReadResults_3_valid;
  wire [31:0]      vrfReadQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire             vrfReadQueueVec_4_enq_valid = vrfReadResults_4_valid;
  wire [31:0]      vrfReadQueueVec_4_enq_bits = vrfReadResults_4_bits;
  wire             vrfReadQueueVec_5_enq_valid = vrfReadResults_5_valid;
  wire [31:0]      vrfReadQueueVec_5_enq_bits = vrfReadResults_5_bits;
  wire             vrfReadQueueVec_6_enq_valid = vrfReadResults_6_valid;
  wire [31:0]      vrfReadQueueVec_6_enq_bits = vrfReadResults_6_bits;
  wire             vrfReadQueueVec_7_enq_valid = vrfReadResults_7_valid;
  wire [31:0]      vrfReadQueueVec_7_enq_bits = vrfReadResults_7_bits;
  wire             addressQueue_deq_ready = storeResponse;
  wire [1:0]       accessStateCheck_lo_lo = 2'h0;
  wire [1:0]       accessStateCheck_lo_hi = 2'h0;
  wire [1:0]       accessStateCheck_hi_lo = 2'h0;
  wire [1:0]       accessStateCheck_hi_hi = 2'h0;
  wire [3:0]       accessStateCheck_lo = 4'h0;
  wire [3:0]       accessStateCheck_hi = 4'h0;
  wire             accessStateCheck = 1'h1;
  wire             accessStateUpdate_0 = 1'h0;
  wire             accessStateUpdate_1 = 1'h0;
  wire             accessStateUpdate_2 = 1'h0;
  wire             accessStateUpdate_3 = 1'h0;
  wire             accessStateUpdate_4 = 1'h0;
  wire             accessStateUpdate_5 = 1'h0;
  wire             accessStateUpdate_6 = 1'h0;
  wire             accessStateUpdate_7 = 1'h0;
  wire [1023:0]    hi = 1024'h0;
  wire [1023:0]    hi_1 = 1024'h0;
  wire [1023:0]    hi_2 = 1024'h0;
  wire [1023:0]    hi_3 = 1024'h0;
  wire [1023:0]    hi_8 = 1024'h0;
  wire [1023:0]    hi_9 = 1024'h0;
  wire [1023:0]    hi_10 = 1024'h0;
  wire [1023:0]    hi_11 = 1024'h0;
  wire [1023:0]    hi_16 = 1024'h0;
  wire [1023:0]    hi_17 = 1024'h0;
  wire [1023:0]    hi_18 = 1024'h0;
  wire [1023:0]    hi_19 = 1024'h0;
  wire [511:0]     lo_hi = 512'h0;
  wire [511:0]     hi_lo = 512'h0;
  wire [511:0]     hi_hi = 512'h0;
  wire [511:0]     lo_hi_1 = 512'h0;
  wire [511:0]     hi_lo_1 = 512'h0;
  wire [511:0]     hi_hi_1 = 512'h0;
  wire [511:0]     hi_lo_2 = 512'h0;
  wire [511:0]     hi_hi_2 = 512'h0;
  wire [511:0]     hi_lo_3 = 512'h0;
  wire [511:0]     hi_hi_3 = 512'h0;
  wire [511:0]     hi_hi_4 = 512'h0;
  wire [511:0]     hi_hi_5 = 512'h0;
  wire [511:0]     lo_hi_8 = 512'h0;
  wire [511:0]     hi_lo_8 = 512'h0;
  wire [511:0]     hi_hi_8 = 512'h0;
  wire [511:0]     lo_hi_9 = 512'h0;
  wire [511:0]     hi_lo_9 = 512'h0;
  wire [511:0]     hi_hi_9 = 512'h0;
  wire [511:0]     hi_lo_10 = 512'h0;
  wire [511:0]     hi_hi_10 = 512'h0;
  wire [511:0]     hi_lo_11 = 512'h0;
  wire [511:0]     hi_hi_11 = 512'h0;
  wire [511:0]     hi_hi_12 = 512'h0;
  wire [511:0]     hi_hi_13 = 512'h0;
  wire [511:0]     lo_hi_16 = 512'h0;
  wire [511:0]     hi_lo_16 = 512'h0;
  wire [511:0]     hi_hi_16 = 512'h0;
  wire [511:0]     lo_hi_17 = 512'h0;
  wire [511:0]     hi_lo_17 = 512'h0;
  wire [511:0]     hi_hi_17 = 512'h0;
  wire [511:0]     hi_lo_18 = 512'h0;
  wire [511:0]     hi_hi_18 = 512'h0;
  wire [511:0]     hi_lo_19 = 512'h0;
  wire [511:0]     hi_hi_19 = 512'h0;
  wire [511:0]     hi_hi_20 = 512'h0;
  wire [511:0]     hi_hi_21 = 512'h0;
  wire [255:0]     res_1 = 256'h0;
  wire [255:0]     res_2 = 256'h0;
  wire [255:0]     res_3 = 256'h0;
  wire [255:0]     res_4 = 256'h0;
  wire [255:0]     res_5 = 256'h0;
  wire [255:0]     res_6 = 256'h0;
  wire [255:0]     res_7 = 256'h0;
  wire [255:0]     res_10 = 256'h0;
  wire [255:0]     res_11 = 256'h0;
  wire [255:0]     res_12 = 256'h0;
  wire [255:0]     res_13 = 256'h0;
  wire [255:0]     res_14 = 256'h0;
  wire [255:0]     res_15 = 256'h0;
  wire [255:0]     res_19 = 256'h0;
  wire [255:0]     res_20 = 256'h0;
  wire [255:0]     res_21 = 256'h0;
  wire [255:0]     res_22 = 256'h0;
  wire [255:0]     res_23 = 256'h0;
  wire [255:0]     res_28 = 256'h0;
  wire [255:0]     res_29 = 256'h0;
  wire [255:0]     res_30 = 256'h0;
  wire [255:0]     res_31 = 256'h0;
  wire [255:0]     res_37 = 256'h0;
  wire [255:0]     res_38 = 256'h0;
  wire [255:0]     res_39 = 256'h0;
  wire [255:0]     res_46 = 256'h0;
  wire [255:0]     res_47 = 256'h0;
  wire [255:0]     res_55 = 256'h0;
  wire [255:0]     res_65 = 256'h0;
  wire [255:0]     res_66 = 256'h0;
  wire [255:0]     res_67 = 256'h0;
  wire [255:0]     res_68 = 256'h0;
  wire [255:0]     res_69 = 256'h0;
  wire [255:0]     res_70 = 256'h0;
  wire [255:0]     res_71 = 256'h0;
  wire [255:0]     res_74 = 256'h0;
  wire [255:0]     res_75 = 256'h0;
  wire [255:0]     res_76 = 256'h0;
  wire [255:0]     res_77 = 256'h0;
  wire [255:0]     res_78 = 256'h0;
  wire [255:0]     res_79 = 256'h0;
  wire [255:0]     res_83 = 256'h0;
  wire [255:0]     res_84 = 256'h0;
  wire [255:0]     res_85 = 256'h0;
  wire [255:0]     res_86 = 256'h0;
  wire [255:0]     res_87 = 256'h0;
  wire [255:0]     res_92 = 256'h0;
  wire [255:0]     res_93 = 256'h0;
  wire [255:0]     res_94 = 256'h0;
  wire [255:0]     res_95 = 256'h0;
  wire [255:0]     res_101 = 256'h0;
  wire [255:0]     res_102 = 256'h0;
  wire [255:0]     res_103 = 256'h0;
  wire [255:0]     res_110 = 256'h0;
  wire [255:0]     res_111 = 256'h0;
  wire [255:0]     res_119 = 256'h0;
  wire [255:0]     res_129 = 256'h0;
  wire [255:0]     res_130 = 256'h0;
  wire [255:0]     res_131 = 256'h0;
  wire [255:0]     res_132 = 256'h0;
  wire [255:0]     res_133 = 256'h0;
  wire [255:0]     res_134 = 256'h0;
  wire [255:0]     res_135 = 256'h0;
  wire [255:0]     res_138 = 256'h0;
  wire [255:0]     res_139 = 256'h0;
  wire [255:0]     res_140 = 256'h0;
  wire [255:0]     res_141 = 256'h0;
  wire [255:0]     res_142 = 256'h0;
  wire [255:0]     res_143 = 256'h0;
  wire [255:0]     res_147 = 256'h0;
  wire [255:0]     res_148 = 256'h0;
  wire [255:0]     res_149 = 256'h0;
  wire [255:0]     res_150 = 256'h0;
  wire [255:0]     res_151 = 256'h0;
  wire [255:0]     res_156 = 256'h0;
  wire [255:0]     res_157 = 256'h0;
  wire [255:0]     res_158 = 256'h0;
  wire [255:0]     res_159 = 256'h0;
  wire [255:0]     res_165 = 256'h0;
  wire [255:0]     res_166 = 256'h0;
  wire [255:0]     res_167 = 256'h0;
  wire [255:0]     res_174 = 256'h0;
  wire [255:0]     res_175 = 256'h0;
  wire [255:0]     res_183 = 256'h0;
  wire [1:0]       vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_4_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_5_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_6_bits_readSource = 2'h2;
  wire [1:0]       vrfReadDataPorts_7_bits_readSource = 2'h2;
  wire [31:0]      alignedDequeueAddress;
  reg  [2:0]       lsuRequestReg_instructionInformation_nf;
  reg              lsuRequestReg_instructionInformation_mew;
  reg  [1:0]       lsuRequestReg_instructionInformation_mop;
  reg  [4:0]       lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]       lsuRequestReg_instructionInformation_eew;
  reg  [4:0]       lsuRequestReg_instructionInformation_vs3;
  reg              lsuRequestReg_instructionInformation_isStore;
  reg              lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]      lsuRequestReg_rs1Data;
  reg  [31:0]      lsuRequestReg_rs2Data;
  reg  [2:0]       lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_0_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_1_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_2_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_3_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_4_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_5_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_6_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]       vrfReadDataPorts_7_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [11:0]      csrInterfaceReg_vl;
  reg  [11:0]      csrInterfaceReg_vStart;
  reg  [2:0]       csrInterfaceReg_vlmul;
  reg  [1:0]       csrInterfaceReg_vSew;
  reg  [1:0]       csrInterfaceReg_vxrm;
  reg              csrInterfaceReg_vta;
  reg              csrInterfaceReg_vma;
  reg              requestFireNext;
  reg  [1:0]       dataEEW;
  wire [3:0]       _dataEEWOH_T = 4'h1 << dataEEW;
  wire [2:0]       dataEEWOH = _dataEEWOH_T[2:0];
  wire             isMaskType = lsuRequest_valid ? lsuRequest_bits_instructionInformation_maskedLoadStore : lsuRequestReg_instructionInformation_maskedLoadStore;
  wire [31:0]      maskAmend = isMaskType ? maskInput : 32'hFFFFFFFF;
  reg  [31:0]      maskReg;
  wire [31:0]      _lastMaskAmend_T_1 = 32'h1 << csrInterface_vl[4:0];
  wire [29:0]      _GEN = _lastMaskAmend_T_1[30:1] | _lastMaskAmend_T_1[31:2];
  wire [28:0]      _GEN_0 = _GEN[28:0] | {_lastMaskAmend_T_1[31], _GEN[29:2]};
  wire [26:0]      _GEN_1 = _GEN_0[26:0] | {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:4]};
  wire [22:0]      _GEN_2 = _GEN_1[22:0] | {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:27], _GEN_1[26:8]};
  wire [30:0]      lastMaskAmend = {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:27], _GEN_1[26:23], _GEN_2[22:15], _GEN_2[14:0] | {_lastMaskAmend_T_1[31], _GEN[29], _GEN_0[28:27], _GEN_1[26:23], _GEN_2[22:16]}};
  reg              needAmend;
  reg  [30:0]      lastMaskAmendReg;
  wire [1:0]       countEndForGroup = {1'h0, dataEEWOH[1]} | {2{dataEEWOH[2]}};
  reg  [5:0]       maskGroupCounter;
  wire [5:0]       nextMaskGroup = maskGroupCounter + 6'h1;
  reg  [1:0]       maskCounterInGroup;
  wire [1:0]       nextMaskCount = maskCounterInGroup + 2'h1;
  wire             isLastDataGroup = maskCounterInGroup == countEndForGroup;
  wire [5:0]       _maskSelect_bits_output = lsuRequest_valid ? 6'h0 : nextMaskGroup;
  reg              isLastMaskGroup;
  wire [31:0]      maskWire = maskReg & (needAmend & isLastMaskGroup ? {1'h0, lastMaskAmendReg} : 32'hFFFFFFFF);
  wire [3:0]       maskForGroupWire_lo_lo_lo_lo = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]       maskForGroupWire_lo_lo_lo_hi = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo = {maskForGroupWire_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo};
  wire [3:0]       maskForGroupWire_lo_lo_hi_lo = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi_hi = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi = {maskForGroupWire_lo_lo_hi_hi, maskForGroupWire_lo_lo_hi_lo};
  wire [15:0]      maskForGroupWire_lo_lo = {maskForGroupWire_lo_lo_hi, maskForGroupWire_lo_lo_lo};
  wire [3:0]       maskForGroupWire_lo_hi_lo_lo = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]       maskForGroupWire_lo_hi_lo_hi = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo = {maskForGroupWire_lo_hi_lo_hi, maskForGroupWire_lo_hi_lo_lo};
  wire [3:0]       maskForGroupWire_lo_hi_hi_lo = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi_hi = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi = {maskForGroupWire_lo_hi_hi_hi, maskForGroupWire_lo_hi_hi_lo};
  wire [15:0]      maskForGroupWire_lo_hi = {maskForGroupWire_lo_hi_hi, maskForGroupWire_lo_hi_lo};
  wire [31:0]      maskForGroupWire_lo = {maskForGroupWire_lo_hi, maskForGroupWire_lo_lo};
  wire [3:0]       maskForGroupWire_hi_lo_lo_lo = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]       maskForGroupWire_hi_lo_lo_hi = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo = {maskForGroupWire_hi_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo};
  wire [3:0]       maskForGroupWire_hi_lo_hi_lo = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi_hi = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi = {maskForGroupWire_hi_lo_hi_hi, maskForGroupWire_hi_lo_hi_lo};
  wire [15:0]      maskForGroupWire_hi_lo = {maskForGroupWire_hi_lo_hi, maskForGroupWire_hi_lo_lo};
  wire [3:0]       maskForGroupWire_hi_hi_lo_lo = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]       maskForGroupWire_hi_hi_lo_hi = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo = {maskForGroupWire_hi_hi_lo_hi, maskForGroupWire_hi_hi_lo_lo};
  wire [3:0]       maskForGroupWire_hi_hi_hi_lo = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi_hi = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_lo};
  wire [15:0]      maskForGroupWire_hi_hi = {maskForGroupWire_hi_hi_hi, maskForGroupWire_hi_hi_lo};
  wire [31:0]      maskForGroupWire_hi = {maskForGroupWire_hi_hi, maskForGroupWire_hi_lo};
  wire [3:0]       maskForGroupWire_lo_lo_lo_lo_1 = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]       maskForGroupWire_lo_lo_lo_hi_1 = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_lo_hi_lo_1 = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]       maskForGroupWire_lo_lo_hi_hi_1 = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_1 = {maskForGroupWire_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_hi_lo_1};
  wire [15:0]      maskForGroupWire_lo_lo_1 = {maskForGroupWire_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_hi_lo_lo_1 = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]       maskForGroupWire_lo_hi_lo_hi_1 = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_1 = {maskForGroupWire_lo_hi_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_lo_hi_hi_lo_1 = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]       maskForGroupWire_lo_hi_hi_hi_1 = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_lo_1};
  wire [15:0]      maskForGroupWire_lo_hi_1 = {maskForGroupWire_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_1};
  wire [31:0]      maskForGroupWire_lo_1 = {maskForGroupWire_lo_hi_1, maskForGroupWire_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_lo_lo_lo_1 = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]       maskForGroupWire_hi_lo_lo_hi_1 = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_1 = {maskForGroupWire_hi_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_lo_hi_lo_1 = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]       maskForGroupWire_hi_lo_hi_hi_1 = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_1 = {maskForGroupWire_hi_lo_hi_hi_1, maskForGroupWire_hi_lo_hi_lo_1};
  wire [15:0]      maskForGroupWire_hi_lo_1 = {maskForGroupWire_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_hi_lo_lo_1 = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]       maskForGroupWire_hi_hi_lo_hi_1 = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_1 = {maskForGroupWire_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_1};
  wire [3:0]       maskForGroupWire_hi_hi_hi_lo_1 = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]       maskForGroupWire_hi_hi_hi_hi_1 = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_lo_1};
  wire [15:0]      maskForGroupWire_hi_hi_1 = {maskForGroupWire_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_1};
  wire [31:0]      maskForGroupWire_hi_1 = {maskForGroupWire_hi_hi_1, maskForGroupWire_hi_lo_1};
  wire [3:0]       _maskForGroupWire_T_133 = 4'h1 << maskCounterInGroup;
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_2 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_2 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_2 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_2 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_2 = {maskForGroupWire_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_hi_lo_2};
  wire [31:0]      maskForGroupWire_lo_lo_2 = {maskForGroupWire_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_2 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_2 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_2 = {maskForGroupWire_lo_hi_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_2 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_2 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_lo_2};
  wire [31:0]      maskForGroupWire_lo_hi_2 = {maskForGroupWire_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_2};
  wire [63:0]      maskForGroupWire_lo_2 = {maskForGroupWire_lo_hi_2, maskForGroupWire_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_2 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_2 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_2 = {maskForGroupWire_hi_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_2 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_2 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_2 = {maskForGroupWire_hi_lo_hi_hi_2, maskForGroupWire_hi_lo_hi_lo_2};
  wire [31:0]      maskForGroupWire_hi_lo_2 = {maskForGroupWire_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_2 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_2 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_2 = {maskForGroupWire_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_2};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_2 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_2 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_lo_2};
  wire [31:0]      maskForGroupWire_hi_hi_2 = {maskForGroupWire_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_2};
  wire [63:0]      maskForGroupWire_hi_2 = {maskForGroupWire_hi_hi_2, maskForGroupWire_hi_lo_2};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_3 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_3 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_3 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_3 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_3 = {maskForGroupWire_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_hi_lo_3};
  wire [31:0]      maskForGroupWire_lo_lo_3 = {maskForGroupWire_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_3 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_3 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_3 = {maskForGroupWire_lo_hi_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_3 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_3 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_lo_3};
  wire [31:0]      maskForGroupWire_lo_hi_3 = {maskForGroupWire_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_3};
  wire [63:0]      maskForGroupWire_lo_3 = {maskForGroupWire_lo_hi_3, maskForGroupWire_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_3 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_3 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_3 = {maskForGroupWire_hi_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_3 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_3 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_3 = {maskForGroupWire_hi_lo_hi_hi_3, maskForGroupWire_hi_lo_hi_lo_3};
  wire [31:0]      maskForGroupWire_hi_lo_3 = {maskForGroupWire_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_3 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_3 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_3 = {maskForGroupWire_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_3};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_3 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_3 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_lo_3};
  wire [31:0]      maskForGroupWire_hi_hi_3 = {maskForGroupWire_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_3};
  wire [63:0]      maskForGroupWire_hi_3 = {maskForGroupWire_hi_hi_3, maskForGroupWire_hi_lo_3};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_4 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_4 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_4 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_4 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_4 = {maskForGroupWire_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_hi_lo_4};
  wire [31:0]      maskForGroupWire_lo_lo_4 = {maskForGroupWire_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_4 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_4 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_4 = {maskForGroupWire_lo_hi_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_4 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_4 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_lo_4};
  wire [31:0]      maskForGroupWire_lo_hi_4 = {maskForGroupWire_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_4};
  wire [63:0]      maskForGroupWire_lo_4 = {maskForGroupWire_lo_hi_4, maskForGroupWire_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_4 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_4 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_4 = {maskForGroupWire_hi_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_4 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_4 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_4 = {maskForGroupWire_hi_lo_hi_hi_4, maskForGroupWire_hi_lo_hi_lo_4};
  wire [31:0]      maskForGroupWire_hi_lo_4 = {maskForGroupWire_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_4 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_4 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_4 = {maskForGroupWire_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_4};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_4 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_4 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_lo_4};
  wire [31:0]      maskForGroupWire_hi_hi_4 = {maskForGroupWire_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_4};
  wire [63:0]      maskForGroupWire_hi_4 = {maskForGroupWire_hi_hi_4, maskForGroupWire_hi_lo_4};
  wire [7:0]       maskForGroupWire_lo_lo_lo_lo_5 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]       maskForGroupWire_lo_lo_lo_hi_5 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]      maskForGroupWire_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_lo_hi_lo_5 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]       maskForGroupWire_lo_lo_hi_hi_5 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]      maskForGroupWire_lo_lo_hi_5 = {maskForGroupWire_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_hi_lo_5};
  wire [31:0]      maskForGroupWire_lo_lo_5 = {maskForGroupWire_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_hi_lo_lo_5 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]       maskForGroupWire_lo_hi_lo_hi_5 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]      maskForGroupWire_lo_hi_lo_5 = {maskForGroupWire_lo_hi_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_lo_hi_hi_lo_5 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]       maskForGroupWire_lo_hi_hi_hi_5 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]      maskForGroupWire_lo_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_lo_5};
  wire [31:0]      maskForGroupWire_lo_hi_5 = {maskForGroupWire_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_5};
  wire [63:0]      maskForGroupWire_lo_5 = {maskForGroupWire_lo_hi_5, maskForGroupWire_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_lo_lo_lo_5 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]       maskForGroupWire_hi_lo_lo_hi_5 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]      maskForGroupWire_hi_lo_lo_5 = {maskForGroupWire_hi_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_lo_hi_lo_5 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]       maskForGroupWire_hi_lo_hi_hi_5 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]      maskForGroupWire_hi_lo_hi_5 = {maskForGroupWire_hi_lo_hi_hi_5, maskForGroupWire_hi_lo_hi_lo_5};
  wire [31:0]      maskForGroupWire_hi_lo_5 = {maskForGroupWire_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_hi_lo_lo_5 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]       maskForGroupWire_hi_hi_lo_hi_5 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]      maskForGroupWire_hi_hi_lo_5 = {maskForGroupWire_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_5};
  wire [7:0]       maskForGroupWire_hi_hi_hi_lo_5 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]       maskForGroupWire_hi_hi_hi_hi_5 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]      maskForGroupWire_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_lo_5};
  wire [31:0]      maskForGroupWire_hi_hi_5 = {maskForGroupWire_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_5};
  wire [63:0]      maskForGroupWire_hi_5 = {maskForGroupWire_hi_hi_5, maskForGroupWire_hi_lo_5};
  wire [31:0]      maskForGroupWire =
    (dataEEWOH[0] ? maskWire : 32'h0) | (dataEEWOH[1] ? (maskCounterInGroup[0] ? maskForGroupWire_hi : maskForGroupWire_lo_1) : 32'h0)
    | (dataEEWOH[2]
         ? (_maskForGroupWire_T_133[0] ? maskForGroupWire_lo_2[31:0] : 32'h0) | (_maskForGroupWire_T_133[1] ? maskForGroupWire_lo_3[63:32] : 32'h0) | (_maskForGroupWire_T_133[2] ? maskForGroupWire_hi_4[31:0] : 32'h0)
           | (_maskForGroupWire_T_133[3] ? maskForGroupWire_hi_5[63:32] : 32'h0)
         : 32'h0);
  wire [1:0]       initSendState_lo = maskForGroupWire[1:0];
  wire [1:0]       fillBySeg_lo_lo_lo_lo = maskForGroupWire[1:0];
  wire [1:0]       initSendState_hi = maskForGroupWire[3:2];
  wire [1:0]       fillBySeg_lo_lo_lo_hi = maskForGroupWire[3:2];
  wire             initSendState_0 = |{initSendState_hi, initSendState_lo};
  wire [1:0]       initSendState_lo_1 = maskForGroupWire[5:4];
  wire [1:0]       fillBySeg_lo_lo_hi_lo = maskForGroupWire[5:4];
  wire [1:0]       initSendState_hi_1 = maskForGroupWire[7:6];
  wire [1:0]       fillBySeg_lo_lo_hi_hi = maskForGroupWire[7:6];
  wire             initSendState_1 = |{initSendState_hi_1, initSendState_lo_1};
  wire [1:0]       initSendState_lo_2 = maskForGroupWire[9:8];
  wire [1:0]       fillBySeg_lo_hi_lo_lo = maskForGroupWire[9:8];
  wire [1:0]       initSendState_hi_2 = maskForGroupWire[11:10];
  wire [1:0]       fillBySeg_lo_hi_lo_hi = maskForGroupWire[11:10];
  wire             initSendState_2 = |{initSendState_hi_2, initSendState_lo_2};
  wire [1:0]       initSendState_lo_3 = maskForGroupWire[13:12];
  wire [1:0]       fillBySeg_lo_hi_hi_lo = maskForGroupWire[13:12];
  wire [1:0]       initSendState_hi_3 = maskForGroupWire[15:14];
  wire [1:0]       fillBySeg_lo_hi_hi_hi = maskForGroupWire[15:14];
  wire             initSendState_3 = |{initSendState_hi_3, initSendState_lo_3};
  wire [1:0]       initSendState_lo_4 = maskForGroupWire[17:16];
  wire [1:0]       fillBySeg_hi_lo_lo_lo = maskForGroupWire[17:16];
  wire [1:0]       initSendState_hi_4 = maskForGroupWire[19:18];
  wire [1:0]       fillBySeg_hi_lo_lo_hi = maskForGroupWire[19:18];
  wire             initSendState_4 = |{initSendState_hi_4, initSendState_lo_4};
  wire [1:0]       initSendState_lo_5 = maskForGroupWire[21:20];
  wire [1:0]       fillBySeg_hi_lo_hi_lo = maskForGroupWire[21:20];
  wire [1:0]       initSendState_hi_5 = maskForGroupWire[23:22];
  wire [1:0]       fillBySeg_hi_lo_hi_hi = maskForGroupWire[23:22];
  wire             initSendState_5 = |{initSendState_hi_5, initSendState_lo_5};
  wire [1:0]       initSendState_lo_6 = maskForGroupWire[25:24];
  wire [1:0]       fillBySeg_hi_hi_lo_lo = maskForGroupWire[25:24];
  wire [1:0]       initSendState_hi_6 = maskForGroupWire[27:26];
  wire [1:0]       fillBySeg_hi_hi_lo_hi = maskForGroupWire[27:26];
  wire             initSendState_6 = |{initSendState_hi_6, initSendState_lo_6};
  wire [1:0]       initSendState_lo_7 = maskForGroupWire[29:28];
  wire [1:0]       fillBySeg_hi_hi_hi_lo = maskForGroupWire[29:28];
  wire [1:0]       initSendState_hi_7 = maskForGroupWire[31:30];
  wire [1:0]       fillBySeg_hi_hi_hi_hi = maskForGroupWire[31:30];
  wire             initSendState_7 = |{initSendState_hi_7, initSendState_lo_7};
  reg  [255:0]     accessData_0;
  wire [255:0]     accessDataUpdate_1 = accessData_0;
  reg  [255:0]     accessData_1;
  wire [255:0]     accessDataUpdate_2 = accessData_1;
  reg  [255:0]     accessData_2;
  wire [255:0]     accessDataUpdate_3 = accessData_2;
  reg  [255:0]     accessData_3;
  wire [255:0]     accessDataUpdate_4 = accessData_3;
  reg  [255:0]     accessData_4;
  wire [255:0]     accessDataUpdate_5 = accessData_4;
  reg  [255:0]     accessData_5;
  wire [255:0]     accessDataUpdate_6 = accessData_5;
  reg  [255:0]     accessData_6;
  wire [255:0]     accessDataUpdate_7 = accessData_6;
  reg  [255:0]     accessData_7;
  reg  [2:0]       accessPtr;
  reg  [5:0]       dataGroup;
  reg  [255:0]     dataBuffer_0;
  reg  [255:0]     dataBuffer_1;
  reg  [255:0]     dataBuffer_2;
  reg  [255:0]     dataBuffer_3;
  reg  [255:0]     dataBuffer_4;
  reg  [255:0]     dataBuffer_5;
  reg  [255:0]     dataBuffer_6;
  reg  [255:0]     dataBuffer_7;
  reg  [6:0]       bufferBaseCacheLineIndex;
  wire [6:0]       memRequest_bits_index_0 = bufferBaseCacheLineIndex;
  reg  [2:0]       cacheLineIndexInBuffer;
  wire [4:0]       initOffset = lsuRequestReg_rs1Data[4:0];
  wire             invalidInstruction = csrInterface_vl == 12'h0;
  reg              invalidInstructionNext;
  wire             wholeType = lsuRequest_bits_instructionInformation_lumop[3];
  wire [2:0]       nfCorrection = wholeType ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [3:0]       segmentInstructionIndexInterval;
  wire [18:0]      bytePerInstruction = {3'h0, {12'h0, {1'h0, nfCorrection} + 4'h1} * {4'h0, csrInterface_vl}} << lsuRequest_bits_instructionInformation_eew;
  wire [18:0]      accessMemSize = bytePerInstruction + {14'h0, lsuRequest_bits_rs1Data[4:0]};
  wire [13:0]      lastCacheLineIndex = accessMemSize[18:5] - {13'h0, accessMemSize[4:0] == 5'h0};
  wire [13:0]      lastWriteVrfIndex = bytePerInstruction[18:5] - {13'h0, bytePerInstruction[4:0] == 5'h0};
  reg  [13:0]      lastWriteVrfIndexReg;
  reg              lastCacheNeedPush;
  reg  [13:0]      cacheLineNumberReg;
  wire [14:0]      dataByteSize = {3'h0, csrInterface_vl} << lsuRequest_bits_instructionInformation_eew;
  wire [9:0]       lastDataGroupForInstruction = dataByteSize[14:5] - {9'h0, dataByteSize[4:0] == 5'h0};
  reg  [9:0]       lastDataGroupReg;
  wire [5:0]       nextDataGroup = lsuRequest_valid ? 6'h0 : dataGroup + 6'h1;
  wire             isLastRead = {4'h0, dataGroup} == lastDataGroupReg;
  reg              hazardCheck;
  wire             accessBufferEnqueueFire;
  wire             vrfReadQueueVec_0_deq_ready;
  wire             vrfReadQueueVec_0_enq_ready = ~_vrfReadQueueVec_fifo_full | vrfReadQueueVec_0_deq_ready;
  wire             vrfReadQueueVec_0_deq_valid = ~_vrfReadQueueVec_fifo_empty | vrfReadQueueVec_0_enq_valid;
  wire [31:0]      vrfReadQueueVec_0_deq_bits = _vrfReadQueueVec_fifo_empty ? vrfReadQueueVec_0_enq_bits : _vrfReadQueueVec_fifo_data_out;
  wire             vrfReadQueueVec_1_deq_ready;
  wire             vrfReadQueueVec_1_enq_ready = ~_vrfReadQueueVec_fifo_1_full | vrfReadQueueVec_1_deq_ready;
  wire             vrfReadQueueVec_1_deq_valid = ~_vrfReadQueueVec_fifo_1_empty | vrfReadQueueVec_1_enq_valid;
  wire [31:0]      vrfReadQueueVec_1_deq_bits = _vrfReadQueueVec_fifo_1_empty ? vrfReadQueueVec_1_enq_bits : _vrfReadQueueVec_fifo_1_data_out;
  wire             vrfReadQueueVec_2_deq_ready;
  wire             vrfReadQueueVec_2_enq_ready = ~_vrfReadQueueVec_fifo_2_full | vrfReadQueueVec_2_deq_ready;
  wire             vrfReadQueueVec_2_deq_valid = ~_vrfReadQueueVec_fifo_2_empty | vrfReadQueueVec_2_enq_valid;
  wire [31:0]      vrfReadQueueVec_2_deq_bits = _vrfReadQueueVec_fifo_2_empty ? vrfReadQueueVec_2_enq_bits : _vrfReadQueueVec_fifo_2_data_out;
  wire             vrfReadQueueVec_3_deq_ready;
  wire             vrfReadQueueVec_3_enq_ready = ~_vrfReadQueueVec_fifo_3_full | vrfReadQueueVec_3_deq_ready;
  wire             vrfReadQueueVec_3_deq_valid = ~_vrfReadQueueVec_fifo_3_empty | vrfReadQueueVec_3_enq_valid;
  wire [31:0]      vrfReadQueueVec_3_deq_bits = _vrfReadQueueVec_fifo_3_empty ? vrfReadQueueVec_3_enq_bits : _vrfReadQueueVec_fifo_3_data_out;
  wire             vrfReadQueueVec_4_deq_ready;
  wire             vrfReadQueueVec_4_enq_ready = ~_vrfReadQueueVec_fifo_4_full | vrfReadQueueVec_4_deq_ready;
  wire             vrfReadQueueVec_4_deq_valid = ~_vrfReadQueueVec_fifo_4_empty | vrfReadQueueVec_4_enq_valid;
  wire [31:0]      vrfReadQueueVec_4_deq_bits = _vrfReadQueueVec_fifo_4_empty ? vrfReadQueueVec_4_enq_bits : _vrfReadQueueVec_fifo_4_data_out;
  wire             vrfReadQueueVec_5_deq_ready;
  wire             vrfReadQueueVec_5_enq_ready = ~_vrfReadQueueVec_fifo_5_full | vrfReadQueueVec_5_deq_ready;
  wire             vrfReadQueueVec_5_deq_valid = ~_vrfReadQueueVec_fifo_5_empty | vrfReadQueueVec_5_enq_valid;
  wire [31:0]      vrfReadQueueVec_5_deq_bits = _vrfReadQueueVec_fifo_5_empty ? vrfReadQueueVec_5_enq_bits : _vrfReadQueueVec_fifo_5_data_out;
  wire             vrfReadQueueVec_6_deq_ready;
  wire             vrfReadQueueVec_6_enq_ready = ~_vrfReadQueueVec_fifo_6_full | vrfReadQueueVec_6_deq_ready;
  wire             vrfReadQueueVec_6_deq_valid = ~_vrfReadQueueVec_fifo_6_empty | vrfReadQueueVec_6_enq_valid;
  wire [31:0]      vrfReadQueueVec_6_deq_bits = _vrfReadQueueVec_fifo_6_empty ? vrfReadQueueVec_6_enq_bits : _vrfReadQueueVec_fifo_6_data_out;
  wire             vrfReadQueueVec_7_deq_ready;
  wire             vrfReadQueueVec_7_enq_ready = ~_vrfReadQueueVec_fifo_7_full | vrfReadQueueVec_7_deq_ready;
  wire             vrfReadQueueVec_7_deq_valid = ~_vrfReadQueueVec_fifo_7_empty | vrfReadQueueVec_7_enq_valid;
  wire [31:0]      vrfReadQueueVec_7_deq_bits = _vrfReadQueueVec_fifo_7_empty ? vrfReadQueueVec_7_enq_bits : _vrfReadQueueVec_fifo_7_data_out;
  reg  [2:0]       readStageValid_segPtr;
  reg  [5:0]       readStageValid_readCount;
  reg              readStageValid_stageValid;
  wire             readStageValid_lastReadPtr = readStageValid_segPtr == 3'h0;
  wire [5:0]       readStageValid_nextReadCount = lsuRequest_valid ? 6'h0 : readStageValid_readCount + 6'h1;
  wire             readStageValid_lastReadGroup = {4'h0, readStageValid_readCount} == lastDataGroupReg;
  wire             vrfReadDataPorts_0_valid_0;
  wire             _readStageValid_T_11 = vrfReadDataPorts_0_ready_0 & vrfReadDataPorts_0_valid_0;
  reg  [3:0]       readStageValid_readCounter;
  wire [3:0]       readStageValid_counterChange = _readStageValid_T_11 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_0_valid_0 = readStageValid_stageValid & ~(readStageValid_readCounter[3]);
  wire [4:0]       _GEN_3 = {1'h0, segmentInstructionIndexInterval};
  wire [4:0]       vrfReadDataPorts_0_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr} * _GEN_3 + {2'h0, readStageValid_readCount[5:3]};
  wire [2:0]       vrfReadDataPorts_0_bits_offset_0 = readStageValid_readCount[2:0];
  reg  [2:0]       readStageValid_segPtr_1;
  reg  [5:0]       readStageValid_readCount_1;
  reg              readStageValid_stageValid_1;
  wire             readStageValid_lastReadPtr_1 = readStageValid_segPtr_1 == 3'h0;
  wire [5:0]       readStageValid_nextReadCount_1 = lsuRequest_valid ? 6'h0 : readStageValid_readCount_1 + 6'h1;
  wire             readStageValid_lastReadGroup_1 = {4'h0, readStageValid_readCount_1} == lastDataGroupReg;
  wire             vrfReadDataPorts_1_valid_0;
  wire             _readStageValid_T_30 = vrfReadDataPorts_1_ready_0 & vrfReadDataPorts_1_valid_0;
  reg  [3:0]       readStageValid_readCounter_1;
  wire [3:0]       readStageValid_counterChange_1 = _readStageValid_T_30 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_1_valid_0 = readStageValid_stageValid_1 & ~(readStageValid_readCounter_1[3]);
  wire [4:0]       vrfReadDataPorts_1_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_1} * _GEN_3 + {2'h0, readStageValid_readCount_1[5:3]};
  wire [2:0]       vrfReadDataPorts_1_bits_offset_0 = readStageValid_readCount_1[2:0];
  reg  [2:0]       readStageValid_segPtr_2;
  reg  [5:0]       readStageValid_readCount_2;
  reg              readStageValid_stageValid_2;
  wire             readStageValid_lastReadPtr_2 = readStageValid_segPtr_2 == 3'h0;
  wire [5:0]       readStageValid_nextReadCount_2 = lsuRequest_valid ? 6'h0 : readStageValid_readCount_2 + 6'h1;
  wire             readStageValid_lastReadGroup_2 = {4'h0, readStageValid_readCount_2} == lastDataGroupReg;
  wire             vrfReadDataPorts_2_valid_0;
  wire             _readStageValid_T_49 = vrfReadDataPorts_2_ready_0 & vrfReadDataPorts_2_valid_0;
  reg  [3:0]       readStageValid_readCounter_2;
  wire [3:0]       readStageValid_counterChange_2 = _readStageValid_T_49 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_2_valid_0 = readStageValid_stageValid_2 & ~(readStageValid_readCounter_2[3]);
  wire [4:0]       vrfReadDataPorts_2_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_2} * _GEN_3 + {2'h0, readStageValid_readCount_2[5:3]};
  wire [2:0]       vrfReadDataPorts_2_bits_offset_0 = readStageValid_readCount_2[2:0];
  reg  [2:0]       readStageValid_segPtr_3;
  reg  [5:0]       readStageValid_readCount_3;
  reg              readStageValid_stageValid_3;
  wire             readStageValid_lastReadPtr_3 = readStageValid_segPtr_3 == 3'h0;
  wire [5:0]       readStageValid_nextReadCount_3 = lsuRequest_valid ? 6'h0 : readStageValid_readCount_3 + 6'h1;
  wire             readStageValid_lastReadGroup_3 = {4'h0, readStageValid_readCount_3} == lastDataGroupReg;
  wire             vrfReadDataPorts_3_valid_0;
  wire             _readStageValid_T_68 = vrfReadDataPorts_3_ready_0 & vrfReadDataPorts_3_valid_0;
  reg  [3:0]       readStageValid_readCounter_3;
  wire [3:0]       readStageValid_counterChange_3 = _readStageValid_T_68 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_3_valid_0 = readStageValid_stageValid_3 & ~(readStageValid_readCounter_3[3]);
  wire [4:0]       vrfReadDataPorts_3_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_3} * _GEN_3 + {2'h0, readStageValid_readCount_3[5:3]};
  wire [2:0]       vrfReadDataPorts_3_bits_offset_0 = readStageValid_readCount_3[2:0];
  reg  [2:0]       readStageValid_segPtr_4;
  reg  [5:0]       readStageValid_readCount_4;
  reg              readStageValid_stageValid_4;
  wire             readStageValid_lastReadPtr_4 = readStageValid_segPtr_4 == 3'h0;
  wire [5:0]       readStageValid_nextReadCount_4 = lsuRequest_valid ? 6'h0 : readStageValid_readCount_4 + 6'h1;
  wire             readStageValid_lastReadGroup_4 = {4'h0, readStageValid_readCount_4} == lastDataGroupReg;
  wire             vrfReadDataPorts_4_valid_0;
  wire             _readStageValid_T_87 = vrfReadDataPorts_4_ready_0 & vrfReadDataPorts_4_valid_0;
  reg  [3:0]       readStageValid_readCounter_4;
  wire [3:0]       readStageValid_counterChange_4 = _readStageValid_T_87 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_4_valid_0 = readStageValid_stageValid_4 & ~(readStageValid_readCounter_4[3]);
  wire [4:0]       vrfReadDataPorts_4_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_4} * _GEN_3 + {2'h0, readStageValid_readCount_4[5:3]};
  wire [2:0]       vrfReadDataPorts_4_bits_offset_0 = readStageValid_readCount_4[2:0];
  reg  [2:0]       readStageValid_segPtr_5;
  reg  [5:0]       readStageValid_readCount_5;
  reg              readStageValid_stageValid_5;
  wire             readStageValid_lastReadPtr_5 = readStageValid_segPtr_5 == 3'h0;
  wire [5:0]       readStageValid_nextReadCount_5 = lsuRequest_valid ? 6'h0 : readStageValid_readCount_5 + 6'h1;
  wire             readStageValid_lastReadGroup_5 = {4'h0, readStageValid_readCount_5} == lastDataGroupReg;
  wire             vrfReadDataPorts_5_valid_0;
  wire             _readStageValid_T_106 = vrfReadDataPorts_5_ready_0 & vrfReadDataPorts_5_valid_0;
  reg  [3:0]       readStageValid_readCounter_5;
  wire [3:0]       readStageValid_counterChange_5 = _readStageValid_T_106 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_5_valid_0 = readStageValid_stageValid_5 & ~(readStageValid_readCounter_5[3]);
  wire [4:0]       vrfReadDataPorts_5_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_5} * _GEN_3 + {2'h0, readStageValid_readCount_5[5:3]};
  wire [2:0]       vrfReadDataPorts_5_bits_offset_0 = readStageValid_readCount_5[2:0];
  reg  [2:0]       readStageValid_segPtr_6;
  reg  [5:0]       readStageValid_readCount_6;
  reg              readStageValid_stageValid_6;
  wire             readStageValid_lastReadPtr_6 = readStageValid_segPtr_6 == 3'h0;
  wire [5:0]       readStageValid_nextReadCount_6 = lsuRequest_valid ? 6'h0 : readStageValid_readCount_6 + 6'h1;
  wire             readStageValid_lastReadGroup_6 = {4'h0, readStageValid_readCount_6} == lastDataGroupReg;
  wire             vrfReadDataPorts_6_valid_0;
  wire             _readStageValid_T_125 = vrfReadDataPorts_6_ready_0 & vrfReadDataPorts_6_valid_0;
  reg  [3:0]       readStageValid_readCounter_6;
  wire [3:0]       readStageValid_counterChange_6 = _readStageValid_T_125 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_6_valid_0 = readStageValid_stageValid_6 & ~(readStageValid_readCounter_6[3]);
  wire [4:0]       vrfReadDataPorts_6_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_6} * _GEN_3 + {2'h0, readStageValid_readCount_6[5:3]};
  wire [2:0]       vrfReadDataPorts_6_bits_offset_0 = readStageValid_readCount_6[2:0];
  reg  [2:0]       readStageValid_segPtr_7;
  reg  [5:0]       readStageValid_readCount_7;
  reg              readStageValid_stageValid_7;
  wire             readStageValid_lastReadPtr_7 = readStageValid_segPtr_7 == 3'h0;
  wire [5:0]       readStageValid_nextReadCount_7 = lsuRequest_valid ? 6'h0 : readStageValid_readCount_7 + 6'h1;
  wire             readStageValid_lastReadGroup_7 = {4'h0, readStageValid_readCount_7} == lastDataGroupReg;
  wire             vrfReadDataPorts_7_valid_0;
  wire             _readStageValid_T_144 = vrfReadDataPorts_7_ready_0 & vrfReadDataPorts_7_valid_0;
  reg  [3:0]       readStageValid_readCounter_7;
  wire [3:0]       readStageValid_counterChange_7 = _readStageValid_T_144 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_7_valid_0 = readStageValid_stageValid_7 & ~(readStageValid_readCounter_7[3]);
  wire [4:0]       vrfReadDataPorts_7_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_7} * _GEN_3 + {2'h0, readStageValid_readCount_7[5:3]};
  wire [2:0]       vrfReadDataPorts_7_bits_offset_0 = readStageValid_readCount_7[2:0];
  wire             readStageValid =
    |{readStageValid_stageValid,
      readStageValid_readCounter,
      readStageValid_stageValid_1,
      readStageValid_readCounter_1,
      readStageValid_stageValid_2,
      readStageValid_readCounter_2,
      readStageValid_stageValid_3,
      readStageValid_readCounter_3,
      readStageValid_stageValid_4,
      readStageValid_readCounter_4,
      readStageValid_stageValid_5,
      readStageValid_readCounter_5,
      readStageValid_stageValid_6,
      readStageValid_readCounter_6,
      readStageValid_stageValid_7,
      readStageValid_readCounter_7};
  reg              bufferFull;
  wire             accessBufferDequeueReady;
  wire             accessBufferEnqueueReady = ~bufferFull | accessBufferDequeueReady;
  wire             accessBufferEnqueueValid =
    vrfReadQueueVec_0_deq_valid & vrfReadQueueVec_1_deq_valid & vrfReadQueueVec_2_deq_valid & vrfReadQueueVec_3_deq_valid & vrfReadQueueVec_4_deq_valid & vrfReadQueueVec_5_deq_valid & vrfReadQueueVec_6_deq_valid
    & vrfReadQueueVec_7_deq_valid;
  wire             readQueueClear =
    ~(vrfReadQueueVec_0_deq_valid | vrfReadQueueVec_1_deq_valid | vrfReadQueueVec_2_deq_valid | vrfReadQueueVec_3_deq_valid | vrfReadQueueVec_4_deq_valid | vrfReadQueueVec_5_deq_valid | vrfReadQueueVec_6_deq_valid
      | vrfReadQueueVec_7_deq_valid);
  assign accessBufferEnqueueFire = accessBufferEnqueueValid & accessBufferEnqueueReady;
  assign vrfReadQueueVec_0_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_1_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_2_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_3_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_4_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_5_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_6_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_7_deq_ready = accessBufferEnqueueFire;
  wire             lastPtr = accessPtr == 3'h0;
  wire             lastPtrEnq = lastPtr & accessBufferEnqueueFire;
  wire             accessBufferDequeueValid = bufferFull | lastPtrEnq;
  wire             accessBufferDequeueFire = accessBufferDequeueValid & accessBufferDequeueReady;
  wire [63:0]      accessDataUpdate_lo_lo = {vrfReadQueueVec_1_deq_bits, vrfReadQueueVec_0_deq_bits};
  wire [63:0]      accessDataUpdate_lo_hi = {vrfReadQueueVec_3_deq_bits, vrfReadQueueVec_2_deq_bits};
  wire [127:0]     accessDataUpdate_lo = {accessDataUpdate_lo_hi, accessDataUpdate_lo_lo};
  wire [63:0]      accessDataUpdate_hi_lo = {vrfReadQueueVec_5_deq_bits, vrfReadQueueVec_4_deq_bits};
  wire [63:0]      accessDataUpdate_hi_hi = {vrfReadQueueVec_7_deq_bits, vrfReadQueueVec_6_deq_bits};
  wire [127:0]     accessDataUpdate_hi = {accessDataUpdate_hi_hi, accessDataUpdate_hi_lo};
  wire [255:0]     accessDataUpdate_0 = {accessDataUpdate_hi, accessDataUpdate_lo};
  reg              bufferValid;
  reg  [31:0]      maskForBufferData_0;
  reg  [31:0]      maskForBufferData_1;
  reg  [31:0]      maskForBufferData_2;
  reg  [31:0]      maskForBufferData_3;
  reg  [31:0]      maskForBufferData_4;
  reg  [31:0]      maskForBufferData_5;
  reg  [31:0]      maskForBufferData_6;
  reg  [31:0]      maskForBufferData_7;
  reg              lastDataGroupInDataBuffer;
  wire             memRequest_valid_0;
  wire             _addressQueue_enq_valid_T = memRequest_ready_0 & memRequest_valid_0;
  wire             alignedDequeueFire;
  assign alignedDequeueFire = _addressQueue_enq_valid_T;
  wire             addressQueue_enq_valid;
  assign addressQueue_enq_valid = _addressQueue_enq_valid_T;
  reg  [255:0]     cacheLineTemp;
  reg  [31:0]      maskTemp;
  reg              canSendTail;
  wire             isLastCacheLineInBuffer = cacheLineIndexInBuffer == lsuRequestReg_instructionInformation_nf;
  wire             bufferWillClear = alignedDequeueFire & isLastCacheLineInBuffer;
  wire             addressQueue_enq_ready;
  wire             addressQueueFree;
  assign accessBufferDequeueReady = ~bufferValid | memRequest_ready_0 & isLastCacheLineInBuffer & addressQueueFree;
  wire [255:0]     bufferStageEnqueueData_0 = bufferFull ? accessData_0 : accessDataUpdate_0;
  wire [255:0]     bufferStageEnqueueData_1 = bufferFull ? accessData_1 : accessDataUpdate_1;
  wire [255:0]     bufferStageEnqueueData_2 = bufferFull ? accessData_2 : accessDataUpdate_2;
  wire [255:0]     bufferStageEnqueueData_3 = bufferFull ? accessData_3 : accessDataUpdate_3;
  wire [255:0]     bufferStageEnqueueData_4 = bufferFull ? accessData_4 : accessDataUpdate_4;
  wire [255:0]     bufferStageEnqueueData_5 = bufferFull ? accessData_5 : accessDataUpdate_5;
  wire [255:0]     bufferStageEnqueueData_6 = bufferFull ? accessData_6 : accessDataUpdate_6;
  wire [255:0]     bufferStageEnqueueData_7 = bufferFull ? accessData_7 : accessDataUpdate_7;
  wire [7:0]       _fillBySeg_T = 8'h1 << lsuRequestReg_instructionInformation_nf;
  wire [3:0]       fillBySeg_lo_lo_lo = {fillBySeg_lo_lo_lo_hi, fillBySeg_lo_lo_lo_lo};
  wire [3:0]       fillBySeg_lo_lo_hi = {fillBySeg_lo_lo_hi_hi, fillBySeg_lo_lo_hi_lo};
  wire [7:0]       fillBySeg_lo_lo = {fillBySeg_lo_lo_hi, fillBySeg_lo_lo_lo};
  wire [3:0]       fillBySeg_lo_hi_lo = {fillBySeg_lo_hi_lo_hi, fillBySeg_lo_hi_lo_lo};
  wire [3:0]       fillBySeg_lo_hi_hi = {fillBySeg_lo_hi_hi_hi, fillBySeg_lo_hi_hi_lo};
  wire [7:0]       fillBySeg_lo_hi = {fillBySeg_lo_hi_hi, fillBySeg_lo_hi_lo};
  wire [15:0]      fillBySeg_lo = {fillBySeg_lo_hi, fillBySeg_lo_lo};
  wire [3:0]       fillBySeg_hi_lo_lo = {fillBySeg_hi_lo_lo_hi, fillBySeg_hi_lo_lo_lo};
  wire [3:0]       fillBySeg_hi_lo_hi = {fillBySeg_hi_lo_hi_hi, fillBySeg_hi_lo_hi_lo};
  wire [7:0]       fillBySeg_hi_lo = {fillBySeg_hi_lo_hi, fillBySeg_hi_lo_lo};
  wire [3:0]       fillBySeg_hi_hi_lo = {fillBySeg_hi_hi_lo_hi, fillBySeg_hi_hi_lo_lo};
  wire [3:0]       fillBySeg_hi_hi_hi = {fillBySeg_hi_hi_hi_hi, fillBySeg_hi_hi_hi_lo};
  wire [7:0]       fillBySeg_hi_hi = {fillBySeg_hi_hi_hi, fillBySeg_hi_hi_lo};
  wire [15:0]      fillBySeg_hi = {fillBySeg_hi_hi, fillBySeg_hi_lo};
  wire [3:0]       fillBySeg_lo_lo_lo_lo_1 = {{2{maskForGroupWire[1]}}, {2{maskForGroupWire[0]}}};
  wire [3:0]       fillBySeg_lo_lo_lo_hi_1 = {{2{maskForGroupWire[3]}}, {2{maskForGroupWire[2]}}};
  wire [7:0]       fillBySeg_lo_lo_lo_1 = {fillBySeg_lo_lo_lo_hi_1, fillBySeg_lo_lo_lo_lo_1};
  wire [3:0]       fillBySeg_lo_lo_hi_lo_1 = {{2{maskForGroupWire[5]}}, {2{maskForGroupWire[4]}}};
  wire [3:0]       fillBySeg_lo_lo_hi_hi_1 = {{2{maskForGroupWire[7]}}, {2{maskForGroupWire[6]}}};
  wire [7:0]       fillBySeg_lo_lo_hi_1 = {fillBySeg_lo_lo_hi_hi_1, fillBySeg_lo_lo_hi_lo_1};
  wire [15:0]      fillBySeg_lo_lo_1 = {fillBySeg_lo_lo_hi_1, fillBySeg_lo_lo_lo_1};
  wire [3:0]       fillBySeg_lo_hi_lo_lo_1 = {{2{maskForGroupWire[9]}}, {2{maskForGroupWire[8]}}};
  wire [3:0]       fillBySeg_lo_hi_lo_hi_1 = {{2{maskForGroupWire[11]}}, {2{maskForGroupWire[10]}}};
  wire [7:0]       fillBySeg_lo_hi_lo_1 = {fillBySeg_lo_hi_lo_hi_1, fillBySeg_lo_hi_lo_lo_1};
  wire [3:0]       fillBySeg_lo_hi_hi_lo_1 = {{2{maskForGroupWire[13]}}, {2{maskForGroupWire[12]}}};
  wire [3:0]       fillBySeg_lo_hi_hi_hi_1 = {{2{maskForGroupWire[15]}}, {2{maskForGroupWire[14]}}};
  wire [7:0]       fillBySeg_lo_hi_hi_1 = {fillBySeg_lo_hi_hi_hi_1, fillBySeg_lo_hi_hi_lo_1};
  wire [15:0]      fillBySeg_lo_hi_1 = {fillBySeg_lo_hi_hi_1, fillBySeg_lo_hi_lo_1};
  wire [31:0]      fillBySeg_lo_1 = {fillBySeg_lo_hi_1, fillBySeg_lo_lo_1};
  wire [3:0]       fillBySeg_hi_lo_lo_lo_1 = {{2{maskForGroupWire[17]}}, {2{maskForGroupWire[16]}}};
  wire [3:0]       fillBySeg_hi_lo_lo_hi_1 = {{2{maskForGroupWire[19]}}, {2{maskForGroupWire[18]}}};
  wire [7:0]       fillBySeg_hi_lo_lo_1 = {fillBySeg_hi_lo_lo_hi_1, fillBySeg_hi_lo_lo_lo_1};
  wire [3:0]       fillBySeg_hi_lo_hi_lo_1 = {{2{maskForGroupWire[21]}}, {2{maskForGroupWire[20]}}};
  wire [3:0]       fillBySeg_hi_lo_hi_hi_1 = {{2{maskForGroupWire[23]}}, {2{maskForGroupWire[22]}}};
  wire [7:0]       fillBySeg_hi_lo_hi_1 = {fillBySeg_hi_lo_hi_hi_1, fillBySeg_hi_lo_hi_lo_1};
  wire [15:0]      fillBySeg_hi_lo_1 = {fillBySeg_hi_lo_hi_1, fillBySeg_hi_lo_lo_1};
  wire [3:0]       fillBySeg_hi_hi_lo_lo_1 = {{2{maskForGroupWire[25]}}, {2{maskForGroupWire[24]}}};
  wire [3:0]       fillBySeg_hi_hi_lo_hi_1 = {{2{maskForGroupWire[27]}}, {2{maskForGroupWire[26]}}};
  wire [7:0]       fillBySeg_hi_hi_lo_1 = {fillBySeg_hi_hi_lo_hi_1, fillBySeg_hi_hi_lo_lo_1};
  wire [3:0]       fillBySeg_hi_hi_hi_lo_1 = {{2{maskForGroupWire[29]}}, {2{maskForGroupWire[28]}}};
  wire [3:0]       fillBySeg_hi_hi_hi_hi_1 = {{2{maskForGroupWire[31]}}, {2{maskForGroupWire[30]}}};
  wire [7:0]       fillBySeg_hi_hi_hi_1 = {fillBySeg_hi_hi_hi_hi_1, fillBySeg_hi_hi_hi_lo_1};
  wire [15:0]      fillBySeg_hi_hi_1 = {fillBySeg_hi_hi_hi_1, fillBySeg_hi_hi_lo_1};
  wire [31:0]      fillBySeg_hi_1 = {fillBySeg_hi_hi_1, fillBySeg_hi_lo_1};
  wire [5:0]       fillBySeg_lo_lo_lo_lo_2 = {{3{maskForGroupWire[1]}}, {3{maskForGroupWire[0]}}};
  wire [5:0]       fillBySeg_lo_lo_lo_hi_2 = {{3{maskForGroupWire[3]}}, {3{maskForGroupWire[2]}}};
  wire [11:0]      fillBySeg_lo_lo_lo_2 = {fillBySeg_lo_lo_lo_hi_2, fillBySeg_lo_lo_lo_lo_2};
  wire [5:0]       fillBySeg_lo_lo_hi_lo_2 = {{3{maskForGroupWire[5]}}, {3{maskForGroupWire[4]}}};
  wire [5:0]       fillBySeg_lo_lo_hi_hi_2 = {{3{maskForGroupWire[7]}}, {3{maskForGroupWire[6]}}};
  wire [11:0]      fillBySeg_lo_lo_hi_2 = {fillBySeg_lo_lo_hi_hi_2, fillBySeg_lo_lo_hi_lo_2};
  wire [23:0]      fillBySeg_lo_lo_2 = {fillBySeg_lo_lo_hi_2, fillBySeg_lo_lo_lo_2};
  wire [5:0]       fillBySeg_lo_hi_lo_lo_2 = {{3{maskForGroupWire[9]}}, {3{maskForGroupWire[8]}}};
  wire [5:0]       fillBySeg_lo_hi_lo_hi_2 = {{3{maskForGroupWire[11]}}, {3{maskForGroupWire[10]}}};
  wire [11:0]      fillBySeg_lo_hi_lo_2 = {fillBySeg_lo_hi_lo_hi_2, fillBySeg_lo_hi_lo_lo_2};
  wire [5:0]       fillBySeg_lo_hi_hi_lo_2 = {{3{maskForGroupWire[13]}}, {3{maskForGroupWire[12]}}};
  wire [5:0]       fillBySeg_lo_hi_hi_hi_2 = {{3{maskForGroupWire[15]}}, {3{maskForGroupWire[14]}}};
  wire [11:0]      fillBySeg_lo_hi_hi_2 = {fillBySeg_lo_hi_hi_hi_2, fillBySeg_lo_hi_hi_lo_2};
  wire [23:0]      fillBySeg_lo_hi_2 = {fillBySeg_lo_hi_hi_2, fillBySeg_lo_hi_lo_2};
  wire [47:0]      fillBySeg_lo_2 = {fillBySeg_lo_hi_2, fillBySeg_lo_lo_2};
  wire [5:0]       fillBySeg_hi_lo_lo_lo_2 = {{3{maskForGroupWire[17]}}, {3{maskForGroupWire[16]}}};
  wire [5:0]       fillBySeg_hi_lo_lo_hi_2 = {{3{maskForGroupWire[19]}}, {3{maskForGroupWire[18]}}};
  wire [11:0]      fillBySeg_hi_lo_lo_2 = {fillBySeg_hi_lo_lo_hi_2, fillBySeg_hi_lo_lo_lo_2};
  wire [5:0]       fillBySeg_hi_lo_hi_lo_2 = {{3{maskForGroupWire[21]}}, {3{maskForGroupWire[20]}}};
  wire [5:0]       fillBySeg_hi_lo_hi_hi_2 = {{3{maskForGroupWire[23]}}, {3{maskForGroupWire[22]}}};
  wire [11:0]      fillBySeg_hi_lo_hi_2 = {fillBySeg_hi_lo_hi_hi_2, fillBySeg_hi_lo_hi_lo_2};
  wire [23:0]      fillBySeg_hi_lo_2 = {fillBySeg_hi_lo_hi_2, fillBySeg_hi_lo_lo_2};
  wire [5:0]       fillBySeg_hi_hi_lo_lo_2 = {{3{maskForGroupWire[25]}}, {3{maskForGroupWire[24]}}};
  wire [5:0]       fillBySeg_hi_hi_lo_hi_2 = {{3{maskForGroupWire[27]}}, {3{maskForGroupWire[26]}}};
  wire [11:0]      fillBySeg_hi_hi_lo_2 = {fillBySeg_hi_hi_lo_hi_2, fillBySeg_hi_hi_lo_lo_2};
  wire [5:0]       fillBySeg_hi_hi_hi_lo_2 = {{3{maskForGroupWire[29]}}, {3{maskForGroupWire[28]}}};
  wire [5:0]       fillBySeg_hi_hi_hi_hi_2 = {{3{maskForGroupWire[31]}}, {3{maskForGroupWire[30]}}};
  wire [11:0]      fillBySeg_hi_hi_hi_2 = {fillBySeg_hi_hi_hi_hi_2, fillBySeg_hi_hi_hi_lo_2};
  wire [23:0]      fillBySeg_hi_hi_2 = {fillBySeg_hi_hi_hi_2, fillBySeg_hi_hi_lo_2};
  wire [47:0]      fillBySeg_hi_2 = {fillBySeg_hi_hi_2, fillBySeg_hi_lo_2};
  wire [7:0]       fillBySeg_lo_lo_lo_lo_3 = {{4{maskForGroupWire[1]}}, {4{maskForGroupWire[0]}}};
  wire [7:0]       fillBySeg_lo_lo_lo_hi_3 = {{4{maskForGroupWire[3]}}, {4{maskForGroupWire[2]}}};
  wire [15:0]      fillBySeg_lo_lo_lo_3 = {fillBySeg_lo_lo_lo_hi_3, fillBySeg_lo_lo_lo_lo_3};
  wire [7:0]       fillBySeg_lo_lo_hi_lo_3 = {{4{maskForGroupWire[5]}}, {4{maskForGroupWire[4]}}};
  wire [7:0]       fillBySeg_lo_lo_hi_hi_3 = {{4{maskForGroupWire[7]}}, {4{maskForGroupWire[6]}}};
  wire [15:0]      fillBySeg_lo_lo_hi_3 = {fillBySeg_lo_lo_hi_hi_3, fillBySeg_lo_lo_hi_lo_3};
  wire [31:0]      fillBySeg_lo_lo_3 = {fillBySeg_lo_lo_hi_3, fillBySeg_lo_lo_lo_3};
  wire [7:0]       fillBySeg_lo_hi_lo_lo_3 = {{4{maskForGroupWire[9]}}, {4{maskForGroupWire[8]}}};
  wire [7:0]       fillBySeg_lo_hi_lo_hi_3 = {{4{maskForGroupWire[11]}}, {4{maskForGroupWire[10]}}};
  wire [15:0]      fillBySeg_lo_hi_lo_3 = {fillBySeg_lo_hi_lo_hi_3, fillBySeg_lo_hi_lo_lo_3};
  wire [7:0]       fillBySeg_lo_hi_hi_lo_3 = {{4{maskForGroupWire[13]}}, {4{maskForGroupWire[12]}}};
  wire [7:0]       fillBySeg_lo_hi_hi_hi_3 = {{4{maskForGroupWire[15]}}, {4{maskForGroupWire[14]}}};
  wire [15:0]      fillBySeg_lo_hi_hi_3 = {fillBySeg_lo_hi_hi_hi_3, fillBySeg_lo_hi_hi_lo_3};
  wire [31:0]      fillBySeg_lo_hi_3 = {fillBySeg_lo_hi_hi_3, fillBySeg_lo_hi_lo_3};
  wire [63:0]      fillBySeg_lo_3 = {fillBySeg_lo_hi_3, fillBySeg_lo_lo_3};
  wire [7:0]       fillBySeg_hi_lo_lo_lo_3 = {{4{maskForGroupWire[17]}}, {4{maskForGroupWire[16]}}};
  wire [7:0]       fillBySeg_hi_lo_lo_hi_3 = {{4{maskForGroupWire[19]}}, {4{maskForGroupWire[18]}}};
  wire [15:0]      fillBySeg_hi_lo_lo_3 = {fillBySeg_hi_lo_lo_hi_3, fillBySeg_hi_lo_lo_lo_3};
  wire [7:0]       fillBySeg_hi_lo_hi_lo_3 = {{4{maskForGroupWire[21]}}, {4{maskForGroupWire[20]}}};
  wire [7:0]       fillBySeg_hi_lo_hi_hi_3 = {{4{maskForGroupWire[23]}}, {4{maskForGroupWire[22]}}};
  wire [15:0]      fillBySeg_hi_lo_hi_3 = {fillBySeg_hi_lo_hi_hi_3, fillBySeg_hi_lo_hi_lo_3};
  wire [31:0]      fillBySeg_hi_lo_3 = {fillBySeg_hi_lo_hi_3, fillBySeg_hi_lo_lo_3};
  wire [7:0]       fillBySeg_hi_hi_lo_lo_3 = {{4{maskForGroupWire[25]}}, {4{maskForGroupWire[24]}}};
  wire [7:0]       fillBySeg_hi_hi_lo_hi_3 = {{4{maskForGroupWire[27]}}, {4{maskForGroupWire[26]}}};
  wire [15:0]      fillBySeg_hi_hi_lo_3 = {fillBySeg_hi_hi_lo_hi_3, fillBySeg_hi_hi_lo_lo_3};
  wire [7:0]       fillBySeg_hi_hi_hi_lo_3 = {{4{maskForGroupWire[29]}}, {4{maskForGroupWire[28]}}};
  wire [7:0]       fillBySeg_hi_hi_hi_hi_3 = {{4{maskForGroupWire[31]}}, {4{maskForGroupWire[30]}}};
  wire [15:0]      fillBySeg_hi_hi_hi_3 = {fillBySeg_hi_hi_hi_hi_3, fillBySeg_hi_hi_hi_lo_3};
  wire [31:0]      fillBySeg_hi_hi_3 = {fillBySeg_hi_hi_hi_3, fillBySeg_hi_hi_lo_3};
  wire [63:0]      fillBySeg_hi_3 = {fillBySeg_hi_hi_3, fillBySeg_hi_lo_3};
  wire [9:0]       fillBySeg_lo_lo_lo_lo_4 = {{5{maskForGroupWire[1]}}, {5{maskForGroupWire[0]}}};
  wire [9:0]       fillBySeg_lo_lo_lo_hi_4 = {{5{maskForGroupWire[3]}}, {5{maskForGroupWire[2]}}};
  wire [19:0]      fillBySeg_lo_lo_lo_4 = {fillBySeg_lo_lo_lo_hi_4, fillBySeg_lo_lo_lo_lo_4};
  wire [9:0]       fillBySeg_lo_lo_hi_lo_4 = {{5{maskForGroupWire[5]}}, {5{maskForGroupWire[4]}}};
  wire [9:0]       fillBySeg_lo_lo_hi_hi_4 = {{5{maskForGroupWire[7]}}, {5{maskForGroupWire[6]}}};
  wire [19:0]      fillBySeg_lo_lo_hi_4 = {fillBySeg_lo_lo_hi_hi_4, fillBySeg_lo_lo_hi_lo_4};
  wire [39:0]      fillBySeg_lo_lo_4 = {fillBySeg_lo_lo_hi_4, fillBySeg_lo_lo_lo_4};
  wire [9:0]       fillBySeg_lo_hi_lo_lo_4 = {{5{maskForGroupWire[9]}}, {5{maskForGroupWire[8]}}};
  wire [9:0]       fillBySeg_lo_hi_lo_hi_4 = {{5{maskForGroupWire[11]}}, {5{maskForGroupWire[10]}}};
  wire [19:0]      fillBySeg_lo_hi_lo_4 = {fillBySeg_lo_hi_lo_hi_4, fillBySeg_lo_hi_lo_lo_4};
  wire [9:0]       fillBySeg_lo_hi_hi_lo_4 = {{5{maskForGroupWire[13]}}, {5{maskForGroupWire[12]}}};
  wire [9:0]       fillBySeg_lo_hi_hi_hi_4 = {{5{maskForGroupWire[15]}}, {5{maskForGroupWire[14]}}};
  wire [19:0]      fillBySeg_lo_hi_hi_4 = {fillBySeg_lo_hi_hi_hi_4, fillBySeg_lo_hi_hi_lo_4};
  wire [39:0]      fillBySeg_lo_hi_4 = {fillBySeg_lo_hi_hi_4, fillBySeg_lo_hi_lo_4};
  wire [79:0]      fillBySeg_lo_4 = {fillBySeg_lo_hi_4, fillBySeg_lo_lo_4};
  wire [9:0]       fillBySeg_hi_lo_lo_lo_4 = {{5{maskForGroupWire[17]}}, {5{maskForGroupWire[16]}}};
  wire [9:0]       fillBySeg_hi_lo_lo_hi_4 = {{5{maskForGroupWire[19]}}, {5{maskForGroupWire[18]}}};
  wire [19:0]      fillBySeg_hi_lo_lo_4 = {fillBySeg_hi_lo_lo_hi_4, fillBySeg_hi_lo_lo_lo_4};
  wire [9:0]       fillBySeg_hi_lo_hi_lo_4 = {{5{maskForGroupWire[21]}}, {5{maskForGroupWire[20]}}};
  wire [9:0]       fillBySeg_hi_lo_hi_hi_4 = {{5{maskForGroupWire[23]}}, {5{maskForGroupWire[22]}}};
  wire [19:0]      fillBySeg_hi_lo_hi_4 = {fillBySeg_hi_lo_hi_hi_4, fillBySeg_hi_lo_hi_lo_4};
  wire [39:0]      fillBySeg_hi_lo_4 = {fillBySeg_hi_lo_hi_4, fillBySeg_hi_lo_lo_4};
  wire [9:0]       fillBySeg_hi_hi_lo_lo_4 = {{5{maskForGroupWire[25]}}, {5{maskForGroupWire[24]}}};
  wire [9:0]       fillBySeg_hi_hi_lo_hi_4 = {{5{maskForGroupWire[27]}}, {5{maskForGroupWire[26]}}};
  wire [19:0]      fillBySeg_hi_hi_lo_4 = {fillBySeg_hi_hi_lo_hi_4, fillBySeg_hi_hi_lo_lo_4};
  wire [9:0]       fillBySeg_hi_hi_hi_lo_4 = {{5{maskForGroupWire[29]}}, {5{maskForGroupWire[28]}}};
  wire [9:0]       fillBySeg_hi_hi_hi_hi_4 = {{5{maskForGroupWire[31]}}, {5{maskForGroupWire[30]}}};
  wire [19:0]      fillBySeg_hi_hi_hi_4 = {fillBySeg_hi_hi_hi_hi_4, fillBySeg_hi_hi_hi_lo_4};
  wire [39:0]      fillBySeg_hi_hi_4 = {fillBySeg_hi_hi_hi_4, fillBySeg_hi_hi_lo_4};
  wire [79:0]      fillBySeg_hi_4 = {fillBySeg_hi_hi_4, fillBySeg_hi_lo_4};
  wire [11:0]      fillBySeg_lo_lo_lo_lo_5 = {{6{maskForGroupWire[1]}}, {6{maskForGroupWire[0]}}};
  wire [11:0]      fillBySeg_lo_lo_lo_hi_5 = {{6{maskForGroupWire[3]}}, {6{maskForGroupWire[2]}}};
  wire [23:0]      fillBySeg_lo_lo_lo_5 = {fillBySeg_lo_lo_lo_hi_5, fillBySeg_lo_lo_lo_lo_5};
  wire [11:0]      fillBySeg_lo_lo_hi_lo_5 = {{6{maskForGroupWire[5]}}, {6{maskForGroupWire[4]}}};
  wire [11:0]      fillBySeg_lo_lo_hi_hi_5 = {{6{maskForGroupWire[7]}}, {6{maskForGroupWire[6]}}};
  wire [23:0]      fillBySeg_lo_lo_hi_5 = {fillBySeg_lo_lo_hi_hi_5, fillBySeg_lo_lo_hi_lo_5};
  wire [47:0]      fillBySeg_lo_lo_5 = {fillBySeg_lo_lo_hi_5, fillBySeg_lo_lo_lo_5};
  wire [11:0]      fillBySeg_lo_hi_lo_lo_5 = {{6{maskForGroupWire[9]}}, {6{maskForGroupWire[8]}}};
  wire [11:0]      fillBySeg_lo_hi_lo_hi_5 = {{6{maskForGroupWire[11]}}, {6{maskForGroupWire[10]}}};
  wire [23:0]      fillBySeg_lo_hi_lo_5 = {fillBySeg_lo_hi_lo_hi_5, fillBySeg_lo_hi_lo_lo_5};
  wire [11:0]      fillBySeg_lo_hi_hi_lo_5 = {{6{maskForGroupWire[13]}}, {6{maskForGroupWire[12]}}};
  wire [11:0]      fillBySeg_lo_hi_hi_hi_5 = {{6{maskForGroupWire[15]}}, {6{maskForGroupWire[14]}}};
  wire [23:0]      fillBySeg_lo_hi_hi_5 = {fillBySeg_lo_hi_hi_hi_5, fillBySeg_lo_hi_hi_lo_5};
  wire [47:0]      fillBySeg_lo_hi_5 = {fillBySeg_lo_hi_hi_5, fillBySeg_lo_hi_lo_5};
  wire [95:0]      fillBySeg_lo_5 = {fillBySeg_lo_hi_5, fillBySeg_lo_lo_5};
  wire [11:0]      fillBySeg_hi_lo_lo_lo_5 = {{6{maskForGroupWire[17]}}, {6{maskForGroupWire[16]}}};
  wire [11:0]      fillBySeg_hi_lo_lo_hi_5 = {{6{maskForGroupWire[19]}}, {6{maskForGroupWire[18]}}};
  wire [23:0]      fillBySeg_hi_lo_lo_5 = {fillBySeg_hi_lo_lo_hi_5, fillBySeg_hi_lo_lo_lo_5};
  wire [11:0]      fillBySeg_hi_lo_hi_lo_5 = {{6{maskForGroupWire[21]}}, {6{maskForGroupWire[20]}}};
  wire [11:0]      fillBySeg_hi_lo_hi_hi_5 = {{6{maskForGroupWire[23]}}, {6{maskForGroupWire[22]}}};
  wire [23:0]      fillBySeg_hi_lo_hi_5 = {fillBySeg_hi_lo_hi_hi_5, fillBySeg_hi_lo_hi_lo_5};
  wire [47:0]      fillBySeg_hi_lo_5 = {fillBySeg_hi_lo_hi_5, fillBySeg_hi_lo_lo_5};
  wire [11:0]      fillBySeg_hi_hi_lo_lo_5 = {{6{maskForGroupWire[25]}}, {6{maskForGroupWire[24]}}};
  wire [11:0]      fillBySeg_hi_hi_lo_hi_5 = {{6{maskForGroupWire[27]}}, {6{maskForGroupWire[26]}}};
  wire [23:0]      fillBySeg_hi_hi_lo_5 = {fillBySeg_hi_hi_lo_hi_5, fillBySeg_hi_hi_lo_lo_5};
  wire [11:0]      fillBySeg_hi_hi_hi_lo_5 = {{6{maskForGroupWire[29]}}, {6{maskForGroupWire[28]}}};
  wire [11:0]      fillBySeg_hi_hi_hi_hi_5 = {{6{maskForGroupWire[31]}}, {6{maskForGroupWire[30]}}};
  wire [23:0]      fillBySeg_hi_hi_hi_5 = {fillBySeg_hi_hi_hi_hi_5, fillBySeg_hi_hi_hi_lo_5};
  wire [47:0]      fillBySeg_hi_hi_5 = {fillBySeg_hi_hi_hi_5, fillBySeg_hi_hi_lo_5};
  wire [95:0]      fillBySeg_hi_5 = {fillBySeg_hi_hi_5, fillBySeg_hi_lo_5};
  wire [13:0]      fillBySeg_lo_lo_lo_lo_6 = {{7{maskForGroupWire[1]}}, {7{maskForGroupWire[0]}}};
  wire [13:0]      fillBySeg_lo_lo_lo_hi_6 = {{7{maskForGroupWire[3]}}, {7{maskForGroupWire[2]}}};
  wire [27:0]      fillBySeg_lo_lo_lo_6 = {fillBySeg_lo_lo_lo_hi_6, fillBySeg_lo_lo_lo_lo_6};
  wire [13:0]      fillBySeg_lo_lo_hi_lo_6 = {{7{maskForGroupWire[5]}}, {7{maskForGroupWire[4]}}};
  wire [13:0]      fillBySeg_lo_lo_hi_hi_6 = {{7{maskForGroupWire[7]}}, {7{maskForGroupWire[6]}}};
  wire [27:0]      fillBySeg_lo_lo_hi_6 = {fillBySeg_lo_lo_hi_hi_6, fillBySeg_lo_lo_hi_lo_6};
  wire [55:0]      fillBySeg_lo_lo_6 = {fillBySeg_lo_lo_hi_6, fillBySeg_lo_lo_lo_6};
  wire [13:0]      fillBySeg_lo_hi_lo_lo_6 = {{7{maskForGroupWire[9]}}, {7{maskForGroupWire[8]}}};
  wire [13:0]      fillBySeg_lo_hi_lo_hi_6 = {{7{maskForGroupWire[11]}}, {7{maskForGroupWire[10]}}};
  wire [27:0]      fillBySeg_lo_hi_lo_6 = {fillBySeg_lo_hi_lo_hi_6, fillBySeg_lo_hi_lo_lo_6};
  wire [13:0]      fillBySeg_lo_hi_hi_lo_6 = {{7{maskForGroupWire[13]}}, {7{maskForGroupWire[12]}}};
  wire [13:0]      fillBySeg_lo_hi_hi_hi_6 = {{7{maskForGroupWire[15]}}, {7{maskForGroupWire[14]}}};
  wire [27:0]      fillBySeg_lo_hi_hi_6 = {fillBySeg_lo_hi_hi_hi_6, fillBySeg_lo_hi_hi_lo_6};
  wire [55:0]      fillBySeg_lo_hi_6 = {fillBySeg_lo_hi_hi_6, fillBySeg_lo_hi_lo_6};
  wire [111:0]     fillBySeg_lo_6 = {fillBySeg_lo_hi_6, fillBySeg_lo_lo_6};
  wire [13:0]      fillBySeg_hi_lo_lo_lo_6 = {{7{maskForGroupWire[17]}}, {7{maskForGroupWire[16]}}};
  wire [13:0]      fillBySeg_hi_lo_lo_hi_6 = {{7{maskForGroupWire[19]}}, {7{maskForGroupWire[18]}}};
  wire [27:0]      fillBySeg_hi_lo_lo_6 = {fillBySeg_hi_lo_lo_hi_6, fillBySeg_hi_lo_lo_lo_6};
  wire [13:0]      fillBySeg_hi_lo_hi_lo_6 = {{7{maskForGroupWire[21]}}, {7{maskForGroupWire[20]}}};
  wire [13:0]      fillBySeg_hi_lo_hi_hi_6 = {{7{maskForGroupWire[23]}}, {7{maskForGroupWire[22]}}};
  wire [27:0]      fillBySeg_hi_lo_hi_6 = {fillBySeg_hi_lo_hi_hi_6, fillBySeg_hi_lo_hi_lo_6};
  wire [55:0]      fillBySeg_hi_lo_6 = {fillBySeg_hi_lo_hi_6, fillBySeg_hi_lo_lo_6};
  wire [13:0]      fillBySeg_hi_hi_lo_lo_6 = {{7{maskForGroupWire[25]}}, {7{maskForGroupWire[24]}}};
  wire [13:0]      fillBySeg_hi_hi_lo_hi_6 = {{7{maskForGroupWire[27]}}, {7{maskForGroupWire[26]}}};
  wire [27:0]      fillBySeg_hi_hi_lo_6 = {fillBySeg_hi_hi_lo_hi_6, fillBySeg_hi_hi_lo_lo_6};
  wire [13:0]      fillBySeg_hi_hi_hi_lo_6 = {{7{maskForGroupWire[29]}}, {7{maskForGroupWire[28]}}};
  wire [13:0]      fillBySeg_hi_hi_hi_hi_6 = {{7{maskForGroupWire[31]}}, {7{maskForGroupWire[30]}}};
  wire [27:0]      fillBySeg_hi_hi_hi_6 = {fillBySeg_hi_hi_hi_hi_6, fillBySeg_hi_hi_hi_lo_6};
  wire [55:0]      fillBySeg_hi_hi_6 = {fillBySeg_hi_hi_hi_6, fillBySeg_hi_hi_lo_6};
  wire [111:0]     fillBySeg_hi_6 = {fillBySeg_hi_hi_6, fillBySeg_hi_lo_6};
  wire [15:0]      fillBySeg_lo_lo_lo_lo_7 = {{8{maskForGroupWire[1]}}, {8{maskForGroupWire[0]}}};
  wire [15:0]      fillBySeg_lo_lo_lo_hi_7 = {{8{maskForGroupWire[3]}}, {8{maskForGroupWire[2]}}};
  wire [31:0]      fillBySeg_lo_lo_lo_7 = {fillBySeg_lo_lo_lo_hi_7, fillBySeg_lo_lo_lo_lo_7};
  wire [15:0]      fillBySeg_lo_lo_hi_lo_7 = {{8{maskForGroupWire[5]}}, {8{maskForGroupWire[4]}}};
  wire [15:0]      fillBySeg_lo_lo_hi_hi_7 = {{8{maskForGroupWire[7]}}, {8{maskForGroupWire[6]}}};
  wire [31:0]      fillBySeg_lo_lo_hi_7 = {fillBySeg_lo_lo_hi_hi_7, fillBySeg_lo_lo_hi_lo_7};
  wire [63:0]      fillBySeg_lo_lo_7 = {fillBySeg_lo_lo_hi_7, fillBySeg_lo_lo_lo_7};
  wire [15:0]      fillBySeg_lo_hi_lo_lo_7 = {{8{maskForGroupWire[9]}}, {8{maskForGroupWire[8]}}};
  wire [15:0]      fillBySeg_lo_hi_lo_hi_7 = {{8{maskForGroupWire[11]}}, {8{maskForGroupWire[10]}}};
  wire [31:0]      fillBySeg_lo_hi_lo_7 = {fillBySeg_lo_hi_lo_hi_7, fillBySeg_lo_hi_lo_lo_7};
  wire [15:0]      fillBySeg_lo_hi_hi_lo_7 = {{8{maskForGroupWire[13]}}, {8{maskForGroupWire[12]}}};
  wire [15:0]      fillBySeg_lo_hi_hi_hi_7 = {{8{maskForGroupWire[15]}}, {8{maskForGroupWire[14]}}};
  wire [31:0]      fillBySeg_lo_hi_hi_7 = {fillBySeg_lo_hi_hi_hi_7, fillBySeg_lo_hi_hi_lo_7};
  wire [63:0]      fillBySeg_lo_hi_7 = {fillBySeg_lo_hi_hi_7, fillBySeg_lo_hi_lo_7};
  wire [127:0]     fillBySeg_lo_7 = {fillBySeg_lo_hi_7, fillBySeg_lo_lo_7};
  wire [15:0]      fillBySeg_hi_lo_lo_lo_7 = {{8{maskForGroupWire[17]}}, {8{maskForGroupWire[16]}}};
  wire [15:0]      fillBySeg_hi_lo_lo_hi_7 = {{8{maskForGroupWire[19]}}, {8{maskForGroupWire[18]}}};
  wire [31:0]      fillBySeg_hi_lo_lo_7 = {fillBySeg_hi_lo_lo_hi_7, fillBySeg_hi_lo_lo_lo_7};
  wire [15:0]      fillBySeg_hi_lo_hi_lo_7 = {{8{maskForGroupWire[21]}}, {8{maskForGroupWire[20]}}};
  wire [15:0]      fillBySeg_hi_lo_hi_hi_7 = {{8{maskForGroupWire[23]}}, {8{maskForGroupWire[22]}}};
  wire [31:0]      fillBySeg_hi_lo_hi_7 = {fillBySeg_hi_lo_hi_hi_7, fillBySeg_hi_lo_hi_lo_7};
  wire [63:0]      fillBySeg_hi_lo_7 = {fillBySeg_hi_lo_hi_7, fillBySeg_hi_lo_lo_7};
  wire [15:0]      fillBySeg_hi_hi_lo_lo_7 = {{8{maskForGroupWire[25]}}, {8{maskForGroupWire[24]}}};
  wire [15:0]      fillBySeg_hi_hi_lo_hi_7 = {{8{maskForGroupWire[27]}}, {8{maskForGroupWire[26]}}};
  wire [31:0]      fillBySeg_hi_hi_lo_7 = {fillBySeg_hi_hi_lo_hi_7, fillBySeg_hi_hi_lo_lo_7};
  wire [15:0]      fillBySeg_hi_hi_hi_lo_7 = {{8{maskForGroupWire[29]}}, {8{maskForGroupWire[28]}}};
  wire [15:0]      fillBySeg_hi_hi_hi_hi_7 = {{8{maskForGroupWire[31]}}, {8{maskForGroupWire[30]}}};
  wire [31:0]      fillBySeg_hi_hi_hi_7 = {fillBySeg_hi_hi_hi_hi_7, fillBySeg_hi_hi_hi_lo_7};
  wire [63:0]      fillBySeg_hi_hi_7 = {fillBySeg_hi_hi_hi_7, fillBySeg_hi_hi_lo_7};
  wire [127:0]     fillBySeg_hi_7 = {fillBySeg_hi_hi_7, fillBySeg_hi_lo_7};
  wire [255:0]     fillBySeg =
    {32'h0,
     {32'h0,
      {32'h0,
       {32'h0,
        {32'h0, {32'h0, {32'h0, _fillBySeg_T[0] ? {fillBySeg_hi, fillBySeg_lo} : 32'h0} | (_fillBySeg_T[1] ? {fillBySeg_hi_1, fillBySeg_lo_1} : 64'h0)} | (_fillBySeg_T[2] ? {fillBySeg_hi_2, fillBySeg_lo_2} : 96'h0)}
          | (_fillBySeg_T[3] ? {fillBySeg_hi_3, fillBySeg_lo_3} : 128'h0)} | (_fillBySeg_T[4] ? {fillBySeg_hi_4, fillBySeg_lo_4} : 160'h0)} | (_fillBySeg_T[5] ? {fillBySeg_hi_5, fillBySeg_lo_5} : 192'h0)}
       | (_fillBySeg_T[6] ? {fillBySeg_hi_6, fillBySeg_lo_6} : 224'h0)} | (_fillBySeg_T[7] ? {fillBySeg_hi_7, fillBySeg_lo_7} : 256'h0);
  wire [7:0]       dataRegroupBySew_0_0 = bufferStageEnqueueData_0[7:0];
  wire [7:0]       dataRegroupBySew_0_1 = bufferStageEnqueueData_0[15:8];
  wire [7:0]       dataRegroupBySew_0_2 = bufferStageEnqueueData_0[23:16];
  wire [7:0]       dataRegroupBySew_0_3 = bufferStageEnqueueData_0[31:24];
  wire [7:0]       dataRegroupBySew_0_4 = bufferStageEnqueueData_0[39:32];
  wire [7:0]       dataRegroupBySew_0_5 = bufferStageEnqueueData_0[47:40];
  wire [7:0]       dataRegroupBySew_0_6 = bufferStageEnqueueData_0[55:48];
  wire [7:0]       dataRegroupBySew_0_7 = bufferStageEnqueueData_0[63:56];
  wire [7:0]       dataRegroupBySew_0_8 = bufferStageEnqueueData_0[71:64];
  wire [7:0]       dataRegroupBySew_0_9 = bufferStageEnqueueData_0[79:72];
  wire [7:0]       dataRegroupBySew_0_10 = bufferStageEnqueueData_0[87:80];
  wire [7:0]       dataRegroupBySew_0_11 = bufferStageEnqueueData_0[95:88];
  wire [7:0]       dataRegroupBySew_0_12 = bufferStageEnqueueData_0[103:96];
  wire [7:0]       dataRegroupBySew_0_13 = bufferStageEnqueueData_0[111:104];
  wire [7:0]       dataRegroupBySew_0_14 = bufferStageEnqueueData_0[119:112];
  wire [7:0]       dataRegroupBySew_0_15 = bufferStageEnqueueData_0[127:120];
  wire [7:0]       dataRegroupBySew_0_16 = bufferStageEnqueueData_0[135:128];
  wire [7:0]       dataRegroupBySew_0_17 = bufferStageEnqueueData_0[143:136];
  wire [7:0]       dataRegroupBySew_0_18 = bufferStageEnqueueData_0[151:144];
  wire [7:0]       dataRegroupBySew_0_19 = bufferStageEnqueueData_0[159:152];
  wire [7:0]       dataRegroupBySew_0_20 = bufferStageEnqueueData_0[167:160];
  wire [7:0]       dataRegroupBySew_0_21 = bufferStageEnqueueData_0[175:168];
  wire [7:0]       dataRegroupBySew_0_22 = bufferStageEnqueueData_0[183:176];
  wire [7:0]       dataRegroupBySew_0_23 = bufferStageEnqueueData_0[191:184];
  wire [7:0]       dataRegroupBySew_0_24 = bufferStageEnqueueData_0[199:192];
  wire [7:0]       dataRegroupBySew_0_25 = bufferStageEnqueueData_0[207:200];
  wire [7:0]       dataRegroupBySew_0_26 = bufferStageEnqueueData_0[215:208];
  wire [7:0]       dataRegroupBySew_0_27 = bufferStageEnqueueData_0[223:216];
  wire [7:0]       dataRegroupBySew_0_28 = bufferStageEnqueueData_0[231:224];
  wire [7:0]       dataRegroupBySew_0_29 = bufferStageEnqueueData_0[239:232];
  wire [7:0]       dataRegroupBySew_0_30 = bufferStageEnqueueData_0[247:240];
  wire [7:0]       dataRegroupBySew_0_31 = bufferStageEnqueueData_0[255:248];
  wire [7:0]       dataRegroupBySew_1_0 = bufferStageEnqueueData_1[7:0];
  wire [7:0]       dataRegroupBySew_1_1 = bufferStageEnqueueData_1[15:8];
  wire [7:0]       dataRegroupBySew_1_2 = bufferStageEnqueueData_1[23:16];
  wire [7:0]       dataRegroupBySew_1_3 = bufferStageEnqueueData_1[31:24];
  wire [7:0]       dataRegroupBySew_1_4 = bufferStageEnqueueData_1[39:32];
  wire [7:0]       dataRegroupBySew_1_5 = bufferStageEnqueueData_1[47:40];
  wire [7:0]       dataRegroupBySew_1_6 = bufferStageEnqueueData_1[55:48];
  wire [7:0]       dataRegroupBySew_1_7 = bufferStageEnqueueData_1[63:56];
  wire [7:0]       dataRegroupBySew_1_8 = bufferStageEnqueueData_1[71:64];
  wire [7:0]       dataRegroupBySew_1_9 = bufferStageEnqueueData_1[79:72];
  wire [7:0]       dataRegroupBySew_1_10 = bufferStageEnqueueData_1[87:80];
  wire [7:0]       dataRegroupBySew_1_11 = bufferStageEnqueueData_1[95:88];
  wire [7:0]       dataRegroupBySew_1_12 = bufferStageEnqueueData_1[103:96];
  wire [7:0]       dataRegroupBySew_1_13 = bufferStageEnqueueData_1[111:104];
  wire [7:0]       dataRegroupBySew_1_14 = bufferStageEnqueueData_1[119:112];
  wire [7:0]       dataRegroupBySew_1_15 = bufferStageEnqueueData_1[127:120];
  wire [7:0]       dataRegroupBySew_1_16 = bufferStageEnqueueData_1[135:128];
  wire [7:0]       dataRegroupBySew_1_17 = bufferStageEnqueueData_1[143:136];
  wire [7:0]       dataRegroupBySew_1_18 = bufferStageEnqueueData_1[151:144];
  wire [7:0]       dataRegroupBySew_1_19 = bufferStageEnqueueData_1[159:152];
  wire [7:0]       dataRegroupBySew_1_20 = bufferStageEnqueueData_1[167:160];
  wire [7:0]       dataRegroupBySew_1_21 = bufferStageEnqueueData_1[175:168];
  wire [7:0]       dataRegroupBySew_1_22 = bufferStageEnqueueData_1[183:176];
  wire [7:0]       dataRegroupBySew_1_23 = bufferStageEnqueueData_1[191:184];
  wire [7:0]       dataRegroupBySew_1_24 = bufferStageEnqueueData_1[199:192];
  wire [7:0]       dataRegroupBySew_1_25 = bufferStageEnqueueData_1[207:200];
  wire [7:0]       dataRegroupBySew_1_26 = bufferStageEnqueueData_1[215:208];
  wire [7:0]       dataRegroupBySew_1_27 = bufferStageEnqueueData_1[223:216];
  wire [7:0]       dataRegroupBySew_1_28 = bufferStageEnqueueData_1[231:224];
  wire [7:0]       dataRegroupBySew_1_29 = bufferStageEnqueueData_1[239:232];
  wire [7:0]       dataRegroupBySew_1_30 = bufferStageEnqueueData_1[247:240];
  wire [7:0]       dataRegroupBySew_1_31 = bufferStageEnqueueData_1[255:248];
  wire [7:0]       dataRegroupBySew_2_0 = bufferStageEnqueueData_2[7:0];
  wire [7:0]       dataRegroupBySew_2_1 = bufferStageEnqueueData_2[15:8];
  wire [7:0]       dataRegroupBySew_2_2 = bufferStageEnqueueData_2[23:16];
  wire [7:0]       dataRegroupBySew_2_3 = bufferStageEnqueueData_2[31:24];
  wire [7:0]       dataRegroupBySew_2_4 = bufferStageEnqueueData_2[39:32];
  wire [7:0]       dataRegroupBySew_2_5 = bufferStageEnqueueData_2[47:40];
  wire [7:0]       dataRegroupBySew_2_6 = bufferStageEnqueueData_2[55:48];
  wire [7:0]       dataRegroupBySew_2_7 = bufferStageEnqueueData_2[63:56];
  wire [7:0]       dataRegroupBySew_2_8 = bufferStageEnqueueData_2[71:64];
  wire [7:0]       dataRegroupBySew_2_9 = bufferStageEnqueueData_2[79:72];
  wire [7:0]       dataRegroupBySew_2_10 = bufferStageEnqueueData_2[87:80];
  wire [7:0]       dataRegroupBySew_2_11 = bufferStageEnqueueData_2[95:88];
  wire [7:0]       dataRegroupBySew_2_12 = bufferStageEnqueueData_2[103:96];
  wire [7:0]       dataRegroupBySew_2_13 = bufferStageEnqueueData_2[111:104];
  wire [7:0]       dataRegroupBySew_2_14 = bufferStageEnqueueData_2[119:112];
  wire [7:0]       dataRegroupBySew_2_15 = bufferStageEnqueueData_2[127:120];
  wire [7:0]       dataRegroupBySew_2_16 = bufferStageEnqueueData_2[135:128];
  wire [7:0]       dataRegroupBySew_2_17 = bufferStageEnqueueData_2[143:136];
  wire [7:0]       dataRegroupBySew_2_18 = bufferStageEnqueueData_2[151:144];
  wire [7:0]       dataRegroupBySew_2_19 = bufferStageEnqueueData_2[159:152];
  wire [7:0]       dataRegroupBySew_2_20 = bufferStageEnqueueData_2[167:160];
  wire [7:0]       dataRegroupBySew_2_21 = bufferStageEnqueueData_2[175:168];
  wire [7:0]       dataRegroupBySew_2_22 = bufferStageEnqueueData_2[183:176];
  wire [7:0]       dataRegroupBySew_2_23 = bufferStageEnqueueData_2[191:184];
  wire [7:0]       dataRegroupBySew_2_24 = bufferStageEnqueueData_2[199:192];
  wire [7:0]       dataRegroupBySew_2_25 = bufferStageEnqueueData_2[207:200];
  wire [7:0]       dataRegroupBySew_2_26 = bufferStageEnqueueData_2[215:208];
  wire [7:0]       dataRegroupBySew_2_27 = bufferStageEnqueueData_2[223:216];
  wire [7:0]       dataRegroupBySew_2_28 = bufferStageEnqueueData_2[231:224];
  wire [7:0]       dataRegroupBySew_2_29 = bufferStageEnqueueData_2[239:232];
  wire [7:0]       dataRegroupBySew_2_30 = bufferStageEnqueueData_2[247:240];
  wire [7:0]       dataRegroupBySew_2_31 = bufferStageEnqueueData_2[255:248];
  wire [7:0]       dataRegroupBySew_3_0 = bufferStageEnqueueData_3[7:0];
  wire [7:0]       dataRegroupBySew_3_1 = bufferStageEnqueueData_3[15:8];
  wire [7:0]       dataRegroupBySew_3_2 = bufferStageEnqueueData_3[23:16];
  wire [7:0]       dataRegroupBySew_3_3 = bufferStageEnqueueData_3[31:24];
  wire [7:0]       dataRegroupBySew_3_4 = bufferStageEnqueueData_3[39:32];
  wire [7:0]       dataRegroupBySew_3_5 = bufferStageEnqueueData_3[47:40];
  wire [7:0]       dataRegroupBySew_3_6 = bufferStageEnqueueData_3[55:48];
  wire [7:0]       dataRegroupBySew_3_7 = bufferStageEnqueueData_3[63:56];
  wire [7:0]       dataRegroupBySew_3_8 = bufferStageEnqueueData_3[71:64];
  wire [7:0]       dataRegroupBySew_3_9 = bufferStageEnqueueData_3[79:72];
  wire [7:0]       dataRegroupBySew_3_10 = bufferStageEnqueueData_3[87:80];
  wire [7:0]       dataRegroupBySew_3_11 = bufferStageEnqueueData_3[95:88];
  wire [7:0]       dataRegroupBySew_3_12 = bufferStageEnqueueData_3[103:96];
  wire [7:0]       dataRegroupBySew_3_13 = bufferStageEnqueueData_3[111:104];
  wire [7:0]       dataRegroupBySew_3_14 = bufferStageEnqueueData_3[119:112];
  wire [7:0]       dataRegroupBySew_3_15 = bufferStageEnqueueData_3[127:120];
  wire [7:0]       dataRegroupBySew_3_16 = bufferStageEnqueueData_3[135:128];
  wire [7:0]       dataRegroupBySew_3_17 = bufferStageEnqueueData_3[143:136];
  wire [7:0]       dataRegroupBySew_3_18 = bufferStageEnqueueData_3[151:144];
  wire [7:0]       dataRegroupBySew_3_19 = bufferStageEnqueueData_3[159:152];
  wire [7:0]       dataRegroupBySew_3_20 = bufferStageEnqueueData_3[167:160];
  wire [7:0]       dataRegroupBySew_3_21 = bufferStageEnqueueData_3[175:168];
  wire [7:0]       dataRegroupBySew_3_22 = bufferStageEnqueueData_3[183:176];
  wire [7:0]       dataRegroupBySew_3_23 = bufferStageEnqueueData_3[191:184];
  wire [7:0]       dataRegroupBySew_3_24 = bufferStageEnqueueData_3[199:192];
  wire [7:0]       dataRegroupBySew_3_25 = bufferStageEnqueueData_3[207:200];
  wire [7:0]       dataRegroupBySew_3_26 = bufferStageEnqueueData_3[215:208];
  wire [7:0]       dataRegroupBySew_3_27 = bufferStageEnqueueData_3[223:216];
  wire [7:0]       dataRegroupBySew_3_28 = bufferStageEnqueueData_3[231:224];
  wire [7:0]       dataRegroupBySew_3_29 = bufferStageEnqueueData_3[239:232];
  wire [7:0]       dataRegroupBySew_3_30 = bufferStageEnqueueData_3[247:240];
  wire [7:0]       dataRegroupBySew_3_31 = bufferStageEnqueueData_3[255:248];
  wire [7:0]       dataRegroupBySew_4_0 = bufferStageEnqueueData_4[7:0];
  wire [7:0]       dataRegroupBySew_4_1 = bufferStageEnqueueData_4[15:8];
  wire [7:0]       dataRegroupBySew_4_2 = bufferStageEnqueueData_4[23:16];
  wire [7:0]       dataRegroupBySew_4_3 = bufferStageEnqueueData_4[31:24];
  wire [7:0]       dataRegroupBySew_4_4 = bufferStageEnqueueData_4[39:32];
  wire [7:0]       dataRegroupBySew_4_5 = bufferStageEnqueueData_4[47:40];
  wire [7:0]       dataRegroupBySew_4_6 = bufferStageEnqueueData_4[55:48];
  wire [7:0]       dataRegroupBySew_4_7 = bufferStageEnqueueData_4[63:56];
  wire [7:0]       dataRegroupBySew_4_8 = bufferStageEnqueueData_4[71:64];
  wire [7:0]       dataRegroupBySew_4_9 = bufferStageEnqueueData_4[79:72];
  wire [7:0]       dataRegroupBySew_4_10 = bufferStageEnqueueData_4[87:80];
  wire [7:0]       dataRegroupBySew_4_11 = bufferStageEnqueueData_4[95:88];
  wire [7:0]       dataRegroupBySew_4_12 = bufferStageEnqueueData_4[103:96];
  wire [7:0]       dataRegroupBySew_4_13 = bufferStageEnqueueData_4[111:104];
  wire [7:0]       dataRegroupBySew_4_14 = bufferStageEnqueueData_4[119:112];
  wire [7:0]       dataRegroupBySew_4_15 = bufferStageEnqueueData_4[127:120];
  wire [7:0]       dataRegroupBySew_4_16 = bufferStageEnqueueData_4[135:128];
  wire [7:0]       dataRegroupBySew_4_17 = bufferStageEnqueueData_4[143:136];
  wire [7:0]       dataRegroupBySew_4_18 = bufferStageEnqueueData_4[151:144];
  wire [7:0]       dataRegroupBySew_4_19 = bufferStageEnqueueData_4[159:152];
  wire [7:0]       dataRegroupBySew_4_20 = bufferStageEnqueueData_4[167:160];
  wire [7:0]       dataRegroupBySew_4_21 = bufferStageEnqueueData_4[175:168];
  wire [7:0]       dataRegroupBySew_4_22 = bufferStageEnqueueData_4[183:176];
  wire [7:0]       dataRegroupBySew_4_23 = bufferStageEnqueueData_4[191:184];
  wire [7:0]       dataRegroupBySew_4_24 = bufferStageEnqueueData_4[199:192];
  wire [7:0]       dataRegroupBySew_4_25 = bufferStageEnqueueData_4[207:200];
  wire [7:0]       dataRegroupBySew_4_26 = bufferStageEnqueueData_4[215:208];
  wire [7:0]       dataRegroupBySew_4_27 = bufferStageEnqueueData_4[223:216];
  wire [7:0]       dataRegroupBySew_4_28 = bufferStageEnqueueData_4[231:224];
  wire [7:0]       dataRegroupBySew_4_29 = bufferStageEnqueueData_4[239:232];
  wire [7:0]       dataRegroupBySew_4_30 = bufferStageEnqueueData_4[247:240];
  wire [7:0]       dataRegroupBySew_4_31 = bufferStageEnqueueData_4[255:248];
  wire [7:0]       dataRegroupBySew_5_0 = bufferStageEnqueueData_5[7:0];
  wire [7:0]       dataRegroupBySew_5_1 = bufferStageEnqueueData_5[15:8];
  wire [7:0]       dataRegroupBySew_5_2 = bufferStageEnqueueData_5[23:16];
  wire [7:0]       dataRegroupBySew_5_3 = bufferStageEnqueueData_5[31:24];
  wire [7:0]       dataRegroupBySew_5_4 = bufferStageEnqueueData_5[39:32];
  wire [7:0]       dataRegroupBySew_5_5 = bufferStageEnqueueData_5[47:40];
  wire [7:0]       dataRegroupBySew_5_6 = bufferStageEnqueueData_5[55:48];
  wire [7:0]       dataRegroupBySew_5_7 = bufferStageEnqueueData_5[63:56];
  wire [7:0]       dataRegroupBySew_5_8 = bufferStageEnqueueData_5[71:64];
  wire [7:0]       dataRegroupBySew_5_9 = bufferStageEnqueueData_5[79:72];
  wire [7:0]       dataRegroupBySew_5_10 = bufferStageEnqueueData_5[87:80];
  wire [7:0]       dataRegroupBySew_5_11 = bufferStageEnqueueData_5[95:88];
  wire [7:0]       dataRegroupBySew_5_12 = bufferStageEnqueueData_5[103:96];
  wire [7:0]       dataRegroupBySew_5_13 = bufferStageEnqueueData_5[111:104];
  wire [7:0]       dataRegroupBySew_5_14 = bufferStageEnqueueData_5[119:112];
  wire [7:0]       dataRegroupBySew_5_15 = bufferStageEnqueueData_5[127:120];
  wire [7:0]       dataRegroupBySew_5_16 = bufferStageEnqueueData_5[135:128];
  wire [7:0]       dataRegroupBySew_5_17 = bufferStageEnqueueData_5[143:136];
  wire [7:0]       dataRegroupBySew_5_18 = bufferStageEnqueueData_5[151:144];
  wire [7:0]       dataRegroupBySew_5_19 = bufferStageEnqueueData_5[159:152];
  wire [7:0]       dataRegroupBySew_5_20 = bufferStageEnqueueData_5[167:160];
  wire [7:0]       dataRegroupBySew_5_21 = bufferStageEnqueueData_5[175:168];
  wire [7:0]       dataRegroupBySew_5_22 = bufferStageEnqueueData_5[183:176];
  wire [7:0]       dataRegroupBySew_5_23 = bufferStageEnqueueData_5[191:184];
  wire [7:0]       dataRegroupBySew_5_24 = bufferStageEnqueueData_5[199:192];
  wire [7:0]       dataRegroupBySew_5_25 = bufferStageEnqueueData_5[207:200];
  wire [7:0]       dataRegroupBySew_5_26 = bufferStageEnqueueData_5[215:208];
  wire [7:0]       dataRegroupBySew_5_27 = bufferStageEnqueueData_5[223:216];
  wire [7:0]       dataRegroupBySew_5_28 = bufferStageEnqueueData_5[231:224];
  wire [7:0]       dataRegroupBySew_5_29 = bufferStageEnqueueData_5[239:232];
  wire [7:0]       dataRegroupBySew_5_30 = bufferStageEnqueueData_5[247:240];
  wire [7:0]       dataRegroupBySew_5_31 = bufferStageEnqueueData_5[255:248];
  wire [7:0]       dataRegroupBySew_6_0 = bufferStageEnqueueData_6[7:0];
  wire [7:0]       dataRegroupBySew_6_1 = bufferStageEnqueueData_6[15:8];
  wire [7:0]       dataRegroupBySew_6_2 = bufferStageEnqueueData_6[23:16];
  wire [7:0]       dataRegroupBySew_6_3 = bufferStageEnqueueData_6[31:24];
  wire [7:0]       dataRegroupBySew_6_4 = bufferStageEnqueueData_6[39:32];
  wire [7:0]       dataRegroupBySew_6_5 = bufferStageEnqueueData_6[47:40];
  wire [7:0]       dataRegroupBySew_6_6 = bufferStageEnqueueData_6[55:48];
  wire [7:0]       dataRegroupBySew_6_7 = bufferStageEnqueueData_6[63:56];
  wire [7:0]       dataRegroupBySew_6_8 = bufferStageEnqueueData_6[71:64];
  wire [7:0]       dataRegroupBySew_6_9 = bufferStageEnqueueData_6[79:72];
  wire [7:0]       dataRegroupBySew_6_10 = bufferStageEnqueueData_6[87:80];
  wire [7:0]       dataRegroupBySew_6_11 = bufferStageEnqueueData_6[95:88];
  wire [7:0]       dataRegroupBySew_6_12 = bufferStageEnqueueData_6[103:96];
  wire [7:0]       dataRegroupBySew_6_13 = bufferStageEnqueueData_6[111:104];
  wire [7:0]       dataRegroupBySew_6_14 = bufferStageEnqueueData_6[119:112];
  wire [7:0]       dataRegroupBySew_6_15 = bufferStageEnqueueData_6[127:120];
  wire [7:0]       dataRegroupBySew_6_16 = bufferStageEnqueueData_6[135:128];
  wire [7:0]       dataRegroupBySew_6_17 = bufferStageEnqueueData_6[143:136];
  wire [7:0]       dataRegroupBySew_6_18 = bufferStageEnqueueData_6[151:144];
  wire [7:0]       dataRegroupBySew_6_19 = bufferStageEnqueueData_6[159:152];
  wire [7:0]       dataRegroupBySew_6_20 = bufferStageEnqueueData_6[167:160];
  wire [7:0]       dataRegroupBySew_6_21 = bufferStageEnqueueData_6[175:168];
  wire [7:0]       dataRegroupBySew_6_22 = bufferStageEnqueueData_6[183:176];
  wire [7:0]       dataRegroupBySew_6_23 = bufferStageEnqueueData_6[191:184];
  wire [7:0]       dataRegroupBySew_6_24 = bufferStageEnqueueData_6[199:192];
  wire [7:0]       dataRegroupBySew_6_25 = bufferStageEnqueueData_6[207:200];
  wire [7:0]       dataRegroupBySew_6_26 = bufferStageEnqueueData_6[215:208];
  wire [7:0]       dataRegroupBySew_6_27 = bufferStageEnqueueData_6[223:216];
  wire [7:0]       dataRegroupBySew_6_28 = bufferStageEnqueueData_6[231:224];
  wire [7:0]       dataRegroupBySew_6_29 = bufferStageEnqueueData_6[239:232];
  wire [7:0]       dataRegroupBySew_6_30 = bufferStageEnqueueData_6[247:240];
  wire [7:0]       dataRegroupBySew_6_31 = bufferStageEnqueueData_6[255:248];
  wire [7:0]       dataRegroupBySew_7_0 = bufferStageEnqueueData_7[7:0];
  wire [7:0]       dataRegroupBySew_7_1 = bufferStageEnqueueData_7[15:8];
  wire [7:0]       dataRegroupBySew_7_2 = bufferStageEnqueueData_7[23:16];
  wire [7:0]       dataRegroupBySew_7_3 = bufferStageEnqueueData_7[31:24];
  wire [7:0]       dataRegroupBySew_7_4 = bufferStageEnqueueData_7[39:32];
  wire [7:0]       dataRegroupBySew_7_5 = bufferStageEnqueueData_7[47:40];
  wire [7:0]       dataRegroupBySew_7_6 = bufferStageEnqueueData_7[55:48];
  wire [7:0]       dataRegroupBySew_7_7 = bufferStageEnqueueData_7[63:56];
  wire [7:0]       dataRegroupBySew_7_8 = bufferStageEnqueueData_7[71:64];
  wire [7:0]       dataRegroupBySew_7_9 = bufferStageEnqueueData_7[79:72];
  wire [7:0]       dataRegroupBySew_7_10 = bufferStageEnqueueData_7[87:80];
  wire [7:0]       dataRegroupBySew_7_11 = bufferStageEnqueueData_7[95:88];
  wire [7:0]       dataRegroupBySew_7_12 = bufferStageEnqueueData_7[103:96];
  wire [7:0]       dataRegroupBySew_7_13 = bufferStageEnqueueData_7[111:104];
  wire [7:0]       dataRegroupBySew_7_14 = bufferStageEnqueueData_7[119:112];
  wire [7:0]       dataRegroupBySew_7_15 = bufferStageEnqueueData_7[127:120];
  wire [7:0]       dataRegroupBySew_7_16 = bufferStageEnqueueData_7[135:128];
  wire [7:0]       dataRegroupBySew_7_17 = bufferStageEnqueueData_7[143:136];
  wire [7:0]       dataRegroupBySew_7_18 = bufferStageEnqueueData_7[151:144];
  wire [7:0]       dataRegroupBySew_7_19 = bufferStageEnqueueData_7[159:152];
  wire [7:0]       dataRegroupBySew_7_20 = bufferStageEnqueueData_7[167:160];
  wire [7:0]       dataRegroupBySew_7_21 = bufferStageEnqueueData_7[175:168];
  wire [7:0]       dataRegroupBySew_7_22 = bufferStageEnqueueData_7[183:176];
  wire [7:0]       dataRegroupBySew_7_23 = bufferStageEnqueueData_7[191:184];
  wire [7:0]       dataRegroupBySew_7_24 = bufferStageEnqueueData_7[199:192];
  wire [7:0]       dataRegroupBySew_7_25 = bufferStageEnqueueData_7[207:200];
  wire [7:0]       dataRegroupBySew_7_26 = bufferStageEnqueueData_7[215:208];
  wire [7:0]       dataRegroupBySew_7_27 = bufferStageEnqueueData_7[223:216];
  wire [7:0]       dataRegroupBySew_7_28 = bufferStageEnqueueData_7[231:224];
  wire [7:0]       dataRegroupBySew_7_29 = bufferStageEnqueueData_7[239:232];
  wire [7:0]       dataRegroupBySew_7_30 = bufferStageEnqueueData_7[247:240];
  wire [7:0]       dataRegroupBySew_7_31 = bufferStageEnqueueData_7[255:248];
  wire [15:0]      dataInMem_lo_lo_lo_lo = {dataRegroupBySew_0_1, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_lo_lo_lo_hi = {dataRegroupBySew_0_3, dataRegroupBySew_0_2};
  wire [31:0]      dataInMem_lo_lo_lo = {dataInMem_lo_lo_lo_hi, dataInMem_lo_lo_lo_lo};
  wire [15:0]      dataInMem_lo_lo_hi_lo = {dataRegroupBySew_0_5, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_lo_lo_hi_hi = {dataRegroupBySew_0_7, dataRegroupBySew_0_6};
  wire [31:0]      dataInMem_lo_lo_hi = {dataInMem_lo_lo_hi_hi, dataInMem_lo_lo_hi_lo};
  wire [63:0]      dataInMem_lo_lo = {dataInMem_lo_lo_hi, dataInMem_lo_lo_lo};
  wire [15:0]      dataInMem_lo_hi_lo_lo = {dataRegroupBySew_0_9, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_lo_hi_lo_hi = {dataRegroupBySew_0_11, dataRegroupBySew_0_10};
  wire [31:0]      dataInMem_lo_hi_lo = {dataInMem_lo_hi_lo_hi, dataInMem_lo_hi_lo_lo};
  wire [15:0]      dataInMem_lo_hi_hi_lo = {dataRegroupBySew_0_13, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_lo_hi_hi_hi = {dataRegroupBySew_0_15, dataRegroupBySew_0_14};
  wire [31:0]      dataInMem_lo_hi_hi = {dataInMem_lo_hi_hi_hi, dataInMem_lo_hi_hi_lo};
  wire [63:0]      dataInMem_lo_hi = {dataInMem_lo_hi_hi, dataInMem_lo_hi_lo};
  wire [127:0]     dataInMem_lo = {dataInMem_lo_hi, dataInMem_lo_lo};
  wire [15:0]      dataInMem_hi_lo_lo_lo = {dataRegroupBySew_0_17, dataRegroupBySew_0_16};
  wire [15:0]      dataInMem_hi_lo_lo_hi = {dataRegroupBySew_0_19, dataRegroupBySew_0_18};
  wire [31:0]      dataInMem_hi_lo_lo = {dataInMem_hi_lo_lo_hi, dataInMem_hi_lo_lo_lo};
  wire [15:0]      dataInMem_hi_lo_hi_lo = {dataRegroupBySew_0_21, dataRegroupBySew_0_20};
  wire [15:0]      dataInMem_hi_lo_hi_hi = {dataRegroupBySew_0_23, dataRegroupBySew_0_22};
  wire [31:0]      dataInMem_hi_lo_hi = {dataInMem_hi_lo_hi_hi, dataInMem_hi_lo_hi_lo};
  wire [63:0]      dataInMem_hi_lo = {dataInMem_hi_lo_hi, dataInMem_hi_lo_lo};
  wire [15:0]      dataInMem_hi_hi_lo_lo = {dataRegroupBySew_0_25, dataRegroupBySew_0_24};
  wire [15:0]      dataInMem_hi_hi_lo_hi = {dataRegroupBySew_0_27, dataRegroupBySew_0_26};
  wire [31:0]      dataInMem_hi_hi_lo = {dataInMem_hi_hi_lo_hi, dataInMem_hi_hi_lo_lo};
  wire [15:0]      dataInMem_hi_hi_hi_lo = {dataRegroupBySew_0_29, dataRegroupBySew_0_28};
  wire [15:0]      dataInMem_hi_hi_hi_hi = {dataRegroupBySew_0_31, dataRegroupBySew_0_30};
  wire [31:0]      dataInMem_hi_hi_hi = {dataInMem_hi_hi_hi_hi, dataInMem_hi_hi_hi_lo};
  wire [63:0]      dataInMem_hi_hi = {dataInMem_hi_hi_hi, dataInMem_hi_hi_lo};
  wire [127:0]     dataInMem_hi = {dataInMem_hi_hi, dataInMem_hi_lo};
  wire [255:0]     dataInMem = {dataInMem_hi, dataInMem_lo};
  wire [255:0]     regroupCacheLine_0 = dataInMem;
  wire [255:0]     res = regroupCacheLine_0;
  wire [511:0]     lo_lo = {256'h0, res};
  wire [1023:0]    lo = {512'h0, lo_lo};
  wire [2047:0]    regroupLoadData_0_0 = {1024'h0, lo};
  wire [31:0]      dataInMem_lo_lo_lo_lo_1 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1, dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [31:0]      dataInMem_lo_lo_lo_hi_1 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3, dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [63:0]      dataInMem_lo_lo_lo_1 = {dataInMem_lo_lo_lo_hi_1, dataInMem_lo_lo_lo_lo_1};
  wire [31:0]      dataInMem_lo_lo_hi_lo_1 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5, dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [31:0]      dataInMem_lo_lo_hi_hi_1 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7, dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [63:0]      dataInMem_lo_lo_hi_1 = {dataInMem_lo_lo_hi_hi_1, dataInMem_lo_lo_hi_lo_1};
  wire [127:0]     dataInMem_lo_lo_1 = {dataInMem_lo_lo_hi_1, dataInMem_lo_lo_lo_1};
  wire [31:0]      dataInMem_lo_hi_lo_lo_1 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9, dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [31:0]      dataInMem_lo_hi_lo_hi_1 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11, dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [63:0]      dataInMem_lo_hi_lo_1 = {dataInMem_lo_hi_lo_hi_1, dataInMem_lo_hi_lo_lo_1};
  wire [31:0]      dataInMem_lo_hi_hi_lo_1 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13, dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [31:0]      dataInMem_lo_hi_hi_hi_1 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15, dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [63:0]      dataInMem_lo_hi_hi_1 = {dataInMem_lo_hi_hi_hi_1, dataInMem_lo_hi_hi_lo_1};
  wire [127:0]     dataInMem_lo_hi_1 = {dataInMem_lo_hi_hi_1, dataInMem_lo_hi_lo_1};
  wire [255:0]     dataInMem_lo_1 = {dataInMem_lo_hi_1, dataInMem_lo_lo_1};
  wire [31:0]      dataInMem_hi_lo_lo_lo_1 = {dataRegroupBySew_1_17, dataRegroupBySew_0_17, dataRegroupBySew_1_16, dataRegroupBySew_0_16};
  wire [31:0]      dataInMem_hi_lo_lo_hi_1 = {dataRegroupBySew_1_19, dataRegroupBySew_0_19, dataRegroupBySew_1_18, dataRegroupBySew_0_18};
  wire [63:0]      dataInMem_hi_lo_lo_1 = {dataInMem_hi_lo_lo_hi_1, dataInMem_hi_lo_lo_lo_1};
  wire [31:0]      dataInMem_hi_lo_hi_lo_1 = {dataRegroupBySew_1_21, dataRegroupBySew_0_21, dataRegroupBySew_1_20, dataRegroupBySew_0_20};
  wire [31:0]      dataInMem_hi_lo_hi_hi_1 = {dataRegroupBySew_1_23, dataRegroupBySew_0_23, dataRegroupBySew_1_22, dataRegroupBySew_0_22};
  wire [63:0]      dataInMem_hi_lo_hi_1 = {dataInMem_hi_lo_hi_hi_1, dataInMem_hi_lo_hi_lo_1};
  wire [127:0]     dataInMem_hi_lo_1 = {dataInMem_hi_lo_hi_1, dataInMem_hi_lo_lo_1};
  wire [31:0]      dataInMem_hi_hi_lo_lo_1 = {dataRegroupBySew_1_25, dataRegroupBySew_0_25, dataRegroupBySew_1_24, dataRegroupBySew_0_24};
  wire [31:0]      dataInMem_hi_hi_lo_hi_1 = {dataRegroupBySew_1_27, dataRegroupBySew_0_27, dataRegroupBySew_1_26, dataRegroupBySew_0_26};
  wire [63:0]      dataInMem_hi_hi_lo_1 = {dataInMem_hi_hi_lo_hi_1, dataInMem_hi_hi_lo_lo_1};
  wire [31:0]      dataInMem_hi_hi_hi_lo_1 = {dataRegroupBySew_1_29, dataRegroupBySew_0_29, dataRegroupBySew_1_28, dataRegroupBySew_0_28};
  wire [31:0]      dataInMem_hi_hi_hi_hi_1 = {dataRegroupBySew_1_31, dataRegroupBySew_0_31, dataRegroupBySew_1_30, dataRegroupBySew_0_30};
  wire [63:0]      dataInMem_hi_hi_hi_1 = {dataInMem_hi_hi_hi_hi_1, dataInMem_hi_hi_hi_lo_1};
  wire [127:0]     dataInMem_hi_hi_1 = {dataInMem_hi_hi_hi_1, dataInMem_hi_hi_lo_1};
  wire [255:0]     dataInMem_hi_1 = {dataInMem_hi_hi_1, dataInMem_hi_lo_1};
  wire [511:0]     dataInMem_1 = {dataInMem_hi_1, dataInMem_lo_1};
  wire [255:0]     regroupCacheLine_1_0 = dataInMem_1[255:0];
  wire [255:0]     regroupCacheLine_1_1 = dataInMem_1[511:256];
  wire [255:0]     res_8 = regroupCacheLine_1_0;
  wire [255:0]     res_9 = regroupCacheLine_1_1;
  wire [511:0]     lo_lo_1 = {res_9, res_8};
  wire [1023:0]    lo_1 = {512'h0, lo_lo_1};
  wire [2047:0]    regroupLoadData_0_1 = {1024'h0, lo_1};
  wire [15:0]      _GEN_4 = {dataRegroupBySew_2_0, dataRegroupBySew_1_0};
  wire [15:0]      dataInMem_hi_2;
  assign dataInMem_hi_2 = _GEN_4;
  wire [15:0]      dataInMem_lo_hi_5;
  assign dataInMem_lo_hi_5 = _GEN_4;
  wire [15:0]      dataInMem_lo_hi_38;
  assign dataInMem_lo_hi_38 = _GEN_4;
  wire [15:0]      _GEN_5 = {dataRegroupBySew_2_1, dataRegroupBySew_1_1};
  wire [15:0]      dataInMem_hi_3;
  assign dataInMem_hi_3 = _GEN_5;
  wire [15:0]      dataInMem_lo_hi_6;
  assign dataInMem_lo_hi_6 = _GEN_5;
  wire [15:0]      dataInMem_lo_hi_39;
  assign dataInMem_lo_hi_39 = _GEN_5;
  wire [15:0]      _GEN_6 = {dataRegroupBySew_2_2, dataRegroupBySew_1_2};
  wire [15:0]      dataInMem_hi_4;
  assign dataInMem_hi_4 = _GEN_6;
  wire [15:0]      dataInMem_lo_hi_7;
  assign dataInMem_lo_hi_7 = _GEN_6;
  wire [15:0]      dataInMem_lo_hi_40;
  assign dataInMem_lo_hi_40 = _GEN_6;
  wire [15:0]      _GEN_7 = {dataRegroupBySew_2_3, dataRegroupBySew_1_3};
  wire [15:0]      dataInMem_hi_5;
  assign dataInMem_hi_5 = _GEN_7;
  wire [15:0]      dataInMem_lo_hi_8;
  assign dataInMem_lo_hi_8 = _GEN_7;
  wire [15:0]      dataInMem_lo_hi_41;
  assign dataInMem_lo_hi_41 = _GEN_7;
  wire [15:0]      _GEN_8 = {dataRegroupBySew_2_4, dataRegroupBySew_1_4};
  wire [15:0]      dataInMem_hi_6;
  assign dataInMem_hi_6 = _GEN_8;
  wire [15:0]      dataInMem_lo_hi_9;
  assign dataInMem_lo_hi_9 = _GEN_8;
  wire [15:0]      dataInMem_lo_hi_42;
  assign dataInMem_lo_hi_42 = _GEN_8;
  wire [15:0]      _GEN_9 = {dataRegroupBySew_2_5, dataRegroupBySew_1_5};
  wire [15:0]      dataInMem_hi_7;
  assign dataInMem_hi_7 = _GEN_9;
  wire [15:0]      dataInMem_lo_hi_10;
  assign dataInMem_lo_hi_10 = _GEN_9;
  wire [15:0]      dataInMem_lo_hi_43;
  assign dataInMem_lo_hi_43 = _GEN_9;
  wire [15:0]      _GEN_10 = {dataRegroupBySew_2_6, dataRegroupBySew_1_6};
  wire [15:0]      dataInMem_hi_8;
  assign dataInMem_hi_8 = _GEN_10;
  wire [15:0]      dataInMem_lo_hi_11;
  assign dataInMem_lo_hi_11 = _GEN_10;
  wire [15:0]      dataInMem_lo_hi_44;
  assign dataInMem_lo_hi_44 = _GEN_10;
  wire [15:0]      _GEN_11 = {dataRegroupBySew_2_7, dataRegroupBySew_1_7};
  wire [15:0]      dataInMem_hi_9;
  assign dataInMem_hi_9 = _GEN_11;
  wire [15:0]      dataInMem_lo_hi_12;
  assign dataInMem_lo_hi_12 = _GEN_11;
  wire [15:0]      dataInMem_lo_hi_45;
  assign dataInMem_lo_hi_45 = _GEN_11;
  wire [15:0]      _GEN_12 = {dataRegroupBySew_2_8, dataRegroupBySew_1_8};
  wire [15:0]      dataInMem_hi_10;
  assign dataInMem_hi_10 = _GEN_12;
  wire [15:0]      dataInMem_lo_hi_13;
  assign dataInMem_lo_hi_13 = _GEN_12;
  wire [15:0]      dataInMem_lo_hi_46;
  assign dataInMem_lo_hi_46 = _GEN_12;
  wire [15:0]      _GEN_13 = {dataRegroupBySew_2_9, dataRegroupBySew_1_9};
  wire [15:0]      dataInMem_hi_11;
  assign dataInMem_hi_11 = _GEN_13;
  wire [15:0]      dataInMem_lo_hi_14;
  assign dataInMem_lo_hi_14 = _GEN_13;
  wire [15:0]      dataInMem_lo_hi_47;
  assign dataInMem_lo_hi_47 = _GEN_13;
  wire [15:0]      _GEN_14 = {dataRegroupBySew_2_10, dataRegroupBySew_1_10};
  wire [15:0]      dataInMem_hi_12;
  assign dataInMem_hi_12 = _GEN_14;
  wire [15:0]      dataInMem_lo_hi_15;
  assign dataInMem_lo_hi_15 = _GEN_14;
  wire [15:0]      dataInMem_lo_hi_48;
  assign dataInMem_lo_hi_48 = _GEN_14;
  wire [15:0]      _GEN_15 = {dataRegroupBySew_2_11, dataRegroupBySew_1_11};
  wire [15:0]      dataInMem_hi_13;
  assign dataInMem_hi_13 = _GEN_15;
  wire [15:0]      dataInMem_lo_hi_16;
  assign dataInMem_lo_hi_16 = _GEN_15;
  wire [15:0]      dataInMem_lo_hi_49;
  assign dataInMem_lo_hi_49 = _GEN_15;
  wire [15:0]      _GEN_16 = {dataRegroupBySew_2_12, dataRegroupBySew_1_12};
  wire [15:0]      dataInMem_hi_14;
  assign dataInMem_hi_14 = _GEN_16;
  wire [15:0]      dataInMem_lo_hi_17;
  assign dataInMem_lo_hi_17 = _GEN_16;
  wire [15:0]      dataInMem_lo_hi_50;
  assign dataInMem_lo_hi_50 = _GEN_16;
  wire [15:0]      _GEN_17 = {dataRegroupBySew_2_13, dataRegroupBySew_1_13};
  wire [15:0]      dataInMem_hi_15;
  assign dataInMem_hi_15 = _GEN_17;
  wire [15:0]      dataInMem_lo_hi_18;
  assign dataInMem_lo_hi_18 = _GEN_17;
  wire [15:0]      dataInMem_lo_hi_51;
  assign dataInMem_lo_hi_51 = _GEN_17;
  wire [15:0]      _GEN_18 = {dataRegroupBySew_2_14, dataRegroupBySew_1_14};
  wire [15:0]      dataInMem_hi_16;
  assign dataInMem_hi_16 = _GEN_18;
  wire [15:0]      dataInMem_lo_hi_19;
  assign dataInMem_lo_hi_19 = _GEN_18;
  wire [15:0]      dataInMem_lo_hi_52;
  assign dataInMem_lo_hi_52 = _GEN_18;
  wire [15:0]      _GEN_19 = {dataRegroupBySew_2_15, dataRegroupBySew_1_15};
  wire [15:0]      dataInMem_hi_17;
  assign dataInMem_hi_17 = _GEN_19;
  wire [15:0]      dataInMem_lo_hi_20;
  assign dataInMem_lo_hi_20 = _GEN_19;
  wire [15:0]      dataInMem_lo_hi_53;
  assign dataInMem_lo_hi_53 = _GEN_19;
  wire [15:0]      _GEN_20 = {dataRegroupBySew_2_16, dataRegroupBySew_1_16};
  wire [15:0]      dataInMem_hi_18;
  assign dataInMem_hi_18 = _GEN_20;
  wire [15:0]      dataInMem_lo_hi_21;
  assign dataInMem_lo_hi_21 = _GEN_20;
  wire [15:0]      dataInMem_lo_hi_54;
  assign dataInMem_lo_hi_54 = _GEN_20;
  wire [15:0]      _GEN_21 = {dataRegroupBySew_2_17, dataRegroupBySew_1_17};
  wire [15:0]      dataInMem_hi_19;
  assign dataInMem_hi_19 = _GEN_21;
  wire [15:0]      dataInMem_lo_hi_22;
  assign dataInMem_lo_hi_22 = _GEN_21;
  wire [15:0]      dataInMem_lo_hi_55;
  assign dataInMem_lo_hi_55 = _GEN_21;
  wire [15:0]      _GEN_22 = {dataRegroupBySew_2_18, dataRegroupBySew_1_18};
  wire [15:0]      dataInMem_hi_20;
  assign dataInMem_hi_20 = _GEN_22;
  wire [15:0]      dataInMem_lo_hi_23;
  assign dataInMem_lo_hi_23 = _GEN_22;
  wire [15:0]      dataInMem_lo_hi_56;
  assign dataInMem_lo_hi_56 = _GEN_22;
  wire [15:0]      _GEN_23 = {dataRegroupBySew_2_19, dataRegroupBySew_1_19};
  wire [15:0]      dataInMem_hi_21;
  assign dataInMem_hi_21 = _GEN_23;
  wire [15:0]      dataInMem_lo_hi_24;
  assign dataInMem_lo_hi_24 = _GEN_23;
  wire [15:0]      dataInMem_lo_hi_57;
  assign dataInMem_lo_hi_57 = _GEN_23;
  wire [15:0]      _GEN_24 = {dataRegroupBySew_2_20, dataRegroupBySew_1_20};
  wire [15:0]      dataInMem_hi_22;
  assign dataInMem_hi_22 = _GEN_24;
  wire [15:0]      dataInMem_lo_hi_25;
  assign dataInMem_lo_hi_25 = _GEN_24;
  wire [15:0]      dataInMem_lo_hi_58;
  assign dataInMem_lo_hi_58 = _GEN_24;
  wire [15:0]      _GEN_25 = {dataRegroupBySew_2_21, dataRegroupBySew_1_21};
  wire [15:0]      dataInMem_hi_23;
  assign dataInMem_hi_23 = _GEN_25;
  wire [15:0]      dataInMem_lo_hi_26;
  assign dataInMem_lo_hi_26 = _GEN_25;
  wire [15:0]      dataInMem_lo_hi_59;
  assign dataInMem_lo_hi_59 = _GEN_25;
  wire [15:0]      _GEN_26 = {dataRegroupBySew_2_22, dataRegroupBySew_1_22};
  wire [15:0]      dataInMem_hi_24;
  assign dataInMem_hi_24 = _GEN_26;
  wire [15:0]      dataInMem_lo_hi_27;
  assign dataInMem_lo_hi_27 = _GEN_26;
  wire [15:0]      dataInMem_lo_hi_60;
  assign dataInMem_lo_hi_60 = _GEN_26;
  wire [15:0]      _GEN_27 = {dataRegroupBySew_2_23, dataRegroupBySew_1_23};
  wire [15:0]      dataInMem_hi_25;
  assign dataInMem_hi_25 = _GEN_27;
  wire [15:0]      dataInMem_lo_hi_28;
  assign dataInMem_lo_hi_28 = _GEN_27;
  wire [15:0]      dataInMem_lo_hi_61;
  assign dataInMem_lo_hi_61 = _GEN_27;
  wire [15:0]      _GEN_28 = {dataRegroupBySew_2_24, dataRegroupBySew_1_24};
  wire [15:0]      dataInMem_hi_26;
  assign dataInMem_hi_26 = _GEN_28;
  wire [15:0]      dataInMem_lo_hi_29;
  assign dataInMem_lo_hi_29 = _GEN_28;
  wire [15:0]      dataInMem_lo_hi_62;
  assign dataInMem_lo_hi_62 = _GEN_28;
  wire [15:0]      _GEN_29 = {dataRegroupBySew_2_25, dataRegroupBySew_1_25};
  wire [15:0]      dataInMem_hi_27;
  assign dataInMem_hi_27 = _GEN_29;
  wire [15:0]      dataInMem_lo_hi_30;
  assign dataInMem_lo_hi_30 = _GEN_29;
  wire [15:0]      dataInMem_lo_hi_63;
  assign dataInMem_lo_hi_63 = _GEN_29;
  wire [15:0]      _GEN_30 = {dataRegroupBySew_2_26, dataRegroupBySew_1_26};
  wire [15:0]      dataInMem_hi_28;
  assign dataInMem_hi_28 = _GEN_30;
  wire [15:0]      dataInMem_lo_hi_31;
  assign dataInMem_lo_hi_31 = _GEN_30;
  wire [15:0]      dataInMem_lo_hi_64;
  assign dataInMem_lo_hi_64 = _GEN_30;
  wire [15:0]      _GEN_31 = {dataRegroupBySew_2_27, dataRegroupBySew_1_27};
  wire [15:0]      dataInMem_hi_29;
  assign dataInMem_hi_29 = _GEN_31;
  wire [15:0]      dataInMem_lo_hi_32;
  assign dataInMem_lo_hi_32 = _GEN_31;
  wire [15:0]      dataInMem_lo_hi_65;
  assign dataInMem_lo_hi_65 = _GEN_31;
  wire [15:0]      _GEN_32 = {dataRegroupBySew_2_28, dataRegroupBySew_1_28};
  wire [15:0]      dataInMem_hi_30;
  assign dataInMem_hi_30 = _GEN_32;
  wire [15:0]      dataInMem_lo_hi_33;
  assign dataInMem_lo_hi_33 = _GEN_32;
  wire [15:0]      dataInMem_lo_hi_66;
  assign dataInMem_lo_hi_66 = _GEN_32;
  wire [15:0]      _GEN_33 = {dataRegroupBySew_2_29, dataRegroupBySew_1_29};
  wire [15:0]      dataInMem_hi_31;
  assign dataInMem_hi_31 = _GEN_33;
  wire [15:0]      dataInMem_lo_hi_34;
  assign dataInMem_lo_hi_34 = _GEN_33;
  wire [15:0]      dataInMem_lo_hi_67;
  assign dataInMem_lo_hi_67 = _GEN_33;
  wire [15:0]      _GEN_34 = {dataRegroupBySew_2_30, dataRegroupBySew_1_30};
  wire [15:0]      dataInMem_hi_32;
  assign dataInMem_hi_32 = _GEN_34;
  wire [15:0]      dataInMem_lo_hi_35;
  assign dataInMem_lo_hi_35 = _GEN_34;
  wire [15:0]      dataInMem_lo_hi_68;
  assign dataInMem_lo_hi_68 = _GEN_34;
  wire [15:0]      _GEN_35 = {dataRegroupBySew_2_31, dataRegroupBySew_1_31};
  wire [15:0]      dataInMem_hi_33;
  assign dataInMem_hi_33 = _GEN_35;
  wire [15:0]      dataInMem_lo_hi_36;
  assign dataInMem_lo_hi_36 = _GEN_35;
  wire [15:0]      dataInMem_lo_hi_69;
  assign dataInMem_lo_hi_69 = _GEN_35;
  wire [47:0]      dataInMem_lo_lo_lo_lo_2 = {dataInMem_hi_3, dataRegroupBySew_0_1, dataInMem_hi_2, dataRegroupBySew_0_0};
  wire [47:0]      dataInMem_lo_lo_lo_hi_2 = {dataInMem_hi_5, dataRegroupBySew_0_3, dataInMem_hi_4, dataRegroupBySew_0_2};
  wire [95:0]      dataInMem_lo_lo_lo_2 = {dataInMem_lo_lo_lo_hi_2, dataInMem_lo_lo_lo_lo_2};
  wire [47:0]      dataInMem_lo_lo_hi_lo_2 = {dataInMem_hi_7, dataRegroupBySew_0_5, dataInMem_hi_6, dataRegroupBySew_0_4};
  wire [47:0]      dataInMem_lo_lo_hi_hi_2 = {dataInMem_hi_9, dataRegroupBySew_0_7, dataInMem_hi_8, dataRegroupBySew_0_6};
  wire [95:0]      dataInMem_lo_lo_hi_2 = {dataInMem_lo_lo_hi_hi_2, dataInMem_lo_lo_hi_lo_2};
  wire [191:0]     dataInMem_lo_lo_2 = {dataInMem_lo_lo_hi_2, dataInMem_lo_lo_lo_2};
  wire [47:0]      dataInMem_lo_hi_lo_lo_2 = {dataInMem_hi_11, dataRegroupBySew_0_9, dataInMem_hi_10, dataRegroupBySew_0_8};
  wire [47:0]      dataInMem_lo_hi_lo_hi_2 = {dataInMem_hi_13, dataRegroupBySew_0_11, dataInMem_hi_12, dataRegroupBySew_0_10};
  wire [95:0]      dataInMem_lo_hi_lo_2 = {dataInMem_lo_hi_lo_hi_2, dataInMem_lo_hi_lo_lo_2};
  wire [47:0]      dataInMem_lo_hi_hi_lo_2 = {dataInMem_hi_15, dataRegroupBySew_0_13, dataInMem_hi_14, dataRegroupBySew_0_12};
  wire [47:0]      dataInMem_lo_hi_hi_hi_2 = {dataInMem_hi_17, dataRegroupBySew_0_15, dataInMem_hi_16, dataRegroupBySew_0_14};
  wire [95:0]      dataInMem_lo_hi_hi_2 = {dataInMem_lo_hi_hi_hi_2, dataInMem_lo_hi_hi_lo_2};
  wire [191:0]     dataInMem_lo_hi_2 = {dataInMem_lo_hi_hi_2, dataInMem_lo_hi_lo_2};
  wire [383:0]     dataInMem_lo_2 = {dataInMem_lo_hi_2, dataInMem_lo_lo_2};
  wire [47:0]      dataInMem_hi_lo_lo_lo_2 = {dataInMem_hi_19, dataRegroupBySew_0_17, dataInMem_hi_18, dataRegroupBySew_0_16};
  wire [47:0]      dataInMem_hi_lo_lo_hi_2 = {dataInMem_hi_21, dataRegroupBySew_0_19, dataInMem_hi_20, dataRegroupBySew_0_18};
  wire [95:0]      dataInMem_hi_lo_lo_2 = {dataInMem_hi_lo_lo_hi_2, dataInMem_hi_lo_lo_lo_2};
  wire [47:0]      dataInMem_hi_lo_hi_lo_2 = {dataInMem_hi_23, dataRegroupBySew_0_21, dataInMem_hi_22, dataRegroupBySew_0_20};
  wire [47:0]      dataInMem_hi_lo_hi_hi_2 = {dataInMem_hi_25, dataRegroupBySew_0_23, dataInMem_hi_24, dataRegroupBySew_0_22};
  wire [95:0]      dataInMem_hi_lo_hi_2 = {dataInMem_hi_lo_hi_hi_2, dataInMem_hi_lo_hi_lo_2};
  wire [191:0]     dataInMem_hi_lo_2 = {dataInMem_hi_lo_hi_2, dataInMem_hi_lo_lo_2};
  wire [47:0]      dataInMem_hi_hi_lo_lo_2 = {dataInMem_hi_27, dataRegroupBySew_0_25, dataInMem_hi_26, dataRegroupBySew_0_24};
  wire [47:0]      dataInMem_hi_hi_lo_hi_2 = {dataInMem_hi_29, dataRegroupBySew_0_27, dataInMem_hi_28, dataRegroupBySew_0_26};
  wire [95:0]      dataInMem_hi_hi_lo_2 = {dataInMem_hi_hi_lo_hi_2, dataInMem_hi_hi_lo_lo_2};
  wire [47:0]      dataInMem_hi_hi_hi_lo_2 = {dataInMem_hi_31, dataRegroupBySew_0_29, dataInMem_hi_30, dataRegroupBySew_0_28};
  wire [47:0]      dataInMem_hi_hi_hi_hi_2 = {dataInMem_hi_33, dataRegroupBySew_0_31, dataInMem_hi_32, dataRegroupBySew_0_30};
  wire [95:0]      dataInMem_hi_hi_hi_2 = {dataInMem_hi_hi_hi_hi_2, dataInMem_hi_hi_hi_lo_2};
  wire [191:0]     dataInMem_hi_hi_2 = {dataInMem_hi_hi_hi_2, dataInMem_hi_hi_lo_2};
  wire [383:0]     dataInMem_hi_34 = {dataInMem_hi_hi_2, dataInMem_hi_lo_2};
  wire [767:0]     dataInMem_2 = {dataInMem_hi_34, dataInMem_lo_2};
  wire [255:0]     regroupCacheLine_2_0 = dataInMem_2[255:0];
  wire [255:0]     regroupCacheLine_2_1 = dataInMem_2[511:256];
  wire [255:0]     regroupCacheLine_2_2 = dataInMem_2[767:512];
  wire [255:0]     res_16 = regroupCacheLine_2_0;
  wire [255:0]     res_17 = regroupCacheLine_2_1;
  wire [255:0]     res_18 = regroupCacheLine_2_2;
  wire [511:0]     lo_lo_2 = {res_17, res_16};
  wire [511:0]     lo_hi_2 = {256'h0, res_18};
  wire [1023:0]    lo_2 = {lo_hi_2, lo_lo_2};
  wire [2047:0]    regroupLoadData_0_2 = {1024'h0, lo_2};
  wire [15:0]      _GEN_36 = {dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_lo_3;
  assign dataInMem_lo_3 = _GEN_36;
  wire [15:0]      dataInMem_lo_36;
  assign dataInMem_lo_36 = _GEN_36;
  wire [15:0]      dataInMem_lo_lo_7;
  assign dataInMem_lo_lo_7 = _GEN_36;
  wire [15:0]      _GEN_37 = {dataRegroupBySew_3_0, dataRegroupBySew_2_0};
  wire [15:0]      dataInMem_hi_35;
  assign dataInMem_hi_35 = _GEN_37;
  wire [15:0]      dataInMem_lo_hi_71;
  assign dataInMem_lo_hi_71 = _GEN_37;
  wire [15:0]      _GEN_38 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1};
  wire [15:0]      dataInMem_lo_4;
  assign dataInMem_lo_4 = _GEN_38;
  wire [15:0]      dataInMem_lo_37;
  assign dataInMem_lo_37 = _GEN_38;
  wire [15:0]      dataInMem_lo_lo_8;
  assign dataInMem_lo_lo_8 = _GEN_38;
  wire [15:0]      _GEN_39 = {dataRegroupBySew_3_1, dataRegroupBySew_2_1};
  wire [15:0]      dataInMem_hi_36;
  assign dataInMem_hi_36 = _GEN_39;
  wire [15:0]      dataInMem_lo_hi_72;
  assign dataInMem_lo_hi_72 = _GEN_39;
  wire [15:0]      _GEN_40 = {dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [15:0]      dataInMem_lo_5;
  assign dataInMem_lo_5 = _GEN_40;
  wire [15:0]      dataInMem_lo_38;
  assign dataInMem_lo_38 = _GEN_40;
  wire [15:0]      dataInMem_lo_lo_9;
  assign dataInMem_lo_lo_9 = _GEN_40;
  wire [15:0]      _GEN_41 = {dataRegroupBySew_3_2, dataRegroupBySew_2_2};
  wire [15:0]      dataInMem_hi_37;
  assign dataInMem_hi_37 = _GEN_41;
  wire [15:0]      dataInMem_lo_hi_73;
  assign dataInMem_lo_hi_73 = _GEN_41;
  wire [15:0]      _GEN_42 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3};
  wire [15:0]      dataInMem_lo_6;
  assign dataInMem_lo_6 = _GEN_42;
  wire [15:0]      dataInMem_lo_39;
  assign dataInMem_lo_39 = _GEN_42;
  wire [15:0]      dataInMem_lo_lo_10;
  assign dataInMem_lo_lo_10 = _GEN_42;
  wire [15:0]      _GEN_43 = {dataRegroupBySew_3_3, dataRegroupBySew_2_3};
  wire [15:0]      dataInMem_hi_38;
  assign dataInMem_hi_38 = _GEN_43;
  wire [15:0]      dataInMem_lo_hi_74;
  assign dataInMem_lo_hi_74 = _GEN_43;
  wire [15:0]      _GEN_44 = {dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_lo_7;
  assign dataInMem_lo_7 = _GEN_44;
  wire [15:0]      dataInMem_lo_40;
  assign dataInMem_lo_40 = _GEN_44;
  wire [15:0]      dataInMem_lo_lo_11;
  assign dataInMem_lo_lo_11 = _GEN_44;
  wire [15:0]      _GEN_45 = {dataRegroupBySew_3_4, dataRegroupBySew_2_4};
  wire [15:0]      dataInMem_hi_39;
  assign dataInMem_hi_39 = _GEN_45;
  wire [15:0]      dataInMem_lo_hi_75;
  assign dataInMem_lo_hi_75 = _GEN_45;
  wire [15:0]      _GEN_46 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5};
  wire [15:0]      dataInMem_lo_8;
  assign dataInMem_lo_8 = _GEN_46;
  wire [15:0]      dataInMem_lo_41;
  assign dataInMem_lo_41 = _GEN_46;
  wire [15:0]      dataInMem_lo_lo_12;
  assign dataInMem_lo_lo_12 = _GEN_46;
  wire [15:0]      _GEN_47 = {dataRegroupBySew_3_5, dataRegroupBySew_2_5};
  wire [15:0]      dataInMem_hi_40;
  assign dataInMem_hi_40 = _GEN_47;
  wire [15:0]      dataInMem_lo_hi_76;
  assign dataInMem_lo_hi_76 = _GEN_47;
  wire [15:0]      _GEN_48 = {dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [15:0]      dataInMem_lo_9;
  assign dataInMem_lo_9 = _GEN_48;
  wire [15:0]      dataInMem_lo_42;
  assign dataInMem_lo_42 = _GEN_48;
  wire [15:0]      dataInMem_lo_lo_13;
  assign dataInMem_lo_lo_13 = _GEN_48;
  wire [15:0]      _GEN_49 = {dataRegroupBySew_3_6, dataRegroupBySew_2_6};
  wire [15:0]      dataInMem_hi_41;
  assign dataInMem_hi_41 = _GEN_49;
  wire [15:0]      dataInMem_lo_hi_77;
  assign dataInMem_lo_hi_77 = _GEN_49;
  wire [15:0]      _GEN_50 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7};
  wire [15:0]      dataInMem_lo_10;
  assign dataInMem_lo_10 = _GEN_50;
  wire [15:0]      dataInMem_lo_43;
  assign dataInMem_lo_43 = _GEN_50;
  wire [15:0]      dataInMem_lo_lo_14;
  assign dataInMem_lo_lo_14 = _GEN_50;
  wire [15:0]      _GEN_51 = {dataRegroupBySew_3_7, dataRegroupBySew_2_7};
  wire [15:0]      dataInMem_hi_42;
  assign dataInMem_hi_42 = _GEN_51;
  wire [15:0]      dataInMem_lo_hi_78;
  assign dataInMem_lo_hi_78 = _GEN_51;
  wire [15:0]      _GEN_52 = {dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_lo_11;
  assign dataInMem_lo_11 = _GEN_52;
  wire [15:0]      dataInMem_lo_44;
  assign dataInMem_lo_44 = _GEN_52;
  wire [15:0]      dataInMem_lo_lo_15;
  assign dataInMem_lo_lo_15 = _GEN_52;
  wire [15:0]      _GEN_53 = {dataRegroupBySew_3_8, dataRegroupBySew_2_8};
  wire [15:0]      dataInMem_hi_43;
  assign dataInMem_hi_43 = _GEN_53;
  wire [15:0]      dataInMem_lo_hi_79;
  assign dataInMem_lo_hi_79 = _GEN_53;
  wire [15:0]      _GEN_54 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9};
  wire [15:0]      dataInMem_lo_12;
  assign dataInMem_lo_12 = _GEN_54;
  wire [15:0]      dataInMem_lo_45;
  assign dataInMem_lo_45 = _GEN_54;
  wire [15:0]      dataInMem_lo_lo_16;
  assign dataInMem_lo_lo_16 = _GEN_54;
  wire [15:0]      _GEN_55 = {dataRegroupBySew_3_9, dataRegroupBySew_2_9};
  wire [15:0]      dataInMem_hi_44;
  assign dataInMem_hi_44 = _GEN_55;
  wire [15:0]      dataInMem_lo_hi_80;
  assign dataInMem_lo_hi_80 = _GEN_55;
  wire [15:0]      _GEN_56 = {dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [15:0]      dataInMem_lo_13;
  assign dataInMem_lo_13 = _GEN_56;
  wire [15:0]      dataInMem_lo_46;
  assign dataInMem_lo_46 = _GEN_56;
  wire [15:0]      dataInMem_lo_lo_17;
  assign dataInMem_lo_lo_17 = _GEN_56;
  wire [15:0]      _GEN_57 = {dataRegroupBySew_3_10, dataRegroupBySew_2_10};
  wire [15:0]      dataInMem_hi_45;
  assign dataInMem_hi_45 = _GEN_57;
  wire [15:0]      dataInMem_lo_hi_81;
  assign dataInMem_lo_hi_81 = _GEN_57;
  wire [15:0]      _GEN_58 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11};
  wire [15:0]      dataInMem_lo_14;
  assign dataInMem_lo_14 = _GEN_58;
  wire [15:0]      dataInMem_lo_47;
  assign dataInMem_lo_47 = _GEN_58;
  wire [15:0]      dataInMem_lo_lo_18;
  assign dataInMem_lo_lo_18 = _GEN_58;
  wire [15:0]      _GEN_59 = {dataRegroupBySew_3_11, dataRegroupBySew_2_11};
  wire [15:0]      dataInMem_hi_46;
  assign dataInMem_hi_46 = _GEN_59;
  wire [15:0]      dataInMem_lo_hi_82;
  assign dataInMem_lo_hi_82 = _GEN_59;
  wire [15:0]      _GEN_60 = {dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_lo_15;
  assign dataInMem_lo_15 = _GEN_60;
  wire [15:0]      dataInMem_lo_48;
  assign dataInMem_lo_48 = _GEN_60;
  wire [15:0]      dataInMem_lo_lo_19;
  assign dataInMem_lo_lo_19 = _GEN_60;
  wire [15:0]      _GEN_61 = {dataRegroupBySew_3_12, dataRegroupBySew_2_12};
  wire [15:0]      dataInMem_hi_47;
  assign dataInMem_hi_47 = _GEN_61;
  wire [15:0]      dataInMem_lo_hi_83;
  assign dataInMem_lo_hi_83 = _GEN_61;
  wire [15:0]      _GEN_62 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13};
  wire [15:0]      dataInMem_lo_16;
  assign dataInMem_lo_16 = _GEN_62;
  wire [15:0]      dataInMem_lo_49;
  assign dataInMem_lo_49 = _GEN_62;
  wire [15:0]      dataInMem_lo_lo_20;
  assign dataInMem_lo_lo_20 = _GEN_62;
  wire [15:0]      _GEN_63 = {dataRegroupBySew_3_13, dataRegroupBySew_2_13};
  wire [15:0]      dataInMem_hi_48;
  assign dataInMem_hi_48 = _GEN_63;
  wire [15:0]      dataInMem_lo_hi_84;
  assign dataInMem_lo_hi_84 = _GEN_63;
  wire [15:0]      _GEN_64 = {dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [15:0]      dataInMem_lo_17;
  assign dataInMem_lo_17 = _GEN_64;
  wire [15:0]      dataInMem_lo_50;
  assign dataInMem_lo_50 = _GEN_64;
  wire [15:0]      dataInMem_lo_lo_21;
  assign dataInMem_lo_lo_21 = _GEN_64;
  wire [15:0]      _GEN_65 = {dataRegroupBySew_3_14, dataRegroupBySew_2_14};
  wire [15:0]      dataInMem_hi_49;
  assign dataInMem_hi_49 = _GEN_65;
  wire [15:0]      dataInMem_lo_hi_85;
  assign dataInMem_lo_hi_85 = _GEN_65;
  wire [15:0]      _GEN_66 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15};
  wire [15:0]      dataInMem_lo_18;
  assign dataInMem_lo_18 = _GEN_66;
  wire [15:0]      dataInMem_lo_51;
  assign dataInMem_lo_51 = _GEN_66;
  wire [15:0]      dataInMem_lo_lo_22;
  assign dataInMem_lo_lo_22 = _GEN_66;
  wire [15:0]      _GEN_67 = {dataRegroupBySew_3_15, dataRegroupBySew_2_15};
  wire [15:0]      dataInMem_hi_50;
  assign dataInMem_hi_50 = _GEN_67;
  wire [15:0]      dataInMem_lo_hi_86;
  assign dataInMem_lo_hi_86 = _GEN_67;
  wire [15:0]      _GEN_68 = {dataRegroupBySew_1_16, dataRegroupBySew_0_16};
  wire [15:0]      dataInMem_lo_19;
  assign dataInMem_lo_19 = _GEN_68;
  wire [15:0]      dataInMem_lo_52;
  assign dataInMem_lo_52 = _GEN_68;
  wire [15:0]      dataInMem_lo_lo_23;
  assign dataInMem_lo_lo_23 = _GEN_68;
  wire [15:0]      _GEN_69 = {dataRegroupBySew_3_16, dataRegroupBySew_2_16};
  wire [15:0]      dataInMem_hi_51;
  assign dataInMem_hi_51 = _GEN_69;
  wire [15:0]      dataInMem_lo_hi_87;
  assign dataInMem_lo_hi_87 = _GEN_69;
  wire [15:0]      _GEN_70 = {dataRegroupBySew_1_17, dataRegroupBySew_0_17};
  wire [15:0]      dataInMem_lo_20;
  assign dataInMem_lo_20 = _GEN_70;
  wire [15:0]      dataInMem_lo_53;
  assign dataInMem_lo_53 = _GEN_70;
  wire [15:0]      dataInMem_lo_lo_24;
  assign dataInMem_lo_lo_24 = _GEN_70;
  wire [15:0]      _GEN_71 = {dataRegroupBySew_3_17, dataRegroupBySew_2_17};
  wire [15:0]      dataInMem_hi_52;
  assign dataInMem_hi_52 = _GEN_71;
  wire [15:0]      dataInMem_lo_hi_88;
  assign dataInMem_lo_hi_88 = _GEN_71;
  wire [15:0]      _GEN_72 = {dataRegroupBySew_1_18, dataRegroupBySew_0_18};
  wire [15:0]      dataInMem_lo_21;
  assign dataInMem_lo_21 = _GEN_72;
  wire [15:0]      dataInMem_lo_54;
  assign dataInMem_lo_54 = _GEN_72;
  wire [15:0]      dataInMem_lo_lo_25;
  assign dataInMem_lo_lo_25 = _GEN_72;
  wire [15:0]      _GEN_73 = {dataRegroupBySew_3_18, dataRegroupBySew_2_18};
  wire [15:0]      dataInMem_hi_53;
  assign dataInMem_hi_53 = _GEN_73;
  wire [15:0]      dataInMem_lo_hi_89;
  assign dataInMem_lo_hi_89 = _GEN_73;
  wire [15:0]      _GEN_74 = {dataRegroupBySew_1_19, dataRegroupBySew_0_19};
  wire [15:0]      dataInMem_lo_22;
  assign dataInMem_lo_22 = _GEN_74;
  wire [15:0]      dataInMem_lo_55;
  assign dataInMem_lo_55 = _GEN_74;
  wire [15:0]      dataInMem_lo_lo_26;
  assign dataInMem_lo_lo_26 = _GEN_74;
  wire [15:0]      _GEN_75 = {dataRegroupBySew_3_19, dataRegroupBySew_2_19};
  wire [15:0]      dataInMem_hi_54;
  assign dataInMem_hi_54 = _GEN_75;
  wire [15:0]      dataInMem_lo_hi_90;
  assign dataInMem_lo_hi_90 = _GEN_75;
  wire [15:0]      _GEN_76 = {dataRegroupBySew_1_20, dataRegroupBySew_0_20};
  wire [15:0]      dataInMem_lo_23;
  assign dataInMem_lo_23 = _GEN_76;
  wire [15:0]      dataInMem_lo_56;
  assign dataInMem_lo_56 = _GEN_76;
  wire [15:0]      dataInMem_lo_lo_27;
  assign dataInMem_lo_lo_27 = _GEN_76;
  wire [15:0]      _GEN_77 = {dataRegroupBySew_3_20, dataRegroupBySew_2_20};
  wire [15:0]      dataInMem_hi_55;
  assign dataInMem_hi_55 = _GEN_77;
  wire [15:0]      dataInMem_lo_hi_91;
  assign dataInMem_lo_hi_91 = _GEN_77;
  wire [15:0]      _GEN_78 = {dataRegroupBySew_1_21, dataRegroupBySew_0_21};
  wire [15:0]      dataInMem_lo_24;
  assign dataInMem_lo_24 = _GEN_78;
  wire [15:0]      dataInMem_lo_57;
  assign dataInMem_lo_57 = _GEN_78;
  wire [15:0]      dataInMem_lo_lo_28;
  assign dataInMem_lo_lo_28 = _GEN_78;
  wire [15:0]      _GEN_79 = {dataRegroupBySew_3_21, dataRegroupBySew_2_21};
  wire [15:0]      dataInMem_hi_56;
  assign dataInMem_hi_56 = _GEN_79;
  wire [15:0]      dataInMem_lo_hi_92;
  assign dataInMem_lo_hi_92 = _GEN_79;
  wire [15:0]      _GEN_80 = {dataRegroupBySew_1_22, dataRegroupBySew_0_22};
  wire [15:0]      dataInMem_lo_25;
  assign dataInMem_lo_25 = _GEN_80;
  wire [15:0]      dataInMem_lo_58;
  assign dataInMem_lo_58 = _GEN_80;
  wire [15:0]      dataInMem_lo_lo_29;
  assign dataInMem_lo_lo_29 = _GEN_80;
  wire [15:0]      _GEN_81 = {dataRegroupBySew_3_22, dataRegroupBySew_2_22};
  wire [15:0]      dataInMem_hi_57;
  assign dataInMem_hi_57 = _GEN_81;
  wire [15:0]      dataInMem_lo_hi_93;
  assign dataInMem_lo_hi_93 = _GEN_81;
  wire [15:0]      _GEN_82 = {dataRegroupBySew_1_23, dataRegroupBySew_0_23};
  wire [15:0]      dataInMem_lo_26;
  assign dataInMem_lo_26 = _GEN_82;
  wire [15:0]      dataInMem_lo_59;
  assign dataInMem_lo_59 = _GEN_82;
  wire [15:0]      dataInMem_lo_lo_30;
  assign dataInMem_lo_lo_30 = _GEN_82;
  wire [15:0]      _GEN_83 = {dataRegroupBySew_3_23, dataRegroupBySew_2_23};
  wire [15:0]      dataInMem_hi_58;
  assign dataInMem_hi_58 = _GEN_83;
  wire [15:0]      dataInMem_lo_hi_94;
  assign dataInMem_lo_hi_94 = _GEN_83;
  wire [15:0]      _GEN_84 = {dataRegroupBySew_1_24, dataRegroupBySew_0_24};
  wire [15:0]      dataInMem_lo_27;
  assign dataInMem_lo_27 = _GEN_84;
  wire [15:0]      dataInMem_lo_60;
  assign dataInMem_lo_60 = _GEN_84;
  wire [15:0]      dataInMem_lo_lo_31;
  assign dataInMem_lo_lo_31 = _GEN_84;
  wire [15:0]      _GEN_85 = {dataRegroupBySew_3_24, dataRegroupBySew_2_24};
  wire [15:0]      dataInMem_hi_59;
  assign dataInMem_hi_59 = _GEN_85;
  wire [15:0]      dataInMem_lo_hi_95;
  assign dataInMem_lo_hi_95 = _GEN_85;
  wire [15:0]      _GEN_86 = {dataRegroupBySew_1_25, dataRegroupBySew_0_25};
  wire [15:0]      dataInMem_lo_28;
  assign dataInMem_lo_28 = _GEN_86;
  wire [15:0]      dataInMem_lo_61;
  assign dataInMem_lo_61 = _GEN_86;
  wire [15:0]      dataInMem_lo_lo_32;
  assign dataInMem_lo_lo_32 = _GEN_86;
  wire [15:0]      _GEN_87 = {dataRegroupBySew_3_25, dataRegroupBySew_2_25};
  wire [15:0]      dataInMem_hi_60;
  assign dataInMem_hi_60 = _GEN_87;
  wire [15:0]      dataInMem_lo_hi_96;
  assign dataInMem_lo_hi_96 = _GEN_87;
  wire [15:0]      _GEN_88 = {dataRegroupBySew_1_26, dataRegroupBySew_0_26};
  wire [15:0]      dataInMem_lo_29;
  assign dataInMem_lo_29 = _GEN_88;
  wire [15:0]      dataInMem_lo_62;
  assign dataInMem_lo_62 = _GEN_88;
  wire [15:0]      dataInMem_lo_lo_33;
  assign dataInMem_lo_lo_33 = _GEN_88;
  wire [15:0]      _GEN_89 = {dataRegroupBySew_3_26, dataRegroupBySew_2_26};
  wire [15:0]      dataInMem_hi_61;
  assign dataInMem_hi_61 = _GEN_89;
  wire [15:0]      dataInMem_lo_hi_97;
  assign dataInMem_lo_hi_97 = _GEN_89;
  wire [15:0]      _GEN_90 = {dataRegroupBySew_1_27, dataRegroupBySew_0_27};
  wire [15:0]      dataInMem_lo_30;
  assign dataInMem_lo_30 = _GEN_90;
  wire [15:0]      dataInMem_lo_63;
  assign dataInMem_lo_63 = _GEN_90;
  wire [15:0]      dataInMem_lo_lo_34;
  assign dataInMem_lo_lo_34 = _GEN_90;
  wire [15:0]      _GEN_91 = {dataRegroupBySew_3_27, dataRegroupBySew_2_27};
  wire [15:0]      dataInMem_hi_62;
  assign dataInMem_hi_62 = _GEN_91;
  wire [15:0]      dataInMem_lo_hi_98;
  assign dataInMem_lo_hi_98 = _GEN_91;
  wire [15:0]      _GEN_92 = {dataRegroupBySew_1_28, dataRegroupBySew_0_28};
  wire [15:0]      dataInMem_lo_31;
  assign dataInMem_lo_31 = _GEN_92;
  wire [15:0]      dataInMem_lo_64;
  assign dataInMem_lo_64 = _GEN_92;
  wire [15:0]      dataInMem_lo_lo_35;
  assign dataInMem_lo_lo_35 = _GEN_92;
  wire [15:0]      _GEN_93 = {dataRegroupBySew_3_28, dataRegroupBySew_2_28};
  wire [15:0]      dataInMem_hi_63;
  assign dataInMem_hi_63 = _GEN_93;
  wire [15:0]      dataInMem_lo_hi_99;
  assign dataInMem_lo_hi_99 = _GEN_93;
  wire [15:0]      _GEN_94 = {dataRegroupBySew_1_29, dataRegroupBySew_0_29};
  wire [15:0]      dataInMem_lo_32;
  assign dataInMem_lo_32 = _GEN_94;
  wire [15:0]      dataInMem_lo_65;
  assign dataInMem_lo_65 = _GEN_94;
  wire [15:0]      dataInMem_lo_lo_36;
  assign dataInMem_lo_lo_36 = _GEN_94;
  wire [15:0]      _GEN_95 = {dataRegroupBySew_3_29, dataRegroupBySew_2_29};
  wire [15:0]      dataInMem_hi_64;
  assign dataInMem_hi_64 = _GEN_95;
  wire [15:0]      dataInMem_lo_hi_100;
  assign dataInMem_lo_hi_100 = _GEN_95;
  wire [15:0]      _GEN_96 = {dataRegroupBySew_1_30, dataRegroupBySew_0_30};
  wire [15:0]      dataInMem_lo_33;
  assign dataInMem_lo_33 = _GEN_96;
  wire [15:0]      dataInMem_lo_66;
  assign dataInMem_lo_66 = _GEN_96;
  wire [15:0]      dataInMem_lo_lo_37;
  assign dataInMem_lo_lo_37 = _GEN_96;
  wire [15:0]      _GEN_97 = {dataRegroupBySew_3_30, dataRegroupBySew_2_30};
  wire [15:0]      dataInMem_hi_65;
  assign dataInMem_hi_65 = _GEN_97;
  wire [15:0]      dataInMem_lo_hi_101;
  assign dataInMem_lo_hi_101 = _GEN_97;
  wire [15:0]      _GEN_98 = {dataRegroupBySew_1_31, dataRegroupBySew_0_31};
  wire [15:0]      dataInMem_lo_34;
  assign dataInMem_lo_34 = _GEN_98;
  wire [15:0]      dataInMem_lo_67;
  assign dataInMem_lo_67 = _GEN_98;
  wire [15:0]      dataInMem_lo_lo_38;
  assign dataInMem_lo_lo_38 = _GEN_98;
  wire [15:0]      _GEN_99 = {dataRegroupBySew_3_31, dataRegroupBySew_2_31};
  wire [15:0]      dataInMem_hi_66;
  assign dataInMem_hi_66 = _GEN_99;
  wire [15:0]      dataInMem_lo_hi_102;
  assign dataInMem_lo_hi_102 = _GEN_99;
  wire [63:0]      dataInMem_lo_lo_lo_lo_3 = {dataInMem_hi_36, dataInMem_lo_4, dataInMem_hi_35, dataInMem_lo_3};
  wire [63:0]      dataInMem_lo_lo_lo_hi_3 = {dataInMem_hi_38, dataInMem_lo_6, dataInMem_hi_37, dataInMem_lo_5};
  wire [127:0]     dataInMem_lo_lo_lo_3 = {dataInMem_lo_lo_lo_hi_3, dataInMem_lo_lo_lo_lo_3};
  wire [63:0]      dataInMem_lo_lo_hi_lo_3 = {dataInMem_hi_40, dataInMem_lo_8, dataInMem_hi_39, dataInMem_lo_7};
  wire [63:0]      dataInMem_lo_lo_hi_hi_3 = {dataInMem_hi_42, dataInMem_lo_10, dataInMem_hi_41, dataInMem_lo_9};
  wire [127:0]     dataInMem_lo_lo_hi_3 = {dataInMem_lo_lo_hi_hi_3, dataInMem_lo_lo_hi_lo_3};
  wire [255:0]     dataInMem_lo_lo_3 = {dataInMem_lo_lo_hi_3, dataInMem_lo_lo_lo_3};
  wire [63:0]      dataInMem_lo_hi_lo_lo_3 = {dataInMem_hi_44, dataInMem_lo_12, dataInMem_hi_43, dataInMem_lo_11};
  wire [63:0]      dataInMem_lo_hi_lo_hi_3 = {dataInMem_hi_46, dataInMem_lo_14, dataInMem_hi_45, dataInMem_lo_13};
  wire [127:0]     dataInMem_lo_hi_lo_3 = {dataInMem_lo_hi_lo_hi_3, dataInMem_lo_hi_lo_lo_3};
  wire [63:0]      dataInMem_lo_hi_hi_lo_3 = {dataInMem_hi_48, dataInMem_lo_16, dataInMem_hi_47, dataInMem_lo_15};
  wire [63:0]      dataInMem_lo_hi_hi_hi_3 = {dataInMem_hi_50, dataInMem_lo_18, dataInMem_hi_49, dataInMem_lo_17};
  wire [127:0]     dataInMem_lo_hi_hi_3 = {dataInMem_lo_hi_hi_hi_3, dataInMem_lo_hi_hi_lo_3};
  wire [255:0]     dataInMem_lo_hi_3 = {dataInMem_lo_hi_hi_3, dataInMem_lo_hi_lo_3};
  wire [511:0]     dataInMem_lo_35 = {dataInMem_lo_hi_3, dataInMem_lo_lo_3};
  wire [63:0]      dataInMem_hi_lo_lo_lo_3 = {dataInMem_hi_52, dataInMem_lo_20, dataInMem_hi_51, dataInMem_lo_19};
  wire [63:0]      dataInMem_hi_lo_lo_hi_3 = {dataInMem_hi_54, dataInMem_lo_22, dataInMem_hi_53, dataInMem_lo_21};
  wire [127:0]     dataInMem_hi_lo_lo_3 = {dataInMem_hi_lo_lo_hi_3, dataInMem_hi_lo_lo_lo_3};
  wire [63:0]      dataInMem_hi_lo_hi_lo_3 = {dataInMem_hi_56, dataInMem_lo_24, dataInMem_hi_55, dataInMem_lo_23};
  wire [63:0]      dataInMem_hi_lo_hi_hi_3 = {dataInMem_hi_58, dataInMem_lo_26, dataInMem_hi_57, dataInMem_lo_25};
  wire [127:0]     dataInMem_hi_lo_hi_3 = {dataInMem_hi_lo_hi_hi_3, dataInMem_hi_lo_hi_lo_3};
  wire [255:0]     dataInMem_hi_lo_3 = {dataInMem_hi_lo_hi_3, dataInMem_hi_lo_lo_3};
  wire [63:0]      dataInMem_hi_hi_lo_lo_3 = {dataInMem_hi_60, dataInMem_lo_28, dataInMem_hi_59, dataInMem_lo_27};
  wire [63:0]      dataInMem_hi_hi_lo_hi_3 = {dataInMem_hi_62, dataInMem_lo_30, dataInMem_hi_61, dataInMem_lo_29};
  wire [127:0]     dataInMem_hi_hi_lo_3 = {dataInMem_hi_hi_lo_hi_3, dataInMem_hi_hi_lo_lo_3};
  wire [63:0]      dataInMem_hi_hi_hi_lo_3 = {dataInMem_hi_64, dataInMem_lo_32, dataInMem_hi_63, dataInMem_lo_31};
  wire [63:0]      dataInMem_hi_hi_hi_hi_3 = {dataInMem_hi_66, dataInMem_lo_34, dataInMem_hi_65, dataInMem_lo_33};
  wire [127:0]     dataInMem_hi_hi_hi_3 = {dataInMem_hi_hi_hi_hi_3, dataInMem_hi_hi_hi_lo_3};
  wire [255:0]     dataInMem_hi_hi_3 = {dataInMem_hi_hi_hi_3, dataInMem_hi_hi_lo_3};
  wire [511:0]     dataInMem_hi_67 = {dataInMem_hi_hi_3, dataInMem_hi_lo_3};
  wire [1023:0]    dataInMem_3 = {dataInMem_hi_67, dataInMem_lo_35};
  wire [255:0]     regroupCacheLine_3_0 = dataInMem_3[255:0];
  wire [255:0]     regroupCacheLine_3_1 = dataInMem_3[511:256];
  wire [255:0]     regroupCacheLine_3_2 = dataInMem_3[767:512];
  wire [255:0]     regroupCacheLine_3_3 = dataInMem_3[1023:768];
  wire [255:0]     res_24 = regroupCacheLine_3_0;
  wire [255:0]     res_25 = regroupCacheLine_3_1;
  wire [255:0]     res_26 = regroupCacheLine_3_2;
  wire [255:0]     res_27 = regroupCacheLine_3_3;
  wire [511:0]     lo_lo_3 = {res_25, res_24};
  wire [511:0]     lo_hi_3 = {res_27, res_26};
  wire [1023:0]    lo_3 = {lo_hi_3, lo_lo_3};
  wire [2047:0]    regroupLoadData_0_3 = {1024'h0, lo_3};
  wire [15:0]      _GEN_100 = {dataRegroupBySew_4_0, dataRegroupBySew_3_0};
  wire [15:0]      dataInMem_hi_hi_4;
  assign dataInMem_hi_hi_4 = _GEN_100;
  wire [15:0]      dataInMem_hi_lo_6;
  assign dataInMem_hi_lo_6 = _GEN_100;
  wire [23:0]      dataInMem_hi_68 = {dataInMem_hi_hi_4, dataRegroupBySew_2_0};
  wire [15:0]      _GEN_101 = {dataRegroupBySew_4_1, dataRegroupBySew_3_1};
  wire [15:0]      dataInMem_hi_hi_5;
  assign dataInMem_hi_hi_5 = _GEN_101;
  wire [15:0]      dataInMem_hi_lo_7;
  assign dataInMem_hi_lo_7 = _GEN_101;
  wire [23:0]      dataInMem_hi_69 = {dataInMem_hi_hi_5, dataRegroupBySew_2_1};
  wire [15:0]      _GEN_102 = {dataRegroupBySew_4_2, dataRegroupBySew_3_2};
  wire [15:0]      dataInMem_hi_hi_6;
  assign dataInMem_hi_hi_6 = _GEN_102;
  wire [15:0]      dataInMem_hi_lo_8;
  assign dataInMem_hi_lo_8 = _GEN_102;
  wire [23:0]      dataInMem_hi_70 = {dataInMem_hi_hi_6, dataRegroupBySew_2_2};
  wire [15:0]      _GEN_103 = {dataRegroupBySew_4_3, dataRegroupBySew_3_3};
  wire [15:0]      dataInMem_hi_hi_7;
  assign dataInMem_hi_hi_7 = _GEN_103;
  wire [15:0]      dataInMem_hi_lo_9;
  assign dataInMem_hi_lo_9 = _GEN_103;
  wire [23:0]      dataInMem_hi_71 = {dataInMem_hi_hi_7, dataRegroupBySew_2_3};
  wire [15:0]      _GEN_104 = {dataRegroupBySew_4_4, dataRegroupBySew_3_4};
  wire [15:0]      dataInMem_hi_hi_8;
  assign dataInMem_hi_hi_8 = _GEN_104;
  wire [15:0]      dataInMem_hi_lo_10;
  assign dataInMem_hi_lo_10 = _GEN_104;
  wire [23:0]      dataInMem_hi_72 = {dataInMem_hi_hi_8, dataRegroupBySew_2_4};
  wire [15:0]      _GEN_105 = {dataRegroupBySew_4_5, dataRegroupBySew_3_5};
  wire [15:0]      dataInMem_hi_hi_9;
  assign dataInMem_hi_hi_9 = _GEN_105;
  wire [15:0]      dataInMem_hi_lo_11;
  assign dataInMem_hi_lo_11 = _GEN_105;
  wire [23:0]      dataInMem_hi_73 = {dataInMem_hi_hi_9, dataRegroupBySew_2_5};
  wire [15:0]      _GEN_106 = {dataRegroupBySew_4_6, dataRegroupBySew_3_6};
  wire [15:0]      dataInMem_hi_hi_10;
  assign dataInMem_hi_hi_10 = _GEN_106;
  wire [15:0]      dataInMem_hi_lo_12;
  assign dataInMem_hi_lo_12 = _GEN_106;
  wire [23:0]      dataInMem_hi_74 = {dataInMem_hi_hi_10, dataRegroupBySew_2_6};
  wire [15:0]      _GEN_107 = {dataRegroupBySew_4_7, dataRegroupBySew_3_7};
  wire [15:0]      dataInMem_hi_hi_11;
  assign dataInMem_hi_hi_11 = _GEN_107;
  wire [15:0]      dataInMem_hi_lo_13;
  assign dataInMem_hi_lo_13 = _GEN_107;
  wire [23:0]      dataInMem_hi_75 = {dataInMem_hi_hi_11, dataRegroupBySew_2_7};
  wire [15:0]      _GEN_108 = {dataRegroupBySew_4_8, dataRegroupBySew_3_8};
  wire [15:0]      dataInMem_hi_hi_12;
  assign dataInMem_hi_hi_12 = _GEN_108;
  wire [15:0]      dataInMem_hi_lo_14;
  assign dataInMem_hi_lo_14 = _GEN_108;
  wire [23:0]      dataInMem_hi_76 = {dataInMem_hi_hi_12, dataRegroupBySew_2_8};
  wire [15:0]      _GEN_109 = {dataRegroupBySew_4_9, dataRegroupBySew_3_9};
  wire [15:0]      dataInMem_hi_hi_13;
  assign dataInMem_hi_hi_13 = _GEN_109;
  wire [15:0]      dataInMem_hi_lo_15;
  assign dataInMem_hi_lo_15 = _GEN_109;
  wire [23:0]      dataInMem_hi_77 = {dataInMem_hi_hi_13, dataRegroupBySew_2_9};
  wire [15:0]      _GEN_110 = {dataRegroupBySew_4_10, dataRegroupBySew_3_10};
  wire [15:0]      dataInMem_hi_hi_14;
  assign dataInMem_hi_hi_14 = _GEN_110;
  wire [15:0]      dataInMem_hi_lo_16;
  assign dataInMem_hi_lo_16 = _GEN_110;
  wire [23:0]      dataInMem_hi_78 = {dataInMem_hi_hi_14, dataRegroupBySew_2_10};
  wire [15:0]      _GEN_111 = {dataRegroupBySew_4_11, dataRegroupBySew_3_11};
  wire [15:0]      dataInMem_hi_hi_15;
  assign dataInMem_hi_hi_15 = _GEN_111;
  wire [15:0]      dataInMem_hi_lo_17;
  assign dataInMem_hi_lo_17 = _GEN_111;
  wire [23:0]      dataInMem_hi_79 = {dataInMem_hi_hi_15, dataRegroupBySew_2_11};
  wire [15:0]      _GEN_112 = {dataRegroupBySew_4_12, dataRegroupBySew_3_12};
  wire [15:0]      dataInMem_hi_hi_16;
  assign dataInMem_hi_hi_16 = _GEN_112;
  wire [15:0]      dataInMem_hi_lo_18;
  assign dataInMem_hi_lo_18 = _GEN_112;
  wire [23:0]      dataInMem_hi_80 = {dataInMem_hi_hi_16, dataRegroupBySew_2_12};
  wire [15:0]      _GEN_113 = {dataRegroupBySew_4_13, dataRegroupBySew_3_13};
  wire [15:0]      dataInMem_hi_hi_17;
  assign dataInMem_hi_hi_17 = _GEN_113;
  wire [15:0]      dataInMem_hi_lo_19;
  assign dataInMem_hi_lo_19 = _GEN_113;
  wire [23:0]      dataInMem_hi_81 = {dataInMem_hi_hi_17, dataRegroupBySew_2_13};
  wire [15:0]      _GEN_114 = {dataRegroupBySew_4_14, dataRegroupBySew_3_14};
  wire [15:0]      dataInMem_hi_hi_18;
  assign dataInMem_hi_hi_18 = _GEN_114;
  wire [15:0]      dataInMem_hi_lo_20;
  assign dataInMem_hi_lo_20 = _GEN_114;
  wire [23:0]      dataInMem_hi_82 = {dataInMem_hi_hi_18, dataRegroupBySew_2_14};
  wire [15:0]      _GEN_115 = {dataRegroupBySew_4_15, dataRegroupBySew_3_15};
  wire [15:0]      dataInMem_hi_hi_19;
  assign dataInMem_hi_hi_19 = _GEN_115;
  wire [15:0]      dataInMem_hi_lo_21;
  assign dataInMem_hi_lo_21 = _GEN_115;
  wire [23:0]      dataInMem_hi_83 = {dataInMem_hi_hi_19, dataRegroupBySew_2_15};
  wire [15:0]      _GEN_116 = {dataRegroupBySew_4_16, dataRegroupBySew_3_16};
  wire [15:0]      dataInMem_hi_hi_20;
  assign dataInMem_hi_hi_20 = _GEN_116;
  wire [15:0]      dataInMem_hi_lo_22;
  assign dataInMem_hi_lo_22 = _GEN_116;
  wire [23:0]      dataInMem_hi_84 = {dataInMem_hi_hi_20, dataRegroupBySew_2_16};
  wire [15:0]      _GEN_117 = {dataRegroupBySew_4_17, dataRegroupBySew_3_17};
  wire [15:0]      dataInMem_hi_hi_21;
  assign dataInMem_hi_hi_21 = _GEN_117;
  wire [15:0]      dataInMem_hi_lo_23;
  assign dataInMem_hi_lo_23 = _GEN_117;
  wire [23:0]      dataInMem_hi_85 = {dataInMem_hi_hi_21, dataRegroupBySew_2_17};
  wire [15:0]      _GEN_118 = {dataRegroupBySew_4_18, dataRegroupBySew_3_18};
  wire [15:0]      dataInMem_hi_hi_22;
  assign dataInMem_hi_hi_22 = _GEN_118;
  wire [15:0]      dataInMem_hi_lo_24;
  assign dataInMem_hi_lo_24 = _GEN_118;
  wire [23:0]      dataInMem_hi_86 = {dataInMem_hi_hi_22, dataRegroupBySew_2_18};
  wire [15:0]      _GEN_119 = {dataRegroupBySew_4_19, dataRegroupBySew_3_19};
  wire [15:0]      dataInMem_hi_hi_23;
  assign dataInMem_hi_hi_23 = _GEN_119;
  wire [15:0]      dataInMem_hi_lo_25;
  assign dataInMem_hi_lo_25 = _GEN_119;
  wire [23:0]      dataInMem_hi_87 = {dataInMem_hi_hi_23, dataRegroupBySew_2_19};
  wire [15:0]      _GEN_120 = {dataRegroupBySew_4_20, dataRegroupBySew_3_20};
  wire [15:0]      dataInMem_hi_hi_24;
  assign dataInMem_hi_hi_24 = _GEN_120;
  wire [15:0]      dataInMem_hi_lo_26;
  assign dataInMem_hi_lo_26 = _GEN_120;
  wire [23:0]      dataInMem_hi_88 = {dataInMem_hi_hi_24, dataRegroupBySew_2_20};
  wire [15:0]      _GEN_121 = {dataRegroupBySew_4_21, dataRegroupBySew_3_21};
  wire [15:0]      dataInMem_hi_hi_25;
  assign dataInMem_hi_hi_25 = _GEN_121;
  wire [15:0]      dataInMem_hi_lo_27;
  assign dataInMem_hi_lo_27 = _GEN_121;
  wire [23:0]      dataInMem_hi_89 = {dataInMem_hi_hi_25, dataRegroupBySew_2_21};
  wire [15:0]      _GEN_122 = {dataRegroupBySew_4_22, dataRegroupBySew_3_22};
  wire [15:0]      dataInMem_hi_hi_26;
  assign dataInMem_hi_hi_26 = _GEN_122;
  wire [15:0]      dataInMem_hi_lo_28;
  assign dataInMem_hi_lo_28 = _GEN_122;
  wire [23:0]      dataInMem_hi_90 = {dataInMem_hi_hi_26, dataRegroupBySew_2_22};
  wire [15:0]      _GEN_123 = {dataRegroupBySew_4_23, dataRegroupBySew_3_23};
  wire [15:0]      dataInMem_hi_hi_27;
  assign dataInMem_hi_hi_27 = _GEN_123;
  wire [15:0]      dataInMem_hi_lo_29;
  assign dataInMem_hi_lo_29 = _GEN_123;
  wire [23:0]      dataInMem_hi_91 = {dataInMem_hi_hi_27, dataRegroupBySew_2_23};
  wire [15:0]      _GEN_124 = {dataRegroupBySew_4_24, dataRegroupBySew_3_24};
  wire [15:0]      dataInMem_hi_hi_28;
  assign dataInMem_hi_hi_28 = _GEN_124;
  wire [15:0]      dataInMem_hi_lo_30;
  assign dataInMem_hi_lo_30 = _GEN_124;
  wire [23:0]      dataInMem_hi_92 = {dataInMem_hi_hi_28, dataRegroupBySew_2_24};
  wire [15:0]      _GEN_125 = {dataRegroupBySew_4_25, dataRegroupBySew_3_25};
  wire [15:0]      dataInMem_hi_hi_29;
  assign dataInMem_hi_hi_29 = _GEN_125;
  wire [15:0]      dataInMem_hi_lo_31;
  assign dataInMem_hi_lo_31 = _GEN_125;
  wire [23:0]      dataInMem_hi_93 = {dataInMem_hi_hi_29, dataRegroupBySew_2_25};
  wire [15:0]      _GEN_126 = {dataRegroupBySew_4_26, dataRegroupBySew_3_26};
  wire [15:0]      dataInMem_hi_hi_30;
  assign dataInMem_hi_hi_30 = _GEN_126;
  wire [15:0]      dataInMem_hi_lo_32;
  assign dataInMem_hi_lo_32 = _GEN_126;
  wire [23:0]      dataInMem_hi_94 = {dataInMem_hi_hi_30, dataRegroupBySew_2_26};
  wire [15:0]      _GEN_127 = {dataRegroupBySew_4_27, dataRegroupBySew_3_27};
  wire [15:0]      dataInMem_hi_hi_31;
  assign dataInMem_hi_hi_31 = _GEN_127;
  wire [15:0]      dataInMem_hi_lo_33;
  assign dataInMem_hi_lo_33 = _GEN_127;
  wire [23:0]      dataInMem_hi_95 = {dataInMem_hi_hi_31, dataRegroupBySew_2_27};
  wire [15:0]      _GEN_128 = {dataRegroupBySew_4_28, dataRegroupBySew_3_28};
  wire [15:0]      dataInMem_hi_hi_32;
  assign dataInMem_hi_hi_32 = _GEN_128;
  wire [15:0]      dataInMem_hi_lo_34;
  assign dataInMem_hi_lo_34 = _GEN_128;
  wire [23:0]      dataInMem_hi_96 = {dataInMem_hi_hi_32, dataRegroupBySew_2_28};
  wire [15:0]      _GEN_129 = {dataRegroupBySew_4_29, dataRegroupBySew_3_29};
  wire [15:0]      dataInMem_hi_hi_33;
  assign dataInMem_hi_hi_33 = _GEN_129;
  wire [15:0]      dataInMem_hi_lo_35;
  assign dataInMem_hi_lo_35 = _GEN_129;
  wire [23:0]      dataInMem_hi_97 = {dataInMem_hi_hi_33, dataRegroupBySew_2_29};
  wire [15:0]      _GEN_130 = {dataRegroupBySew_4_30, dataRegroupBySew_3_30};
  wire [15:0]      dataInMem_hi_hi_34;
  assign dataInMem_hi_hi_34 = _GEN_130;
  wire [15:0]      dataInMem_hi_lo_36;
  assign dataInMem_hi_lo_36 = _GEN_130;
  wire [23:0]      dataInMem_hi_98 = {dataInMem_hi_hi_34, dataRegroupBySew_2_30};
  wire [15:0]      _GEN_131 = {dataRegroupBySew_4_31, dataRegroupBySew_3_31};
  wire [15:0]      dataInMem_hi_hi_35;
  assign dataInMem_hi_hi_35 = _GEN_131;
  wire [15:0]      dataInMem_hi_lo_37;
  assign dataInMem_hi_lo_37 = _GEN_131;
  wire [23:0]      dataInMem_hi_99 = {dataInMem_hi_hi_35, dataRegroupBySew_2_31};
  wire [79:0]      dataInMem_lo_lo_lo_lo_4 = {dataInMem_hi_69, dataInMem_lo_37, dataInMem_hi_68, dataInMem_lo_36};
  wire [79:0]      dataInMem_lo_lo_lo_hi_4 = {dataInMem_hi_71, dataInMem_lo_39, dataInMem_hi_70, dataInMem_lo_38};
  wire [159:0]     dataInMem_lo_lo_lo_4 = {dataInMem_lo_lo_lo_hi_4, dataInMem_lo_lo_lo_lo_4};
  wire [79:0]      dataInMem_lo_lo_hi_lo_4 = {dataInMem_hi_73, dataInMem_lo_41, dataInMem_hi_72, dataInMem_lo_40};
  wire [79:0]      dataInMem_lo_lo_hi_hi_4 = {dataInMem_hi_75, dataInMem_lo_43, dataInMem_hi_74, dataInMem_lo_42};
  wire [159:0]     dataInMem_lo_lo_hi_4 = {dataInMem_lo_lo_hi_hi_4, dataInMem_lo_lo_hi_lo_4};
  wire [319:0]     dataInMem_lo_lo_4 = {dataInMem_lo_lo_hi_4, dataInMem_lo_lo_lo_4};
  wire [79:0]      dataInMem_lo_hi_lo_lo_4 = {dataInMem_hi_77, dataInMem_lo_45, dataInMem_hi_76, dataInMem_lo_44};
  wire [79:0]      dataInMem_lo_hi_lo_hi_4 = {dataInMem_hi_79, dataInMem_lo_47, dataInMem_hi_78, dataInMem_lo_46};
  wire [159:0]     dataInMem_lo_hi_lo_4 = {dataInMem_lo_hi_lo_hi_4, dataInMem_lo_hi_lo_lo_4};
  wire [79:0]      dataInMem_lo_hi_hi_lo_4 = {dataInMem_hi_81, dataInMem_lo_49, dataInMem_hi_80, dataInMem_lo_48};
  wire [79:0]      dataInMem_lo_hi_hi_hi_4 = {dataInMem_hi_83, dataInMem_lo_51, dataInMem_hi_82, dataInMem_lo_50};
  wire [159:0]     dataInMem_lo_hi_hi_4 = {dataInMem_lo_hi_hi_hi_4, dataInMem_lo_hi_hi_lo_4};
  wire [319:0]     dataInMem_lo_hi_4 = {dataInMem_lo_hi_hi_4, dataInMem_lo_hi_lo_4};
  wire [639:0]     dataInMem_lo_68 = {dataInMem_lo_hi_4, dataInMem_lo_lo_4};
  wire [79:0]      dataInMem_hi_lo_lo_lo_4 = {dataInMem_hi_85, dataInMem_lo_53, dataInMem_hi_84, dataInMem_lo_52};
  wire [79:0]      dataInMem_hi_lo_lo_hi_4 = {dataInMem_hi_87, dataInMem_lo_55, dataInMem_hi_86, dataInMem_lo_54};
  wire [159:0]     dataInMem_hi_lo_lo_4 = {dataInMem_hi_lo_lo_hi_4, dataInMem_hi_lo_lo_lo_4};
  wire [79:0]      dataInMem_hi_lo_hi_lo_4 = {dataInMem_hi_89, dataInMem_lo_57, dataInMem_hi_88, dataInMem_lo_56};
  wire [79:0]      dataInMem_hi_lo_hi_hi_4 = {dataInMem_hi_91, dataInMem_lo_59, dataInMem_hi_90, dataInMem_lo_58};
  wire [159:0]     dataInMem_hi_lo_hi_4 = {dataInMem_hi_lo_hi_hi_4, dataInMem_hi_lo_hi_lo_4};
  wire [319:0]     dataInMem_hi_lo_4 = {dataInMem_hi_lo_hi_4, dataInMem_hi_lo_lo_4};
  wire [79:0]      dataInMem_hi_hi_lo_lo_4 = {dataInMem_hi_93, dataInMem_lo_61, dataInMem_hi_92, dataInMem_lo_60};
  wire [79:0]      dataInMem_hi_hi_lo_hi_4 = {dataInMem_hi_95, dataInMem_lo_63, dataInMem_hi_94, dataInMem_lo_62};
  wire [159:0]     dataInMem_hi_hi_lo_4 = {dataInMem_hi_hi_lo_hi_4, dataInMem_hi_hi_lo_lo_4};
  wire [79:0]      dataInMem_hi_hi_hi_lo_4 = {dataInMem_hi_97, dataInMem_lo_65, dataInMem_hi_96, dataInMem_lo_64};
  wire [79:0]      dataInMem_hi_hi_hi_hi_4 = {dataInMem_hi_99, dataInMem_lo_67, dataInMem_hi_98, dataInMem_lo_66};
  wire [159:0]     dataInMem_hi_hi_hi_4 = {dataInMem_hi_hi_hi_hi_4, dataInMem_hi_hi_hi_lo_4};
  wire [319:0]     dataInMem_hi_hi_36 = {dataInMem_hi_hi_hi_4, dataInMem_hi_hi_lo_4};
  wire [639:0]     dataInMem_hi_100 = {dataInMem_hi_hi_36, dataInMem_hi_lo_4};
  wire [1279:0]    dataInMem_4 = {dataInMem_hi_100, dataInMem_lo_68};
  wire [255:0]     regroupCacheLine_4_0 = dataInMem_4[255:0];
  wire [255:0]     regroupCacheLine_4_1 = dataInMem_4[511:256];
  wire [255:0]     regroupCacheLine_4_2 = dataInMem_4[767:512];
  wire [255:0]     regroupCacheLine_4_3 = dataInMem_4[1023:768];
  wire [255:0]     regroupCacheLine_4_4 = dataInMem_4[1279:1024];
  wire [255:0]     res_32 = regroupCacheLine_4_0;
  wire [255:0]     res_33 = regroupCacheLine_4_1;
  wire [255:0]     res_34 = regroupCacheLine_4_2;
  wire [255:0]     res_35 = regroupCacheLine_4_3;
  wire [255:0]     res_36 = regroupCacheLine_4_4;
  wire [511:0]     lo_lo_4 = {res_33, res_32};
  wire [511:0]     lo_hi_4 = {res_35, res_34};
  wire [1023:0]    lo_4 = {lo_hi_4, lo_lo_4};
  wire [511:0]     hi_lo_4 = {256'h0, res_36};
  wire [1023:0]    hi_4 = {512'h0, hi_lo_4};
  wire [2047:0]    regroupLoadData_0_4 = {hi_4, lo_4};
  wire [23:0]      dataInMem_lo_69 = {dataInMem_lo_hi_5, dataRegroupBySew_0_0};
  wire [15:0]      _GEN_132 = {dataRegroupBySew_5_0, dataRegroupBySew_4_0};
  wire [15:0]      dataInMem_hi_hi_37;
  assign dataInMem_hi_hi_37 = _GEN_132;
  wire [15:0]      dataInMem_hi_lo_39;
  assign dataInMem_hi_lo_39 = _GEN_132;
  wire [23:0]      dataInMem_hi_101 = {dataInMem_hi_hi_37, dataRegroupBySew_3_0};
  wire [23:0]      dataInMem_lo_70 = {dataInMem_lo_hi_6, dataRegroupBySew_0_1};
  wire [15:0]      _GEN_133 = {dataRegroupBySew_5_1, dataRegroupBySew_4_1};
  wire [15:0]      dataInMem_hi_hi_38;
  assign dataInMem_hi_hi_38 = _GEN_133;
  wire [15:0]      dataInMem_hi_lo_40;
  assign dataInMem_hi_lo_40 = _GEN_133;
  wire [23:0]      dataInMem_hi_102 = {dataInMem_hi_hi_38, dataRegroupBySew_3_1};
  wire [23:0]      dataInMem_lo_71 = {dataInMem_lo_hi_7, dataRegroupBySew_0_2};
  wire [15:0]      _GEN_134 = {dataRegroupBySew_5_2, dataRegroupBySew_4_2};
  wire [15:0]      dataInMem_hi_hi_39;
  assign dataInMem_hi_hi_39 = _GEN_134;
  wire [15:0]      dataInMem_hi_lo_41;
  assign dataInMem_hi_lo_41 = _GEN_134;
  wire [23:0]      dataInMem_hi_103 = {dataInMem_hi_hi_39, dataRegroupBySew_3_2};
  wire [23:0]      dataInMem_lo_72 = {dataInMem_lo_hi_8, dataRegroupBySew_0_3};
  wire [15:0]      _GEN_135 = {dataRegroupBySew_5_3, dataRegroupBySew_4_3};
  wire [15:0]      dataInMem_hi_hi_40;
  assign dataInMem_hi_hi_40 = _GEN_135;
  wire [15:0]      dataInMem_hi_lo_42;
  assign dataInMem_hi_lo_42 = _GEN_135;
  wire [23:0]      dataInMem_hi_104 = {dataInMem_hi_hi_40, dataRegroupBySew_3_3};
  wire [23:0]      dataInMem_lo_73 = {dataInMem_lo_hi_9, dataRegroupBySew_0_4};
  wire [15:0]      _GEN_136 = {dataRegroupBySew_5_4, dataRegroupBySew_4_4};
  wire [15:0]      dataInMem_hi_hi_41;
  assign dataInMem_hi_hi_41 = _GEN_136;
  wire [15:0]      dataInMem_hi_lo_43;
  assign dataInMem_hi_lo_43 = _GEN_136;
  wire [23:0]      dataInMem_hi_105 = {dataInMem_hi_hi_41, dataRegroupBySew_3_4};
  wire [23:0]      dataInMem_lo_74 = {dataInMem_lo_hi_10, dataRegroupBySew_0_5};
  wire [15:0]      _GEN_137 = {dataRegroupBySew_5_5, dataRegroupBySew_4_5};
  wire [15:0]      dataInMem_hi_hi_42;
  assign dataInMem_hi_hi_42 = _GEN_137;
  wire [15:0]      dataInMem_hi_lo_44;
  assign dataInMem_hi_lo_44 = _GEN_137;
  wire [23:0]      dataInMem_hi_106 = {dataInMem_hi_hi_42, dataRegroupBySew_3_5};
  wire [23:0]      dataInMem_lo_75 = {dataInMem_lo_hi_11, dataRegroupBySew_0_6};
  wire [15:0]      _GEN_138 = {dataRegroupBySew_5_6, dataRegroupBySew_4_6};
  wire [15:0]      dataInMem_hi_hi_43;
  assign dataInMem_hi_hi_43 = _GEN_138;
  wire [15:0]      dataInMem_hi_lo_45;
  assign dataInMem_hi_lo_45 = _GEN_138;
  wire [23:0]      dataInMem_hi_107 = {dataInMem_hi_hi_43, dataRegroupBySew_3_6};
  wire [23:0]      dataInMem_lo_76 = {dataInMem_lo_hi_12, dataRegroupBySew_0_7};
  wire [15:0]      _GEN_139 = {dataRegroupBySew_5_7, dataRegroupBySew_4_7};
  wire [15:0]      dataInMem_hi_hi_44;
  assign dataInMem_hi_hi_44 = _GEN_139;
  wire [15:0]      dataInMem_hi_lo_46;
  assign dataInMem_hi_lo_46 = _GEN_139;
  wire [23:0]      dataInMem_hi_108 = {dataInMem_hi_hi_44, dataRegroupBySew_3_7};
  wire [23:0]      dataInMem_lo_77 = {dataInMem_lo_hi_13, dataRegroupBySew_0_8};
  wire [15:0]      _GEN_140 = {dataRegroupBySew_5_8, dataRegroupBySew_4_8};
  wire [15:0]      dataInMem_hi_hi_45;
  assign dataInMem_hi_hi_45 = _GEN_140;
  wire [15:0]      dataInMem_hi_lo_47;
  assign dataInMem_hi_lo_47 = _GEN_140;
  wire [23:0]      dataInMem_hi_109 = {dataInMem_hi_hi_45, dataRegroupBySew_3_8};
  wire [23:0]      dataInMem_lo_78 = {dataInMem_lo_hi_14, dataRegroupBySew_0_9};
  wire [15:0]      _GEN_141 = {dataRegroupBySew_5_9, dataRegroupBySew_4_9};
  wire [15:0]      dataInMem_hi_hi_46;
  assign dataInMem_hi_hi_46 = _GEN_141;
  wire [15:0]      dataInMem_hi_lo_48;
  assign dataInMem_hi_lo_48 = _GEN_141;
  wire [23:0]      dataInMem_hi_110 = {dataInMem_hi_hi_46, dataRegroupBySew_3_9};
  wire [23:0]      dataInMem_lo_79 = {dataInMem_lo_hi_15, dataRegroupBySew_0_10};
  wire [15:0]      _GEN_142 = {dataRegroupBySew_5_10, dataRegroupBySew_4_10};
  wire [15:0]      dataInMem_hi_hi_47;
  assign dataInMem_hi_hi_47 = _GEN_142;
  wire [15:0]      dataInMem_hi_lo_49;
  assign dataInMem_hi_lo_49 = _GEN_142;
  wire [23:0]      dataInMem_hi_111 = {dataInMem_hi_hi_47, dataRegroupBySew_3_10};
  wire [23:0]      dataInMem_lo_80 = {dataInMem_lo_hi_16, dataRegroupBySew_0_11};
  wire [15:0]      _GEN_143 = {dataRegroupBySew_5_11, dataRegroupBySew_4_11};
  wire [15:0]      dataInMem_hi_hi_48;
  assign dataInMem_hi_hi_48 = _GEN_143;
  wire [15:0]      dataInMem_hi_lo_50;
  assign dataInMem_hi_lo_50 = _GEN_143;
  wire [23:0]      dataInMem_hi_112 = {dataInMem_hi_hi_48, dataRegroupBySew_3_11};
  wire [23:0]      dataInMem_lo_81 = {dataInMem_lo_hi_17, dataRegroupBySew_0_12};
  wire [15:0]      _GEN_144 = {dataRegroupBySew_5_12, dataRegroupBySew_4_12};
  wire [15:0]      dataInMem_hi_hi_49;
  assign dataInMem_hi_hi_49 = _GEN_144;
  wire [15:0]      dataInMem_hi_lo_51;
  assign dataInMem_hi_lo_51 = _GEN_144;
  wire [23:0]      dataInMem_hi_113 = {dataInMem_hi_hi_49, dataRegroupBySew_3_12};
  wire [23:0]      dataInMem_lo_82 = {dataInMem_lo_hi_18, dataRegroupBySew_0_13};
  wire [15:0]      _GEN_145 = {dataRegroupBySew_5_13, dataRegroupBySew_4_13};
  wire [15:0]      dataInMem_hi_hi_50;
  assign dataInMem_hi_hi_50 = _GEN_145;
  wire [15:0]      dataInMem_hi_lo_52;
  assign dataInMem_hi_lo_52 = _GEN_145;
  wire [23:0]      dataInMem_hi_114 = {dataInMem_hi_hi_50, dataRegroupBySew_3_13};
  wire [23:0]      dataInMem_lo_83 = {dataInMem_lo_hi_19, dataRegroupBySew_0_14};
  wire [15:0]      _GEN_146 = {dataRegroupBySew_5_14, dataRegroupBySew_4_14};
  wire [15:0]      dataInMem_hi_hi_51;
  assign dataInMem_hi_hi_51 = _GEN_146;
  wire [15:0]      dataInMem_hi_lo_53;
  assign dataInMem_hi_lo_53 = _GEN_146;
  wire [23:0]      dataInMem_hi_115 = {dataInMem_hi_hi_51, dataRegroupBySew_3_14};
  wire [23:0]      dataInMem_lo_84 = {dataInMem_lo_hi_20, dataRegroupBySew_0_15};
  wire [15:0]      _GEN_147 = {dataRegroupBySew_5_15, dataRegroupBySew_4_15};
  wire [15:0]      dataInMem_hi_hi_52;
  assign dataInMem_hi_hi_52 = _GEN_147;
  wire [15:0]      dataInMem_hi_lo_54;
  assign dataInMem_hi_lo_54 = _GEN_147;
  wire [23:0]      dataInMem_hi_116 = {dataInMem_hi_hi_52, dataRegroupBySew_3_15};
  wire [23:0]      dataInMem_lo_85 = {dataInMem_lo_hi_21, dataRegroupBySew_0_16};
  wire [15:0]      _GEN_148 = {dataRegroupBySew_5_16, dataRegroupBySew_4_16};
  wire [15:0]      dataInMem_hi_hi_53;
  assign dataInMem_hi_hi_53 = _GEN_148;
  wire [15:0]      dataInMem_hi_lo_55;
  assign dataInMem_hi_lo_55 = _GEN_148;
  wire [23:0]      dataInMem_hi_117 = {dataInMem_hi_hi_53, dataRegroupBySew_3_16};
  wire [23:0]      dataInMem_lo_86 = {dataInMem_lo_hi_22, dataRegroupBySew_0_17};
  wire [15:0]      _GEN_149 = {dataRegroupBySew_5_17, dataRegroupBySew_4_17};
  wire [15:0]      dataInMem_hi_hi_54;
  assign dataInMem_hi_hi_54 = _GEN_149;
  wire [15:0]      dataInMem_hi_lo_56;
  assign dataInMem_hi_lo_56 = _GEN_149;
  wire [23:0]      dataInMem_hi_118 = {dataInMem_hi_hi_54, dataRegroupBySew_3_17};
  wire [23:0]      dataInMem_lo_87 = {dataInMem_lo_hi_23, dataRegroupBySew_0_18};
  wire [15:0]      _GEN_150 = {dataRegroupBySew_5_18, dataRegroupBySew_4_18};
  wire [15:0]      dataInMem_hi_hi_55;
  assign dataInMem_hi_hi_55 = _GEN_150;
  wire [15:0]      dataInMem_hi_lo_57;
  assign dataInMem_hi_lo_57 = _GEN_150;
  wire [23:0]      dataInMem_hi_119 = {dataInMem_hi_hi_55, dataRegroupBySew_3_18};
  wire [23:0]      dataInMem_lo_88 = {dataInMem_lo_hi_24, dataRegroupBySew_0_19};
  wire [15:0]      _GEN_151 = {dataRegroupBySew_5_19, dataRegroupBySew_4_19};
  wire [15:0]      dataInMem_hi_hi_56;
  assign dataInMem_hi_hi_56 = _GEN_151;
  wire [15:0]      dataInMem_hi_lo_58;
  assign dataInMem_hi_lo_58 = _GEN_151;
  wire [23:0]      dataInMem_hi_120 = {dataInMem_hi_hi_56, dataRegroupBySew_3_19};
  wire [23:0]      dataInMem_lo_89 = {dataInMem_lo_hi_25, dataRegroupBySew_0_20};
  wire [15:0]      _GEN_152 = {dataRegroupBySew_5_20, dataRegroupBySew_4_20};
  wire [15:0]      dataInMem_hi_hi_57;
  assign dataInMem_hi_hi_57 = _GEN_152;
  wire [15:0]      dataInMem_hi_lo_59;
  assign dataInMem_hi_lo_59 = _GEN_152;
  wire [23:0]      dataInMem_hi_121 = {dataInMem_hi_hi_57, dataRegroupBySew_3_20};
  wire [23:0]      dataInMem_lo_90 = {dataInMem_lo_hi_26, dataRegroupBySew_0_21};
  wire [15:0]      _GEN_153 = {dataRegroupBySew_5_21, dataRegroupBySew_4_21};
  wire [15:0]      dataInMem_hi_hi_58;
  assign dataInMem_hi_hi_58 = _GEN_153;
  wire [15:0]      dataInMem_hi_lo_60;
  assign dataInMem_hi_lo_60 = _GEN_153;
  wire [23:0]      dataInMem_hi_122 = {dataInMem_hi_hi_58, dataRegroupBySew_3_21};
  wire [23:0]      dataInMem_lo_91 = {dataInMem_lo_hi_27, dataRegroupBySew_0_22};
  wire [15:0]      _GEN_154 = {dataRegroupBySew_5_22, dataRegroupBySew_4_22};
  wire [15:0]      dataInMem_hi_hi_59;
  assign dataInMem_hi_hi_59 = _GEN_154;
  wire [15:0]      dataInMem_hi_lo_61;
  assign dataInMem_hi_lo_61 = _GEN_154;
  wire [23:0]      dataInMem_hi_123 = {dataInMem_hi_hi_59, dataRegroupBySew_3_22};
  wire [23:0]      dataInMem_lo_92 = {dataInMem_lo_hi_28, dataRegroupBySew_0_23};
  wire [15:0]      _GEN_155 = {dataRegroupBySew_5_23, dataRegroupBySew_4_23};
  wire [15:0]      dataInMem_hi_hi_60;
  assign dataInMem_hi_hi_60 = _GEN_155;
  wire [15:0]      dataInMem_hi_lo_62;
  assign dataInMem_hi_lo_62 = _GEN_155;
  wire [23:0]      dataInMem_hi_124 = {dataInMem_hi_hi_60, dataRegroupBySew_3_23};
  wire [23:0]      dataInMem_lo_93 = {dataInMem_lo_hi_29, dataRegroupBySew_0_24};
  wire [15:0]      _GEN_156 = {dataRegroupBySew_5_24, dataRegroupBySew_4_24};
  wire [15:0]      dataInMem_hi_hi_61;
  assign dataInMem_hi_hi_61 = _GEN_156;
  wire [15:0]      dataInMem_hi_lo_63;
  assign dataInMem_hi_lo_63 = _GEN_156;
  wire [23:0]      dataInMem_hi_125 = {dataInMem_hi_hi_61, dataRegroupBySew_3_24};
  wire [23:0]      dataInMem_lo_94 = {dataInMem_lo_hi_30, dataRegroupBySew_0_25};
  wire [15:0]      _GEN_157 = {dataRegroupBySew_5_25, dataRegroupBySew_4_25};
  wire [15:0]      dataInMem_hi_hi_62;
  assign dataInMem_hi_hi_62 = _GEN_157;
  wire [15:0]      dataInMem_hi_lo_64;
  assign dataInMem_hi_lo_64 = _GEN_157;
  wire [23:0]      dataInMem_hi_126 = {dataInMem_hi_hi_62, dataRegroupBySew_3_25};
  wire [23:0]      dataInMem_lo_95 = {dataInMem_lo_hi_31, dataRegroupBySew_0_26};
  wire [15:0]      _GEN_158 = {dataRegroupBySew_5_26, dataRegroupBySew_4_26};
  wire [15:0]      dataInMem_hi_hi_63;
  assign dataInMem_hi_hi_63 = _GEN_158;
  wire [15:0]      dataInMem_hi_lo_65;
  assign dataInMem_hi_lo_65 = _GEN_158;
  wire [23:0]      dataInMem_hi_127 = {dataInMem_hi_hi_63, dataRegroupBySew_3_26};
  wire [23:0]      dataInMem_lo_96 = {dataInMem_lo_hi_32, dataRegroupBySew_0_27};
  wire [15:0]      _GEN_159 = {dataRegroupBySew_5_27, dataRegroupBySew_4_27};
  wire [15:0]      dataInMem_hi_hi_64;
  assign dataInMem_hi_hi_64 = _GEN_159;
  wire [15:0]      dataInMem_hi_lo_66;
  assign dataInMem_hi_lo_66 = _GEN_159;
  wire [23:0]      dataInMem_hi_128 = {dataInMem_hi_hi_64, dataRegroupBySew_3_27};
  wire [23:0]      dataInMem_lo_97 = {dataInMem_lo_hi_33, dataRegroupBySew_0_28};
  wire [15:0]      _GEN_160 = {dataRegroupBySew_5_28, dataRegroupBySew_4_28};
  wire [15:0]      dataInMem_hi_hi_65;
  assign dataInMem_hi_hi_65 = _GEN_160;
  wire [15:0]      dataInMem_hi_lo_67;
  assign dataInMem_hi_lo_67 = _GEN_160;
  wire [23:0]      dataInMem_hi_129 = {dataInMem_hi_hi_65, dataRegroupBySew_3_28};
  wire [23:0]      dataInMem_lo_98 = {dataInMem_lo_hi_34, dataRegroupBySew_0_29};
  wire [15:0]      _GEN_161 = {dataRegroupBySew_5_29, dataRegroupBySew_4_29};
  wire [15:0]      dataInMem_hi_hi_66;
  assign dataInMem_hi_hi_66 = _GEN_161;
  wire [15:0]      dataInMem_hi_lo_68;
  assign dataInMem_hi_lo_68 = _GEN_161;
  wire [23:0]      dataInMem_hi_130 = {dataInMem_hi_hi_66, dataRegroupBySew_3_29};
  wire [23:0]      dataInMem_lo_99 = {dataInMem_lo_hi_35, dataRegroupBySew_0_30};
  wire [15:0]      _GEN_162 = {dataRegroupBySew_5_30, dataRegroupBySew_4_30};
  wire [15:0]      dataInMem_hi_hi_67;
  assign dataInMem_hi_hi_67 = _GEN_162;
  wire [15:0]      dataInMem_hi_lo_69;
  assign dataInMem_hi_lo_69 = _GEN_162;
  wire [23:0]      dataInMem_hi_131 = {dataInMem_hi_hi_67, dataRegroupBySew_3_30};
  wire [23:0]      dataInMem_lo_100 = {dataInMem_lo_hi_36, dataRegroupBySew_0_31};
  wire [15:0]      _GEN_163 = {dataRegroupBySew_5_31, dataRegroupBySew_4_31};
  wire [15:0]      dataInMem_hi_hi_68;
  assign dataInMem_hi_hi_68 = _GEN_163;
  wire [15:0]      dataInMem_hi_lo_70;
  assign dataInMem_hi_lo_70 = _GEN_163;
  wire [23:0]      dataInMem_hi_132 = {dataInMem_hi_hi_68, dataRegroupBySew_3_31};
  wire [95:0]      dataInMem_lo_lo_lo_lo_5 = {dataInMem_hi_102, dataInMem_lo_70, dataInMem_hi_101, dataInMem_lo_69};
  wire [95:0]      dataInMem_lo_lo_lo_hi_5 = {dataInMem_hi_104, dataInMem_lo_72, dataInMem_hi_103, dataInMem_lo_71};
  wire [191:0]     dataInMem_lo_lo_lo_5 = {dataInMem_lo_lo_lo_hi_5, dataInMem_lo_lo_lo_lo_5};
  wire [95:0]      dataInMem_lo_lo_hi_lo_5 = {dataInMem_hi_106, dataInMem_lo_74, dataInMem_hi_105, dataInMem_lo_73};
  wire [95:0]      dataInMem_lo_lo_hi_hi_5 = {dataInMem_hi_108, dataInMem_lo_76, dataInMem_hi_107, dataInMem_lo_75};
  wire [191:0]     dataInMem_lo_lo_hi_5 = {dataInMem_lo_lo_hi_hi_5, dataInMem_lo_lo_hi_lo_5};
  wire [383:0]     dataInMem_lo_lo_5 = {dataInMem_lo_lo_hi_5, dataInMem_lo_lo_lo_5};
  wire [95:0]      dataInMem_lo_hi_lo_lo_5 = {dataInMem_hi_110, dataInMem_lo_78, dataInMem_hi_109, dataInMem_lo_77};
  wire [95:0]      dataInMem_lo_hi_lo_hi_5 = {dataInMem_hi_112, dataInMem_lo_80, dataInMem_hi_111, dataInMem_lo_79};
  wire [191:0]     dataInMem_lo_hi_lo_5 = {dataInMem_lo_hi_lo_hi_5, dataInMem_lo_hi_lo_lo_5};
  wire [95:0]      dataInMem_lo_hi_hi_lo_5 = {dataInMem_hi_114, dataInMem_lo_82, dataInMem_hi_113, dataInMem_lo_81};
  wire [95:0]      dataInMem_lo_hi_hi_hi_5 = {dataInMem_hi_116, dataInMem_lo_84, dataInMem_hi_115, dataInMem_lo_83};
  wire [191:0]     dataInMem_lo_hi_hi_5 = {dataInMem_lo_hi_hi_hi_5, dataInMem_lo_hi_hi_lo_5};
  wire [383:0]     dataInMem_lo_hi_37 = {dataInMem_lo_hi_hi_5, dataInMem_lo_hi_lo_5};
  wire [767:0]     dataInMem_lo_101 = {dataInMem_lo_hi_37, dataInMem_lo_lo_5};
  wire [95:0]      dataInMem_hi_lo_lo_lo_5 = {dataInMem_hi_118, dataInMem_lo_86, dataInMem_hi_117, dataInMem_lo_85};
  wire [95:0]      dataInMem_hi_lo_lo_hi_5 = {dataInMem_hi_120, dataInMem_lo_88, dataInMem_hi_119, dataInMem_lo_87};
  wire [191:0]     dataInMem_hi_lo_lo_5 = {dataInMem_hi_lo_lo_hi_5, dataInMem_hi_lo_lo_lo_5};
  wire [95:0]      dataInMem_hi_lo_hi_lo_5 = {dataInMem_hi_122, dataInMem_lo_90, dataInMem_hi_121, dataInMem_lo_89};
  wire [95:0]      dataInMem_hi_lo_hi_hi_5 = {dataInMem_hi_124, dataInMem_lo_92, dataInMem_hi_123, dataInMem_lo_91};
  wire [191:0]     dataInMem_hi_lo_hi_5 = {dataInMem_hi_lo_hi_hi_5, dataInMem_hi_lo_hi_lo_5};
  wire [383:0]     dataInMem_hi_lo_5 = {dataInMem_hi_lo_hi_5, dataInMem_hi_lo_lo_5};
  wire [95:0]      dataInMem_hi_hi_lo_lo_5 = {dataInMem_hi_126, dataInMem_lo_94, dataInMem_hi_125, dataInMem_lo_93};
  wire [95:0]      dataInMem_hi_hi_lo_hi_5 = {dataInMem_hi_128, dataInMem_lo_96, dataInMem_hi_127, dataInMem_lo_95};
  wire [191:0]     dataInMem_hi_hi_lo_5 = {dataInMem_hi_hi_lo_hi_5, dataInMem_hi_hi_lo_lo_5};
  wire [95:0]      dataInMem_hi_hi_hi_lo_5 = {dataInMem_hi_130, dataInMem_lo_98, dataInMem_hi_129, dataInMem_lo_97};
  wire [95:0]      dataInMem_hi_hi_hi_hi_5 = {dataInMem_hi_132, dataInMem_lo_100, dataInMem_hi_131, dataInMem_lo_99};
  wire [191:0]     dataInMem_hi_hi_hi_5 = {dataInMem_hi_hi_hi_hi_5, dataInMem_hi_hi_hi_lo_5};
  wire [383:0]     dataInMem_hi_hi_69 = {dataInMem_hi_hi_hi_5, dataInMem_hi_hi_lo_5};
  wire [767:0]     dataInMem_hi_133 = {dataInMem_hi_hi_69, dataInMem_hi_lo_5};
  wire [1535:0]    dataInMem_5 = {dataInMem_hi_133, dataInMem_lo_101};
  wire [255:0]     regroupCacheLine_5_0 = dataInMem_5[255:0];
  wire [255:0]     regroupCacheLine_5_1 = dataInMem_5[511:256];
  wire [255:0]     regroupCacheLine_5_2 = dataInMem_5[767:512];
  wire [255:0]     regroupCacheLine_5_3 = dataInMem_5[1023:768];
  wire [255:0]     regroupCacheLine_5_4 = dataInMem_5[1279:1024];
  wire [255:0]     regroupCacheLine_5_5 = dataInMem_5[1535:1280];
  wire [255:0]     res_40 = regroupCacheLine_5_0;
  wire [255:0]     res_41 = regroupCacheLine_5_1;
  wire [255:0]     res_42 = regroupCacheLine_5_2;
  wire [255:0]     res_43 = regroupCacheLine_5_3;
  wire [255:0]     res_44 = regroupCacheLine_5_4;
  wire [255:0]     res_45 = regroupCacheLine_5_5;
  wire [511:0]     lo_lo_5 = {res_41, res_40};
  wire [511:0]     lo_hi_5 = {res_43, res_42};
  wire [1023:0]    lo_5 = {lo_hi_5, lo_lo_5};
  wire [511:0]     hi_lo_5 = {res_45, res_44};
  wire [1023:0]    hi_5 = {512'h0, hi_lo_5};
  wire [2047:0]    regroupLoadData_0_5 = {hi_5, lo_5};
  wire [23:0]      dataInMem_lo_102 = {dataInMem_lo_hi_38, dataRegroupBySew_0_0};
  wire [15:0]      dataInMem_hi_hi_70 = {dataRegroupBySew_6_0, dataRegroupBySew_5_0};
  wire [31:0]      dataInMem_hi_134 = {dataInMem_hi_hi_70, dataInMem_hi_lo_6};
  wire [23:0]      dataInMem_lo_103 = {dataInMem_lo_hi_39, dataRegroupBySew_0_1};
  wire [15:0]      dataInMem_hi_hi_71 = {dataRegroupBySew_6_1, dataRegroupBySew_5_1};
  wire [31:0]      dataInMem_hi_135 = {dataInMem_hi_hi_71, dataInMem_hi_lo_7};
  wire [23:0]      dataInMem_lo_104 = {dataInMem_lo_hi_40, dataRegroupBySew_0_2};
  wire [15:0]      dataInMem_hi_hi_72 = {dataRegroupBySew_6_2, dataRegroupBySew_5_2};
  wire [31:0]      dataInMem_hi_136 = {dataInMem_hi_hi_72, dataInMem_hi_lo_8};
  wire [23:0]      dataInMem_lo_105 = {dataInMem_lo_hi_41, dataRegroupBySew_0_3};
  wire [15:0]      dataInMem_hi_hi_73 = {dataRegroupBySew_6_3, dataRegroupBySew_5_3};
  wire [31:0]      dataInMem_hi_137 = {dataInMem_hi_hi_73, dataInMem_hi_lo_9};
  wire [23:0]      dataInMem_lo_106 = {dataInMem_lo_hi_42, dataRegroupBySew_0_4};
  wire [15:0]      dataInMem_hi_hi_74 = {dataRegroupBySew_6_4, dataRegroupBySew_5_4};
  wire [31:0]      dataInMem_hi_138 = {dataInMem_hi_hi_74, dataInMem_hi_lo_10};
  wire [23:0]      dataInMem_lo_107 = {dataInMem_lo_hi_43, dataRegroupBySew_0_5};
  wire [15:0]      dataInMem_hi_hi_75 = {dataRegroupBySew_6_5, dataRegroupBySew_5_5};
  wire [31:0]      dataInMem_hi_139 = {dataInMem_hi_hi_75, dataInMem_hi_lo_11};
  wire [23:0]      dataInMem_lo_108 = {dataInMem_lo_hi_44, dataRegroupBySew_0_6};
  wire [15:0]      dataInMem_hi_hi_76 = {dataRegroupBySew_6_6, dataRegroupBySew_5_6};
  wire [31:0]      dataInMem_hi_140 = {dataInMem_hi_hi_76, dataInMem_hi_lo_12};
  wire [23:0]      dataInMem_lo_109 = {dataInMem_lo_hi_45, dataRegroupBySew_0_7};
  wire [15:0]      dataInMem_hi_hi_77 = {dataRegroupBySew_6_7, dataRegroupBySew_5_7};
  wire [31:0]      dataInMem_hi_141 = {dataInMem_hi_hi_77, dataInMem_hi_lo_13};
  wire [23:0]      dataInMem_lo_110 = {dataInMem_lo_hi_46, dataRegroupBySew_0_8};
  wire [15:0]      dataInMem_hi_hi_78 = {dataRegroupBySew_6_8, dataRegroupBySew_5_8};
  wire [31:0]      dataInMem_hi_142 = {dataInMem_hi_hi_78, dataInMem_hi_lo_14};
  wire [23:0]      dataInMem_lo_111 = {dataInMem_lo_hi_47, dataRegroupBySew_0_9};
  wire [15:0]      dataInMem_hi_hi_79 = {dataRegroupBySew_6_9, dataRegroupBySew_5_9};
  wire [31:0]      dataInMem_hi_143 = {dataInMem_hi_hi_79, dataInMem_hi_lo_15};
  wire [23:0]      dataInMem_lo_112 = {dataInMem_lo_hi_48, dataRegroupBySew_0_10};
  wire [15:0]      dataInMem_hi_hi_80 = {dataRegroupBySew_6_10, dataRegroupBySew_5_10};
  wire [31:0]      dataInMem_hi_144 = {dataInMem_hi_hi_80, dataInMem_hi_lo_16};
  wire [23:0]      dataInMem_lo_113 = {dataInMem_lo_hi_49, dataRegroupBySew_0_11};
  wire [15:0]      dataInMem_hi_hi_81 = {dataRegroupBySew_6_11, dataRegroupBySew_5_11};
  wire [31:0]      dataInMem_hi_145 = {dataInMem_hi_hi_81, dataInMem_hi_lo_17};
  wire [23:0]      dataInMem_lo_114 = {dataInMem_lo_hi_50, dataRegroupBySew_0_12};
  wire [15:0]      dataInMem_hi_hi_82 = {dataRegroupBySew_6_12, dataRegroupBySew_5_12};
  wire [31:0]      dataInMem_hi_146 = {dataInMem_hi_hi_82, dataInMem_hi_lo_18};
  wire [23:0]      dataInMem_lo_115 = {dataInMem_lo_hi_51, dataRegroupBySew_0_13};
  wire [15:0]      dataInMem_hi_hi_83 = {dataRegroupBySew_6_13, dataRegroupBySew_5_13};
  wire [31:0]      dataInMem_hi_147 = {dataInMem_hi_hi_83, dataInMem_hi_lo_19};
  wire [23:0]      dataInMem_lo_116 = {dataInMem_lo_hi_52, dataRegroupBySew_0_14};
  wire [15:0]      dataInMem_hi_hi_84 = {dataRegroupBySew_6_14, dataRegroupBySew_5_14};
  wire [31:0]      dataInMem_hi_148 = {dataInMem_hi_hi_84, dataInMem_hi_lo_20};
  wire [23:0]      dataInMem_lo_117 = {dataInMem_lo_hi_53, dataRegroupBySew_0_15};
  wire [15:0]      dataInMem_hi_hi_85 = {dataRegroupBySew_6_15, dataRegroupBySew_5_15};
  wire [31:0]      dataInMem_hi_149 = {dataInMem_hi_hi_85, dataInMem_hi_lo_21};
  wire [23:0]      dataInMem_lo_118 = {dataInMem_lo_hi_54, dataRegroupBySew_0_16};
  wire [15:0]      dataInMem_hi_hi_86 = {dataRegroupBySew_6_16, dataRegroupBySew_5_16};
  wire [31:0]      dataInMem_hi_150 = {dataInMem_hi_hi_86, dataInMem_hi_lo_22};
  wire [23:0]      dataInMem_lo_119 = {dataInMem_lo_hi_55, dataRegroupBySew_0_17};
  wire [15:0]      dataInMem_hi_hi_87 = {dataRegroupBySew_6_17, dataRegroupBySew_5_17};
  wire [31:0]      dataInMem_hi_151 = {dataInMem_hi_hi_87, dataInMem_hi_lo_23};
  wire [23:0]      dataInMem_lo_120 = {dataInMem_lo_hi_56, dataRegroupBySew_0_18};
  wire [15:0]      dataInMem_hi_hi_88 = {dataRegroupBySew_6_18, dataRegroupBySew_5_18};
  wire [31:0]      dataInMem_hi_152 = {dataInMem_hi_hi_88, dataInMem_hi_lo_24};
  wire [23:0]      dataInMem_lo_121 = {dataInMem_lo_hi_57, dataRegroupBySew_0_19};
  wire [15:0]      dataInMem_hi_hi_89 = {dataRegroupBySew_6_19, dataRegroupBySew_5_19};
  wire [31:0]      dataInMem_hi_153 = {dataInMem_hi_hi_89, dataInMem_hi_lo_25};
  wire [23:0]      dataInMem_lo_122 = {dataInMem_lo_hi_58, dataRegroupBySew_0_20};
  wire [15:0]      dataInMem_hi_hi_90 = {dataRegroupBySew_6_20, dataRegroupBySew_5_20};
  wire [31:0]      dataInMem_hi_154 = {dataInMem_hi_hi_90, dataInMem_hi_lo_26};
  wire [23:0]      dataInMem_lo_123 = {dataInMem_lo_hi_59, dataRegroupBySew_0_21};
  wire [15:0]      dataInMem_hi_hi_91 = {dataRegroupBySew_6_21, dataRegroupBySew_5_21};
  wire [31:0]      dataInMem_hi_155 = {dataInMem_hi_hi_91, dataInMem_hi_lo_27};
  wire [23:0]      dataInMem_lo_124 = {dataInMem_lo_hi_60, dataRegroupBySew_0_22};
  wire [15:0]      dataInMem_hi_hi_92 = {dataRegroupBySew_6_22, dataRegroupBySew_5_22};
  wire [31:0]      dataInMem_hi_156 = {dataInMem_hi_hi_92, dataInMem_hi_lo_28};
  wire [23:0]      dataInMem_lo_125 = {dataInMem_lo_hi_61, dataRegroupBySew_0_23};
  wire [15:0]      dataInMem_hi_hi_93 = {dataRegroupBySew_6_23, dataRegroupBySew_5_23};
  wire [31:0]      dataInMem_hi_157 = {dataInMem_hi_hi_93, dataInMem_hi_lo_29};
  wire [23:0]      dataInMem_lo_126 = {dataInMem_lo_hi_62, dataRegroupBySew_0_24};
  wire [15:0]      dataInMem_hi_hi_94 = {dataRegroupBySew_6_24, dataRegroupBySew_5_24};
  wire [31:0]      dataInMem_hi_158 = {dataInMem_hi_hi_94, dataInMem_hi_lo_30};
  wire [23:0]      dataInMem_lo_127 = {dataInMem_lo_hi_63, dataRegroupBySew_0_25};
  wire [15:0]      dataInMem_hi_hi_95 = {dataRegroupBySew_6_25, dataRegroupBySew_5_25};
  wire [31:0]      dataInMem_hi_159 = {dataInMem_hi_hi_95, dataInMem_hi_lo_31};
  wire [23:0]      dataInMem_lo_128 = {dataInMem_lo_hi_64, dataRegroupBySew_0_26};
  wire [15:0]      dataInMem_hi_hi_96 = {dataRegroupBySew_6_26, dataRegroupBySew_5_26};
  wire [31:0]      dataInMem_hi_160 = {dataInMem_hi_hi_96, dataInMem_hi_lo_32};
  wire [23:0]      dataInMem_lo_129 = {dataInMem_lo_hi_65, dataRegroupBySew_0_27};
  wire [15:0]      dataInMem_hi_hi_97 = {dataRegroupBySew_6_27, dataRegroupBySew_5_27};
  wire [31:0]      dataInMem_hi_161 = {dataInMem_hi_hi_97, dataInMem_hi_lo_33};
  wire [23:0]      dataInMem_lo_130 = {dataInMem_lo_hi_66, dataRegroupBySew_0_28};
  wire [15:0]      dataInMem_hi_hi_98 = {dataRegroupBySew_6_28, dataRegroupBySew_5_28};
  wire [31:0]      dataInMem_hi_162 = {dataInMem_hi_hi_98, dataInMem_hi_lo_34};
  wire [23:0]      dataInMem_lo_131 = {dataInMem_lo_hi_67, dataRegroupBySew_0_29};
  wire [15:0]      dataInMem_hi_hi_99 = {dataRegroupBySew_6_29, dataRegroupBySew_5_29};
  wire [31:0]      dataInMem_hi_163 = {dataInMem_hi_hi_99, dataInMem_hi_lo_35};
  wire [23:0]      dataInMem_lo_132 = {dataInMem_lo_hi_68, dataRegroupBySew_0_30};
  wire [15:0]      dataInMem_hi_hi_100 = {dataRegroupBySew_6_30, dataRegroupBySew_5_30};
  wire [31:0]      dataInMem_hi_164 = {dataInMem_hi_hi_100, dataInMem_hi_lo_36};
  wire [23:0]      dataInMem_lo_133 = {dataInMem_lo_hi_69, dataRegroupBySew_0_31};
  wire [15:0]      dataInMem_hi_hi_101 = {dataRegroupBySew_6_31, dataRegroupBySew_5_31};
  wire [31:0]      dataInMem_hi_165 = {dataInMem_hi_hi_101, dataInMem_hi_lo_37};
  wire [111:0]     dataInMem_lo_lo_lo_lo_6 = {dataInMem_hi_135, dataInMem_lo_103, dataInMem_hi_134, dataInMem_lo_102};
  wire [111:0]     dataInMem_lo_lo_lo_hi_6 = {dataInMem_hi_137, dataInMem_lo_105, dataInMem_hi_136, dataInMem_lo_104};
  wire [223:0]     dataInMem_lo_lo_lo_6 = {dataInMem_lo_lo_lo_hi_6, dataInMem_lo_lo_lo_lo_6};
  wire [111:0]     dataInMem_lo_lo_hi_lo_6 = {dataInMem_hi_139, dataInMem_lo_107, dataInMem_hi_138, dataInMem_lo_106};
  wire [111:0]     dataInMem_lo_lo_hi_hi_6 = {dataInMem_hi_141, dataInMem_lo_109, dataInMem_hi_140, dataInMem_lo_108};
  wire [223:0]     dataInMem_lo_lo_hi_6 = {dataInMem_lo_lo_hi_hi_6, dataInMem_lo_lo_hi_lo_6};
  wire [447:0]     dataInMem_lo_lo_6 = {dataInMem_lo_lo_hi_6, dataInMem_lo_lo_lo_6};
  wire [111:0]     dataInMem_lo_hi_lo_lo_6 = {dataInMem_hi_143, dataInMem_lo_111, dataInMem_hi_142, dataInMem_lo_110};
  wire [111:0]     dataInMem_lo_hi_lo_hi_6 = {dataInMem_hi_145, dataInMem_lo_113, dataInMem_hi_144, dataInMem_lo_112};
  wire [223:0]     dataInMem_lo_hi_lo_6 = {dataInMem_lo_hi_lo_hi_6, dataInMem_lo_hi_lo_lo_6};
  wire [111:0]     dataInMem_lo_hi_hi_lo_6 = {dataInMem_hi_147, dataInMem_lo_115, dataInMem_hi_146, dataInMem_lo_114};
  wire [111:0]     dataInMem_lo_hi_hi_hi_6 = {dataInMem_hi_149, dataInMem_lo_117, dataInMem_hi_148, dataInMem_lo_116};
  wire [223:0]     dataInMem_lo_hi_hi_6 = {dataInMem_lo_hi_hi_hi_6, dataInMem_lo_hi_hi_lo_6};
  wire [447:0]     dataInMem_lo_hi_70 = {dataInMem_lo_hi_hi_6, dataInMem_lo_hi_lo_6};
  wire [895:0]     dataInMem_lo_134 = {dataInMem_lo_hi_70, dataInMem_lo_lo_6};
  wire [111:0]     dataInMem_hi_lo_lo_lo_6 = {dataInMem_hi_151, dataInMem_lo_119, dataInMem_hi_150, dataInMem_lo_118};
  wire [111:0]     dataInMem_hi_lo_lo_hi_6 = {dataInMem_hi_153, dataInMem_lo_121, dataInMem_hi_152, dataInMem_lo_120};
  wire [223:0]     dataInMem_hi_lo_lo_6 = {dataInMem_hi_lo_lo_hi_6, dataInMem_hi_lo_lo_lo_6};
  wire [111:0]     dataInMem_hi_lo_hi_lo_6 = {dataInMem_hi_155, dataInMem_lo_123, dataInMem_hi_154, dataInMem_lo_122};
  wire [111:0]     dataInMem_hi_lo_hi_hi_6 = {dataInMem_hi_157, dataInMem_lo_125, dataInMem_hi_156, dataInMem_lo_124};
  wire [223:0]     dataInMem_hi_lo_hi_6 = {dataInMem_hi_lo_hi_hi_6, dataInMem_hi_lo_hi_lo_6};
  wire [447:0]     dataInMem_hi_lo_38 = {dataInMem_hi_lo_hi_6, dataInMem_hi_lo_lo_6};
  wire [111:0]     dataInMem_hi_hi_lo_lo_6 = {dataInMem_hi_159, dataInMem_lo_127, dataInMem_hi_158, dataInMem_lo_126};
  wire [111:0]     dataInMem_hi_hi_lo_hi_6 = {dataInMem_hi_161, dataInMem_lo_129, dataInMem_hi_160, dataInMem_lo_128};
  wire [223:0]     dataInMem_hi_hi_lo_6 = {dataInMem_hi_hi_lo_hi_6, dataInMem_hi_hi_lo_lo_6};
  wire [111:0]     dataInMem_hi_hi_hi_lo_6 = {dataInMem_hi_163, dataInMem_lo_131, dataInMem_hi_162, dataInMem_lo_130};
  wire [111:0]     dataInMem_hi_hi_hi_hi_6 = {dataInMem_hi_165, dataInMem_lo_133, dataInMem_hi_164, dataInMem_lo_132};
  wire [223:0]     dataInMem_hi_hi_hi_6 = {dataInMem_hi_hi_hi_hi_6, dataInMem_hi_hi_hi_lo_6};
  wire [447:0]     dataInMem_hi_hi_102 = {dataInMem_hi_hi_hi_6, dataInMem_hi_hi_lo_6};
  wire [895:0]     dataInMem_hi_166 = {dataInMem_hi_hi_102, dataInMem_hi_lo_38};
  wire [1791:0]    dataInMem_6 = {dataInMem_hi_166, dataInMem_lo_134};
  wire [255:0]     regroupCacheLine_6_0 = dataInMem_6[255:0];
  wire [255:0]     regroupCacheLine_6_1 = dataInMem_6[511:256];
  wire [255:0]     regroupCacheLine_6_2 = dataInMem_6[767:512];
  wire [255:0]     regroupCacheLine_6_3 = dataInMem_6[1023:768];
  wire [255:0]     regroupCacheLine_6_4 = dataInMem_6[1279:1024];
  wire [255:0]     regroupCacheLine_6_5 = dataInMem_6[1535:1280];
  wire [255:0]     regroupCacheLine_6_6 = dataInMem_6[1791:1536];
  wire [255:0]     res_48 = regroupCacheLine_6_0;
  wire [255:0]     res_49 = regroupCacheLine_6_1;
  wire [255:0]     res_50 = regroupCacheLine_6_2;
  wire [255:0]     res_51 = regroupCacheLine_6_3;
  wire [255:0]     res_52 = regroupCacheLine_6_4;
  wire [255:0]     res_53 = regroupCacheLine_6_5;
  wire [255:0]     res_54 = regroupCacheLine_6_6;
  wire [511:0]     lo_lo_6 = {res_49, res_48};
  wire [511:0]     lo_hi_6 = {res_51, res_50};
  wire [1023:0]    lo_6 = {lo_hi_6, lo_lo_6};
  wire [511:0]     hi_lo_6 = {res_53, res_52};
  wire [511:0]     hi_hi_6 = {256'h0, res_54};
  wire [1023:0]    hi_6 = {hi_hi_6, hi_lo_6};
  wire [2047:0]    regroupLoadData_0_6 = {hi_6, lo_6};
  wire [31:0]      dataInMem_lo_135 = {dataInMem_lo_hi_71, dataInMem_lo_lo_7};
  wire [15:0]      dataInMem_hi_hi_103 = {dataRegroupBySew_7_0, dataRegroupBySew_6_0};
  wire [31:0]      dataInMem_hi_167 = {dataInMem_hi_hi_103, dataInMem_hi_lo_39};
  wire [31:0]      dataInMem_lo_136 = {dataInMem_lo_hi_72, dataInMem_lo_lo_8};
  wire [15:0]      dataInMem_hi_hi_104 = {dataRegroupBySew_7_1, dataRegroupBySew_6_1};
  wire [31:0]      dataInMem_hi_168 = {dataInMem_hi_hi_104, dataInMem_hi_lo_40};
  wire [31:0]      dataInMem_lo_137 = {dataInMem_lo_hi_73, dataInMem_lo_lo_9};
  wire [15:0]      dataInMem_hi_hi_105 = {dataRegroupBySew_7_2, dataRegroupBySew_6_2};
  wire [31:0]      dataInMem_hi_169 = {dataInMem_hi_hi_105, dataInMem_hi_lo_41};
  wire [31:0]      dataInMem_lo_138 = {dataInMem_lo_hi_74, dataInMem_lo_lo_10};
  wire [15:0]      dataInMem_hi_hi_106 = {dataRegroupBySew_7_3, dataRegroupBySew_6_3};
  wire [31:0]      dataInMem_hi_170 = {dataInMem_hi_hi_106, dataInMem_hi_lo_42};
  wire [31:0]      dataInMem_lo_139 = {dataInMem_lo_hi_75, dataInMem_lo_lo_11};
  wire [15:0]      dataInMem_hi_hi_107 = {dataRegroupBySew_7_4, dataRegroupBySew_6_4};
  wire [31:0]      dataInMem_hi_171 = {dataInMem_hi_hi_107, dataInMem_hi_lo_43};
  wire [31:0]      dataInMem_lo_140 = {dataInMem_lo_hi_76, dataInMem_lo_lo_12};
  wire [15:0]      dataInMem_hi_hi_108 = {dataRegroupBySew_7_5, dataRegroupBySew_6_5};
  wire [31:0]      dataInMem_hi_172 = {dataInMem_hi_hi_108, dataInMem_hi_lo_44};
  wire [31:0]      dataInMem_lo_141 = {dataInMem_lo_hi_77, dataInMem_lo_lo_13};
  wire [15:0]      dataInMem_hi_hi_109 = {dataRegroupBySew_7_6, dataRegroupBySew_6_6};
  wire [31:0]      dataInMem_hi_173 = {dataInMem_hi_hi_109, dataInMem_hi_lo_45};
  wire [31:0]      dataInMem_lo_142 = {dataInMem_lo_hi_78, dataInMem_lo_lo_14};
  wire [15:0]      dataInMem_hi_hi_110 = {dataRegroupBySew_7_7, dataRegroupBySew_6_7};
  wire [31:0]      dataInMem_hi_174 = {dataInMem_hi_hi_110, dataInMem_hi_lo_46};
  wire [31:0]      dataInMem_lo_143 = {dataInMem_lo_hi_79, dataInMem_lo_lo_15};
  wire [15:0]      dataInMem_hi_hi_111 = {dataRegroupBySew_7_8, dataRegroupBySew_6_8};
  wire [31:0]      dataInMem_hi_175 = {dataInMem_hi_hi_111, dataInMem_hi_lo_47};
  wire [31:0]      dataInMem_lo_144 = {dataInMem_lo_hi_80, dataInMem_lo_lo_16};
  wire [15:0]      dataInMem_hi_hi_112 = {dataRegroupBySew_7_9, dataRegroupBySew_6_9};
  wire [31:0]      dataInMem_hi_176 = {dataInMem_hi_hi_112, dataInMem_hi_lo_48};
  wire [31:0]      dataInMem_lo_145 = {dataInMem_lo_hi_81, dataInMem_lo_lo_17};
  wire [15:0]      dataInMem_hi_hi_113 = {dataRegroupBySew_7_10, dataRegroupBySew_6_10};
  wire [31:0]      dataInMem_hi_177 = {dataInMem_hi_hi_113, dataInMem_hi_lo_49};
  wire [31:0]      dataInMem_lo_146 = {dataInMem_lo_hi_82, dataInMem_lo_lo_18};
  wire [15:0]      dataInMem_hi_hi_114 = {dataRegroupBySew_7_11, dataRegroupBySew_6_11};
  wire [31:0]      dataInMem_hi_178 = {dataInMem_hi_hi_114, dataInMem_hi_lo_50};
  wire [31:0]      dataInMem_lo_147 = {dataInMem_lo_hi_83, dataInMem_lo_lo_19};
  wire [15:0]      dataInMem_hi_hi_115 = {dataRegroupBySew_7_12, dataRegroupBySew_6_12};
  wire [31:0]      dataInMem_hi_179 = {dataInMem_hi_hi_115, dataInMem_hi_lo_51};
  wire [31:0]      dataInMem_lo_148 = {dataInMem_lo_hi_84, dataInMem_lo_lo_20};
  wire [15:0]      dataInMem_hi_hi_116 = {dataRegroupBySew_7_13, dataRegroupBySew_6_13};
  wire [31:0]      dataInMem_hi_180 = {dataInMem_hi_hi_116, dataInMem_hi_lo_52};
  wire [31:0]      dataInMem_lo_149 = {dataInMem_lo_hi_85, dataInMem_lo_lo_21};
  wire [15:0]      dataInMem_hi_hi_117 = {dataRegroupBySew_7_14, dataRegroupBySew_6_14};
  wire [31:0]      dataInMem_hi_181 = {dataInMem_hi_hi_117, dataInMem_hi_lo_53};
  wire [31:0]      dataInMem_lo_150 = {dataInMem_lo_hi_86, dataInMem_lo_lo_22};
  wire [15:0]      dataInMem_hi_hi_118 = {dataRegroupBySew_7_15, dataRegroupBySew_6_15};
  wire [31:0]      dataInMem_hi_182 = {dataInMem_hi_hi_118, dataInMem_hi_lo_54};
  wire [31:0]      dataInMem_lo_151 = {dataInMem_lo_hi_87, dataInMem_lo_lo_23};
  wire [15:0]      dataInMem_hi_hi_119 = {dataRegroupBySew_7_16, dataRegroupBySew_6_16};
  wire [31:0]      dataInMem_hi_183 = {dataInMem_hi_hi_119, dataInMem_hi_lo_55};
  wire [31:0]      dataInMem_lo_152 = {dataInMem_lo_hi_88, dataInMem_lo_lo_24};
  wire [15:0]      dataInMem_hi_hi_120 = {dataRegroupBySew_7_17, dataRegroupBySew_6_17};
  wire [31:0]      dataInMem_hi_184 = {dataInMem_hi_hi_120, dataInMem_hi_lo_56};
  wire [31:0]      dataInMem_lo_153 = {dataInMem_lo_hi_89, dataInMem_lo_lo_25};
  wire [15:0]      dataInMem_hi_hi_121 = {dataRegroupBySew_7_18, dataRegroupBySew_6_18};
  wire [31:0]      dataInMem_hi_185 = {dataInMem_hi_hi_121, dataInMem_hi_lo_57};
  wire [31:0]      dataInMem_lo_154 = {dataInMem_lo_hi_90, dataInMem_lo_lo_26};
  wire [15:0]      dataInMem_hi_hi_122 = {dataRegroupBySew_7_19, dataRegroupBySew_6_19};
  wire [31:0]      dataInMem_hi_186 = {dataInMem_hi_hi_122, dataInMem_hi_lo_58};
  wire [31:0]      dataInMem_lo_155 = {dataInMem_lo_hi_91, dataInMem_lo_lo_27};
  wire [15:0]      dataInMem_hi_hi_123 = {dataRegroupBySew_7_20, dataRegroupBySew_6_20};
  wire [31:0]      dataInMem_hi_187 = {dataInMem_hi_hi_123, dataInMem_hi_lo_59};
  wire [31:0]      dataInMem_lo_156 = {dataInMem_lo_hi_92, dataInMem_lo_lo_28};
  wire [15:0]      dataInMem_hi_hi_124 = {dataRegroupBySew_7_21, dataRegroupBySew_6_21};
  wire [31:0]      dataInMem_hi_188 = {dataInMem_hi_hi_124, dataInMem_hi_lo_60};
  wire [31:0]      dataInMem_lo_157 = {dataInMem_lo_hi_93, dataInMem_lo_lo_29};
  wire [15:0]      dataInMem_hi_hi_125 = {dataRegroupBySew_7_22, dataRegroupBySew_6_22};
  wire [31:0]      dataInMem_hi_189 = {dataInMem_hi_hi_125, dataInMem_hi_lo_61};
  wire [31:0]      dataInMem_lo_158 = {dataInMem_lo_hi_94, dataInMem_lo_lo_30};
  wire [15:0]      dataInMem_hi_hi_126 = {dataRegroupBySew_7_23, dataRegroupBySew_6_23};
  wire [31:0]      dataInMem_hi_190 = {dataInMem_hi_hi_126, dataInMem_hi_lo_62};
  wire [31:0]      dataInMem_lo_159 = {dataInMem_lo_hi_95, dataInMem_lo_lo_31};
  wire [15:0]      dataInMem_hi_hi_127 = {dataRegroupBySew_7_24, dataRegroupBySew_6_24};
  wire [31:0]      dataInMem_hi_191 = {dataInMem_hi_hi_127, dataInMem_hi_lo_63};
  wire [31:0]      dataInMem_lo_160 = {dataInMem_lo_hi_96, dataInMem_lo_lo_32};
  wire [15:0]      dataInMem_hi_hi_128 = {dataRegroupBySew_7_25, dataRegroupBySew_6_25};
  wire [31:0]      dataInMem_hi_192 = {dataInMem_hi_hi_128, dataInMem_hi_lo_64};
  wire [31:0]      dataInMem_lo_161 = {dataInMem_lo_hi_97, dataInMem_lo_lo_33};
  wire [15:0]      dataInMem_hi_hi_129 = {dataRegroupBySew_7_26, dataRegroupBySew_6_26};
  wire [31:0]      dataInMem_hi_193 = {dataInMem_hi_hi_129, dataInMem_hi_lo_65};
  wire [31:0]      dataInMem_lo_162 = {dataInMem_lo_hi_98, dataInMem_lo_lo_34};
  wire [15:0]      dataInMem_hi_hi_130 = {dataRegroupBySew_7_27, dataRegroupBySew_6_27};
  wire [31:0]      dataInMem_hi_194 = {dataInMem_hi_hi_130, dataInMem_hi_lo_66};
  wire [31:0]      dataInMem_lo_163 = {dataInMem_lo_hi_99, dataInMem_lo_lo_35};
  wire [15:0]      dataInMem_hi_hi_131 = {dataRegroupBySew_7_28, dataRegroupBySew_6_28};
  wire [31:0]      dataInMem_hi_195 = {dataInMem_hi_hi_131, dataInMem_hi_lo_67};
  wire [31:0]      dataInMem_lo_164 = {dataInMem_lo_hi_100, dataInMem_lo_lo_36};
  wire [15:0]      dataInMem_hi_hi_132 = {dataRegroupBySew_7_29, dataRegroupBySew_6_29};
  wire [31:0]      dataInMem_hi_196 = {dataInMem_hi_hi_132, dataInMem_hi_lo_68};
  wire [31:0]      dataInMem_lo_165 = {dataInMem_lo_hi_101, dataInMem_lo_lo_37};
  wire [15:0]      dataInMem_hi_hi_133 = {dataRegroupBySew_7_30, dataRegroupBySew_6_30};
  wire [31:0]      dataInMem_hi_197 = {dataInMem_hi_hi_133, dataInMem_hi_lo_69};
  wire [31:0]      dataInMem_lo_166 = {dataInMem_lo_hi_102, dataInMem_lo_lo_38};
  wire [15:0]      dataInMem_hi_hi_134 = {dataRegroupBySew_7_31, dataRegroupBySew_6_31};
  wire [31:0]      dataInMem_hi_198 = {dataInMem_hi_hi_134, dataInMem_hi_lo_70};
  wire [127:0]     dataInMem_lo_lo_lo_lo_7 = {dataInMem_hi_168, dataInMem_lo_136, dataInMem_hi_167, dataInMem_lo_135};
  wire [127:0]     dataInMem_lo_lo_lo_hi_7 = {dataInMem_hi_170, dataInMem_lo_138, dataInMem_hi_169, dataInMem_lo_137};
  wire [255:0]     dataInMem_lo_lo_lo_7 = {dataInMem_lo_lo_lo_hi_7, dataInMem_lo_lo_lo_lo_7};
  wire [127:0]     dataInMem_lo_lo_hi_lo_7 = {dataInMem_hi_172, dataInMem_lo_140, dataInMem_hi_171, dataInMem_lo_139};
  wire [127:0]     dataInMem_lo_lo_hi_hi_7 = {dataInMem_hi_174, dataInMem_lo_142, dataInMem_hi_173, dataInMem_lo_141};
  wire [255:0]     dataInMem_lo_lo_hi_7 = {dataInMem_lo_lo_hi_hi_7, dataInMem_lo_lo_hi_lo_7};
  wire [511:0]     dataInMem_lo_lo_39 = {dataInMem_lo_lo_hi_7, dataInMem_lo_lo_lo_7};
  wire [127:0]     dataInMem_lo_hi_lo_lo_7 = {dataInMem_hi_176, dataInMem_lo_144, dataInMem_hi_175, dataInMem_lo_143};
  wire [127:0]     dataInMem_lo_hi_lo_hi_7 = {dataInMem_hi_178, dataInMem_lo_146, dataInMem_hi_177, dataInMem_lo_145};
  wire [255:0]     dataInMem_lo_hi_lo_7 = {dataInMem_lo_hi_lo_hi_7, dataInMem_lo_hi_lo_lo_7};
  wire [127:0]     dataInMem_lo_hi_hi_lo_7 = {dataInMem_hi_180, dataInMem_lo_148, dataInMem_hi_179, dataInMem_lo_147};
  wire [127:0]     dataInMem_lo_hi_hi_hi_7 = {dataInMem_hi_182, dataInMem_lo_150, dataInMem_hi_181, dataInMem_lo_149};
  wire [255:0]     dataInMem_lo_hi_hi_7 = {dataInMem_lo_hi_hi_hi_7, dataInMem_lo_hi_hi_lo_7};
  wire [511:0]     dataInMem_lo_hi_103 = {dataInMem_lo_hi_hi_7, dataInMem_lo_hi_lo_7};
  wire [1023:0]    dataInMem_lo_167 = {dataInMem_lo_hi_103, dataInMem_lo_lo_39};
  wire [127:0]     dataInMem_hi_lo_lo_lo_7 = {dataInMem_hi_184, dataInMem_lo_152, dataInMem_hi_183, dataInMem_lo_151};
  wire [127:0]     dataInMem_hi_lo_lo_hi_7 = {dataInMem_hi_186, dataInMem_lo_154, dataInMem_hi_185, dataInMem_lo_153};
  wire [255:0]     dataInMem_hi_lo_lo_7 = {dataInMem_hi_lo_lo_hi_7, dataInMem_hi_lo_lo_lo_7};
  wire [127:0]     dataInMem_hi_lo_hi_lo_7 = {dataInMem_hi_188, dataInMem_lo_156, dataInMem_hi_187, dataInMem_lo_155};
  wire [127:0]     dataInMem_hi_lo_hi_hi_7 = {dataInMem_hi_190, dataInMem_lo_158, dataInMem_hi_189, dataInMem_lo_157};
  wire [255:0]     dataInMem_hi_lo_hi_7 = {dataInMem_hi_lo_hi_hi_7, dataInMem_hi_lo_hi_lo_7};
  wire [511:0]     dataInMem_hi_lo_71 = {dataInMem_hi_lo_hi_7, dataInMem_hi_lo_lo_7};
  wire [127:0]     dataInMem_hi_hi_lo_lo_7 = {dataInMem_hi_192, dataInMem_lo_160, dataInMem_hi_191, dataInMem_lo_159};
  wire [127:0]     dataInMem_hi_hi_lo_hi_7 = {dataInMem_hi_194, dataInMem_lo_162, dataInMem_hi_193, dataInMem_lo_161};
  wire [255:0]     dataInMem_hi_hi_lo_7 = {dataInMem_hi_hi_lo_hi_7, dataInMem_hi_hi_lo_lo_7};
  wire [127:0]     dataInMem_hi_hi_hi_lo_7 = {dataInMem_hi_196, dataInMem_lo_164, dataInMem_hi_195, dataInMem_lo_163};
  wire [127:0]     dataInMem_hi_hi_hi_hi_7 = {dataInMem_hi_198, dataInMem_lo_166, dataInMem_hi_197, dataInMem_lo_165};
  wire [255:0]     dataInMem_hi_hi_hi_7 = {dataInMem_hi_hi_hi_hi_7, dataInMem_hi_hi_hi_lo_7};
  wire [511:0]     dataInMem_hi_hi_135 = {dataInMem_hi_hi_hi_7, dataInMem_hi_hi_lo_7};
  wire [1023:0]    dataInMem_hi_199 = {dataInMem_hi_hi_135, dataInMem_hi_lo_71};
  wire [2047:0]    dataInMem_7 = {dataInMem_hi_199, dataInMem_lo_167};
  wire [255:0]     regroupCacheLine_7_0 = dataInMem_7[255:0];
  wire [255:0]     regroupCacheLine_7_1 = dataInMem_7[511:256];
  wire [255:0]     regroupCacheLine_7_2 = dataInMem_7[767:512];
  wire [255:0]     regroupCacheLine_7_3 = dataInMem_7[1023:768];
  wire [255:0]     regroupCacheLine_7_4 = dataInMem_7[1279:1024];
  wire [255:0]     regroupCacheLine_7_5 = dataInMem_7[1535:1280];
  wire [255:0]     regroupCacheLine_7_6 = dataInMem_7[1791:1536];
  wire [255:0]     regroupCacheLine_7_7 = dataInMem_7[2047:1792];
  wire [255:0]     res_56 = regroupCacheLine_7_0;
  wire [255:0]     res_57 = regroupCacheLine_7_1;
  wire [255:0]     res_58 = regroupCacheLine_7_2;
  wire [255:0]     res_59 = regroupCacheLine_7_3;
  wire [255:0]     res_60 = regroupCacheLine_7_4;
  wire [255:0]     res_61 = regroupCacheLine_7_5;
  wire [255:0]     res_62 = regroupCacheLine_7_6;
  wire [255:0]     res_63 = regroupCacheLine_7_7;
  wire [511:0]     lo_lo_7 = {res_57, res_56};
  wire [511:0]     lo_hi_7 = {res_59, res_58};
  wire [1023:0]    lo_7 = {lo_hi_7, lo_lo_7};
  wire [511:0]     hi_lo_7 = {res_61, res_60};
  wire [511:0]     hi_hi_7 = {res_63, res_62};
  wire [1023:0]    hi_7 = {hi_hi_7, hi_lo_7};
  wire [2047:0]    regroupLoadData_0_7 = {hi_7, lo_7};
  wire [15:0]      dataRegroupBySew_0_1_0 = bufferStageEnqueueData_0[15:0];
  wire [15:0]      dataRegroupBySew_0_1_1 = bufferStageEnqueueData_0[31:16];
  wire [15:0]      dataRegroupBySew_0_1_2 = bufferStageEnqueueData_0[47:32];
  wire [15:0]      dataRegroupBySew_0_1_3 = bufferStageEnqueueData_0[63:48];
  wire [15:0]      dataRegroupBySew_0_1_4 = bufferStageEnqueueData_0[79:64];
  wire [15:0]      dataRegroupBySew_0_1_5 = bufferStageEnqueueData_0[95:80];
  wire [15:0]      dataRegroupBySew_0_1_6 = bufferStageEnqueueData_0[111:96];
  wire [15:0]      dataRegroupBySew_0_1_7 = bufferStageEnqueueData_0[127:112];
  wire [15:0]      dataRegroupBySew_0_1_8 = bufferStageEnqueueData_0[143:128];
  wire [15:0]      dataRegroupBySew_0_1_9 = bufferStageEnqueueData_0[159:144];
  wire [15:0]      dataRegroupBySew_0_1_10 = bufferStageEnqueueData_0[175:160];
  wire [15:0]      dataRegroupBySew_0_1_11 = bufferStageEnqueueData_0[191:176];
  wire [15:0]      dataRegroupBySew_0_1_12 = bufferStageEnqueueData_0[207:192];
  wire [15:0]      dataRegroupBySew_0_1_13 = bufferStageEnqueueData_0[223:208];
  wire [15:0]      dataRegroupBySew_0_1_14 = bufferStageEnqueueData_0[239:224];
  wire [15:0]      dataRegroupBySew_0_1_15 = bufferStageEnqueueData_0[255:240];
  wire [15:0]      dataRegroupBySew_1_1_0 = bufferStageEnqueueData_1[15:0];
  wire [15:0]      dataRegroupBySew_1_1_1 = bufferStageEnqueueData_1[31:16];
  wire [15:0]      dataRegroupBySew_1_1_2 = bufferStageEnqueueData_1[47:32];
  wire [15:0]      dataRegroupBySew_1_1_3 = bufferStageEnqueueData_1[63:48];
  wire [15:0]      dataRegroupBySew_1_1_4 = bufferStageEnqueueData_1[79:64];
  wire [15:0]      dataRegroupBySew_1_1_5 = bufferStageEnqueueData_1[95:80];
  wire [15:0]      dataRegroupBySew_1_1_6 = bufferStageEnqueueData_1[111:96];
  wire [15:0]      dataRegroupBySew_1_1_7 = bufferStageEnqueueData_1[127:112];
  wire [15:0]      dataRegroupBySew_1_1_8 = bufferStageEnqueueData_1[143:128];
  wire [15:0]      dataRegroupBySew_1_1_9 = bufferStageEnqueueData_1[159:144];
  wire [15:0]      dataRegroupBySew_1_1_10 = bufferStageEnqueueData_1[175:160];
  wire [15:0]      dataRegroupBySew_1_1_11 = bufferStageEnqueueData_1[191:176];
  wire [15:0]      dataRegroupBySew_1_1_12 = bufferStageEnqueueData_1[207:192];
  wire [15:0]      dataRegroupBySew_1_1_13 = bufferStageEnqueueData_1[223:208];
  wire [15:0]      dataRegroupBySew_1_1_14 = bufferStageEnqueueData_1[239:224];
  wire [15:0]      dataRegroupBySew_1_1_15 = bufferStageEnqueueData_1[255:240];
  wire [15:0]      dataRegroupBySew_2_1_0 = bufferStageEnqueueData_2[15:0];
  wire [15:0]      dataRegroupBySew_2_1_1 = bufferStageEnqueueData_2[31:16];
  wire [15:0]      dataRegroupBySew_2_1_2 = bufferStageEnqueueData_2[47:32];
  wire [15:0]      dataRegroupBySew_2_1_3 = bufferStageEnqueueData_2[63:48];
  wire [15:0]      dataRegroupBySew_2_1_4 = bufferStageEnqueueData_2[79:64];
  wire [15:0]      dataRegroupBySew_2_1_5 = bufferStageEnqueueData_2[95:80];
  wire [15:0]      dataRegroupBySew_2_1_6 = bufferStageEnqueueData_2[111:96];
  wire [15:0]      dataRegroupBySew_2_1_7 = bufferStageEnqueueData_2[127:112];
  wire [15:0]      dataRegroupBySew_2_1_8 = bufferStageEnqueueData_2[143:128];
  wire [15:0]      dataRegroupBySew_2_1_9 = bufferStageEnqueueData_2[159:144];
  wire [15:0]      dataRegroupBySew_2_1_10 = bufferStageEnqueueData_2[175:160];
  wire [15:0]      dataRegroupBySew_2_1_11 = bufferStageEnqueueData_2[191:176];
  wire [15:0]      dataRegroupBySew_2_1_12 = bufferStageEnqueueData_2[207:192];
  wire [15:0]      dataRegroupBySew_2_1_13 = bufferStageEnqueueData_2[223:208];
  wire [15:0]      dataRegroupBySew_2_1_14 = bufferStageEnqueueData_2[239:224];
  wire [15:0]      dataRegroupBySew_2_1_15 = bufferStageEnqueueData_2[255:240];
  wire [15:0]      dataRegroupBySew_3_1_0 = bufferStageEnqueueData_3[15:0];
  wire [15:0]      dataRegroupBySew_3_1_1 = bufferStageEnqueueData_3[31:16];
  wire [15:0]      dataRegroupBySew_3_1_2 = bufferStageEnqueueData_3[47:32];
  wire [15:0]      dataRegroupBySew_3_1_3 = bufferStageEnqueueData_3[63:48];
  wire [15:0]      dataRegroupBySew_3_1_4 = bufferStageEnqueueData_3[79:64];
  wire [15:0]      dataRegroupBySew_3_1_5 = bufferStageEnqueueData_3[95:80];
  wire [15:0]      dataRegroupBySew_3_1_6 = bufferStageEnqueueData_3[111:96];
  wire [15:0]      dataRegroupBySew_3_1_7 = bufferStageEnqueueData_3[127:112];
  wire [15:0]      dataRegroupBySew_3_1_8 = bufferStageEnqueueData_3[143:128];
  wire [15:0]      dataRegroupBySew_3_1_9 = bufferStageEnqueueData_3[159:144];
  wire [15:0]      dataRegroupBySew_3_1_10 = bufferStageEnqueueData_3[175:160];
  wire [15:0]      dataRegroupBySew_3_1_11 = bufferStageEnqueueData_3[191:176];
  wire [15:0]      dataRegroupBySew_3_1_12 = bufferStageEnqueueData_3[207:192];
  wire [15:0]      dataRegroupBySew_3_1_13 = bufferStageEnqueueData_3[223:208];
  wire [15:0]      dataRegroupBySew_3_1_14 = bufferStageEnqueueData_3[239:224];
  wire [15:0]      dataRegroupBySew_3_1_15 = bufferStageEnqueueData_3[255:240];
  wire [15:0]      dataRegroupBySew_4_1_0 = bufferStageEnqueueData_4[15:0];
  wire [15:0]      dataRegroupBySew_4_1_1 = bufferStageEnqueueData_4[31:16];
  wire [15:0]      dataRegroupBySew_4_1_2 = bufferStageEnqueueData_4[47:32];
  wire [15:0]      dataRegroupBySew_4_1_3 = bufferStageEnqueueData_4[63:48];
  wire [15:0]      dataRegroupBySew_4_1_4 = bufferStageEnqueueData_4[79:64];
  wire [15:0]      dataRegroupBySew_4_1_5 = bufferStageEnqueueData_4[95:80];
  wire [15:0]      dataRegroupBySew_4_1_6 = bufferStageEnqueueData_4[111:96];
  wire [15:0]      dataRegroupBySew_4_1_7 = bufferStageEnqueueData_4[127:112];
  wire [15:0]      dataRegroupBySew_4_1_8 = bufferStageEnqueueData_4[143:128];
  wire [15:0]      dataRegroupBySew_4_1_9 = bufferStageEnqueueData_4[159:144];
  wire [15:0]      dataRegroupBySew_4_1_10 = bufferStageEnqueueData_4[175:160];
  wire [15:0]      dataRegroupBySew_4_1_11 = bufferStageEnqueueData_4[191:176];
  wire [15:0]      dataRegroupBySew_4_1_12 = bufferStageEnqueueData_4[207:192];
  wire [15:0]      dataRegroupBySew_4_1_13 = bufferStageEnqueueData_4[223:208];
  wire [15:0]      dataRegroupBySew_4_1_14 = bufferStageEnqueueData_4[239:224];
  wire [15:0]      dataRegroupBySew_4_1_15 = bufferStageEnqueueData_4[255:240];
  wire [15:0]      dataRegroupBySew_5_1_0 = bufferStageEnqueueData_5[15:0];
  wire [15:0]      dataRegroupBySew_5_1_1 = bufferStageEnqueueData_5[31:16];
  wire [15:0]      dataRegroupBySew_5_1_2 = bufferStageEnqueueData_5[47:32];
  wire [15:0]      dataRegroupBySew_5_1_3 = bufferStageEnqueueData_5[63:48];
  wire [15:0]      dataRegroupBySew_5_1_4 = bufferStageEnqueueData_5[79:64];
  wire [15:0]      dataRegroupBySew_5_1_5 = bufferStageEnqueueData_5[95:80];
  wire [15:0]      dataRegroupBySew_5_1_6 = bufferStageEnqueueData_5[111:96];
  wire [15:0]      dataRegroupBySew_5_1_7 = bufferStageEnqueueData_5[127:112];
  wire [15:0]      dataRegroupBySew_5_1_8 = bufferStageEnqueueData_5[143:128];
  wire [15:0]      dataRegroupBySew_5_1_9 = bufferStageEnqueueData_5[159:144];
  wire [15:0]      dataRegroupBySew_5_1_10 = bufferStageEnqueueData_5[175:160];
  wire [15:0]      dataRegroupBySew_5_1_11 = bufferStageEnqueueData_5[191:176];
  wire [15:0]      dataRegroupBySew_5_1_12 = bufferStageEnqueueData_5[207:192];
  wire [15:0]      dataRegroupBySew_5_1_13 = bufferStageEnqueueData_5[223:208];
  wire [15:0]      dataRegroupBySew_5_1_14 = bufferStageEnqueueData_5[239:224];
  wire [15:0]      dataRegroupBySew_5_1_15 = bufferStageEnqueueData_5[255:240];
  wire [15:0]      dataRegroupBySew_6_1_0 = bufferStageEnqueueData_6[15:0];
  wire [15:0]      dataRegroupBySew_6_1_1 = bufferStageEnqueueData_6[31:16];
  wire [15:0]      dataRegroupBySew_6_1_2 = bufferStageEnqueueData_6[47:32];
  wire [15:0]      dataRegroupBySew_6_1_3 = bufferStageEnqueueData_6[63:48];
  wire [15:0]      dataRegroupBySew_6_1_4 = bufferStageEnqueueData_6[79:64];
  wire [15:0]      dataRegroupBySew_6_1_5 = bufferStageEnqueueData_6[95:80];
  wire [15:0]      dataRegroupBySew_6_1_6 = bufferStageEnqueueData_6[111:96];
  wire [15:0]      dataRegroupBySew_6_1_7 = bufferStageEnqueueData_6[127:112];
  wire [15:0]      dataRegroupBySew_6_1_8 = bufferStageEnqueueData_6[143:128];
  wire [15:0]      dataRegroupBySew_6_1_9 = bufferStageEnqueueData_6[159:144];
  wire [15:0]      dataRegroupBySew_6_1_10 = bufferStageEnqueueData_6[175:160];
  wire [15:0]      dataRegroupBySew_6_1_11 = bufferStageEnqueueData_6[191:176];
  wire [15:0]      dataRegroupBySew_6_1_12 = bufferStageEnqueueData_6[207:192];
  wire [15:0]      dataRegroupBySew_6_1_13 = bufferStageEnqueueData_6[223:208];
  wire [15:0]      dataRegroupBySew_6_1_14 = bufferStageEnqueueData_6[239:224];
  wire [15:0]      dataRegroupBySew_6_1_15 = bufferStageEnqueueData_6[255:240];
  wire [15:0]      dataRegroupBySew_7_1_0 = bufferStageEnqueueData_7[15:0];
  wire [15:0]      dataRegroupBySew_7_1_1 = bufferStageEnqueueData_7[31:16];
  wire [15:0]      dataRegroupBySew_7_1_2 = bufferStageEnqueueData_7[47:32];
  wire [15:0]      dataRegroupBySew_7_1_3 = bufferStageEnqueueData_7[63:48];
  wire [15:0]      dataRegroupBySew_7_1_4 = bufferStageEnqueueData_7[79:64];
  wire [15:0]      dataRegroupBySew_7_1_5 = bufferStageEnqueueData_7[95:80];
  wire [15:0]      dataRegroupBySew_7_1_6 = bufferStageEnqueueData_7[111:96];
  wire [15:0]      dataRegroupBySew_7_1_7 = bufferStageEnqueueData_7[127:112];
  wire [15:0]      dataRegroupBySew_7_1_8 = bufferStageEnqueueData_7[143:128];
  wire [15:0]      dataRegroupBySew_7_1_9 = bufferStageEnqueueData_7[159:144];
  wire [15:0]      dataRegroupBySew_7_1_10 = bufferStageEnqueueData_7[175:160];
  wire [15:0]      dataRegroupBySew_7_1_11 = bufferStageEnqueueData_7[191:176];
  wire [15:0]      dataRegroupBySew_7_1_12 = bufferStageEnqueueData_7[207:192];
  wire [15:0]      dataRegroupBySew_7_1_13 = bufferStageEnqueueData_7[223:208];
  wire [15:0]      dataRegroupBySew_7_1_14 = bufferStageEnqueueData_7[239:224];
  wire [15:0]      dataRegroupBySew_7_1_15 = bufferStageEnqueueData_7[255:240];
  wire [31:0]      dataInMem_lo_lo_lo_8 = {dataRegroupBySew_0_1_1, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_lo_lo_hi_8 = {dataRegroupBySew_0_1_3, dataRegroupBySew_0_1_2};
  wire [63:0]      dataInMem_lo_lo_40 = {dataInMem_lo_lo_hi_8, dataInMem_lo_lo_lo_8};
  wire [31:0]      dataInMem_lo_hi_lo_8 = {dataRegroupBySew_0_1_5, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_lo_hi_hi_8 = {dataRegroupBySew_0_1_7, dataRegroupBySew_0_1_6};
  wire [63:0]      dataInMem_lo_hi_104 = {dataInMem_lo_hi_hi_8, dataInMem_lo_hi_lo_8};
  wire [127:0]     dataInMem_lo_168 = {dataInMem_lo_hi_104, dataInMem_lo_lo_40};
  wire [31:0]      dataInMem_hi_lo_lo_8 = {dataRegroupBySew_0_1_9, dataRegroupBySew_0_1_8};
  wire [31:0]      dataInMem_hi_lo_hi_8 = {dataRegroupBySew_0_1_11, dataRegroupBySew_0_1_10};
  wire [63:0]      dataInMem_hi_lo_72 = {dataInMem_hi_lo_hi_8, dataInMem_hi_lo_lo_8};
  wire [31:0]      dataInMem_hi_hi_lo_8 = {dataRegroupBySew_0_1_13, dataRegroupBySew_0_1_12};
  wire [31:0]      dataInMem_hi_hi_hi_8 = {dataRegroupBySew_0_1_15, dataRegroupBySew_0_1_14};
  wire [63:0]      dataInMem_hi_hi_136 = {dataInMem_hi_hi_hi_8, dataInMem_hi_hi_lo_8};
  wire [127:0]     dataInMem_hi_200 = {dataInMem_hi_hi_136, dataInMem_hi_lo_72};
  wire [255:0]     dataInMem_8 = {dataInMem_hi_200, dataInMem_lo_168};
  wire [255:0]     regroupCacheLine_8_0 = dataInMem_8;
  wire [255:0]     res_64 = regroupCacheLine_8_0;
  wire [511:0]     lo_lo_8 = {256'h0, res_64};
  wire [1023:0]    lo_8 = {512'h0, lo_lo_8};
  wire [2047:0]    regroupLoadData_1_0 = {1024'h0, lo_8};
  wire [63:0]      dataInMem_lo_lo_lo_9 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1, dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [63:0]      dataInMem_lo_lo_hi_9 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3, dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [127:0]     dataInMem_lo_lo_41 = {dataInMem_lo_lo_hi_9, dataInMem_lo_lo_lo_9};
  wire [63:0]      dataInMem_lo_hi_lo_9 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5, dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [63:0]      dataInMem_lo_hi_hi_9 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7, dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [127:0]     dataInMem_lo_hi_105 = {dataInMem_lo_hi_hi_9, dataInMem_lo_hi_lo_9};
  wire [255:0]     dataInMem_lo_169 = {dataInMem_lo_hi_105, dataInMem_lo_lo_41};
  wire [63:0]      dataInMem_hi_lo_lo_9 = {dataRegroupBySew_1_1_9, dataRegroupBySew_0_1_9, dataRegroupBySew_1_1_8, dataRegroupBySew_0_1_8};
  wire [63:0]      dataInMem_hi_lo_hi_9 = {dataRegroupBySew_1_1_11, dataRegroupBySew_0_1_11, dataRegroupBySew_1_1_10, dataRegroupBySew_0_1_10};
  wire [127:0]     dataInMem_hi_lo_73 = {dataInMem_hi_lo_hi_9, dataInMem_hi_lo_lo_9};
  wire [63:0]      dataInMem_hi_hi_lo_9 = {dataRegroupBySew_1_1_13, dataRegroupBySew_0_1_13, dataRegroupBySew_1_1_12, dataRegroupBySew_0_1_12};
  wire [63:0]      dataInMem_hi_hi_hi_9 = {dataRegroupBySew_1_1_15, dataRegroupBySew_0_1_15, dataRegroupBySew_1_1_14, dataRegroupBySew_0_1_14};
  wire [127:0]     dataInMem_hi_hi_137 = {dataInMem_hi_hi_hi_9, dataInMem_hi_hi_lo_9};
  wire [255:0]     dataInMem_hi_201 = {dataInMem_hi_hi_137, dataInMem_hi_lo_73};
  wire [511:0]     dataInMem_9 = {dataInMem_hi_201, dataInMem_lo_169};
  wire [255:0]     regroupCacheLine_9_0 = dataInMem_9[255:0];
  wire [255:0]     regroupCacheLine_9_1 = dataInMem_9[511:256];
  wire [255:0]     res_72 = regroupCacheLine_9_0;
  wire [255:0]     res_73 = regroupCacheLine_9_1;
  wire [511:0]     lo_lo_9 = {res_73, res_72};
  wire [1023:0]    lo_9 = {512'h0, lo_lo_9};
  wire [2047:0]    regroupLoadData_1_1 = {1024'h0, lo_9};
  wire [31:0]      _GEN_164 = {dataRegroupBySew_2_1_0, dataRegroupBySew_1_1_0};
  wire [31:0]      dataInMem_hi_202;
  assign dataInMem_hi_202 = _GEN_164;
  wire [31:0]      dataInMem_lo_hi_109;
  assign dataInMem_lo_hi_109 = _GEN_164;
  wire [31:0]      dataInMem_lo_hi_126;
  assign dataInMem_lo_hi_126 = _GEN_164;
  wire [31:0]      _GEN_165 = {dataRegroupBySew_2_1_1, dataRegroupBySew_1_1_1};
  wire [31:0]      dataInMem_hi_203;
  assign dataInMem_hi_203 = _GEN_165;
  wire [31:0]      dataInMem_lo_hi_110;
  assign dataInMem_lo_hi_110 = _GEN_165;
  wire [31:0]      dataInMem_lo_hi_127;
  assign dataInMem_lo_hi_127 = _GEN_165;
  wire [31:0]      _GEN_166 = {dataRegroupBySew_2_1_2, dataRegroupBySew_1_1_2};
  wire [31:0]      dataInMem_hi_204;
  assign dataInMem_hi_204 = _GEN_166;
  wire [31:0]      dataInMem_lo_hi_111;
  assign dataInMem_lo_hi_111 = _GEN_166;
  wire [31:0]      dataInMem_lo_hi_128;
  assign dataInMem_lo_hi_128 = _GEN_166;
  wire [31:0]      _GEN_167 = {dataRegroupBySew_2_1_3, dataRegroupBySew_1_1_3};
  wire [31:0]      dataInMem_hi_205;
  assign dataInMem_hi_205 = _GEN_167;
  wire [31:0]      dataInMem_lo_hi_112;
  assign dataInMem_lo_hi_112 = _GEN_167;
  wire [31:0]      dataInMem_lo_hi_129;
  assign dataInMem_lo_hi_129 = _GEN_167;
  wire [31:0]      _GEN_168 = {dataRegroupBySew_2_1_4, dataRegroupBySew_1_1_4};
  wire [31:0]      dataInMem_hi_206;
  assign dataInMem_hi_206 = _GEN_168;
  wire [31:0]      dataInMem_lo_hi_113;
  assign dataInMem_lo_hi_113 = _GEN_168;
  wire [31:0]      dataInMem_lo_hi_130;
  assign dataInMem_lo_hi_130 = _GEN_168;
  wire [31:0]      _GEN_169 = {dataRegroupBySew_2_1_5, dataRegroupBySew_1_1_5};
  wire [31:0]      dataInMem_hi_207;
  assign dataInMem_hi_207 = _GEN_169;
  wire [31:0]      dataInMem_lo_hi_114;
  assign dataInMem_lo_hi_114 = _GEN_169;
  wire [31:0]      dataInMem_lo_hi_131;
  assign dataInMem_lo_hi_131 = _GEN_169;
  wire [31:0]      _GEN_170 = {dataRegroupBySew_2_1_6, dataRegroupBySew_1_1_6};
  wire [31:0]      dataInMem_hi_208;
  assign dataInMem_hi_208 = _GEN_170;
  wire [31:0]      dataInMem_lo_hi_115;
  assign dataInMem_lo_hi_115 = _GEN_170;
  wire [31:0]      dataInMem_lo_hi_132;
  assign dataInMem_lo_hi_132 = _GEN_170;
  wire [31:0]      _GEN_171 = {dataRegroupBySew_2_1_7, dataRegroupBySew_1_1_7};
  wire [31:0]      dataInMem_hi_209;
  assign dataInMem_hi_209 = _GEN_171;
  wire [31:0]      dataInMem_lo_hi_116;
  assign dataInMem_lo_hi_116 = _GEN_171;
  wire [31:0]      dataInMem_lo_hi_133;
  assign dataInMem_lo_hi_133 = _GEN_171;
  wire [31:0]      _GEN_172 = {dataRegroupBySew_2_1_8, dataRegroupBySew_1_1_8};
  wire [31:0]      dataInMem_hi_210;
  assign dataInMem_hi_210 = _GEN_172;
  wire [31:0]      dataInMem_lo_hi_117;
  assign dataInMem_lo_hi_117 = _GEN_172;
  wire [31:0]      dataInMem_lo_hi_134;
  assign dataInMem_lo_hi_134 = _GEN_172;
  wire [31:0]      _GEN_173 = {dataRegroupBySew_2_1_9, dataRegroupBySew_1_1_9};
  wire [31:0]      dataInMem_hi_211;
  assign dataInMem_hi_211 = _GEN_173;
  wire [31:0]      dataInMem_lo_hi_118;
  assign dataInMem_lo_hi_118 = _GEN_173;
  wire [31:0]      dataInMem_lo_hi_135;
  assign dataInMem_lo_hi_135 = _GEN_173;
  wire [31:0]      _GEN_174 = {dataRegroupBySew_2_1_10, dataRegroupBySew_1_1_10};
  wire [31:0]      dataInMem_hi_212;
  assign dataInMem_hi_212 = _GEN_174;
  wire [31:0]      dataInMem_lo_hi_119;
  assign dataInMem_lo_hi_119 = _GEN_174;
  wire [31:0]      dataInMem_lo_hi_136;
  assign dataInMem_lo_hi_136 = _GEN_174;
  wire [31:0]      _GEN_175 = {dataRegroupBySew_2_1_11, dataRegroupBySew_1_1_11};
  wire [31:0]      dataInMem_hi_213;
  assign dataInMem_hi_213 = _GEN_175;
  wire [31:0]      dataInMem_lo_hi_120;
  assign dataInMem_lo_hi_120 = _GEN_175;
  wire [31:0]      dataInMem_lo_hi_137;
  assign dataInMem_lo_hi_137 = _GEN_175;
  wire [31:0]      _GEN_176 = {dataRegroupBySew_2_1_12, dataRegroupBySew_1_1_12};
  wire [31:0]      dataInMem_hi_214;
  assign dataInMem_hi_214 = _GEN_176;
  wire [31:0]      dataInMem_lo_hi_121;
  assign dataInMem_lo_hi_121 = _GEN_176;
  wire [31:0]      dataInMem_lo_hi_138;
  assign dataInMem_lo_hi_138 = _GEN_176;
  wire [31:0]      _GEN_177 = {dataRegroupBySew_2_1_13, dataRegroupBySew_1_1_13};
  wire [31:0]      dataInMem_hi_215;
  assign dataInMem_hi_215 = _GEN_177;
  wire [31:0]      dataInMem_lo_hi_122;
  assign dataInMem_lo_hi_122 = _GEN_177;
  wire [31:0]      dataInMem_lo_hi_139;
  assign dataInMem_lo_hi_139 = _GEN_177;
  wire [31:0]      _GEN_178 = {dataRegroupBySew_2_1_14, dataRegroupBySew_1_1_14};
  wire [31:0]      dataInMem_hi_216;
  assign dataInMem_hi_216 = _GEN_178;
  wire [31:0]      dataInMem_lo_hi_123;
  assign dataInMem_lo_hi_123 = _GEN_178;
  wire [31:0]      dataInMem_lo_hi_140;
  assign dataInMem_lo_hi_140 = _GEN_178;
  wire [31:0]      _GEN_179 = {dataRegroupBySew_2_1_15, dataRegroupBySew_1_1_15};
  wire [31:0]      dataInMem_hi_217;
  assign dataInMem_hi_217 = _GEN_179;
  wire [31:0]      dataInMem_lo_hi_124;
  assign dataInMem_lo_hi_124 = _GEN_179;
  wire [31:0]      dataInMem_lo_hi_141;
  assign dataInMem_lo_hi_141 = _GEN_179;
  wire [95:0]      dataInMem_lo_lo_lo_10 = {dataInMem_hi_203, dataRegroupBySew_0_1_1, dataInMem_hi_202, dataRegroupBySew_0_1_0};
  wire [95:0]      dataInMem_lo_lo_hi_10 = {dataInMem_hi_205, dataRegroupBySew_0_1_3, dataInMem_hi_204, dataRegroupBySew_0_1_2};
  wire [191:0]     dataInMem_lo_lo_42 = {dataInMem_lo_lo_hi_10, dataInMem_lo_lo_lo_10};
  wire [95:0]      dataInMem_lo_hi_lo_10 = {dataInMem_hi_207, dataRegroupBySew_0_1_5, dataInMem_hi_206, dataRegroupBySew_0_1_4};
  wire [95:0]      dataInMem_lo_hi_hi_10 = {dataInMem_hi_209, dataRegroupBySew_0_1_7, dataInMem_hi_208, dataRegroupBySew_0_1_6};
  wire [191:0]     dataInMem_lo_hi_106 = {dataInMem_lo_hi_hi_10, dataInMem_lo_hi_lo_10};
  wire [383:0]     dataInMem_lo_170 = {dataInMem_lo_hi_106, dataInMem_lo_lo_42};
  wire [95:0]      dataInMem_hi_lo_lo_10 = {dataInMem_hi_211, dataRegroupBySew_0_1_9, dataInMem_hi_210, dataRegroupBySew_0_1_8};
  wire [95:0]      dataInMem_hi_lo_hi_10 = {dataInMem_hi_213, dataRegroupBySew_0_1_11, dataInMem_hi_212, dataRegroupBySew_0_1_10};
  wire [191:0]     dataInMem_hi_lo_74 = {dataInMem_hi_lo_hi_10, dataInMem_hi_lo_lo_10};
  wire [95:0]      dataInMem_hi_hi_lo_10 = {dataInMem_hi_215, dataRegroupBySew_0_1_13, dataInMem_hi_214, dataRegroupBySew_0_1_12};
  wire [95:0]      dataInMem_hi_hi_hi_10 = {dataInMem_hi_217, dataRegroupBySew_0_1_15, dataInMem_hi_216, dataRegroupBySew_0_1_14};
  wire [191:0]     dataInMem_hi_hi_138 = {dataInMem_hi_hi_hi_10, dataInMem_hi_hi_lo_10};
  wire [383:0]     dataInMem_hi_218 = {dataInMem_hi_hi_138, dataInMem_hi_lo_74};
  wire [767:0]     dataInMem_10 = {dataInMem_hi_218, dataInMem_lo_170};
  wire [255:0]     regroupCacheLine_10_0 = dataInMem_10[255:0];
  wire [255:0]     regroupCacheLine_10_1 = dataInMem_10[511:256];
  wire [255:0]     regroupCacheLine_10_2 = dataInMem_10[767:512];
  wire [255:0]     res_80 = regroupCacheLine_10_0;
  wire [255:0]     res_81 = regroupCacheLine_10_1;
  wire [255:0]     res_82 = regroupCacheLine_10_2;
  wire [511:0]     lo_lo_10 = {res_81, res_80};
  wire [511:0]     lo_hi_10 = {256'h0, res_82};
  wire [1023:0]    lo_10 = {lo_hi_10, lo_lo_10};
  wire [2047:0]    regroupLoadData_1_2 = {1024'h0, lo_10};
  wire [31:0]      _GEN_180 = {dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_lo_171;
  assign dataInMem_lo_171 = _GEN_180;
  wire [31:0]      dataInMem_lo_188;
  assign dataInMem_lo_188 = _GEN_180;
  wire [31:0]      dataInMem_lo_lo_47;
  assign dataInMem_lo_lo_47 = _GEN_180;
  wire [31:0]      _GEN_181 = {dataRegroupBySew_3_1_0, dataRegroupBySew_2_1_0};
  wire [31:0]      dataInMem_hi_219;
  assign dataInMem_hi_219 = _GEN_181;
  wire [31:0]      dataInMem_lo_hi_143;
  assign dataInMem_lo_hi_143 = _GEN_181;
  wire [31:0]      _GEN_182 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1};
  wire [31:0]      dataInMem_lo_172;
  assign dataInMem_lo_172 = _GEN_182;
  wire [31:0]      dataInMem_lo_189;
  assign dataInMem_lo_189 = _GEN_182;
  wire [31:0]      dataInMem_lo_lo_48;
  assign dataInMem_lo_lo_48 = _GEN_182;
  wire [31:0]      _GEN_183 = {dataRegroupBySew_3_1_1, dataRegroupBySew_2_1_1};
  wire [31:0]      dataInMem_hi_220;
  assign dataInMem_hi_220 = _GEN_183;
  wire [31:0]      dataInMem_lo_hi_144;
  assign dataInMem_lo_hi_144 = _GEN_183;
  wire [31:0]      _GEN_184 = {dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [31:0]      dataInMem_lo_173;
  assign dataInMem_lo_173 = _GEN_184;
  wire [31:0]      dataInMem_lo_190;
  assign dataInMem_lo_190 = _GEN_184;
  wire [31:0]      dataInMem_lo_lo_49;
  assign dataInMem_lo_lo_49 = _GEN_184;
  wire [31:0]      _GEN_185 = {dataRegroupBySew_3_1_2, dataRegroupBySew_2_1_2};
  wire [31:0]      dataInMem_hi_221;
  assign dataInMem_hi_221 = _GEN_185;
  wire [31:0]      dataInMem_lo_hi_145;
  assign dataInMem_lo_hi_145 = _GEN_185;
  wire [31:0]      _GEN_186 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3};
  wire [31:0]      dataInMem_lo_174;
  assign dataInMem_lo_174 = _GEN_186;
  wire [31:0]      dataInMem_lo_191;
  assign dataInMem_lo_191 = _GEN_186;
  wire [31:0]      dataInMem_lo_lo_50;
  assign dataInMem_lo_lo_50 = _GEN_186;
  wire [31:0]      _GEN_187 = {dataRegroupBySew_3_1_3, dataRegroupBySew_2_1_3};
  wire [31:0]      dataInMem_hi_222;
  assign dataInMem_hi_222 = _GEN_187;
  wire [31:0]      dataInMem_lo_hi_146;
  assign dataInMem_lo_hi_146 = _GEN_187;
  wire [31:0]      _GEN_188 = {dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_lo_175;
  assign dataInMem_lo_175 = _GEN_188;
  wire [31:0]      dataInMem_lo_192;
  assign dataInMem_lo_192 = _GEN_188;
  wire [31:0]      dataInMem_lo_lo_51;
  assign dataInMem_lo_lo_51 = _GEN_188;
  wire [31:0]      _GEN_189 = {dataRegroupBySew_3_1_4, dataRegroupBySew_2_1_4};
  wire [31:0]      dataInMem_hi_223;
  assign dataInMem_hi_223 = _GEN_189;
  wire [31:0]      dataInMem_lo_hi_147;
  assign dataInMem_lo_hi_147 = _GEN_189;
  wire [31:0]      _GEN_190 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5};
  wire [31:0]      dataInMem_lo_176;
  assign dataInMem_lo_176 = _GEN_190;
  wire [31:0]      dataInMem_lo_193;
  assign dataInMem_lo_193 = _GEN_190;
  wire [31:0]      dataInMem_lo_lo_52;
  assign dataInMem_lo_lo_52 = _GEN_190;
  wire [31:0]      _GEN_191 = {dataRegroupBySew_3_1_5, dataRegroupBySew_2_1_5};
  wire [31:0]      dataInMem_hi_224;
  assign dataInMem_hi_224 = _GEN_191;
  wire [31:0]      dataInMem_lo_hi_148;
  assign dataInMem_lo_hi_148 = _GEN_191;
  wire [31:0]      _GEN_192 = {dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [31:0]      dataInMem_lo_177;
  assign dataInMem_lo_177 = _GEN_192;
  wire [31:0]      dataInMem_lo_194;
  assign dataInMem_lo_194 = _GEN_192;
  wire [31:0]      dataInMem_lo_lo_53;
  assign dataInMem_lo_lo_53 = _GEN_192;
  wire [31:0]      _GEN_193 = {dataRegroupBySew_3_1_6, dataRegroupBySew_2_1_6};
  wire [31:0]      dataInMem_hi_225;
  assign dataInMem_hi_225 = _GEN_193;
  wire [31:0]      dataInMem_lo_hi_149;
  assign dataInMem_lo_hi_149 = _GEN_193;
  wire [31:0]      _GEN_194 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7};
  wire [31:0]      dataInMem_lo_178;
  assign dataInMem_lo_178 = _GEN_194;
  wire [31:0]      dataInMem_lo_195;
  assign dataInMem_lo_195 = _GEN_194;
  wire [31:0]      dataInMem_lo_lo_54;
  assign dataInMem_lo_lo_54 = _GEN_194;
  wire [31:0]      _GEN_195 = {dataRegroupBySew_3_1_7, dataRegroupBySew_2_1_7};
  wire [31:0]      dataInMem_hi_226;
  assign dataInMem_hi_226 = _GEN_195;
  wire [31:0]      dataInMem_lo_hi_150;
  assign dataInMem_lo_hi_150 = _GEN_195;
  wire [31:0]      _GEN_196 = {dataRegroupBySew_1_1_8, dataRegroupBySew_0_1_8};
  wire [31:0]      dataInMem_lo_179;
  assign dataInMem_lo_179 = _GEN_196;
  wire [31:0]      dataInMem_lo_196;
  assign dataInMem_lo_196 = _GEN_196;
  wire [31:0]      dataInMem_lo_lo_55;
  assign dataInMem_lo_lo_55 = _GEN_196;
  wire [31:0]      _GEN_197 = {dataRegroupBySew_3_1_8, dataRegroupBySew_2_1_8};
  wire [31:0]      dataInMem_hi_227;
  assign dataInMem_hi_227 = _GEN_197;
  wire [31:0]      dataInMem_lo_hi_151;
  assign dataInMem_lo_hi_151 = _GEN_197;
  wire [31:0]      _GEN_198 = {dataRegroupBySew_1_1_9, dataRegroupBySew_0_1_9};
  wire [31:0]      dataInMem_lo_180;
  assign dataInMem_lo_180 = _GEN_198;
  wire [31:0]      dataInMem_lo_197;
  assign dataInMem_lo_197 = _GEN_198;
  wire [31:0]      dataInMem_lo_lo_56;
  assign dataInMem_lo_lo_56 = _GEN_198;
  wire [31:0]      _GEN_199 = {dataRegroupBySew_3_1_9, dataRegroupBySew_2_1_9};
  wire [31:0]      dataInMem_hi_228;
  assign dataInMem_hi_228 = _GEN_199;
  wire [31:0]      dataInMem_lo_hi_152;
  assign dataInMem_lo_hi_152 = _GEN_199;
  wire [31:0]      _GEN_200 = {dataRegroupBySew_1_1_10, dataRegroupBySew_0_1_10};
  wire [31:0]      dataInMem_lo_181;
  assign dataInMem_lo_181 = _GEN_200;
  wire [31:0]      dataInMem_lo_198;
  assign dataInMem_lo_198 = _GEN_200;
  wire [31:0]      dataInMem_lo_lo_57;
  assign dataInMem_lo_lo_57 = _GEN_200;
  wire [31:0]      _GEN_201 = {dataRegroupBySew_3_1_10, dataRegroupBySew_2_1_10};
  wire [31:0]      dataInMem_hi_229;
  assign dataInMem_hi_229 = _GEN_201;
  wire [31:0]      dataInMem_lo_hi_153;
  assign dataInMem_lo_hi_153 = _GEN_201;
  wire [31:0]      _GEN_202 = {dataRegroupBySew_1_1_11, dataRegroupBySew_0_1_11};
  wire [31:0]      dataInMem_lo_182;
  assign dataInMem_lo_182 = _GEN_202;
  wire [31:0]      dataInMem_lo_199;
  assign dataInMem_lo_199 = _GEN_202;
  wire [31:0]      dataInMem_lo_lo_58;
  assign dataInMem_lo_lo_58 = _GEN_202;
  wire [31:0]      _GEN_203 = {dataRegroupBySew_3_1_11, dataRegroupBySew_2_1_11};
  wire [31:0]      dataInMem_hi_230;
  assign dataInMem_hi_230 = _GEN_203;
  wire [31:0]      dataInMem_lo_hi_154;
  assign dataInMem_lo_hi_154 = _GEN_203;
  wire [31:0]      _GEN_204 = {dataRegroupBySew_1_1_12, dataRegroupBySew_0_1_12};
  wire [31:0]      dataInMem_lo_183;
  assign dataInMem_lo_183 = _GEN_204;
  wire [31:0]      dataInMem_lo_200;
  assign dataInMem_lo_200 = _GEN_204;
  wire [31:0]      dataInMem_lo_lo_59;
  assign dataInMem_lo_lo_59 = _GEN_204;
  wire [31:0]      _GEN_205 = {dataRegroupBySew_3_1_12, dataRegroupBySew_2_1_12};
  wire [31:0]      dataInMem_hi_231;
  assign dataInMem_hi_231 = _GEN_205;
  wire [31:0]      dataInMem_lo_hi_155;
  assign dataInMem_lo_hi_155 = _GEN_205;
  wire [31:0]      _GEN_206 = {dataRegroupBySew_1_1_13, dataRegroupBySew_0_1_13};
  wire [31:0]      dataInMem_lo_184;
  assign dataInMem_lo_184 = _GEN_206;
  wire [31:0]      dataInMem_lo_201;
  assign dataInMem_lo_201 = _GEN_206;
  wire [31:0]      dataInMem_lo_lo_60;
  assign dataInMem_lo_lo_60 = _GEN_206;
  wire [31:0]      _GEN_207 = {dataRegroupBySew_3_1_13, dataRegroupBySew_2_1_13};
  wire [31:0]      dataInMem_hi_232;
  assign dataInMem_hi_232 = _GEN_207;
  wire [31:0]      dataInMem_lo_hi_156;
  assign dataInMem_lo_hi_156 = _GEN_207;
  wire [31:0]      _GEN_208 = {dataRegroupBySew_1_1_14, dataRegroupBySew_0_1_14};
  wire [31:0]      dataInMem_lo_185;
  assign dataInMem_lo_185 = _GEN_208;
  wire [31:0]      dataInMem_lo_202;
  assign dataInMem_lo_202 = _GEN_208;
  wire [31:0]      dataInMem_lo_lo_61;
  assign dataInMem_lo_lo_61 = _GEN_208;
  wire [31:0]      _GEN_209 = {dataRegroupBySew_3_1_14, dataRegroupBySew_2_1_14};
  wire [31:0]      dataInMem_hi_233;
  assign dataInMem_hi_233 = _GEN_209;
  wire [31:0]      dataInMem_lo_hi_157;
  assign dataInMem_lo_hi_157 = _GEN_209;
  wire [31:0]      _GEN_210 = {dataRegroupBySew_1_1_15, dataRegroupBySew_0_1_15};
  wire [31:0]      dataInMem_lo_186;
  assign dataInMem_lo_186 = _GEN_210;
  wire [31:0]      dataInMem_lo_203;
  assign dataInMem_lo_203 = _GEN_210;
  wire [31:0]      dataInMem_lo_lo_62;
  assign dataInMem_lo_lo_62 = _GEN_210;
  wire [31:0]      _GEN_211 = {dataRegroupBySew_3_1_15, dataRegroupBySew_2_1_15};
  wire [31:0]      dataInMem_hi_234;
  assign dataInMem_hi_234 = _GEN_211;
  wire [31:0]      dataInMem_lo_hi_158;
  assign dataInMem_lo_hi_158 = _GEN_211;
  wire [127:0]     dataInMem_lo_lo_lo_11 = {dataInMem_hi_220, dataInMem_lo_172, dataInMem_hi_219, dataInMem_lo_171};
  wire [127:0]     dataInMem_lo_lo_hi_11 = {dataInMem_hi_222, dataInMem_lo_174, dataInMem_hi_221, dataInMem_lo_173};
  wire [255:0]     dataInMem_lo_lo_43 = {dataInMem_lo_lo_hi_11, dataInMem_lo_lo_lo_11};
  wire [127:0]     dataInMem_lo_hi_lo_11 = {dataInMem_hi_224, dataInMem_lo_176, dataInMem_hi_223, dataInMem_lo_175};
  wire [127:0]     dataInMem_lo_hi_hi_11 = {dataInMem_hi_226, dataInMem_lo_178, dataInMem_hi_225, dataInMem_lo_177};
  wire [255:0]     dataInMem_lo_hi_107 = {dataInMem_lo_hi_hi_11, dataInMem_lo_hi_lo_11};
  wire [511:0]     dataInMem_lo_187 = {dataInMem_lo_hi_107, dataInMem_lo_lo_43};
  wire [127:0]     dataInMem_hi_lo_lo_11 = {dataInMem_hi_228, dataInMem_lo_180, dataInMem_hi_227, dataInMem_lo_179};
  wire [127:0]     dataInMem_hi_lo_hi_11 = {dataInMem_hi_230, dataInMem_lo_182, dataInMem_hi_229, dataInMem_lo_181};
  wire [255:0]     dataInMem_hi_lo_75 = {dataInMem_hi_lo_hi_11, dataInMem_hi_lo_lo_11};
  wire [127:0]     dataInMem_hi_hi_lo_11 = {dataInMem_hi_232, dataInMem_lo_184, dataInMem_hi_231, dataInMem_lo_183};
  wire [127:0]     dataInMem_hi_hi_hi_11 = {dataInMem_hi_234, dataInMem_lo_186, dataInMem_hi_233, dataInMem_lo_185};
  wire [255:0]     dataInMem_hi_hi_139 = {dataInMem_hi_hi_hi_11, dataInMem_hi_hi_lo_11};
  wire [511:0]     dataInMem_hi_235 = {dataInMem_hi_hi_139, dataInMem_hi_lo_75};
  wire [1023:0]    dataInMem_11 = {dataInMem_hi_235, dataInMem_lo_187};
  wire [255:0]     regroupCacheLine_11_0 = dataInMem_11[255:0];
  wire [255:0]     regroupCacheLine_11_1 = dataInMem_11[511:256];
  wire [255:0]     regroupCacheLine_11_2 = dataInMem_11[767:512];
  wire [255:0]     regroupCacheLine_11_3 = dataInMem_11[1023:768];
  wire [255:0]     res_88 = regroupCacheLine_11_0;
  wire [255:0]     res_89 = regroupCacheLine_11_1;
  wire [255:0]     res_90 = regroupCacheLine_11_2;
  wire [255:0]     res_91 = regroupCacheLine_11_3;
  wire [511:0]     lo_lo_11 = {res_89, res_88};
  wire [511:0]     lo_hi_11 = {res_91, res_90};
  wire [1023:0]    lo_11 = {lo_hi_11, lo_lo_11};
  wire [2047:0]    regroupLoadData_1_3 = {1024'h0, lo_11};
  wire [31:0]      _GEN_212 = {dataRegroupBySew_4_1_0, dataRegroupBySew_3_1_0};
  wire [31:0]      dataInMem_hi_hi_140;
  assign dataInMem_hi_hi_140 = _GEN_212;
  wire [31:0]      dataInMem_hi_lo_78;
  assign dataInMem_hi_lo_78 = _GEN_212;
  wire [47:0]      dataInMem_hi_236 = {dataInMem_hi_hi_140, dataRegroupBySew_2_1_0};
  wire [31:0]      _GEN_213 = {dataRegroupBySew_4_1_1, dataRegroupBySew_3_1_1};
  wire [31:0]      dataInMem_hi_hi_141;
  assign dataInMem_hi_hi_141 = _GEN_213;
  wire [31:0]      dataInMem_hi_lo_79;
  assign dataInMem_hi_lo_79 = _GEN_213;
  wire [47:0]      dataInMem_hi_237 = {dataInMem_hi_hi_141, dataRegroupBySew_2_1_1};
  wire [31:0]      _GEN_214 = {dataRegroupBySew_4_1_2, dataRegroupBySew_3_1_2};
  wire [31:0]      dataInMem_hi_hi_142;
  assign dataInMem_hi_hi_142 = _GEN_214;
  wire [31:0]      dataInMem_hi_lo_80;
  assign dataInMem_hi_lo_80 = _GEN_214;
  wire [47:0]      dataInMem_hi_238 = {dataInMem_hi_hi_142, dataRegroupBySew_2_1_2};
  wire [31:0]      _GEN_215 = {dataRegroupBySew_4_1_3, dataRegroupBySew_3_1_3};
  wire [31:0]      dataInMem_hi_hi_143;
  assign dataInMem_hi_hi_143 = _GEN_215;
  wire [31:0]      dataInMem_hi_lo_81;
  assign dataInMem_hi_lo_81 = _GEN_215;
  wire [47:0]      dataInMem_hi_239 = {dataInMem_hi_hi_143, dataRegroupBySew_2_1_3};
  wire [31:0]      _GEN_216 = {dataRegroupBySew_4_1_4, dataRegroupBySew_3_1_4};
  wire [31:0]      dataInMem_hi_hi_144;
  assign dataInMem_hi_hi_144 = _GEN_216;
  wire [31:0]      dataInMem_hi_lo_82;
  assign dataInMem_hi_lo_82 = _GEN_216;
  wire [47:0]      dataInMem_hi_240 = {dataInMem_hi_hi_144, dataRegroupBySew_2_1_4};
  wire [31:0]      _GEN_217 = {dataRegroupBySew_4_1_5, dataRegroupBySew_3_1_5};
  wire [31:0]      dataInMem_hi_hi_145;
  assign dataInMem_hi_hi_145 = _GEN_217;
  wire [31:0]      dataInMem_hi_lo_83;
  assign dataInMem_hi_lo_83 = _GEN_217;
  wire [47:0]      dataInMem_hi_241 = {dataInMem_hi_hi_145, dataRegroupBySew_2_1_5};
  wire [31:0]      _GEN_218 = {dataRegroupBySew_4_1_6, dataRegroupBySew_3_1_6};
  wire [31:0]      dataInMem_hi_hi_146;
  assign dataInMem_hi_hi_146 = _GEN_218;
  wire [31:0]      dataInMem_hi_lo_84;
  assign dataInMem_hi_lo_84 = _GEN_218;
  wire [47:0]      dataInMem_hi_242 = {dataInMem_hi_hi_146, dataRegroupBySew_2_1_6};
  wire [31:0]      _GEN_219 = {dataRegroupBySew_4_1_7, dataRegroupBySew_3_1_7};
  wire [31:0]      dataInMem_hi_hi_147;
  assign dataInMem_hi_hi_147 = _GEN_219;
  wire [31:0]      dataInMem_hi_lo_85;
  assign dataInMem_hi_lo_85 = _GEN_219;
  wire [47:0]      dataInMem_hi_243 = {dataInMem_hi_hi_147, dataRegroupBySew_2_1_7};
  wire [31:0]      _GEN_220 = {dataRegroupBySew_4_1_8, dataRegroupBySew_3_1_8};
  wire [31:0]      dataInMem_hi_hi_148;
  assign dataInMem_hi_hi_148 = _GEN_220;
  wire [31:0]      dataInMem_hi_lo_86;
  assign dataInMem_hi_lo_86 = _GEN_220;
  wire [47:0]      dataInMem_hi_244 = {dataInMem_hi_hi_148, dataRegroupBySew_2_1_8};
  wire [31:0]      _GEN_221 = {dataRegroupBySew_4_1_9, dataRegroupBySew_3_1_9};
  wire [31:0]      dataInMem_hi_hi_149;
  assign dataInMem_hi_hi_149 = _GEN_221;
  wire [31:0]      dataInMem_hi_lo_87;
  assign dataInMem_hi_lo_87 = _GEN_221;
  wire [47:0]      dataInMem_hi_245 = {dataInMem_hi_hi_149, dataRegroupBySew_2_1_9};
  wire [31:0]      _GEN_222 = {dataRegroupBySew_4_1_10, dataRegroupBySew_3_1_10};
  wire [31:0]      dataInMem_hi_hi_150;
  assign dataInMem_hi_hi_150 = _GEN_222;
  wire [31:0]      dataInMem_hi_lo_88;
  assign dataInMem_hi_lo_88 = _GEN_222;
  wire [47:0]      dataInMem_hi_246 = {dataInMem_hi_hi_150, dataRegroupBySew_2_1_10};
  wire [31:0]      _GEN_223 = {dataRegroupBySew_4_1_11, dataRegroupBySew_3_1_11};
  wire [31:0]      dataInMem_hi_hi_151;
  assign dataInMem_hi_hi_151 = _GEN_223;
  wire [31:0]      dataInMem_hi_lo_89;
  assign dataInMem_hi_lo_89 = _GEN_223;
  wire [47:0]      dataInMem_hi_247 = {dataInMem_hi_hi_151, dataRegroupBySew_2_1_11};
  wire [31:0]      _GEN_224 = {dataRegroupBySew_4_1_12, dataRegroupBySew_3_1_12};
  wire [31:0]      dataInMem_hi_hi_152;
  assign dataInMem_hi_hi_152 = _GEN_224;
  wire [31:0]      dataInMem_hi_lo_90;
  assign dataInMem_hi_lo_90 = _GEN_224;
  wire [47:0]      dataInMem_hi_248 = {dataInMem_hi_hi_152, dataRegroupBySew_2_1_12};
  wire [31:0]      _GEN_225 = {dataRegroupBySew_4_1_13, dataRegroupBySew_3_1_13};
  wire [31:0]      dataInMem_hi_hi_153;
  assign dataInMem_hi_hi_153 = _GEN_225;
  wire [31:0]      dataInMem_hi_lo_91;
  assign dataInMem_hi_lo_91 = _GEN_225;
  wire [47:0]      dataInMem_hi_249 = {dataInMem_hi_hi_153, dataRegroupBySew_2_1_13};
  wire [31:0]      _GEN_226 = {dataRegroupBySew_4_1_14, dataRegroupBySew_3_1_14};
  wire [31:0]      dataInMem_hi_hi_154;
  assign dataInMem_hi_hi_154 = _GEN_226;
  wire [31:0]      dataInMem_hi_lo_92;
  assign dataInMem_hi_lo_92 = _GEN_226;
  wire [47:0]      dataInMem_hi_250 = {dataInMem_hi_hi_154, dataRegroupBySew_2_1_14};
  wire [31:0]      _GEN_227 = {dataRegroupBySew_4_1_15, dataRegroupBySew_3_1_15};
  wire [31:0]      dataInMem_hi_hi_155;
  assign dataInMem_hi_hi_155 = _GEN_227;
  wire [31:0]      dataInMem_hi_lo_93;
  assign dataInMem_hi_lo_93 = _GEN_227;
  wire [47:0]      dataInMem_hi_251 = {dataInMem_hi_hi_155, dataRegroupBySew_2_1_15};
  wire [159:0]     dataInMem_lo_lo_lo_12 = {dataInMem_hi_237, dataInMem_lo_189, dataInMem_hi_236, dataInMem_lo_188};
  wire [159:0]     dataInMem_lo_lo_hi_12 = {dataInMem_hi_239, dataInMem_lo_191, dataInMem_hi_238, dataInMem_lo_190};
  wire [319:0]     dataInMem_lo_lo_44 = {dataInMem_lo_lo_hi_12, dataInMem_lo_lo_lo_12};
  wire [159:0]     dataInMem_lo_hi_lo_12 = {dataInMem_hi_241, dataInMem_lo_193, dataInMem_hi_240, dataInMem_lo_192};
  wire [159:0]     dataInMem_lo_hi_hi_12 = {dataInMem_hi_243, dataInMem_lo_195, dataInMem_hi_242, dataInMem_lo_194};
  wire [319:0]     dataInMem_lo_hi_108 = {dataInMem_lo_hi_hi_12, dataInMem_lo_hi_lo_12};
  wire [639:0]     dataInMem_lo_204 = {dataInMem_lo_hi_108, dataInMem_lo_lo_44};
  wire [159:0]     dataInMem_hi_lo_lo_12 = {dataInMem_hi_245, dataInMem_lo_197, dataInMem_hi_244, dataInMem_lo_196};
  wire [159:0]     dataInMem_hi_lo_hi_12 = {dataInMem_hi_247, dataInMem_lo_199, dataInMem_hi_246, dataInMem_lo_198};
  wire [319:0]     dataInMem_hi_lo_76 = {dataInMem_hi_lo_hi_12, dataInMem_hi_lo_lo_12};
  wire [159:0]     dataInMem_hi_hi_lo_12 = {dataInMem_hi_249, dataInMem_lo_201, dataInMem_hi_248, dataInMem_lo_200};
  wire [159:0]     dataInMem_hi_hi_hi_12 = {dataInMem_hi_251, dataInMem_lo_203, dataInMem_hi_250, dataInMem_lo_202};
  wire [319:0]     dataInMem_hi_hi_156 = {dataInMem_hi_hi_hi_12, dataInMem_hi_hi_lo_12};
  wire [639:0]     dataInMem_hi_252 = {dataInMem_hi_hi_156, dataInMem_hi_lo_76};
  wire [1279:0]    dataInMem_12 = {dataInMem_hi_252, dataInMem_lo_204};
  wire [255:0]     regroupCacheLine_12_0 = dataInMem_12[255:0];
  wire [255:0]     regroupCacheLine_12_1 = dataInMem_12[511:256];
  wire [255:0]     regroupCacheLine_12_2 = dataInMem_12[767:512];
  wire [255:0]     regroupCacheLine_12_3 = dataInMem_12[1023:768];
  wire [255:0]     regroupCacheLine_12_4 = dataInMem_12[1279:1024];
  wire [255:0]     res_96 = regroupCacheLine_12_0;
  wire [255:0]     res_97 = regroupCacheLine_12_1;
  wire [255:0]     res_98 = regroupCacheLine_12_2;
  wire [255:0]     res_99 = regroupCacheLine_12_3;
  wire [255:0]     res_100 = regroupCacheLine_12_4;
  wire [511:0]     lo_lo_12 = {res_97, res_96};
  wire [511:0]     lo_hi_12 = {res_99, res_98};
  wire [1023:0]    lo_12 = {lo_hi_12, lo_lo_12};
  wire [511:0]     hi_lo_12 = {256'h0, res_100};
  wire [1023:0]    hi_12 = {512'h0, hi_lo_12};
  wire [2047:0]    regroupLoadData_1_4 = {hi_12, lo_12};
  wire [47:0]      dataInMem_lo_205 = {dataInMem_lo_hi_109, dataRegroupBySew_0_1_0};
  wire [31:0]      _GEN_228 = {dataRegroupBySew_5_1_0, dataRegroupBySew_4_1_0};
  wire [31:0]      dataInMem_hi_hi_157;
  assign dataInMem_hi_hi_157 = _GEN_228;
  wire [31:0]      dataInMem_hi_lo_95;
  assign dataInMem_hi_lo_95 = _GEN_228;
  wire [47:0]      dataInMem_hi_253 = {dataInMem_hi_hi_157, dataRegroupBySew_3_1_0};
  wire [47:0]      dataInMem_lo_206 = {dataInMem_lo_hi_110, dataRegroupBySew_0_1_1};
  wire [31:0]      _GEN_229 = {dataRegroupBySew_5_1_1, dataRegroupBySew_4_1_1};
  wire [31:0]      dataInMem_hi_hi_158;
  assign dataInMem_hi_hi_158 = _GEN_229;
  wire [31:0]      dataInMem_hi_lo_96;
  assign dataInMem_hi_lo_96 = _GEN_229;
  wire [47:0]      dataInMem_hi_254 = {dataInMem_hi_hi_158, dataRegroupBySew_3_1_1};
  wire [47:0]      dataInMem_lo_207 = {dataInMem_lo_hi_111, dataRegroupBySew_0_1_2};
  wire [31:0]      _GEN_230 = {dataRegroupBySew_5_1_2, dataRegroupBySew_4_1_2};
  wire [31:0]      dataInMem_hi_hi_159;
  assign dataInMem_hi_hi_159 = _GEN_230;
  wire [31:0]      dataInMem_hi_lo_97;
  assign dataInMem_hi_lo_97 = _GEN_230;
  wire [47:0]      dataInMem_hi_255 = {dataInMem_hi_hi_159, dataRegroupBySew_3_1_2};
  wire [47:0]      dataInMem_lo_208 = {dataInMem_lo_hi_112, dataRegroupBySew_0_1_3};
  wire [31:0]      _GEN_231 = {dataRegroupBySew_5_1_3, dataRegroupBySew_4_1_3};
  wire [31:0]      dataInMem_hi_hi_160;
  assign dataInMem_hi_hi_160 = _GEN_231;
  wire [31:0]      dataInMem_hi_lo_98;
  assign dataInMem_hi_lo_98 = _GEN_231;
  wire [47:0]      dataInMem_hi_256 = {dataInMem_hi_hi_160, dataRegroupBySew_3_1_3};
  wire [47:0]      dataInMem_lo_209 = {dataInMem_lo_hi_113, dataRegroupBySew_0_1_4};
  wire [31:0]      _GEN_232 = {dataRegroupBySew_5_1_4, dataRegroupBySew_4_1_4};
  wire [31:0]      dataInMem_hi_hi_161;
  assign dataInMem_hi_hi_161 = _GEN_232;
  wire [31:0]      dataInMem_hi_lo_99;
  assign dataInMem_hi_lo_99 = _GEN_232;
  wire [47:0]      dataInMem_hi_257 = {dataInMem_hi_hi_161, dataRegroupBySew_3_1_4};
  wire [47:0]      dataInMem_lo_210 = {dataInMem_lo_hi_114, dataRegroupBySew_0_1_5};
  wire [31:0]      _GEN_233 = {dataRegroupBySew_5_1_5, dataRegroupBySew_4_1_5};
  wire [31:0]      dataInMem_hi_hi_162;
  assign dataInMem_hi_hi_162 = _GEN_233;
  wire [31:0]      dataInMem_hi_lo_100;
  assign dataInMem_hi_lo_100 = _GEN_233;
  wire [47:0]      dataInMem_hi_258 = {dataInMem_hi_hi_162, dataRegroupBySew_3_1_5};
  wire [47:0]      dataInMem_lo_211 = {dataInMem_lo_hi_115, dataRegroupBySew_0_1_6};
  wire [31:0]      _GEN_234 = {dataRegroupBySew_5_1_6, dataRegroupBySew_4_1_6};
  wire [31:0]      dataInMem_hi_hi_163;
  assign dataInMem_hi_hi_163 = _GEN_234;
  wire [31:0]      dataInMem_hi_lo_101;
  assign dataInMem_hi_lo_101 = _GEN_234;
  wire [47:0]      dataInMem_hi_259 = {dataInMem_hi_hi_163, dataRegroupBySew_3_1_6};
  wire [47:0]      dataInMem_lo_212 = {dataInMem_lo_hi_116, dataRegroupBySew_0_1_7};
  wire [31:0]      _GEN_235 = {dataRegroupBySew_5_1_7, dataRegroupBySew_4_1_7};
  wire [31:0]      dataInMem_hi_hi_164;
  assign dataInMem_hi_hi_164 = _GEN_235;
  wire [31:0]      dataInMem_hi_lo_102;
  assign dataInMem_hi_lo_102 = _GEN_235;
  wire [47:0]      dataInMem_hi_260 = {dataInMem_hi_hi_164, dataRegroupBySew_3_1_7};
  wire [47:0]      dataInMem_lo_213 = {dataInMem_lo_hi_117, dataRegroupBySew_0_1_8};
  wire [31:0]      _GEN_236 = {dataRegroupBySew_5_1_8, dataRegroupBySew_4_1_8};
  wire [31:0]      dataInMem_hi_hi_165;
  assign dataInMem_hi_hi_165 = _GEN_236;
  wire [31:0]      dataInMem_hi_lo_103;
  assign dataInMem_hi_lo_103 = _GEN_236;
  wire [47:0]      dataInMem_hi_261 = {dataInMem_hi_hi_165, dataRegroupBySew_3_1_8};
  wire [47:0]      dataInMem_lo_214 = {dataInMem_lo_hi_118, dataRegroupBySew_0_1_9};
  wire [31:0]      _GEN_237 = {dataRegroupBySew_5_1_9, dataRegroupBySew_4_1_9};
  wire [31:0]      dataInMem_hi_hi_166;
  assign dataInMem_hi_hi_166 = _GEN_237;
  wire [31:0]      dataInMem_hi_lo_104;
  assign dataInMem_hi_lo_104 = _GEN_237;
  wire [47:0]      dataInMem_hi_262 = {dataInMem_hi_hi_166, dataRegroupBySew_3_1_9};
  wire [47:0]      dataInMem_lo_215 = {dataInMem_lo_hi_119, dataRegroupBySew_0_1_10};
  wire [31:0]      _GEN_238 = {dataRegroupBySew_5_1_10, dataRegroupBySew_4_1_10};
  wire [31:0]      dataInMem_hi_hi_167;
  assign dataInMem_hi_hi_167 = _GEN_238;
  wire [31:0]      dataInMem_hi_lo_105;
  assign dataInMem_hi_lo_105 = _GEN_238;
  wire [47:0]      dataInMem_hi_263 = {dataInMem_hi_hi_167, dataRegroupBySew_3_1_10};
  wire [47:0]      dataInMem_lo_216 = {dataInMem_lo_hi_120, dataRegroupBySew_0_1_11};
  wire [31:0]      _GEN_239 = {dataRegroupBySew_5_1_11, dataRegroupBySew_4_1_11};
  wire [31:0]      dataInMem_hi_hi_168;
  assign dataInMem_hi_hi_168 = _GEN_239;
  wire [31:0]      dataInMem_hi_lo_106;
  assign dataInMem_hi_lo_106 = _GEN_239;
  wire [47:0]      dataInMem_hi_264 = {dataInMem_hi_hi_168, dataRegroupBySew_3_1_11};
  wire [47:0]      dataInMem_lo_217 = {dataInMem_lo_hi_121, dataRegroupBySew_0_1_12};
  wire [31:0]      _GEN_240 = {dataRegroupBySew_5_1_12, dataRegroupBySew_4_1_12};
  wire [31:0]      dataInMem_hi_hi_169;
  assign dataInMem_hi_hi_169 = _GEN_240;
  wire [31:0]      dataInMem_hi_lo_107;
  assign dataInMem_hi_lo_107 = _GEN_240;
  wire [47:0]      dataInMem_hi_265 = {dataInMem_hi_hi_169, dataRegroupBySew_3_1_12};
  wire [47:0]      dataInMem_lo_218 = {dataInMem_lo_hi_122, dataRegroupBySew_0_1_13};
  wire [31:0]      _GEN_241 = {dataRegroupBySew_5_1_13, dataRegroupBySew_4_1_13};
  wire [31:0]      dataInMem_hi_hi_170;
  assign dataInMem_hi_hi_170 = _GEN_241;
  wire [31:0]      dataInMem_hi_lo_108;
  assign dataInMem_hi_lo_108 = _GEN_241;
  wire [47:0]      dataInMem_hi_266 = {dataInMem_hi_hi_170, dataRegroupBySew_3_1_13};
  wire [47:0]      dataInMem_lo_219 = {dataInMem_lo_hi_123, dataRegroupBySew_0_1_14};
  wire [31:0]      _GEN_242 = {dataRegroupBySew_5_1_14, dataRegroupBySew_4_1_14};
  wire [31:0]      dataInMem_hi_hi_171;
  assign dataInMem_hi_hi_171 = _GEN_242;
  wire [31:0]      dataInMem_hi_lo_109;
  assign dataInMem_hi_lo_109 = _GEN_242;
  wire [47:0]      dataInMem_hi_267 = {dataInMem_hi_hi_171, dataRegroupBySew_3_1_14};
  wire [47:0]      dataInMem_lo_220 = {dataInMem_lo_hi_124, dataRegroupBySew_0_1_15};
  wire [31:0]      _GEN_243 = {dataRegroupBySew_5_1_15, dataRegroupBySew_4_1_15};
  wire [31:0]      dataInMem_hi_hi_172;
  assign dataInMem_hi_hi_172 = _GEN_243;
  wire [31:0]      dataInMem_hi_lo_110;
  assign dataInMem_hi_lo_110 = _GEN_243;
  wire [47:0]      dataInMem_hi_268 = {dataInMem_hi_hi_172, dataRegroupBySew_3_1_15};
  wire [191:0]     dataInMem_lo_lo_lo_13 = {dataInMem_hi_254, dataInMem_lo_206, dataInMem_hi_253, dataInMem_lo_205};
  wire [191:0]     dataInMem_lo_lo_hi_13 = {dataInMem_hi_256, dataInMem_lo_208, dataInMem_hi_255, dataInMem_lo_207};
  wire [383:0]     dataInMem_lo_lo_45 = {dataInMem_lo_lo_hi_13, dataInMem_lo_lo_lo_13};
  wire [191:0]     dataInMem_lo_hi_lo_13 = {dataInMem_hi_258, dataInMem_lo_210, dataInMem_hi_257, dataInMem_lo_209};
  wire [191:0]     dataInMem_lo_hi_hi_13 = {dataInMem_hi_260, dataInMem_lo_212, dataInMem_hi_259, dataInMem_lo_211};
  wire [383:0]     dataInMem_lo_hi_125 = {dataInMem_lo_hi_hi_13, dataInMem_lo_hi_lo_13};
  wire [767:0]     dataInMem_lo_221 = {dataInMem_lo_hi_125, dataInMem_lo_lo_45};
  wire [191:0]     dataInMem_hi_lo_lo_13 = {dataInMem_hi_262, dataInMem_lo_214, dataInMem_hi_261, dataInMem_lo_213};
  wire [191:0]     dataInMem_hi_lo_hi_13 = {dataInMem_hi_264, dataInMem_lo_216, dataInMem_hi_263, dataInMem_lo_215};
  wire [383:0]     dataInMem_hi_lo_77 = {dataInMem_hi_lo_hi_13, dataInMem_hi_lo_lo_13};
  wire [191:0]     dataInMem_hi_hi_lo_13 = {dataInMem_hi_266, dataInMem_lo_218, dataInMem_hi_265, dataInMem_lo_217};
  wire [191:0]     dataInMem_hi_hi_hi_13 = {dataInMem_hi_268, dataInMem_lo_220, dataInMem_hi_267, dataInMem_lo_219};
  wire [383:0]     dataInMem_hi_hi_173 = {dataInMem_hi_hi_hi_13, dataInMem_hi_hi_lo_13};
  wire [767:0]     dataInMem_hi_269 = {dataInMem_hi_hi_173, dataInMem_hi_lo_77};
  wire [1535:0]    dataInMem_13 = {dataInMem_hi_269, dataInMem_lo_221};
  wire [255:0]     regroupCacheLine_13_0 = dataInMem_13[255:0];
  wire [255:0]     regroupCacheLine_13_1 = dataInMem_13[511:256];
  wire [255:0]     regroupCacheLine_13_2 = dataInMem_13[767:512];
  wire [255:0]     regroupCacheLine_13_3 = dataInMem_13[1023:768];
  wire [255:0]     regroupCacheLine_13_4 = dataInMem_13[1279:1024];
  wire [255:0]     regroupCacheLine_13_5 = dataInMem_13[1535:1280];
  wire [255:0]     res_104 = regroupCacheLine_13_0;
  wire [255:0]     res_105 = regroupCacheLine_13_1;
  wire [255:0]     res_106 = regroupCacheLine_13_2;
  wire [255:0]     res_107 = regroupCacheLine_13_3;
  wire [255:0]     res_108 = regroupCacheLine_13_4;
  wire [255:0]     res_109 = regroupCacheLine_13_5;
  wire [511:0]     lo_lo_13 = {res_105, res_104};
  wire [511:0]     lo_hi_13 = {res_107, res_106};
  wire [1023:0]    lo_13 = {lo_hi_13, lo_lo_13};
  wire [511:0]     hi_lo_13 = {res_109, res_108};
  wire [1023:0]    hi_13 = {512'h0, hi_lo_13};
  wire [2047:0]    regroupLoadData_1_5 = {hi_13, lo_13};
  wire [47:0]      dataInMem_lo_222 = {dataInMem_lo_hi_126, dataRegroupBySew_0_1_0};
  wire [31:0]      dataInMem_hi_hi_174 = {dataRegroupBySew_6_1_0, dataRegroupBySew_5_1_0};
  wire [63:0]      dataInMem_hi_270 = {dataInMem_hi_hi_174, dataInMem_hi_lo_78};
  wire [47:0]      dataInMem_lo_223 = {dataInMem_lo_hi_127, dataRegroupBySew_0_1_1};
  wire [31:0]      dataInMem_hi_hi_175 = {dataRegroupBySew_6_1_1, dataRegroupBySew_5_1_1};
  wire [63:0]      dataInMem_hi_271 = {dataInMem_hi_hi_175, dataInMem_hi_lo_79};
  wire [47:0]      dataInMem_lo_224 = {dataInMem_lo_hi_128, dataRegroupBySew_0_1_2};
  wire [31:0]      dataInMem_hi_hi_176 = {dataRegroupBySew_6_1_2, dataRegroupBySew_5_1_2};
  wire [63:0]      dataInMem_hi_272 = {dataInMem_hi_hi_176, dataInMem_hi_lo_80};
  wire [47:0]      dataInMem_lo_225 = {dataInMem_lo_hi_129, dataRegroupBySew_0_1_3};
  wire [31:0]      dataInMem_hi_hi_177 = {dataRegroupBySew_6_1_3, dataRegroupBySew_5_1_3};
  wire [63:0]      dataInMem_hi_273 = {dataInMem_hi_hi_177, dataInMem_hi_lo_81};
  wire [47:0]      dataInMem_lo_226 = {dataInMem_lo_hi_130, dataRegroupBySew_0_1_4};
  wire [31:0]      dataInMem_hi_hi_178 = {dataRegroupBySew_6_1_4, dataRegroupBySew_5_1_4};
  wire [63:0]      dataInMem_hi_274 = {dataInMem_hi_hi_178, dataInMem_hi_lo_82};
  wire [47:0]      dataInMem_lo_227 = {dataInMem_lo_hi_131, dataRegroupBySew_0_1_5};
  wire [31:0]      dataInMem_hi_hi_179 = {dataRegroupBySew_6_1_5, dataRegroupBySew_5_1_5};
  wire [63:0]      dataInMem_hi_275 = {dataInMem_hi_hi_179, dataInMem_hi_lo_83};
  wire [47:0]      dataInMem_lo_228 = {dataInMem_lo_hi_132, dataRegroupBySew_0_1_6};
  wire [31:0]      dataInMem_hi_hi_180 = {dataRegroupBySew_6_1_6, dataRegroupBySew_5_1_6};
  wire [63:0]      dataInMem_hi_276 = {dataInMem_hi_hi_180, dataInMem_hi_lo_84};
  wire [47:0]      dataInMem_lo_229 = {dataInMem_lo_hi_133, dataRegroupBySew_0_1_7};
  wire [31:0]      dataInMem_hi_hi_181 = {dataRegroupBySew_6_1_7, dataRegroupBySew_5_1_7};
  wire [63:0]      dataInMem_hi_277 = {dataInMem_hi_hi_181, dataInMem_hi_lo_85};
  wire [47:0]      dataInMem_lo_230 = {dataInMem_lo_hi_134, dataRegroupBySew_0_1_8};
  wire [31:0]      dataInMem_hi_hi_182 = {dataRegroupBySew_6_1_8, dataRegroupBySew_5_1_8};
  wire [63:0]      dataInMem_hi_278 = {dataInMem_hi_hi_182, dataInMem_hi_lo_86};
  wire [47:0]      dataInMem_lo_231 = {dataInMem_lo_hi_135, dataRegroupBySew_0_1_9};
  wire [31:0]      dataInMem_hi_hi_183 = {dataRegroupBySew_6_1_9, dataRegroupBySew_5_1_9};
  wire [63:0]      dataInMem_hi_279 = {dataInMem_hi_hi_183, dataInMem_hi_lo_87};
  wire [47:0]      dataInMem_lo_232 = {dataInMem_lo_hi_136, dataRegroupBySew_0_1_10};
  wire [31:0]      dataInMem_hi_hi_184 = {dataRegroupBySew_6_1_10, dataRegroupBySew_5_1_10};
  wire [63:0]      dataInMem_hi_280 = {dataInMem_hi_hi_184, dataInMem_hi_lo_88};
  wire [47:0]      dataInMem_lo_233 = {dataInMem_lo_hi_137, dataRegroupBySew_0_1_11};
  wire [31:0]      dataInMem_hi_hi_185 = {dataRegroupBySew_6_1_11, dataRegroupBySew_5_1_11};
  wire [63:0]      dataInMem_hi_281 = {dataInMem_hi_hi_185, dataInMem_hi_lo_89};
  wire [47:0]      dataInMem_lo_234 = {dataInMem_lo_hi_138, dataRegroupBySew_0_1_12};
  wire [31:0]      dataInMem_hi_hi_186 = {dataRegroupBySew_6_1_12, dataRegroupBySew_5_1_12};
  wire [63:0]      dataInMem_hi_282 = {dataInMem_hi_hi_186, dataInMem_hi_lo_90};
  wire [47:0]      dataInMem_lo_235 = {dataInMem_lo_hi_139, dataRegroupBySew_0_1_13};
  wire [31:0]      dataInMem_hi_hi_187 = {dataRegroupBySew_6_1_13, dataRegroupBySew_5_1_13};
  wire [63:0]      dataInMem_hi_283 = {dataInMem_hi_hi_187, dataInMem_hi_lo_91};
  wire [47:0]      dataInMem_lo_236 = {dataInMem_lo_hi_140, dataRegroupBySew_0_1_14};
  wire [31:0]      dataInMem_hi_hi_188 = {dataRegroupBySew_6_1_14, dataRegroupBySew_5_1_14};
  wire [63:0]      dataInMem_hi_284 = {dataInMem_hi_hi_188, dataInMem_hi_lo_92};
  wire [47:0]      dataInMem_lo_237 = {dataInMem_lo_hi_141, dataRegroupBySew_0_1_15};
  wire [31:0]      dataInMem_hi_hi_189 = {dataRegroupBySew_6_1_15, dataRegroupBySew_5_1_15};
  wire [63:0]      dataInMem_hi_285 = {dataInMem_hi_hi_189, dataInMem_hi_lo_93};
  wire [223:0]     dataInMem_lo_lo_lo_14 = {dataInMem_hi_271, dataInMem_lo_223, dataInMem_hi_270, dataInMem_lo_222};
  wire [223:0]     dataInMem_lo_lo_hi_14 = {dataInMem_hi_273, dataInMem_lo_225, dataInMem_hi_272, dataInMem_lo_224};
  wire [447:0]     dataInMem_lo_lo_46 = {dataInMem_lo_lo_hi_14, dataInMem_lo_lo_lo_14};
  wire [223:0]     dataInMem_lo_hi_lo_14 = {dataInMem_hi_275, dataInMem_lo_227, dataInMem_hi_274, dataInMem_lo_226};
  wire [223:0]     dataInMem_lo_hi_hi_14 = {dataInMem_hi_277, dataInMem_lo_229, dataInMem_hi_276, dataInMem_lo_228};
  wire [447:0]     dataInMem_lo_hi_142 = {dataInMem_lo_hi_hi_14, dataInMem_lo_hi_lo_14};
  wire [895:0]     dataInMem_lo_238 = {dataInMem_lo_hi_142, dataInMem_lo_lo_46};
  wire [223:0]     dataInMem_hi_lo_lo_14 = {dataInMem_hi_279, dataInMem_lo_231, dataInMem_hi_278, dataInMem_lo_230};
  wire [223:0]     dataInMem_hi_lo_hi_14 = {dataInMem_hi_281, dataInMem_lo_233, dataInMem_hi_280, dataInMem_lo_232};
  wire [447:0]     dataInMem_hi_lo_94 = {dataInMem_hi_lo_hi_14, dataInMem_hi_lo_lo_14};
  wire [223:0]     dataInMem_hi_hi_lo_14 = {dataInMem_hi_283, dataInMem_lo_235, dataInMem_hi_282, dataInMem_lo_234};
  wire [223:0]     dataInMem_hi_hi_hi_14 = {dataInMem_hi_285, dataInMem_lo_237, dataInMem_hi_284, dataInMem_lo_236};
  wire [447:0]     dataInMem_hi_hi_190 = {dataInMem_hi_hi_hi_14, dataInMem_hi_hi_lo_14};
  wire [895:0]     dataInMem_hi_286 = {dataInMem_hi_hi_190, dataInMem_hi_lo_94};
  wire [1791:0]    dataInMem_14 = {dataInMem_hi_286, dataInMem_lo_238};
  wire [255:0]     regroupCacheLine_14_0 = dataInMem_14[255:0];
  wire [255:0]     regroupCacheLine_14_1 = dataInMem_14[511:256];
  wire [255:0]     regroupCacheLine_14_2 = dataInMem_14[767:512];
  wire [255:0]     regroupCacheLine_14_3 = dataInMem_14[1023:768];
  wire [255:0]     regroupCacheLine_14_4 = dataInMem_14[1279:1024];
  wire [255:0]     regroupCacheLine_14_5 = dataInMem_14[1535:1280];
  wire [255:0]     regroupCacheLine_14_6 = dataInMem_14[1791:1536];
  wire [255:0]     res_112 = regroupCacheLine_14_0;
  wire [255:0]     res_113 = regroupCacheLine_14_1;
  wire [255:0]     res_114 = regroupCacheLine_14_2;
  wire [255:0]     res_115 = regroupCacheLine_14_3;
  wire [255:0]     res_116 = regroupCacheLine_14_4;
  wire [255:0]     res_117 = regroupCacheLine_14_5;
  wire [255:0]     res_118 = regroupCacheLine_14_6;
  wire [511:0]     lo_lo_14 = {res_113, res_112};
  wire [511:0]     lo_hi_14 = {res_115, res_114};
  wire [1023:0]    lo_14 = {lo_hi_14, lo_lo_14};
  wire [511:0]     hi_lo_14 = {res_117, res_116};
  wire [511:0]     hi_hi_14 = {256'h0, res_118};
  wire [1023:0]    hi_14 = {hi_hi_14, hi_lo_14};
  wire [2047:0]    regroupLoadData_1_6 = {hi_14, lo_14};
  wire [63:0]      dataInMem_lo_239 = {dataInMem_lo_hi_143, dataInMem_lo_lo_47};
  wire [31:0]      dataInMem_hi_hi_191 = {dataRegroupBySew_7_1_0, dataRegroupBySew_6_1_0};
  wire [63:0]      dataInMem_hi_287 = {dataInMem_hi_hi_191, dataInMem_hi_lo_95};
  wire [63:0]      dataInMem_lo_240 = {dataInMem_lo_hi_144, dataInMem_lo_lo_48};
  wire [31:0]      dataInMem_hi_hi_192 = {dataRegroupBySew_7_1_1, dataRegroupBySew_6_1_1};
  wire [63:0]      dataInMem_hi_288 = {dataInMem_hi_hi_192, dataInMem_hi_lo_96};
  wire [63:0]      dataInMem_lo_241 = {dataInMem_lo_hi_145, dataInMem_lo_lo_49};
  wire [31:0]      dataInMem_hi_hi_193 = {dataRegroupBySew_7_1_2, dataRegroupBySew_6_1_2};
  wire [63:0]      dataInMem_hi_289 = {dataInMem_hi_hi_193, dataInMem_hi_lo_97};
  wire [63:0]      dataInMem_lo_242 = {dataInMem_lo_hi_146, dataInMem_lo_lo_50};
  wire [31:0]      dataInMem_hi_hi_194 = {dataRegroupBySew_7_1_3, dataRegroupBySew_6_1_3};
  wire [63:0]      dataInMem_hi_290 = {dataInMem_hi_hi_194, dataInMem_hi_lo_98};
  wire [63:0]      dataInMem_lo_243 = {dataInMem_lo_hi_147, dataInMem_lo_lo_51};
  wire [31:0]      dataInMem_hi_hi_195 = {dataRegroupBySew_7_1_4, dataRegroupBySew_6_1_4};
  wire [63:0]      dataInMem_hi_291 = {dataInMem_hi_hi_195, dataInMem_hi_lo_99};
  wire [63:0]      dataInMem_lo_244 = {dataInMem_lo_hi_148, dataInMem_lo_lo_52};
  wire [31:0]      dataInMem_hi_hi_196 = {dataRegroupBySew_7_1_5, dataRegroupBySew_6_1_5};
  wire [63:0]      dataInMem_hi_292 = {dataInMem_hi_hi_196, dataInMem_hi_lo_100};
  wire [63:0]      dataInMem_lo_245 = {dataInMem_lo_hi_149, dataInMem_lo_lo_53};
  wire [31:0]      dataInMem_hi_hi_197 = {dataRegroupBySew_7_1_6, dataRegroupBySew_6_1_6};
  wire [63:0]      dataInMem_hi_293 = {dataInMem_hi_hi_197, dataInMem_hi_lo_101};
  wire [63:0]      dataInMem_lo_246 = {dataInMem_lo_hi_150, dataInMem_lo_lo_54};
  wire [31:0]      dataInMem_hi_hi_198 = {dataRegroupBySew_7_1_7, dataRegroupBySew_6_1_7};
  wire [63:0]      dataInMem_hi_294 = {dataInMem_hi_hi_198, dataInMem_hi_lo_102};
  wire [63:0]      dataInMem_lo_247 = {dataInMem_lo_hi_151, dataInMem_lo_lo_55};
  wire [31:0]      dataInMem_hi_hi_199 = {dataRegroupBySew_7_1_8, dataRegroupBySew_6_1_8};
  wire [63:0]      dataInMem_hi_295 = {dataInMem_hi_hi_199, dataInMem_hi_lo_103};
  wire [63:0]      dataInMem_lo_248 = {dataInMem_lo_hi_152, dataInMem_lo_lo_56};
  wire [31:0]      dataInMem_hi_hi_200 = {dataRegroupBySew_7_1_9, dataRegroupBySew_6_1_9};
  wire [63:0]      dataInMem_hi_296 = {dataInMem_hi_hi_200, dataInMem_hi_lo_104};
  wire [63:0]      dataInMem_lo_249 = {dataInMem_lo_hi_153, dataInMem_lo_lo_57};
  wire [31:0]      dataInMem_hi_hi_201 = {dataRegroupBySew_7_1_10, dataRegroupBySew_6_1_10};
  wire [63:0]      dataInMem_hi_297 = {dataInMem_hi_hi_201, dataInMem_hi_lo_105};
  wire [63:0]      dataInMem_lo_250 = {dataInMem_lo_hi_154, dataInMem_lo_lo_58};
  wire [31:0]      dataInMem_hi_hi_202 = {dataRegroupBySew_7_1_11, dataRegroupBySew_6_1_11};
  wire [63:0]      dataInMem_hi_298 = {dataInMem_hi_hi_202, dataInMem_hi_lo_106};
  wire [63:0]      dataInMem_lo_251 = {dataInMem_lo_hi_155, dataInMem_lo_lo_59};
  wire [31:0]      dataInMem_hi_hi_203 = {dataRegroupBySew_7_1_12, dataRegroupBySew_6_1_12};
  wire [63:0]      dataInMem_hi_299 = {dataInMem_hi_hi_203, dataInMem_hi_lo_107};
  wire [63:0]      dataInMem_lo_252 = {dataInMem_lo_hi_156, dataInMem_lo_lo_60};
  wire [31:0]      dataInMem_hi_hi_204 = {dataRegroupBySew_7_1_13, dataRegroupBySew_6_1_13};
  wire [63:0]      dataInMem_hi_300 = {dataInMem_hi_hi_204, dataInMem_hi_lo_108};
  wire [63:0]      dataInMem_lo_253 = {dataInMem_lo_hi_157, dataInMem_lo_lo_61};
  wire [31:0]      dataInMem_hi_hi_205 = {dataRegroupBySew_7_1_14, dataRegroupBySew_6_1_14};
  wire [63:0]      dataInMem_hi_301 = {dataInMem_hi_hi_205, dataInMem_hi_lo_109};
  wire [63:0]      dataInMem_lo_254 = {dataInMem_lo_hi_158, dataInMem_lo_lo_62};
  wire [31:0]      dataInMem_hi_hi_206 = {dataRegroupBySew_7_1_15, dataRegroupBySew_6_1_15};
  wire [63:0]      dataInMem_hi_302 = {dataInMem_hi_hi_206, dataInMem_hi_lo_110};
  wire [255:0]     dataInMem_lo_lo_lo_15 = {dataInMem_hi_288, dataInMem_lo_240, dataInMem_hi_287, dataInMem_lo_239};
  wire [255:0]     dataInMem_lo_lo_hi_15 = {dataInMem_hi_290, dataInMem_lo_242, dataInMem_hi_289, dataInMem_lo_241};
  wire [511:0]     dataInMem_lo_lo_63 = {dataInMem_lo_lo_hi_15, dataInMem_lo_lo_lo_15};
  wire [255:0]     dataInMem_lo_hi_lo_15 = {dataInMem_hi_292, dataInMem_lo_244, dataInMem_hi_291, dataInMem_lo_243};
  wire [255:0]     dataInMem_lo_hi_hi_15 = {dataInMem_hi_294, dataInMem_lo_246, dataInMem_hi_293, dataInMem_lo_245};
  wire [511:0]     dataInMem_lo_hi_159 = {dataInMem_lo_hi_hi_15, dataInMem_lo_hi_lo_15};
  wire [1023:0]    dataInMem_lo_255 = {dataInMem_lo_hi_159, dataInMem_lo_lo_63};
  wire [255:0]     dataInMem_hi_lo_lo_15 = {dataInMem_hi_296, dataInMem_lo_248, dataInMem_hi_295, dataInMem_lo_247};
  wire [255:0]     dataInMem_hi_lo_hi_15 = {dataInMem_hi_298, dataInMem_lo_250, dataInMem_hi_297, dataInMem_lo_249};
  wire [511:0]     dataInMem_hi_lo_111 = {dataInMem_hi_lo_hi_15, dataInMem_hi_lo_lo_15};
  wire [255:0]     dataInMem_hi_hi_lo_15 = {dataInMem_hi_300, dataInMem_lo_252, dataInMem_hi_299, dataInMem_lo_251};
  wire [255:0]     dataInMem_hi_hi_hi_15 = {dataInMem_hi_302, dataInMem_lo_254, dataInMem_hi_301, dataInMem_lo_253};
  wire [511:0]     dataInMem_hi_hi_207 = {dataInMem_hi_hi_hi_15, dataInMem_hi_hi_lo_15};
  wire [1023:0]    dataInMem_hi_303 = {dataInMem_hi_hi_207, dataInMem_hi_lo_111};
  wire [2047:0]    dataInMem_15 = {dataInMem_hi_303, dataInMem_lo_255};
  wire [255:0]     regroupCacheLine_15_0 = dataInMem_15[255:0];
  wire [255:0]     regroupCacheLine_15_1 = dataInMem_15[511:256];
  wire [255:0]     regroupCacheLine_15_2 = dataInMem_15[767:512];
  wire [255:0]     regroupCacheLine_15_3 = dataInMem_15[1023:768];
  wire [255:0]     regroupCacheLine_15_4 = dataInMem_15[1279:1024];
  wire [255:0]     regroupCacheLine_15_5 = dataInMem_15[1535:1280];
  wire [255:0]     regroupCacheLine_15_6 = dataInMem_15[1791:1536];
  wire [255:0]     regroupCacheLine_15_7 = dataInMem_15[2047:1792];
  wire [255:0]     res_120 = regroupCacheLine_15_0;
  wire [255:0]     res_121 = regroupCacheLine_15_1;
  wire [255:0]     res_122 = regroupCacheLine_15_2;
  wire [255:0]     res_123 = regroupCacheLine_15_3;
  wire [255:0]     res_124 = regroupCacheLine_15_4;
  wire [255:0]     res_125 = regroupCacheLine_15_5;
  wire [255:0]     res_126 = regroupCacheLine_15_6;
  wire [255:0]     res_127 = regroupCacheLine_15_7;
  wire [511:0]     lo_lo_15 = {res_121, res_120};
  wire [511:0]     lo_hi_15 = {res_123, res_122};
  wire [1023:0]    lo_15 = {lo_hi_15, lo_lo_15};
  wire [511:0]     hi_lo_15 = {res_125, res_124};
  wire [511:0]     hi_hi_15 = {res_127, res_126};
  wire [1023:0]    hi_15 = {hi_hi_15, hi_lo_15};
  wire [2047:0]    regroupLoadData_1_7 = {hi_15, lo_15};
  wire [31:0]      dataRegroupBySew_0_2_0 = bufferStageEnqueueData_0[31:0];
  wire [31:0]      dataRegroupBySew_0_2_1 = bufferStageEnqueueData_0[63:32];
  wire [31:0]      dataRegroupBySew_0_2_2 = bufferStageEnqueueData_0[95:64];
  wire [31:0]      dataRegroupBySew_0_2_3 = bufferStageEnqueueData_0[127:96];
  wire [31:0]      dataRegroupBySew_0_2_4 = bufferStageEnqueueData_0[159:128];
  wire [31:0]      dataRegroupBySew_0_2_5 = bufferStageEnqueueData_0[191:160];
  wire [31:0]      dataRegroupBySew_0_2_6 = bufferStageEnqueueData_0[223:192];
  wire [31:0]      dataRegroupBySew_0_2_7 = bufferStageEnqueueData_0[255:224];
  wire [31:0]      dataRegroupBySew_1_2_0 = bufferStageEnqueueData_1[31:0];
  wire [31:0]      dataRegroupBySew_1_2_1 = bufferStageEnqueueData_1[63:32];
  wire [31:0]      dataRegroupBySew_1_2_2 = bufferStageEnqueueData_1[95:64];
  wire [31:0]      dataRegroupBySew_1_2_3 = bufferStageEnqueueData_1[127:96];
  wire [31:0]      dataRegroupBySew_1_2_4 = bufferStageEnqueueData_1[159:128];
  wire [31:0]      dataRegroupBySew_1_2_5 = bufferStageEnqueueData_1[191:160];
  wire [31:0]      dataRegroupBySew_1_2_6 = bufferStageEnqueueData_1[223:192];
  wire [31:0]      dataRegroupBySew_1_2_7 = bufferStageEnqueueData_1[255:224];
  wire [31:0]      dataRegroupBySew_2_2_0 = bufferStageEnqueueData_2[31:0];
  wire [31:0]      dataRegroupBySew_2_2_1 = bufferStageEnqueueData_2[63:32];
  wire [31:0]      dataRegroupBySew_2_2_2 = bufferStageEnqueueData_2[95:64];
  wire [31:0]      dataRegroupBySew_2_2_3 = bufferStageEnqueueData_2[127:96];
  wire [31:0]      dataRegroupBySew_2_2_4 = bufferStageEnqueueData_2[159:128];
  wire [31:0]      dataRegroupBySew_2_2_5 = bufferStageEnqueueData_2[191:160];
  wire [31:0]      dataRegroupBySew_2_2_6 = bufferStageEnqueueData_2[223:192];
  wire [31:0]      dataRegroupBySew_2_2_7 = bufferStageEnqueueData_2[255:224];
  wire [31:0]      dataRegroupBySew_3_2_0 = bufferStageEnqueueData_3[31:0];
  wire [31:0]      dataRegroupBySew_3_2_1 = bufferStageEnqueueData_3[63:32];
  wire [31:0]      dataRegroupBySew_3_2_2 = bufferStageEnqueueData_3[95:64];
  wire [31:0]      dataRegroupBySew_3_2_3 = bufferStageEnqueueData_3[127:96];
  wire [31:0]      dataRegroupBySew_3_2_4 = bufferStageEnqueueData_3[159:128];
  wire [31:0]      dataRegroupBySew_3_2_5 = bufferStageEnqueueData_3[191:160];
  wire [31:0]      dataRegroupBySew_3_2_6 = bufferStageEnqueueData_3[223:192];
  wire [31:0]      dataRegroupBySew_3_2_7 = bufferStageEnqueueData_3[255:224];
  wire [31:0]      dataRegroupBySew_4_2_0 = bufferStageEnqueueData_4[31:0];
  wire [31:0]      dataRegroupBySew_4_2_1 = bufferStageEnqueueData_4[63:32];
  wire [31:0]      dataRegroupBySew_4_2_2 = bufferStageEnqueueData_4[95:64];
  wire [31:0]      dataRegroupBySew_4_2_3 = bufferStageEnqueueData_4[127:96];
  wire [31:0]      dataRegroupBySew_4_2_4 = bufferStageEnqueueData_4[159:128];
  wire [31:0]      dataRegroupBySew_4_2_5 = bufferStageEnqueueData_4[191:160];
  wire [31:0]      dataRegroupBySew_4_2_6 = bufferStageEnqueueData_4[223:192];
  wire [31:0]      dataRegroupBySew_4_2_7 = bufferStageEnqueueData_4[255:224];
  wire [31:0]      dataRegroupBySew_5_2_0 = bufferStageEnqueueData_5[31:0];
  wire [31:0]      dataRegroupBySew_5_2_1 = bufferStageEnqueueData_5[63:32];
  wire [31:0]      dataRegroupBySew_5_2_2 = bufferStageEnqueueData_5[95:64];
  wire [31:0]      dataRegroupBySew_5_2_3 = bufferStageEnqueueData_5[127:96];
  wire [31:0]      dataRegroupBySew_5_2_4 = bufferStageEnqueueData_5[159:128];
  wire [31:0]      dataRegroupBySew_5_2_5 = bufferStageEnqueueData_5[191:160];
  wire [31:0]      dataRegroupBySew_5_2_6 = bufferStageEnqueueData_5[223:192];
  wire [31:0]      dataRegroupBySew_5_2_7 = bufferStageEnqueueData_5[255:224];
  wire [31:0]      dataRegroupBySew_6_2_0 = bufferStageEnqueueData_6[31:0];
  wire [31:0]      dataRegroupBySew_6_2_1 = bufferStageEnqueueData_6[63:32];
  wire [31:0]      dataRegroupBySew_6_2_2 = bufferStageEnqueueData_6[95:64];
  wire [31:0]      dataRegroupBySew_6_2_3 = bufferStageEnqueueData_6[127:96];
  wire [31:0]      dataRegroupBySew_6_2_4 = bufferStageEnqueueData_6[159:128];
  wire [31:0]      dataRegroupBySew_6_2_5 = bufferStageEnqueueData_6[191:160];
  wire [31:0]      dataRegroupBySew_6_2_6 = bufferStageEnqueueData_6[223:192];
  wire [31:0]      dataRegroupBySew_6_2_7 = bufferStageEnqueueData_6[255:224];
  wire [31:0]      dataRegroupBySew_7_2_0 = bufferStageEnqueueData_7[31:0];
  wire [31:0]      dataRegroupBySew_7_2_1 = bufferStageEnqueueData_7[63:32];
  wire [31:0]      dataRegroupBySew_7_2_2 = bufferStageEnqueueData_7[95:64];
  wire [31:0]      dataRegroupBySew_7_2_3 = bufferStageEnqueueData_7[127:96];
  wire [31:0]      dataRegroupBySew_7_2_4 = bufferStageEnqueueData_7[159:128];
  wire [31:0]      dataRegroupBySew_7_2_5 = bufferStageEnqueueData_7[191:160];
  wire [31:0]      dataRegroupBySew_7_2_6 = bufferStageEnqueueData_7[223:192];
  wire [31:0]      dataRegroupBySew_7_2_7 = bufferStageEnqueueData_7[255:224];
  wire [63:0]      dataInMem_lo_lo_64 = {dataRegroupBySew_0_2_1, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_lo_hi_160 = {dataRegroupBySew_0_2_3, dataRegroupBySew_0_2_2};
  wire [127:0]     dataInMem_lo_256 = {dataInMem_lo_hi_160, dataInMem_lo_lo_64};
  wire [63:0]      dataInMem_hi_lo_112 = {dataRegroupBySew_0_2_5, dataRegroupBySew_0_2_4};
  wire [63:0]      dataInMem_hi_hi_208 = {dataRegroupBySew_0_2_7, dataRegroupBySew_0_2_6};
  wire [127:0]     dataInMem_hi_304 = {dataInMem_hi_hi_208, dataInMem_hi_lo_112};
  wire [255:0]     dataInMem_16 = {dataInMem_hi_304, dataInMem_lo_256};
  wire [255:0]     regroupCacheLine_16_0 = dataInMem_16;
  wire [255:0]     res_128 = regroupCacheLine_16_0;
  wire [511:0]     lo_lo_16 = {256'h0, res_128};
  wire [1023:0]    lo_16 = {512'h0, lo_lo_16};
  wire [2047:0]    regroupLoadData_2_0 = {1024'h0, lo_16};
  wire [127:0]     dataInMem_lo_lo_65 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1, dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [127:0]     dataInMem_lo_hi_161 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3, dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [255:0]     dataInMem_lo_257 = {dataInMem_lo_hi_161, dataInMem_lo_lo_65};
  wire [127:0]     dataInMem_hi_lo_113 = {dataRegroupBySew_1_2_5, dataRegroupBySew_0_2_5, dataRegroupBySew_1_2_4, dataRegroupBySew_0_2_4};
  wire [127:0]     dataInMem_hi_hi_209 = {dataRegroupBySew_1_2_7, dataRegroupBySew_0_2_7, dataRegroupBySew_1_2_6, dataRegroupBySew_0_2_6};
  wire [255:0]     dataInMem_hi_305 = {dataInMem_hi_hi_209, dataInMem_hi_lo_113};
  wire [511:0]     dataInMem_17 = {dataInMem_hi_305, dataInMem_lo_257};
  wire [255:0]     regroupCacheLine_17_0 = dataInMem_17[255:0];
  wire [255:0]     regroupCacheLine_17_1 = dataInMem_17[511:256];
  wire [255:0]     res_136 = regroupCacheLine_17_0;
  wire [255:0]     res_137 = regroupCacheLine_17_1;
  wire [511:0]     lo_lo_17 = {res_137, res_136};
  wire [1023:0]    lo_17 = {512'h0, lo_lo_17};
  wire [2047:0]    regroupLoadData_2_1 = {1024'h0, lo_17};
  wire [63:0]      _GEN_244 = {dataRegroupBySew_2_2_0, dataRegroupBySew_1_2_0};
  wire [63:0]      dataInMem_hi_306;
  assign dataInMem_hi_306 = _GEN_244;
  wire [63:0]      dataInMem_lo_hi_165;
  assign dataInMem_lo_hi_165 = _GEN_244;
  wire [63:0]      dataInMem_lo_hi_174;
  assign dataInMem_lo_hi_174 = _GEN_244;
  wire [63:0]      _GEN_245 = {dataRegroupBySew_2_2_1, dataRegroupBySew_1_2_1};
  wire [63:0]      dataInMem_hi_307;
  assign dataInMem_hi_307 = _GEN_245;
  wire [63:0]      dataInMem_lo_hi_166;
  assign dataInMem_lo_hi_166 = _GEN_245;
  wire [63:0]      dataInMem_lo_hi_175;
  assign dataInMem_lo_hi_175 = _GEN_245;
  wire [63:0]      _GEN_246 = {dataRegroupBySew_2_2_2, dataRegroupBySew_1_2_2};
  wire [63:0]      dataInMem_hi_308;
  assign dataInMem_hi_308 = _GEN_246;
  wire [63:0]      dataInMem_lo_hi_167;
  assign dataInMem_lo_hi_167 = _GEN_246;
  wire [63:0]      dataInMem_lo_hi_176;
  assign dataInMem_lo_hi_176 = _GEN_246;
  wire [63:0]      _GEN_247 = {dataRegroupBySew_2_2_3, dataRegroupBySew_1_2_3};
  wire [63:0]      dataInMem_hi_309;
  assign dataInMem_hi_309 = _GEN_247;
  wire [63:0]      dataInMem_lo_hi_168;
  assign dataInMem_lo_hi_168 = _GEN_247;
  wire [63:0]      dataInMem_lo_hi_177;
  assign dataInMem_lo_hi_177 = _GEN_247;
  wire [63:0]      _GEN_248 = {dataRegroupBySew_2_2_4, dataRegroupBySew_1_2_4};
  wire [63:0]      dataInMem_hi_310;
  assign dataInMem_hi_310 = _GEN_248;
  wire [63:0]      dataInMem_lo_hi_169;
  assign dataInMem_lo_hi_169 = _GEN_248;
  wire [63:0]      dataInMem_lo_hi_178;
  assign dataInMem_lo_hi_178 = _GEN_248;
  wire [63:0]      _GEN_249 = {dataRegroupBySew_2_2_5, dataRegroupBySew_1_2_5};
  wire [63:0]      dataInMem_hi_311;
  assign dataInMem_hi_311 = _GEN_249;
  wire [63:0]      dataInMem_lo_hi_170;
  assign dataInMem_lo_hi_170 = _GEN_249;
  wire [63:0]      dataInMem_lo_hi_179;
  assign dataInMem_lo_hi_179 = _GEN_249;
  wire [63:0]      _GEN_250 = {dataRegroupBySew_2_2_6, dataRegroupBySew_1_2_6};
  wire [63:0]      dataInMem_hi_312;
  assign dataInMem_hi_312 = _GEN_250;
  wire [63:0]      dataInMem_lo_hi_171;
  assign dataInMem_lo_hi_171 = _GEN_250;
  wire [63:0]      dataInMem_lo_hi_180;
  assign dataInMem_lo_hi_180 = _GEN_250;
  wire [63:0]      _GEN_251 = {dataRegroupBySew_2_2_7, dataRegroupBySew_1_2_7};
  wire [63:0]      dataInMem_hi_313;
  assign dataInMem_hi_313 = _GEN_251;
  wire [63:0]      dataInMem_lo_hi_172;
  assign dataInMem_lo_hi_172 = _GEN_251;
  wire [63:0]      dataInMem_lo_hi_181;
  assign dataInMem_lo_hi_181 = _GEN_251;
  wire [191:0]     dataInMem_lo_lo_66 = {dataInMem_hi_307, dataRegroupBySew_0_2_1, dataInMem_hi_306, dataRegroupBySew_0_2_0};
  wire [191:0]     dataInMem_lo_hi_162 = {dataInMem_hi_309, dataRegroupBySew_0_2_3, dataInMem_hi_308, dataRegroupBySew_0_2_2};
  wire [383:0]     dataInMem_lo_258 = {dataInMem_lo_hi_162, dataInMem_lo_lo_66};
  wire [191:0]     dataInMem_hi_lo_114 = {dataInMem_hi_311, dataRegroupBySew_0_2_5, dataInMem_hi_310, dataRegroupBySew_0_2_4};
  wire [191:0]     dataInMem_hi_hi_210 = {dataInMem_hi_313, dataRegroupBySew_0_2_7, dataInMem_hi_312, dataRegroupBySew_0_2_6};
  wire [383:0]     dataInMem_hi_314 = {dataInMem_hi_hi_210, dataInMem_hi_lo_114};
  wire [767:0]     dataInMem_18 = {dataInMem_hi_314, dataInMem_lo_258};
  wire [255:0]     regroupCacheLine_18_0 = dataInMem_18[255:0];
  wire [255:0]     regroupCacheLine_18_1 = dataInMem_18[511:256];
  wire [255:0]     regroupCacheLine_18_2 = dataInMem_18[767:512];
  wire [255:0]     res_144 = regroupCacheLine_18_0;
  wire [255:0]     res_145 = regroupCacheLine_18_1;
  wire [255:0]     res_146 = regroupCacheLine_18_2;
  wire [511:0]     lo_lo_18 = {res_145, res_144};
  wire [511:0]     lo_hi_18 = {256'h0, res_146};
  wire [1023:0]    lo_18 = {lo_hi_18, lo_lo_18};
  wire [2047:0]    regroupLoadData_2_2 = {1024'h0, lo_18};
  wire [63:0]      _GEN_252 = {dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_lo_259;
  assign dataInMem_lo_259 = _GEN_252;
  wire [63:0]      dataInMem_lo_268;
  assign dataInMem_lo_268 = _GEN_252;
  wire [63:0]      dataInMem_lo_lo_71;
  assign dataInMem_lo_lo_71 = _GEN_252;
  wire [63:0]      _GEN_253 = {dataRegroupBySew_3_2_0, dataRegroupBySew_2_2_0};
  wire [63:0]      dataInMem_hi_315;
  assign dataInMem_hi_315 = _GEN_253;
  wire [63:0]      dataInMem_lo_hi_183;
  assign dataInMem_lo_hi_183 = _GEN_253;
  wire [63:0]      _GEN_254 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1};
  wire [63:0]      dataInMem_lo_260;
  assign dataInMem_lo_260 = _GEN_254;
  wire [63:0]      dataInMem_lo_269;
  assign dataInMem_lo_269 = _GEN_254;
  wire [63:0]      dataInMem_lo_lo_72;
  assign dataInMem_lo_lo_72 = _GEN_254;
  wire [63:0]      _GEN_255 = {dataRegroupBySew_3_2_1, dataRegroupBySew_2_2_1};
  wire [63:0]      dataInMem_hi_316;
  assign dataInMem_hi_316 = _GEN_255;
  wire [63:0]      dataInMem_lo_hi_184;
  assign dataInMem_lo_hi_184 = _GEN_255;
  wire [63:0]      _GEN_256 = {dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [63:0]      dataInMem_lo_261;
  assign dataInMem_lo_261 = _GEN_256;
  wire [63:0]      dataInMem_lo_270;
  assign dataInMem_lo_270 = _GEN_256;
  wire [63:0]      dataInMem_lo_lo_73;
  assign dataInMem_lo_lo_73 = _GEN_256;
  wire [63:0]      _GEN_257 = {dataRegroupBySew_3_2_2, dataRegroupBySew_2_2_2};
  wire [63:0]      dataInMem_hi_317;
  assign dataInMem_hi_317 = _GEN_257;
  wire [63:0]      dataInMem_lo_hi_185;
  assign dataInMem_lo_hi_185 = _GEN_257;
  wire [63:0]      _GEN_258 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3};
  wire [63:0]      dataInMem_lo_262;
  assign dataInMem_lo_262 = _GEN_258;
  wire [63:0]      dataInMem_lo_271;
  assign dataInMem_lo_271 = _GEN_258;
  wire [63:0]      dataInMem_lo_lo_74;
  assign dataInMem_lo_lo_74 = _GEN_258;
  wire [63:0]      _GEN_259 = {dataRegroupBySew_3_2_3, dataRegroupBySew_2_2_3};
  wire [63:0]      dataInMem_hi_318;
  assign dataInMem_hi_318 = _GEN_259;
  wire [63:0]      dataInMem_lo_hi_186;
  assign dataInMem_lo_hi_186 = _GEN_259;
  wire [63:0]      _GEN_260 = {dataRegroupBySew_1_2_4, dataRegroupBySew_0_2_4};
  wire [63:0]      dataInMem_lo_263;
  assign dataInMem_lo_263 = _GEN_260;
  wire [63:0]      dataInMem_lo_272;
  assign dataInMem_lo_272 = _GEN_260;
  wire [63:0]      dataInMem_lo_lo_75;
  assign dataInMem_lo_lo_75 = _GEN_260;
  wire [63:0]      _GEN_261 = {dataRegroupBySew_3_2_4, dataRegroupBySew_2_2_4};
  wire [63:0]      dataInMem_hi_319;
  assign dataInMem_hi_319 = _GEN_261;
  wire [63:0]      dataInMem_lo_hi_187;
  assign dataInMem_lo_hi_187 = _GEN_261;
  wire [63:0]      _GEN_262 = {dataRegroupBySew_1_2_5, dataRegroupBySew_0_2_5};
  wire [63:0]      dataInMem_lo_264;
  assign dataInMem_lo_264 = _GEN_262;
  wire [63:0]      dataInMem_lo_273;
  assign dataInMem_lo_273 = _GEN_262;
  wire [63:0]      dataInMem_lo_lo_76;
  assign dataInMem_lo_lo_76 = _GEN_262;
  wire [63:0]      _GEN_263 = {dataRegroupBySew_3_2_5, dataRegroupBySew_2_2_5};
  wire [63:0]      dataInMem_hi_320;
  assign dataInMem_hi_320 = _GEN_263;
  wire [63:0]      dataInMem_lo_hi_188;
  assign dataInMem_lo_hi_188 = _GEN_263;
  wire [63:0]      _GEN_264 = {dataRegroupBySew_1_2_6, dataRegroupBySew_0_2_6};
  wire [63:0]      dataInMem_lo_265;
  assign dataInMem_lo_265 = _GEN_264;
  wire [63:0]      dataInMem_lo_274;
  assign dataInMem_lo_274 = _GEN_264;
  wire [63:0]      dataInMem_lo_lo_77;
  assign dataInMem_lo_lo_77 = _GEN_264;
  wire [63:0]      _GEN_265 = {dataRegroupBySew_3_2_6, dataRegroupBySew_2_2_6};
  wire [63:0]      dataInMem_hi_321;
  assign dataInMem_hi_321 = _GEN_265;
  wire [63:0]      dataInMem_lo_hi_189;
  assign dataInMem_lo_hi_189 = _GEN_265;
  wire [63:0]      _GEN_266 = {dataRegroupBySew_1_2_7, dataRegroupBySew_0_2_7};
  wire [63:0]      dataInMem_lo_266;
  assign dataInMem_lo_266 = _GEN_266;
  wire [63:0]      dataInMem_lo_275;
  assign dataInMem_lo_275 = _GEN_266;
  wire [63:0]      dataInMem_lo_lo_78;
  assign dataInMem_lo_lo_78 = _GEN_266;
  wire [63:0]      _GEN_267 = {dataRegroupBySew_3_2_7, dataRegroupBySew_2_2_7};
  wire [63:0]      dataInMem_hi_322;
  assign dataInMem_hi_322 = _GEN_267;
  wire [63:0]      dataInMem_lo_hi_190;
  assign dataInMem_lo_hi_190 = _GEN_267;
  wire [255:0]     dataInMem_lo_lo_67 = {dataInMem_hi_316, dataInMem_lo_260, dataInMem_hi_315, dataInMem_lo_259};
  wire [255:0]     dataInMem_lo_hi_163 = {dataInMem_hi_318, dataInMem_lo_262, dataInMem_hi_317, dataInMem_lo_261};
  wire [511:0]     dataInMem_lo_267 = {dataInMem_lo_hi_163, dataInMem_lo_lo_67};
  wire [255:0]     dataInMem_hi_lo_115 = {dataInMem_hi_320, dataInMem_lo_264, dataInMem_hi_319, dataInMem_lo_263};
  wire [255:0]     dataInMem_hi_hi_211 = {dataInMem_hi_322, dataInMem_lo_266, dataInMem_hi_321, dataInMem_lo_265};
  wire [511:0]     dataInMem_hi_323 = {dataInMem_hi_hi_211, dataInMem_hi_lo_115};
  wire [1023:0]    dataInMem_19 = {dataInMem_hi_323, dataInMem_lo_267};
  wire [255:0]     regroupCacheLine_19_0 = dataInMem_19[255:0];
  wire [255:0]     regroupCacheLine_19_1 = dataInMem_19[511:256];
  wire [255:0]     regroupCacheLine_19_2 = dataInMem_19[767:512];
  wire [255:0]     regroupCacheLine_19_3 = dataInMem_19[1023:768];
  wire [255:0]     res_152 = regroupCacheLine_19_0;
  wire [255:0]     res_153 = regroupCacheLine_19_1;
  wire [255:0]     res_154 = regroupCacheLine_19_2;
  wire [255:0]     res_155 = regroupCacheLine_19_3;
  wire [511:0]     lo_lo_19 = {res_153, res_152};
  wire [511:0]     lo_hi_19 = {res_155, res_154};
  wire [1023:0]    lo_19 = {lo_hi_19, lo_lo_19};
  wire [2047:0]    regroupLoadData_2_3 = {1024'h0, lo_19};
  wire [63:0]      _GEN_268 = {dataRegroupBySew_4_2_0, dataRegroupBySew_3_2_0};
  wire [63:0]      dataInMem_hi_hi_212;
  assign dataInMem_hi_hi_212 = _GEN_268;
  wire [63:0]      dataInMem_hi_lo_118;
  assign dataInMem_hi_lo_118 = _GEN_268;
  wire [95:0]      dataInMem_hi_324 = {dataInMem_hi_hi_212, dataRegroupBySew_2_2_0};
  wire [63:0]      _GEN_269 = {dataRegroupBySew_4_2_1, dataRegroupBySew_3_2_1};
  wire [63:0]      dataInMem_hi_hi_213;
  assign dataInMem_hi_hi_213 = _GEN_269;
  wire [63:0]      dataInMem_hi_lo_119;
  assign dataInMem_hi_lo_119 = _GEN_269;
  wire [95:0]      dataInMem_hi_325 = {dataInMem_hi_hi_213, dataRegroupBySew_2_2_1};
  wire [63:0]      _GEN_270 = {dataRegroupBySew_4_2_2, dataRegroupBySew_3_2_2};
  wire [63:0]      dataInMem_hi_hi_214;
  assign dataInMem_hi_hi_214 = _GEN_270;
  wire [63:0]      dataInMem_hi_lo_120;
  assign dataInMem_hi_lo_120 = _GEN_270;
  wire [95:0]      dataInMem_hi_326 = {dataInMem_hi_hi_214, dataRegroupBySew_2_2_2};
  wire [63:0]      _GEN_271 = {dataRegroupBySew_4_2_3, dataRegroupBySew_3_2_3};
  wire [63:0]      dataInMem_hi_hi_215;
  assign dataInMem_hi_hi_215 = _GEN_271;
  wire [63:0]      dataInMem_hi_lo_121;
  assign dataInMem_hi_lo_121 = _GEN_271;
  wire [95:0]      dataInMem_hi_327 = {dataInMem_hi_hi_215, dataRegroupBySew_2_2_3};
  wire [63:0]      _GEN_272 = {dataRegroupBySew_4_2_4, dataRegroupBySew_3_2_4};
  wire [63:0]      dataInMem_hi_hi_216;
  assign dataInMem_hi_hi_216 = _GEN_272;
  wire [63:0]      dataInMem_hi_lo_122;
  assign dataInMem_hi_lo_122 = _GEN_272;
  wire [95:0]      dataInMem_hi_328 = {dataInMem_hi_hi_216, dataRegroupBySew_2_2_4};
  wire [63:0]      _GEN_273 = {dataRegroupBySew_4_2_5, dataRegroupBySew_3_2_5};
  wire [63:0]      dataInMem_hi_hi_217;
  assign dataInMem_hi_hi_217 = _GEN_273;
  wire [63:0]      dataInMem_hi_lo_123;
  assign dataInMem_hi_lo_123 = _GEN_273;
  wire [95:0]      dataInMem_hi_329 = {dataInMem_hi_hi_217, dataRegroupBySew_2_2_5};
  wire [63:0]      _GEN_274 = {dataRegroupBySew_4_2_6, dataRegroupBySew_3_2_6};
  wire [63:0]      dataInMem_hi_hi_218;
  assign dataInMem_hi_hi_218 = _GEN_274;
  wire [63:0]      dataInMem_hi_lo_124;
  assign dataInMem_hi_lo_124 = _GEN_274;
  wire [95:0]      dataInMem_hi_330 = {dataInMem_hi_hi_218, dataRegroupBySew_2_2_6};
  wire [63:0]      _GEN_275 = {dataRegroupBySew_4_2_7, dataRegroupBySew_3_2_7};
  wire [63:0]      dataInMem_hi_hi_219;
  assign dataInMem_hi_hi_219 = _GEN_275;
  wire [63:0]      dataInMem_hi_lo_125;
  assign dataInMem_hi_lo_125 = _GEN_275;
  wire [95:0]      dataInMem_hi_331 = {dataInMem_hi_hi_219, dataRegroupBySew_2_2_7};
  wire [319:0]     dataInMem_lo_lo_68 = {dataInMem_hi_325, dataInMem_lo_269, dataInMem_hi_324, dataInMem_lo_268};
  wire [319:0]     dataInMem_lo_hi_164 = {dataInMem_hi_327, dataInMem_lo_271, dataInMem_hi_326, dataInMem_lo_270};
  wire [639:0]     dataInMem_lo_276 = {dataInMem_lo_hi_164, dataInMem_lo_lo_68};
  wire [319:0]     dataInMem_hi_lo_116 = {dataInMem_hi_329, dataInMem_lo_273, dataInMem_hi_328, dataInMem_lo_272};
  wire [319:0]     dataInMem_hi_hi_220 = {dataInMem_hi_331, dataInMem_lo_275, dataInMem_hi_330, dataInMem_lo_274};
  wire [639:0]     dataInMem_hi_332 = {dataInMem_hi_hi_220, dataInMem_hi_lo_116};
  wire [1279:0]    dataInMem_20 = {dataInMem_hi_332, dataInMem_lo_276};
  wire [255:0]     regroupCacheLine_20_0 = dataInMem_20[255:0];
  wire [255:0]     regroupCacheLine_20_1 = dataInMem_20[511:256];
  wire [255:0]     regroupCacheLine_20_2 = dataInMem_20[767:512];
  wire [255:0]     regroupCacheLine_20_3 = dataInMem_20[1023:768];
  wire [255:0]     regroupCacheLine_20_4 = dataInMem_20[1279:1024];
  wire [255:0]     res_160 = regroupCacheLine_20_0;
  wire [255:0]     res_161 = regroupCacheLine_20_1;
  wire [255:0]     res_162 = regroupCacheLine_20_2;
  wire [255:0]     res_163 = regroupCacheLine_20_3;
  wire [255:0]     res_164 = regroupCacheLine_20_4;
  wire [511:0]     lo_lo_20 = {res_161, res_160};
  wire [511:0]     lo_hi_20 = {res_163, res_162};
  wire [1023:0]    lo_20 = {lo_hi_20, lo_lo_20};
  wire [511:0]     hi_lo_20 = {256'h0, res_164};
  wire [1023:0]    hi_20 = {512'h0, hi_lo_20};
  wire [2047:0]    regroupLoadData_2_4 = {hi_20, lo_20};
  wire [95:0]      dataInMem_lo_277 = {dataInMem_lo_hi_165, dataRegroupBySew_0_2_0};
  wire [63:0]      _GEN_276 = {dataRegroupBySew_5_2_0, dataRegroupBySew_4_2_0};
  wire [63:0]      dataInMem_hi_hi_221;
  assign dataInMem_hi_hi_221 = _GEN_276;
  wire [63:0]      dataInMem_hi_lo_127;
  assign dataInMem_hi_lo_127 = _GEN_276;
  wire [95:0]      dataInMem_hi_333 = {dataInMem_hi_hi_221, dataRegroupBySew_3_2_0};
  wire [95:0]      dataInMem_lo_278 = {dataInMem_lo_hi_166, dataRegroupBySew_0_2_1};
  wire [63:0]      _GEN_277 = {dataRegroupBySew_5_2_1, dataRegroupBySew_4_2_1};
  wire [63:0]      dataInMem_hi_hi_222;
  assign dataInMem_hi_hi_222 = _GEN_277;
  wire [63:0]      dataInMem_hi_lo_128;
  assign dataInMem_hi_lo_128 = _GEN_277;
  wire [95:0]      dataInMem_hi_334 = {dataInMem_hi_hi_222, dataRegroupBySew_3_2_1};
  wire [95:0]      dataInMem_lo_279 = {dataInMem_lo_hi_167, dataRegroupBySew_0_2_2};
  wire [63:0]      _GEN_278 = {dataRegroupBySew_5_2_2, dataRegroupBySew_4_2_2};
  wire [63:0]      dataInMem_hi_hi_223;
  assign dataInMem_hi_hi_223 = _GEN_278;
  wire [63:0]      dataInMem_hi_lo_129;
  assign dataInMem_hi_lo_129 = _GEN_278;
  wire [95:0]      dataInMem_hi_335 = {dataInMem_hi_hi_223, dataRegroupBySew_3_2_2};
  wire [95:0]      dataInMem_lo_280 = {dataInMem_lo_hi_168, dataRegroupBySew_0_2_3};
  wire [63:0]      _GEN_279 = {dataRegroupBySew_5_2_3, dataRegroupBySew_4_2_3};
  wire [63:0]      dataInMem_hi_hi_224;
  assign dataInMem_hi_hi_224 = _GEN_279;
  wire [63:0]      dataInMem_hi_lo_130;
  assign dataInMem_hi_lo_130 = _GEN_279;
  wire [95:0]      dataInMem_hi_336 = {dataInMem_hi_hi_224, dataRegroupBySew_3_2_3};
  wire [95:0]      dataInMem_lo_281 = {dataInMem_lo_hi_169, dataRegroupBySew_0_2_4};
  wire [63:0]      _GEN_280 = {dataRegroupBySew_5_2_4, dataRegroupBySew_4_2_4};
  wire [63:0]      dataInMem_hi_hi_225;
  assign dataInMem_hi_hi_225 = _GEN_280;
  wire [63:0]      dataInMem_hi_lo_131;
  assign dataInMem_hi_lo_131 = _GEN_280;
  wire [95:0]      dataInMem_hi_337 = {dataInMem_hi_hi_225, dataRegroupBySew_3_2_4};
  wire [95:0]      dataInMem_lo_282 = {dataInMem_lo_hi_170, dataRegroupBySew_0_2_5};
  wire [63:0]      _GEN_281 = {dataRegroupBySew_5_2_5, dataRegroupBySew_4_2_5};
  wire [63:0]      dataInMem_hi_hi_226;
  assign dataInMem_hi_hi_226 = _GEN_281;
  wire [63:0]      dataInMem_hi_lo_132;
  assign dataInMem_hi_lo_132 = _GEN_281;
  wire [95:0]      dataInMem_hi_338 = {dataInMem_hi_hi_226, dataRegroupBySew_3_2_5};
  wire [95:0]      dataInMem_lo_283 = {dataInMem_lo_hi_171, dataRegroupBySew_0_2_6};
  wire [63:0]      _GEN_282 = {dataRegroupBySew_5_2_6, dataRegroupBySew_4_2_6};
  wire [63:0]      dataInMem_hi_hi_227;
  assign dataInMem_hi_hi_227 = _GEN_282;
  wire [63:0]      dataInMem_hi_lo_133;
  assign dataInMem_hi_lo_133 = _GEN_282;
  wire [95:0]      dataInMem_hi_339 = {dataInMem_hi_hi_227, dataRegroupBySew_3_2_6};
  wire [95:0]      dataInMem_lo_284 = {dataInMem_lo_hi_172, dataRegroupBySew_0_2_7};
  wire [63:0]      _GEN_283 = {dataRegroupBySew_5_2_7, dataRegroupBySew_4_2_7};
  wire [63:0]      dataInMem_hi_hi_228;
  assign dataInMem_hi_hi_228 = _GEN_283;
  wire [63:0]      dataInMem_hi_lo_134;
  assign dataInMem_hi_lo_134 = _GEN_283;
  wire [95:0]      dataInMem_hi_340 = {dataInMem_hi_hi_228, dataRegroupBySew_3_2_7};
  wire [383:0]     dataInMem_lo_lo_69 = {dataInMem_hi_334, dataInMem_lo_278, dataInMem_hi_333, dataInMem_lo_277};
  wire [383:0]     dataInMem_lo_hi_173 = {dataInMem_hi_336, dataInMem_lo_280, dataInMem_hi_335, dataInMem_lo_279};
  wire [767:0]     dataInMem_lo_285 = {dataInMem_lo_hi_173, dataInMem_lo_lo_69};
  wire [383:0]     dataInMem_hi_lo_117 = {dataInMem_hi_338, dataInMem_lo_282, dataInMem_hi_337, dataInMem_lo_281};
  wire [383:0]     dataInMem_hi_hi_229 = {dataInMem_hi_340, dataInMem_lo_284, dataInMem_hi_339, dataInMem_lo_283};
  wire [767:0]     dataInMem_hi_341 = {dataInMem_hi_hi_229, dataInMem_hi_lo_117};
  wire [1535:0]    dataInMem_21 = {dataInMem_hi_341, dataInMem_lo_285};
  wire [255:0]     regroupCacheLine_21_0 = dataInMem_21[255:0];
  wire [255:0]     regroupCacheLine_21_1 = dataInMem_21[511:256];
  wire [255:0]     regroupCacheLine_21_2 = dataInMem_21[767:512];
  wire [255:0]     regroupCacheLine_21_3 = dataInMem_21[1023:768];
  wire [255:0]     regroupCacheLine_21_4 = dataInMem_21[1279:1024];
  wire [255:0]     regroupCacheLine_21_5 = dataInMem_21[1535:1280];
  wire [255:0]     res_168 = regroupCacheLine_21_0;
  wire [255:0]     res_169 = regroupCacheLine_21_1;
  wire [255:0]     res_170 = regroupCacheLine_21_2;
  wire [255:0]     res_171 = regroupCacheLine_21_3;
  wire [255:0]     res_172 = regroupCacheLine_21_4;
  wire [255:0]     res_173 = regroupCacheLine_21_5;
  wire [511:0]     lo_lo_21 = {res_169, res_168};
  wire [511:0]     lo_hi_21 = {res_171, res_170};
  wire [1023:0]    lo_21 = {lo_hi_21, lo_lo_21};
  wire [511:0]     hi_lo_21 = {res_173, res_172};
  wire [1023:0]    hi_21 = {512'h0, hi_lo_21};
  wire [2047:0]    regroupLoadData_2_5 = {hi_21, lo_21};
  wire [95:0]      dataInMem_lo_286 = {dataInMem_lo_hi_174, dataRegroupBySew_0_2_0};
  wire [63:0]      dataInMem_hi_hi_230 = {dataRegroupBySew_6_2_0, dataRegroupBySew_5_2_0};
  wire [127:0]     dataInMem_hi_342 = {dataInMem_hi_hi_230, dataInMem_hi_lo_118};
  wire [95:0]      dataInMem_lo_287 = {dataInMem_lo_hi_175, dataRegroupBySew_0_2_1};
  wire [63:0]      dataInMem_hi_hi_231 = {dataRegroupBySew_6_2_1, dataRegroupBySew_5_2_1};
  wire [127:0]     dataInMem_hi_343 = {dataInMem_hi_hi_231, dataInMem_hi_lo_119};
  wire [95:0]      dataInMem_lo_288 = {dataInMem_lo_hi_176, dataRegroupBySew_0_2_2};
  wire [63:0]      dataInMem_hi_hi_232 = {dataRegroupBySew_6_2_2, dataRegroupBySew_5_2_2};
  wire [127:0]     dataInMem_hi_344 = {dataInMem_hi_hi_232, dataInMem_hi_lo_120};
  wire [95:0]      dataInMem_lo_289 = {dataInMem_lo_hi_177, dataRegroupBySew_0_2_3};
  wire [63:0]      dataInMem_hi_hi_233 = {dataRegroupBySew_6_2_3, dataRegroupBySew_5_2_3};
  wire [127:0]     dataInMem_hi_345 = {dataInMem_hi_hi_233, dataInMem_hi_lo_121};
  wire [95:0]      dataInMem_lo_290 = {dataInMem_lo_hi_178, dataRegroupBySew_0_2_4};
  wire [63:0]      dataInMem_hi_hi_234 = {dataRegroupBySew_6_2_4, dataRegroupBySew_5_2_4};
  wire [127:0]     dataInMem_hi_346 = {dataInMem_hi_hi_234, dataInMem_hi_lo_122};
  wire [95:0]      dataInMem_lo_291 = {dataInMem_lo_hi_179, dataRegroupBySew_0_2_5};
  wire [63:0]      dataInMem_hi_hi_235 = {dataRegroupBySew_6_2_5, dataRegroupBySew_5_2_5};
  wire [127:0]     dataInMem_hi_347 = {dataInMem_hi_hi_235, dataInMem_hi_lo_123};
  wire [95:0]      dataInMem_lo_292 = {dataInMem_lo_hi_180, dataRegroupBySew_0_2_6};
  wire [63:0]      dataInMem_hi_hi_236 = {dataRegroupBySew_6_2_6, dataRegroupBySew_5_2_6};
  wire [127:0]     dataInMem_hi_348 = {dataInMem_hi_hi_236, dataInMem_hi_lo_124};
  wire [95:0]      dataInMem_lo_293 = {dataInMem_lo_hi_181, dataRegroupBySew_0_2_7};
  wire [63:0]      dataInMem_hi_hi_237 = {dataRegroupBySew_6_2_7, dataRegroupBySew_5_2_7};
  wire [127:0]     dataInMem_hi_349 = {dataInMem_hi_hi_237, dataInMem_hi_lo_125};
  wire [447:0]     dataInMem_lo_lo_70 = {dataInMem_hi_343, dataInMem_lo_287, dataInMem_hi_342, dataInMem_lo_286};
  wire [447:0]     dataInMem_lo_hi_182 = {dataInMem_hi_345, dataInMem_lo_289, dataInMem_hi_344, dataInMem_lo_288};
  wire [895:0]     dataInMem_lo_294 = {dataInMem_lo_hi_182, dataInMem_lo_lo_70};
  wire [447:0]     dataInMem_hi_lo_126 = {dataInMem_hi_347, dataInMem_lo_291, dataInMem_hi_346, dataInMem_lo_290};
  wire [447:0]     dataInMem_hi_hi_238 = {dataInMem_hi_349, dataInMem_lo_293, dataInMem_hi_348, dataInMem_lo_292};
  wire [895:0]     dataInMem_hi_350 = {dataInMem_hi_hi_238, dataInMem_hi_lo_126};
  wire [1791:0]    dataInMem_22 = {dataInMem_hi_350, dataInMem_lo_294};
  wire [255:0]     regroupCacheLine_22_0 = dataInMem_22[255:0];
  wire [255:0]     regroupCacheLine_22_1 = dataInMem_22[511:256];
  wire [255:0]     regroupCacheLine_22_2 = dataInMem_22[767:512];
  wire [255:0]     regroupCacheLine_22_3 = dataInMem_22[1023:768];
  wire [255:0]     regroupCacheLine_22_4 = dataInMem_22[1279:1024];
  wire [255:0]     regroupCacheLine_22_5 = dataInMem_22[1535:1280];
  wire [255:0]     regroupCacheLine_22_6 = dataInMem_22[1791:1536];
  wire [255:0]     res_176 = regroupCacheLine_22_0;
  wire [255:0]     res_177 = regroupCacheLine_22_1;
  wire [255:0]     res_178 = regroupCacheLine_22_2;
  wire [255:0]     res_179 = regroupCacheLine_22_3;
  wire [255:0]     res_180 = regroupCacheLine_22_4;
  wire [255:0]     res_181 = regroupCacheLine_22_5;
  wire [255:0]     res_182 = regroupCacheLine_22_6;
  wire [511:0]     lo_lo_22 = {res_177, res_176};
  wire [511:0]     lo_hi_22 = {res_179, res_178};
  wire [1023:0]    lo_22 = {lo_hi_22, lo_lo_22};
  wire [511:0]     hi_lo_22 = {res_181, res_180};
  wire [511:0]     hi_hi_22 = {256'h0, res_182};
  wire [1023:0]    hi_22 = {hi_hi_22, hi_lo_22};
  wire [2047:0]    regroupLoadData_2_6 = {hi_22, lo_22};
  wire [127:0]     dataInMem_lo_295 = {dataInMem_lo_hi_183, dataInMem_lo_lo_71};
  wire [63:0]      dataInMem_hi_hi_239 = {dataRegroupBySew_7_2_0, dataRegroupBySew_6_2_0};
  wire [127:0]     dataInMem_hi_351 = {dataInMem_hi_hi_239, dataInMem_hi_lo_127};
  wire [127:0]     dataInMem_lo_296 = {dataInMem_lo_hi_184, dataInMem_lo_lo_72};
  wire [63:0]      dataInMem_hi_hi_240 = {dataRegroupBySew_7_2_1, dataRegroupBySew_6_2_1};
  wire [127:0]     dataInMem_hi_352 = {dataInMem_hi_hi_240, dataInMem_hi_lo_128};
  wire [127:0]     dataInMem_lo_297 = {dataInMem_lo_hi_185, dataInMem_lo_lo_73};
  wire [63:0]      dataInMem_hi_hi_241 = {dataRegroupBySew_7_2_2, dataRegroupBySew_6_2_2};
  wire [127:0]     dataInMem_hi_353 = {dataInMem_hi_hi_241, dataInMem_hi_lo_129};
  wire [127:0]     dataInMem_lo_298 = {dataInMem_lo_hi_186, dataInMem_lo_lo_74};
  wire [63:0]      dataInMem_hi_hi_242 = {dataRegroupBySew_7_2_3, dataRegroupBySew_6_2_3};
  wire [127:0]     dataInMem_hi_354 = {dataInMem_hi_hi_242, dataInMem_hi_lo_130};
  wire [127:0]     dataInMem_lo_299 = {dataInMem_lo_hi_187, dataInMem_lo_lo_75};
  wire [63:0]      dataInMem_hi_hi_243 = {dataRegroupBySew_7_2_4, dataRegroupBySew_6_2_4};
  wire [127:0]     dataInMem_hi_355 = {dataInMem_hi_hi_243, dataInMem_hi_lo_131};
  wire [127:0]     dataInMem_lo_300 = {dataInMem_lo_hi_188, dataInMem_lo_lo_76};
  wire [63:0]      dataInMem_hi_hi_244 = {dataRegroupBySew_7_2_5, dataRegroupBySew_6_2_5};
  wire [127:0]     dataInMem_hi_356 = {dataInMem_hi_hi_244, dataInMem_hi_lo_132};
  wire [127:0]     dataInMem_lo_301 = {dataInMem_lo_hi_189, dataInMem_lo_lo_77};
  wire [63:0]      dataInMem_hi_hi_245 = {dataRegroupBySew_7_2_6, dataRegroupBySew_6_2_6};
  wire [127:0]     dataInMem_hi_357 = {dataInMem_hi_hi_245, dataInMem_hi_lo_133};
  wire [127:0]     dataInMem_lo_302 = {dataInMem_lo_hi_190, dataInMem_lo_lo_78};
  wire [63:0]      dataInMem_hi_hi_246 = {dataRegroupBySew_7_2_7, dataRegroupBySew_6_2_7};
  wire [127:0]     dataInMem_hi_358 = {dataInMem_hi_hi_246, dataInMem_hi_lo_134};
  wire [511:0]     dataInMem_lo_lo_79 = {dataInMem_hi_352, dataInMem_lo_296, dataInMem_hi_351, dataInMem_lo_295};
  wire [511:0]     dataInMem_lo_hi_191 = {dataInMem_hi_354, dataInMem_lo_298, dataInMem_hi_353, dataInMem_lo_297};
  wire [1023:0]    dataInMem_lo_303 = {dataInMem_lo_hi_191, dataInMem_lo_lo_79};
  wire [511:0]     dataInMem_hi_lo_135 = {dataInMem_hi_356, dataInMem_lo_300, dataInMem_hi_355, dataInMem_lo_299};
  wire [511:0]     dataInMem_hi_hi_247 = {dataInMem_hi_358, dataInMem_lo_302, dataInMem_hi_357, dataInMem_lo_301};
  wire [1023:0]    dataInMem_hi_359 = {dataInMem_hi_hi_247, dataInMem_hi_lo_135};
  wire [2047:0]    dataInMem_23 = {dataInMem_hi_359, dataInMem_lo_303};
  wire [255:0]     regroupCacheLine_23_0 = dataInMem_23[255:0];
  wire [255:0]     regroupCacheLine_23_1 = dataInMem_23[511:256];
  wire [255:0]     regroupCacheLine_23_2 = dataInMem_23[767:512];
  wire [255:0]     regroupCacheLine_23_3 = dataInMem_23[1023:768];
  wire [255:0]     regroupCacheLine_23_4 = dataInMem_23[1279:1024];
  wire [255:0]     regroupCacheLine_23_5 = dataInMem_23[1535:1280];
  wire [255:0]     regroupCacheLine_23_6 = dataInMem_23[1791:1536];
  wire [255:0]     regroupCacheLine_23_7 = dataInMem_23[2047:1792];
  wire [255:0]     res_184 = regroupCacheLine_23_0;
  wire [255:0]     res_185 = regroupCacheLine_23_1;
  wire [255:0]     res_186 = regroupCacheLine_23_2;
  wire [255:0]     res_187 = regroupCacheLine_23_3;
  wire [255:0]     res_188 = regroupCacheLine_23_4;
  wire [255:0]     res_189 = regroupCacheLine_23_5;
  wire [255:0]     res_190 = regroupCacheLine_23_6;
  wire [255:0]     res_191 = regroupCacheLine_23_7;
  wire [511:0]     lo_lo_23 = {res_185, res_184};
  wire [511:0]     lo_hi_23 = {res_187, res_186};
  wire [1023:0]    lo_23 = {lo_hi_23, lo_lo_23};
  wire [511:0]     hi_lo_23 = {res_189, res_188};
  wire [511:0]     hi_hi_23 = {res_191, res_190};
  wire [1023:0]    hi_23 = {hi_hi_23, hi_lo_23};
  wire [2047:0]    regroupLoadData_2_7 = {hi_23, lo_23};
  wire             _GEN_284 = lsuRequest_valid | accessBufferDequeueFire;
  wire             _GEN_285 = isLastDataGroup & ~isLastMaskGroup;
  wire             _maskSelect_valid_output = _GEN_284 & _GEN_285;
  wire [7:0][31:0] _GEN_286 = {{maskForBufferData_7}, {maskForBufferData_6}, {maskForBufferData_5}, {maskForBufferData_4}, {maskForBufferData_3}, {maskForBufferData_2}, {maskForBufferData_1}, {maskForBufferData_0}};
  wire [31:0]      _GEN_287 = _GEN_286[cacheLineIndexInBuffer];
  wire             needSendTail = {7'h0, bufferBaseCacheLineIndex} == cacheLineNumberReg;
  assign memRequest_valid_0 = (bufferValid | canSendTail & needSendTail) & addressQueueFree;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo = {cacheLineTemp[8], cacheLineTemp[0]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi = {cacheLineTemp[24], cacheLineTemp[16]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo = {cacheLineTemp[40], cacheLineTemp[32]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi = {cacheLineTemp[56], cacheLineTemp[48]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi = {memRequest_bits_data_lo_lo_lo_hi_hi, memRequest_bits_data_lo_lo_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo = {cacheLineTemp[72], cacheLineTemp[64]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi = {cacheLineTemp[88], cacheLineTemp[80]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo = {memRequest_bits_data_lo_lo_hi_lo_hi, memRequest_bits_data_lo_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo = {cacheLineTemp[104], cacheLineTemp[96]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi = {cacheLineTemp[120], cacheLineTemp[112]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi = {memRequest_bits_data_lo_lo_hi_hi_hi, memRequest_bits_data_lo_lo_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_lo_hi = {memRequest_bits_data_lo_lo_hi_hi, memRequest_bits_data_lo_lo_hi_lo};
  wire [15:0]      memRequest_bits_data_lo_lo = {memRequest_bits_data_lo_lo_hi, memRequest_bits_data_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo = {cacheLineTemp[136], cacheLineTemp[128]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi = {cacheLineTemp[152], cacheLineTemp[144]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo = {memRequest_bits_data_lo_hi_lo_lo_hi, memRequest_bits_data_lo_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo = {cacheLineTemp[168], cacheLineTemp[160]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi = {cacheLineTemp[184], cacheLineTemp[176]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi = {memRequest_bits_data_lo_hi_lo_hi_hi, memRequest_bits_data_lo_hi_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_hi_lo = {memRequest_bits_data_lo_hi_lo_hi, memRequest_bits_data_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo = {cacheLineTemp[200], cacheLineTemp[192]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi = {cacheLineTemp[216], cacheLineTemp[208]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo = {memRequest_bits_data_lo_hi_hi_lo_hi, memRequest_bits_data_lo_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo = {cacheLineTemp[232], cacheLineTemp[224]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi = {cacheLineTemp[248], cacheLineTemp[240]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi = {memRequest_bits_data_lo_hi_hi_hi_hi, memRequest_bits_data_lo_hi_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_lo_hi_hi = {memRequest_bits_data_lo_hi_hi_hi, memRequest_bits_data_lo_hi_hi_lo};
  wire [15:0]      memRequest_bits_data_lo_hi = {memRequest_bits_data_lo_hi_hi, memRequest_bits_data_lo_hi_lo};
  wire [31:0]      memRequest_bits_data_lo = {memRequest_bits_data_lo_hi, memRequest_bits_data_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo = {dataBuffer_0[8], dataBuffer_0[0]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi = {dataBuffer_0[24], dataBuffer_0[16]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo = {memRequest_bits_data_hi_lo_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo = {dataBuffer_0[40], dataBuffer_0[32]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi = {dataBuffer_0[56], dataBuffer_0[48]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi = {memRequest_bits_data_hi_lo_lo_hi_hi, memRequest_bits_data_hi_lo_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_lo_lo = {memRequest_bits_data_hi_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo = {dataBuffer_0[72], dataBuffer_0[64]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi = {dataBuffer_0[88], dataBuffer_0[80]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo = {memRequest_bits_data_hi_lo_hi_lo_hi, memRequest_bits_data_hi_lo_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo = {dataBuffer_0[104], dataBuffer_0[96]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi = {dataBuffer_0[120], dataBuffer_0[112]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi = {memRequest_bits_data_hi_lo_hi_hi_hi, memRequest_bits_data_hi_lo_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_lo_hi = {memRequest_bits_data_hi_lo_hi_hi, memRequest_bits_data_hi_lo_hi_lo};
  wire [15:0]      memRequest_bits_data_hi_lo = {memRequest_bits_data_hi_lo_hi, memRequest_bits_data_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo = {dataBuffer_0[136], dataBuffer_0[128]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi = {dataBuffer_0[152], dataBuffer_0[144]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo = {memRequest_bits_data_hi_hi_lo_lo_hi, memRequest_bits_data_hi_hi_lo_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo = {dataBuffer_0[168], dataBuffer_0[160]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi = {dataBuffer_0[184], dataBuffer_0[176]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi = {memRequest_bits_data_hi_hi_lo_hi_hi, memRequest_bits_data_hi_hi_lo_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_hi_lo = {memRequest_bits_data_hi_hi_lo_hi, memRequest_bits_data_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo = {dataBuffer_0[200], dataBuffer_0[192]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi = {dataBuffer_0[216], dataBuffer_0[208]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo = {memRequest_bits_data_hi_hi_hi_lo_hi, memRequest_bits_data_hi_hi_hi_lo_lo};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo = {dataBuffer_0[232], dataBuffer_0[224]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi = {dataBuffer_0[248], dataBuffer_0[240]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_hi_lo};
  wire [7:0]       memRequest_bits_data_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_lo};
  wire [15:0]      memRequest_bits_data_hi_hi = {memRequest_bits_data_hi_hi_hi, memRequest_bits_data_hi_hi_lo};
  wire [31:0]      memRequest_bits_data_hi = {memRequest_bits_data_hi_hi, memRequest_bits_data_hi_lo};
  wire [94:0]      _GEN_288 = {90'h0, initOffset};
  wire [94:0]      _memRequest_bits_data_T_514 = {31'h0, memRequest_bits_data_hi, memRequest_bits_data_lo} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_1 = {cacheLineTemp[9], cacheLineTemp[1]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_1 = {cacheLineTemp[25], cacheLineTemp[17]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_1 = {cacheLineTemp[41], cacheLineTemp[33]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_1 = {cacheLineTemp[57], cacheLineTemp[49]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_1 = {cacheLineTemp[73], cacheLineTemp[65]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_1 = {cacheLineTemp[89], cacheLineTemp[81]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_1 = {memRequest_bits_data_lo_lo_hi_lo_hi_1, memRequest_bits_data_lo_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_1 = {cacheLineTemp[105], cacheLineTemp[97]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_1 = {cacheLineTemp[121], cacheLineTemp[113]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_hi_1, memRequest_bits_data_lo_lo_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_1};
  wire [15:0]      memRequest_bits_data_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_1 = {cacheLineTemp[137], cacheLineTemp[129]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_1 = {cacheLineTemp[153], cacheLineTemp[145]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_1 = {memRequest_bits_data_lo_hi_lo_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_1 = {cacheLineTemp[169], cacheLineTemp[161]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_1 = {cacheLineTemp[185], cacheLineTemp[177]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_1 = {memRequest_bits_data_lo_hi_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_1 = {cacheLineTemp[201], cacheLineTemp[193]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_1 = {cacheLineTemp[217], cacheLineTemp[209]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_1 = {memRequest_bits_data_lo_hi_hi_lo_hi_1, memRequest_bits_data_lo_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_1 = {cacheLineTemp[233], cacheLineTemp[225]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_1 = {cacheLineTemp[249], cacheLineTemp[241]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_1};
  wire [15:0]      memRequest_bits_data_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_1};
  wire [31:0]      memRequest_bits_data_lo_1 = {memRequest_bits_data_lo_hi_1, memRequest_bits_data_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_1 = {dataBuffer_0[9], dataBuffer_0[1]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_1 = {dataBuffer_0[25], dataBuffer_0[17]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_1 = {dataBuffer_0[41], dataBuffer_0[33]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_1 = {dataBuffer_0[57], dataBuffer_0[49]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_1 = {memRequest_bits_data_hi_lo_lo_hi_hi_1, memRequest_bits_data_hi_lo_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_1 = {dataBuffer_0[73], dataBuffer_0[65]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_1 = {dataBuffer_0[89], dataBuffer_0[81]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_lo_hi_1, memRequest_bits_data_hi_lo_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_1 = {dataBuffer_0[105], dataBuffer_0[97]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_1 = {dataBuffer_0[121], dataBuffer_0[113]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_hi_1, memRequest_bits_data_hi_lo_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_1};
  wire [15:0]      memRequest_bits_data_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_1 = {dataBuffer_0[137], dataBuffer_0[129]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_1 = {dataBuffer_0[153], dataBuffer_0[145]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_1 = {memRequest_bits_data_hi_hi_lo_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_1 = {dataBuffer_0[169], dataBuffer_0[161]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_1 = {dataBuffer_0[185], dataBuffer_0[177]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_1 = {memRequest_bits_data_hi_hi_lo_hi_hi_1, memRequest_bits_data_hi_hi_lo_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_1 = {dataBuffer_0[201], dataBuffer_0[193]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_1 = {dataBuffer_0[217], dataBuffer_0[209]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_hi_lo_lo_1};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_1 = {dataBuffer_0[233], dataBuffer_0[225]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_1 = {dataBuffer_0[249], dataBuffer_0[241]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_hi_lo_1};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_1};
  wire [15:0]      memRequest_bits_data_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_1};
  wire [31:0]      memRequest_bits_data_hi_1 = {memRequest_bits_data_hi_hi_1, memRequest_bits_data_hi_lo_1};
  wire [94:0]      _memRequest_bits_data_T_611 = {31'h0, memRequest_bits_data_hi_1, memRequest_bits_data_lo_1} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_2 = {cacheLineTemp[10], cacheLineTemp[2]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_2 = {cacheLineTemp[26], cacheLineTemp[18]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_2 = {cacheLineTemp[42], cacheLineTemp[34]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_2 = {cacheLineTemp[58], cacheLineTemp[50]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_2 = {cacheLineTemp[74], cacheLineTemp[66]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_2 = {cacheLineTemp[90], cacheLineTemp[82]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_2 = {memRequest_bits_data_lo_lo_hi_lo_hi_2, memRequest_bits_data_lo_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_2 = {cacheLineTemp[106], cacheLineTemp[98]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_2 = {cacheLineTemp[122], cacheLineTemp[114]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_hi_2, memRequest_bits_data_lo_lo_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_2};
  wire [15:0]      memRequest_bits_data_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_2 = {cacheLineTemp[138], cacheLineTemp[130]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_2 = {cacheLineTemp[154], cacheLineTemp[146]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_2 = {memRequest_bits_data_lo_hi_lo_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_2 = {cacheLineTemp[170], cacheLineTemp[162]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_2 = {cacheLineTemp[186], cacheLineTemp[178]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_2 = {memRequest_bits_data_lo_hi_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_2 = {cacheLineTemp[202], cacheLineTemp[194]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_2 = {cacheLineTemp[218], cacheLineTemp[210]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_2 = {memRequest_bits_data_lo_hi_hi_lo_hi_2, memRequest_bits_data_lo_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_2 = {cacheLineTemp[234], cacheLineTemp[226]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_2 = {cacheLineTemp[250], cacheLineTemp[242]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_2};
  wire [15:0]      memRequest_bits_data_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_2};
  wire [31:0]      memRequest_bits_data_lo_2 = {memRequest_bits_data_lo_hi_2, memRequest_bits_data_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_2 = {dataBuffer_0[10], dataBuffer_0[2]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_2 = {dataBuffer_0[26], dataBuffer_0[18]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_2 = {dataBuffer_0[42], dataBuffer_0[34]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_2 = {dataBuffer_0[58], dataBuffer_0[50]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_2 = {memRequest_bits_data_hi_lo_lo_hi_hi_2, memRequest_bits_data_hi_lo_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_2 = {dataBuffer_0[74], dataBuffer_0[66]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_2 = {dataBuffer_0[90], dataBuffer_0[82]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_lo_hi_2, memRequest_bits_data_hi_lo_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_2 = {dataBuffer_0[106], dataBuffer_0[98]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_2 = {dataBuffer_0[122], dataBuffer_0[114]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_hi_2, memRequest_bits_data_hi_lo_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_2};
  wire [15:0]      memRequest_bits_data_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_2 = {dataBuffer_0[138], dataBuffer_0[130]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_2 = {dataBuffer_0[154], dataBuffer_0[146]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_2 = {memRequest_bits_data_hi_hi_lo_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_2 = {dataBuffer_0[170], dataBuffer_0[162]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_2 = {dataBuffer_0[186], dataBuffer_0[178]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_2 = {memRequest_bits_data_hi_hi_lo_hi_hi_2, memRequest_bits_data_hi_hi_lo_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_2 = {dataBuffer_0[202], dataBuffer_0[194]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_2 = {dataBuffer_0[218], dataBuffer_0[210]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_hi_lo_lo_2};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_2 = {dataBuffer_0[234], dataBuffer_0[226]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_2 = {dataBuffer_0[250], dataBuffer_0[242]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_hi_lo_2};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_2};
  wire [15:0]      memRequest_bits_data_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_2};
  wire [31:0]      memRequest_bits_data_hi_2 = {memRequest_bits_data_hi_hi_2, memRequest_bits_data_hi_lo_2};
  wire [94:0]      _memRequest_bits_data_T_708 = {31'h0, memRequest_bits_data_hi_2, memRequest_bits_data_lo_2} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_3 = {cacheLineTemp[11], cacheLineTemp[3]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_3 = {cacheLineTemp[27], cacheLineTemp[19]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_3 = {cacheLineTemp[43], cacheLineTemp[35]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_3 = {cacheLineTemp[59], cacheLineTemp[51]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_3 = {cacheLineTemp[75], cacheLineTemp[67]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_3 = {cacheLineTemp[91], cacheLineTemp[83]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_3 = {memRequest_bits_data_lo_lo_hi_lo_hi_3, memRequest_bits_data_lo_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_3 = {cacheLineTemp[107], cacheLineTemp[99]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_3 = {cacheLineTemp[123], cacheLineTemp[115]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_hi_3, memRequest_bits_data_lo_lo_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_3};
  wire [15:0]      memRequest_bits_data_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_3 = {cacheLineTemp[139], cacheLineTemp[131]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_3 = {cacheLineTemp[155], cacheLineTemp[147]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_3 = {memRequest_bits_data_lo_hi_lo_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_3 = {cacheLineTemp[171], cacheLineTemp[163]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_3 = {cacheLineTemp[187], cacheLineTemp[179]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_3 = {memRequest_bits_data_lo_hi_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_3 = {cacheLineTemp[203], cacheLineTemp[195]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_3 = {cacheLineTemp[219], cacheLineTemp[211]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_3 = {memRequest_bits_data_lo_hi_hi_lo_hi_3, memRequest_bits_data_lo_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_3 = {cacheLineTemp[235], cacheLineTemp[227]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_3 = {cacheLineTemp[251], cacheLineTemp[243]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_3};
  wire [15:0]      memRequest_bits_data_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_3};
  wire [31:0]      memRequest_bits_data_lo_3 = {memRequest_bits_data_lo_hi_3, memRequest_bits_data_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_3 = {dataBuffer_0[11], dataBuffer_0[3]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_3 = {dataBuffer_0[27], dataBuffer_0[19]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_3 = {dataBuffer_0[43], dataBuffer_0[35]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_3 = {dataBuffer_0[59], dataBuffer_0[51]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_3 = {memRequest_bits_data_hi_lo_lo_hi_hi_3, memRequest_bits_data_hi_lo_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_3 = {dataBuffer_0[75], dataBuffer_0[67]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_3 = {dataBuffer_0[91], dataBuffer_0[83]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_lo_hi_3, memRequest_bits_data_hi_lo_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_3 = {dataBuffer_0[107], dataBuffer_0[99]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_3 = {dataBuffer_0[123], dataBuffer_0[115]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_hi_3, memRequest_bits_data_hi_lo_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_3};
  wire [15:0]      memRequest_bits_data_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_3 = {dataBuffer_0[139], dataBuffer_0[131]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_3 = {dataBuffer_0[155], dataBuffer_0[147]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_3 = {memRequest_bits_data_hi_hi_lo_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_3 = {dataBuffer_0[171], dataBuffer_0[163]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_3 = {dataBuffer_0[187], dataBuffer_0[179]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_3 = {memRequest_bits_data_hi_hi_lo_hi_hi_3, memRequest_bits_data_hi_hi_lo_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_3 = {dataBuffer_0[203], dataBuffer_0[195]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_3 = {dataBuffer_0[219], dataBuffer_0[211]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_hi_lo_lo_3};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_3 = {dataBuffer_0[235], dataBuffer_0[227]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_3 = {dataBuffer_0[251], dataBuffer_0[243]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_hi_lo_3};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_3};
  wire [15:0]      memRequest_bits_data_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_3};
  wire [31:0]      memRequest_bits_data_hi_3 = {memRequest_bits_data_hi_hi_3, memRequest_bits_data_hi_lo_3};
  wire [94:0]      _memRequest_bits_data_T_805 = {31'h0, memRequest_bits_data_hi_3, memRequest_bits_data_lo_3} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_4 = {cacheLineTemp[12], cacheLineTemp[4]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_4 = {cacheLineTemp[28], cacheLineTemp[20]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_4 = {cacheLineTemp[44], cacheLineTemp[36]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_4 = {cacheLineTemp[60], cacheLineTemp[52]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_4 = {cacheLineTemp[76], cacheLineTemp[68]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_4 = {cacheLineTemp[92], cacheLineTemp[84]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_4 = {memRequest_bits_data_lo_lo_hi_lo_hi_4, memRequest_bits_data_lo_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_4 = {cacheLineTemp[108], cacheLineTemp[100]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_4 = {cacheLineTemp[124], cacheLineTemp[116]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_hi_4, memRequest_bits_data_lo_lo_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_4};
  wire [15:0]      memRequest_bits_data_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_4 = {cacheLineTemp[140], cacheLineTemp[132]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_4 = {cacheLineTemp[156], cacheLineTemp[148]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_4 = {memRequest_bits_data_lo_hi_lo_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_4 = {cacheLineTemp[172], cacheLineTemp[164]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_4 = {cacheLineTemp[188], cacheLineTemp[180]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_4 = {memRequest_bits_data_lo_hi_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_4 = {cacheLineTemp[204], cacheLineTemp[196]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_4 = {cacheLineTemp[220], cacheLineTemp[212]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_4 = {memRequest_bits_data_lo_hi_hi_lo_hi_4, memRequest_bits_data_lo_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_4 = {cacheLineTemp[236], cacheLineTemp[228]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_4 = {cacheLineTemp[252], cacheLineTemp[244]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_4};
  wire [15:0]      memRequest_bits_data_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_4};
  wire [31:0]      memRequest_bits_data_lo_4 = {memRequest_bits_data_lo_hi_4, memRequest_bits_data_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_4 = {dataBuffer_0[12], dataBuffer_0[4]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_4 = {dataBuffer_0[28], dataBuffer_0[20]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_4 = {dataBuffer_0[44], dataBuffer_0[36]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_4 = {dataBuffer_0[60], dataBuffer_0[52]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_4 = {memRequest_bits_data_hi_lo_lo_hi_hi_4, memRequest_bits_data_hi_lo_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_4 = {dataBuffer_0[76], dataBuffer_0[68]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_4 = {dataBuffer_0[92], dataBuffer_0[84]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_lo_hi_4, memRequest_bits_data_hi_lo_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_4 = {dataBuffer_0[108], dataBuffer_0[100]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_4 = {dataBuffer_0[124], dataBuffer_0[116]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_hi_4, memRequest_bits_data_hi_lo_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_4};
  wire [15:0]      memRequest_bits_data_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_4 = {dataBuffer_0[140], dataBuffer_0[132]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_4 = {dataBuffer_0[156], dataBuffer_0[148]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_4 = {memRequest_bits_data_hi_hi_lo_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_4 = {dataBuffer_0[172], dataBuffer_0[164]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_4 = {dataBuffer_0[188], dataBuffer_0[180]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_4 = {memRequest_bits_data_hi_hi_lo_hi_hi_4, memRequest_bits_data_hi_hi_lo_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_4 = {dataBuffer_0[204], dataBuffer_0[196]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_4 = {dataBuffer_0[220], dataBuffer_0[212]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_hi_lo_lo_4};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_4 = {dataBuffer_0[236], dataBuffer_0[228]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_4 = {dataBuffer_0[252], dataBuffer_0[244]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_hi_lo_4};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_4};
  wire [15:0]      memRequest_bits_data_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_4};
  wire [31:0]      memRequest_bits_data_hi_4 = {memRequest_bits_data_hi_hi_4, memRequest_bits_data_hi_lo_4};
  wire [94:0]      _memRequest_bits_data_T_902 = {31'h0, memRequest_bits_data_hi_4, memRequest_bits_data_lo_4} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_5 = {cacheLineTemp[13], cacheLineTemp[5]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_5 = {cacheLineTemp[29], cacheLineTemp[21]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_5 = {cacheLineTemp[45], cacheLineTemp[37]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_5 = {cacheLineTemp[61], cacheLineTemp[53]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_5 = {cacheLineTemp[77], cacheLineTemp[69]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_5 = {cacheLineTemp[93], cacheLineTemp[85]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_5 = {memRequest_bits_data_lo_lo_hi_lo_hi_5, memRequest_bits_data_lo_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_5 = {cacheLineTemp[109], cacheLineTemp[101]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_5 = {cacheLineTemp[125], cacheLineTemp[117]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_hi_5, memRequest_bits_data_lo_lo_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_5};
  wire [15:0]      memRequest_bits_data_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_5 = {cacheLineTemp[141], cacheLineTemp[133]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_5 = {cacheLineTemp[157], cacheLineTemp[149]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_5 = {memRequest_bits_data_lo_hi_lo_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_5 = {cacheLineTemp[173], cacheLineTemp[165]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_5 = {cacheLineTemp[189], cacheLineTemp[181]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_5 = {memRequest_bits_data_lo_hi_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_5 = {cacheLineTemp[205], cacheLineTemp[197]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_5 = {cacheLineTemp[221], cacheLineTemp[213]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_5 = {memRequest_bits_data_lo_hi_hi_lo_hi_5, memRequest_bits_data_lo_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_5 = {cacheLineTemp[237], cacheLineTemp[229]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_5 = {cacheLineTemp[253], cacheLineTemp[245]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_5};
  wire [15:0]      memRequest_bits_data_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_5};
  wire [31:0]      memRequest_bits_data_lo_5 = {memRequest_bits_data_lo_hi_5, memRequest_bits_data_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_5 = {dataBuffer_0[13], dataBuffer_0[5]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_5 = {dataBuffer_0[29], dataBuffer_0[21]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_5 = {dataBuffer_0[45], dataBuffer_0[37]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_5 = {dataBuffer_0[61], dataBuffer_0[53]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_5 = {memRequest_bits_data_hi_lo_lo_hi_hi_5, memRequest_bits_data_hi_lo_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_5 = {dataBuffer_0[77], dataBuffer_0[69]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_5 = {dataBuffer_0[93], dataBuffer_0[85]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_lo_hi_5, memRequest_bits_data_hi_lo_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_5 = {dataBuffer_0[109], dataBuffer_0[101]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_5 = {dataBuffer_0[125], dataBuffer_0[117]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_hi_5, memRequest_bits_data_hi_lo_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_5};
  wire [15:0]      memRequest_bits_data_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_5 = {dataBuffer_0[141], dataBuffer_0[133]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_5 = {dataBuffer_0[157], dataBuffer_0[149]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_5 = {memRequest_bits_data_hi_hi_lo_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_5 = {dataBuffer_0[173], dataBuffer_0[165]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_5 = {dataBuffer_0[189], dataBuffer_0[181]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_5 = {memRequest_bits_data_hi_hi_lo_hi_hi_5, memRequest_bits_data_hi_hi_lo_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_5 = {dataBuffer_0[205], dataBuffer_0[197]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_5 = {dataBuffer_0[221], dataBuffer_0[213]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_hi_lo_lo_5};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_5 = {dataBuffer_0[237], dataBuffer_0[229]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_5 = {dataBuffer_0[253], dataBuffer_0[245]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_hi_lo_5};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_5};
  wire [15:0]      memRequest_bits_data_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_5};
  wire [31:0]      memRequest_bits_data_hi_5 = {memRequest_bits_data_hi_hi_5, memRequest_bits_data_hi_lo_5};
  wire [94:0]      _memRequest_bits_data_T_999 = {31'h0, memRequest_bits_data_hi_5, memRequest_bits_data_lo_5} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_6 = {cacheLineTemp[14], cacheLineTemp[6]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_6 = {cacheLineTemp[30], cacheLineTemp[22]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_6 = {cacheLineTemp[46], cacheLineTemp[38]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_6 = {cacheLineTemp[62], cacheLineTemp[54]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_6 = {cacheLineTemp[78], cacheLineTemp[70]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_6 = {cacheLineTemp[94], cacheLineTemp[86]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_6 = {memRequest_bits_data_lo_lo_hi_lo_hi_6, memRequest_bits_data_lo_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_6 = {cacheLineTemp[110], cacheLineTemp[102]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_6 = {cacheLineTemp[126], cacheLineTemp[118]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_hi_6, memRequest_bits_data_lo_lo_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_6};
  wire [15:0]      memRequest_bits_data_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_6 = {cacheLineTemp[142], cacheLineTemp[134]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_6 = {cacheLineTemp[158], cacheLineTemp[150]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_6 = {memRequest_bits_data_lo_hi_lo_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_6 = {cacheLineTemp[174], cacheLineTemp[166]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_6 = {cacheLineTemp[190], cacheLineTemp[182]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_6 = {memRequest_bits_data_lo_hi_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_6 = {cacheLineTemp[206], cacheLineTemp[198]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_6 = {cacheLineTemp[222], cacheLineTemp[214]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_6 = {memRequest_bits_data_lo_hi_hi_lo_hi_6, memRequest_bits_data_lo_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_6 = {cacheLineTemp[238], cacheLineTemp[230]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_6 = {cacheLineTemp[254], cacheLineTemp[246]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_6};
  wire [15:0]      memRequest_bits_data_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_6};
  wire [31:0]      memRequest_bits_data_lo_6 = {memRequest_bits_data_lo_hi_6, memRequest_bits_data_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_6 = {dataBuffer_0[14], dataBuffer_0[6]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_6 = {dataBuffer_0[30], dataBuffer_0[22]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_6 = {dataBuffer_0[46], dataBuffer_0[38]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_6 = {dataBuffer_0[62], dataBuffer_0[54]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_6 = {memRequest_bits_data_hi_lo_lo_hi_hi_6, memRequest_bits_data_hi_lo_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_6 = {dataBuffer_0[78], dataBuffer_0[70]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_6 = {dataBuffer_0[94], dataBuffer_0[86]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_lo_hi_6, memRequest_bits_data_hi_lo_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_6 = {dataBuffer_0[110], dataBuffer_0[102]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_6 = {dataBuffer_0[126], dataBuffer_0[118]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_hi_6, memRequest_bits_data_hi_lo_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_6};
  wire [15:0]      memRequest_bits_data_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_6 = {dataBuffer_0[142], dataBuffer_0[134]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_6 = {dataBuffer_0[158], dataBuffer_0[150]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_6 = {memRequest_bits_data_hi_hi_lo_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_6 = {dataBuffer_0[174], dataBuffer_0[166]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_6 = {dataBuffer_0[190], dataBuffer_0[182]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_6 = {memRequest_bits_data_hi_hi_lo_hi_hi_6, memRequest_bits_data_hi_hi_lo_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_6 = {dataBuffer_0[206], dataBuffer_0[198]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_6 = {dataBuffer_0[222], dataBuffer_0[214]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_hi_lo_lo_6};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_6 = {dataBuffer_0[238], dataBuffer_0[230]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_6 = {dataBuffer_0[254], dataBuffer_0[246]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_hi_lo_6};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_6};
  wire [15:0]      memRequest_bits_data_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_6};
  wire [31:0]      memRequest_bits_data_hi_6 = {memRequest_bits_data_hi_hi_6, memRequest_bits_data_hi_lo_6};
  wire [94:0]      _memRequest_bits_data_T_1096 = {31'h0, memRequest_bits_data_hi_6, memRequest_bits_data_lo_6} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_lo_7 = {cacheLineTemp[15], cacheLineTemp[7]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_lo_hi_7 = {cacheLineTemp[31], cacheLineTemp[23]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_lo_7 = {cacheLineTemp[47], cacheLineTemp[39]};
  wire [1:0]       memRequest_bits_data_lo_lo_lo_hi_hi_7 = {cacheLineTemp[63], cacheLineTemp[55]};
  wire [3:0]       memRequest_bits_data_lo_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_lo_7 = {cacheLineTemp[79], cacheLineTemp[71]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_lo_hi_7 = {cacheLineTemp[95], cacheLineTemp[87]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_lo_7 = {memRequest_bits_data_lo_lo_hi_lo_hi_7, memRequest_bits_data_lo_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_lo_7 = {cacheLineTemp[111], cacheLineTemp[103]};
  wire [1:0]       memRequest_bits_data_lo_lo_hi_hi_hi_7 = {cacheLineTemp[127], cacheLineTemp[119]};
  wire [3:0]       memRequest_bits_data_lo_lo_hi_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_hi_7, memRequest_bits_data_lo_lo_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_7};
  wire [15:0]      memRequest_bits_data_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_lo_7 = {cacheLineTemp[143], cacheLineTemp[135]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_lo_hi_7 = {cacheLineTemp[159], cacheLineTemp[151]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_lo_7 = {memRequest_bits_data_lo_hi_lo_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_lo_7 = {cacheLineTemp[175], cacheLineTemp[167]};
  wire [1:0]       memRequest_bits_data_lo_hi_lo_hi_hi_7 = {cacheLineTemp[191], cacheLineTemp[183]};
  wire [3:0]       memRequest_bits_data_lo_hi_lo_hi_7 = {memRequest_bits_data_lo_hi_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_lo_7 = {cacheLineTemp[207], cacheLineTemp[199]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_lo_hi_7 = {cacheLineTemp[223], cacheLineTemp[215]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_lo_7 = {memRequest_bits_data_lo_hi_hi_lo_hi_7, memRequest_bits_data_lo_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_lo_7 = {cacheLineTemp[239], cacheLineTemp[231]};
  wire [1:0]       memRequest_bits_data_lo_hi_hi_hi_hi_7 = {cacheLineTemp[255], cacheLineTemp[247]};
  wire [3:0]       memRequest_bits_data_lo_hi_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_7};
  wire [15:0]      memRequest_bits_data_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_7};
  wire [31:0]      memRequest_bits_data_lo_7 = {memRequest_bits_data_lo_hi_7, memRequest_bits_data_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_lo_7 = {dataBuffer_0[15], dataBuffer_0[7]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_lo_hi_7 = {dataBuffer_0[31], dataBuffer_0[23]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_lo_7 = {dataBuffer_0[47], dataBuffer_0[39]};
  wire [1:0]       memRequest_bits_data_hi_lo_lo_hi_hi_7 = {dataBuffer_0[63], dataBuffer_0[55]};
  wire [3:0]       memRequest_bits_data_hi_lo_lo_hi_7 = {memRequest_bits_data_hi_lo_lo_hi_hi_7, memRequest_bits_data_hi_lo_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_lo_7 = {dataBuffer_0[79], dataBuffer_0[71]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_lo_hi_7 = {dataBuffer_0[95], dataBuffer_0[87]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_lo_hi_7, memRequest_bits_data_hi_lo_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_lo_7 = {dataBuffer_0[111], dataBuffer_0[103]};
  wire [1:0]       memRequest_bits_data_hi_lo_hi_hi_hi_7 = {dataBuffer_0[127], dataBuffer_0[119]};
  wire [3:0]       memRequest_bits_data_hi_lo_hi_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_hi_7, memRequest_bits_data_hi_lo_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_7};
  wire [15:0]      memRequest_bits_data_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_lo_7 = {dataBuffer_0[143], dataBuffer_0[135]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_lo_hi_7 = {dataBuffer_0[159], dataBuffer_0[151]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_lo_7 = {memRequest_bits_data_hi_hi_lo_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_lo_7 = {dataBuffer_0[175], dataBuffer_0[167]};
  wire [1:0]       memRequest_bits_data_hi_hi_lo_hi_hi_7 = {dataBuffer_0[191], dataBuffer_0[183]};
  wire [3:0]       memRequest_bits_data_hi_hi_lo_hi_7 = {memRequest_bits_data_hi_hi_lo_hi_hi_7, memRequest_bits_data_hi_hi_lo_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_lo_7 = {dataBuffer_0[207], dataBuffer_0[199]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_lo_hi_7 = {dataBuffer_0[223], dataBuffer_0[215]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_hi_lo_lo_7};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_lo_7 = {dataBuffer_0[239], dataBuffer_0[231]};
  wire [1:0]       memRequest_bits_data_hi_hi_hi_hi_hi_7 = {dataBuffer_0[255], dataBuffer_0[247]};
  wire [3:0]       memRequest_bits_data_hi_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_hi_lo_7};
  wire [7:0]       memRequest_bits_data_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_7};
  wire [15:0]      memRequest_bits_data_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_7};
  wire [31:0]      memRequest_bits_data_hi_7 = {memRequest_bits_data_hi_hi_7, memRequest_bits_data_hi_lo_7};
  wire [94:0]      _memRequest_bits_data_T_1193 = {31'h0, memRequest_bits_data_hi_7, memRequest_bits_data_lo_7} << _GEN_288;
  wire [1:0]       memRequest_bits_data_lo_lo_8 = {_memRequest_bits_data_T_611[0], _memRequest_bits_data_T_514[0]};
  wire [1:0]       memRequest_bits_data_lo_hi_8 = {_memRequest_bits_data_T_805[0], _memRequest_bits_data_T_708[0]};
  wire [3:0]       memRequest_bits_data_lo_8 = {memRequest_bits_data_lo_hi_8, memRequest_bits_data_lo_lo_8};
  wire [1:0]       memRequest_bits_data_hi_lo_8 = {_memRequest_bits_data_T_999[0], _memRequest_bits_data_T_902[0]};
  wire [1:0]       memRequest_bits_data_hi_hi_8 = {_memRequest_bits_data_T_1193[0], _memRequest_bits_data_T_1096[0]};
  wire [3:0]       memRequest_bits_data_hi_8 = {memRequest_bits_data_hi_hi_8, memRequest_bits_data_hi_lo_8};
  wire [1:0]       memRequest_bits_data_lo_lo_9 = {_memRequest_bits_data_T_611[1], _memRequest_bits_data_T_514[1]};
  wire [1:0]       memRequest_bits_data_lo_hi_9 = {_memRequest_bits_data_T_805[1], _memRequest_bits_data_T_708[1]};
  wire [3:0]       memRequest_bits_data_lo_9 = {memRequest_bits_data_lo_hi_9, memRequest_bits_data_lo_lo_9};
  wire [1:0]       memRequest_bits_data_hi_lo_9 = {_memRequest_bits_data_T_999[1], _memRequest_bits_data_T_902[1]};
  wire [1:0]       memRequest_bits_data_hi_hi_9 = {_memRequest_bits_data_T_1193[1], _memRequest_bits_data_T_1096[1]};
  wire [3:0]       memRequest_bits_data_hi_9 = {memRequest_bits_data_hi_hi_9, memRequest_bits_data_hi_lo_9};
  wire [1:0]       memRequest_bits_data_lo_lo_10 = {_memRequest_bits_data_T_611[2], _memRequest_bits_data_T_514[2]};
  wire [1:0]       memRequest_bits_data_lo_hi_10 = {_memRequest_bits_data_T_805[2], _memRequest_bits_data_T_708[2]};
  wire [3:0]       memRequest_bits_data_lo_10 = {memRequest_bits_data_lo_hi_10, memRequest_bits_data_lo_lo_10};
  wire [1:0]       memRequest_bits_data_hi_lo_10 = {_memRequest_bits_data_T_999[2], _memRequest_bits_data_T_902[2]};
  wire [1:0]       memRequest_bits_data_hi_hi_10 = {_memRequest_bits_data_T_1193[2], _memRequest_bits_data_T_1096[2]};
  wire [3:0]       memRequest_bits_data_hi_10 = {memRequest_bits_data_hi_hi_10, memRequest_bits_data_hi_lo_10};
  wire [1:0]       memRequest_bits_data_lo_lo_11 = {_memRequest_bits_data_T_611[3], _memRequest_bits_data_T_514[3]};
  wire [1:0]       memRequest_bits_data_lo_hi_11 = {_memRequest_bits_data_T_805[3], _memRequest_bits_data_T_708[3]};
  wire [3:0]       memRequest_bits_data_lo_11 = {memRequest_bits_data_lo_hi_11, memRequest_bits_data_lo_lo_11};
  wire [1:0]       memRequest_bits_data_hi_lo_11 = {_memRequest_bits_data_T_999[3], _memRequest_bits_data_T_902[3]};
  wire [1:0]       memRequest_bits_data_hi_hi_11 = {_memRequest_bits_data_T_1193[3], _memRequest_bits_data_T_1096[3]};
  wire [3:0]       memRequest_bits_data_hi_11 = {memRequest_bits_data_hi_hi_11, memRequest_bits_data_hi_lo_11};
  wire [1:0]       memRequest_bits_data_lo_lo_12 = {_memRequest_bits_data_T_611[4], _memRequest_bits_data_T_514[4]};
  wire [1:0]       memRequest_bits_data_lo_hi_12 = {_memRequest_bits_data_T_805[4], _memRequest_bits_data_T_708[4]};
  wire [3:0]       memRequest_bits_data_lo_12 = {memRequest_bits_data_lo_hi_12, memRequest_bits_data_lo_lo_12};
  wire [1:0]       memRequest_bits_data_hi_lo_12 = {_memRequest_bits_data_T_999[4], _memRequest_bits_data_T_902[4]};
  wire [1:0]       memRequest_bits_data_hi_hi_12 = {_memRequest_bits_data_T_1193[4], _memRequest_bits_data_T_1096[4]};
  wire [3:0]       memRequest_bits_data_hi_12 = {memRequest_bits_data_hi_hi_12, memRequest_bits_data_hi_lo_12};
  wire [1:0]       memRequest_bits_data_lo_lo_13 = {_memRequest_bits_data_T_611[5], _memRequest_bits_data_T_514[5]};
  wire [1:0]       memRequest_bits_data_lo_hi_13 = {_memRequest_bits_data_T_805[5], _memRequest_bits_data_T_708[5]};
  wire [3:0]       memRequest_bits_data_lo_13 = {memRequest_bits_data_lo_hi_13, memRequest_bits_data_lo_lo_13};
  wire [1:0]       memRequest_bits_data_hi_lo_13 = {_memRequest_bits_data_T_999[5], _memRequest_bits_data_T_902[5]};
  wire [1:0]       memRequest_bits_data_hi_hi_13 = {_memRequest_bits_data_T_1193[5], _memRequest_bits_data_T_1096[5]};
  wire [3:0]       memRequest_bits_data_hi_13 = {memRequest_bits_data_hi_hi_13, memRequest_bits_data_hi_lo_13};
  wire [1:0]       memRequest_bits_data_lo_lo_14 = {_memRequest_bits_data_T_611[6], _memRequest_bits_data_T_514[6]};
  wire [1:0]       memRequest_bits_data_lo_hi_14 = {_memRequest_bits_data_T_805[6], _memRequest_bits_data_T_708[6]};
  wire [3:0]       memRequest_bits_data_lo_14 = {memRequest_bits_data_lo_hi_14, memRequest_bits_data_lo_lo_14};
  wire [1:0]       memRequest_bits_data_hi_lo_14 = {_memRequest_bits_data_T_999[6], _memRequest_bits_data_T_902[6]};
  wire [1:0]       memRequest_bits_data_hi_hi_14 = {_memRequest_bits_data_T_1193[6], _memRequest_bits_data_T_1096[6]};
  wire [3:0]       memRequest_bits_data_hi_14 = {memRequest_bits_data_hi_hi_14, memRequest_bits_data_hi_lo_14};
  wire [1:0]       memRequest_bits_data_lo_lo_15 = {_memRequest_bits_data_T_611[7], _memRequest_bits_data_T_514[7]};
  wire [1:0]       memRequest_bits_data_lo_hi_15 = {_memRequest_bits_data_T_805[7], _memRequest_bits_data_T_708[7]};
  wire [3:0]       memRequest_bits_data_lo_15 = {memRequest_bits_data_lo_hi_15, memRequest_bits_data_lo_lo_15};
  wire [1:0]       memRequest_bits_data_hi_lo_15 = {_memRequest_bits_data_T_999[7], _memRequest_bits_data_T_902[7]};
  wire [1:0]       memRequest_bits_data_hi_hi_15 = {_memRequest_bits_data_T_1193[7], _memRequest_bits_data_T_1096[7]};
  wire [3:0]       memRequest_bits_data_hi_15 = {memRequest_bits_data_hi_hi_15, memRequest_bits_data_hi_lo_15};
  wire [1:0]       memRequest_bits_data_lo_lo_16 = {_memRequest_bits_data_T_611[8], _memRequest_bits_data_T_514[8]};
  wire [1:0]       memRequest_bits_data_lo_hi_16 = {_memRequest_bits_data_T_805[8], _memRequest_bits_data_T_708[8]};
  wire [3:0]       memRequest_bits_data_lo_16 = {memRequest_bits_data_lo_hi_16, memRequest_bits_data_lo_lo_16};
  wire [1:0]       memRequest_bits_data_hi_lo_16 = {_memRequest_bits_data_T_999[8], _memRequest_bits_data_T_902[8]};
  wire [1:0]       memRequest_bits_data_hi_hi_16 = {_memRequest_bits_data_T_1193[8], _memRequest_bits_data_T_1096[8]};
  wire [3:0]       memRequest_bits_data_hi_16 = {memRequest_bits_data_hi_hi_16, memRequest_bits_data_hi_lo_16};
  wire [1:0]       memRequest_bits_data_lo_lo_17 = {_memRequest_bits_data_T_611[9], _memRequest_bits_data_T_514[9]};
  wire [1:0]       memRequest_bits_data_lo_hi_17 = {_memRequest_bits_data_T_805[9], _memRequest_bits_data_T_708[9]};
  wire [3:0]       memRequest_bits_data_lo_17 = {memRequest_bits_data_lo_hi_17, memRequest_bits_data_lo_lo_17};
  wire [1:0]       memRequest_bits_data_hi_lo_17 = {_memRequest_bits_data_T_999[9], _memRequest_bits_data_T_902[9]};
  wire [1:0]       memRequest_bits_data_hi_hi_17 = {_memRequest_bits_data_T_1193[9], _memRequest_bits_data_T_1096[9]};
  wire [3:0]       memRequest_bits_data_hi_17 = {memRequest_bits_data_hi_hi_17, memRequest_bits_data_hi_lo_17};
  wire [1:0]       memRequest_bits_data_lo_lo_18 = {_memRequest_bits_data_T_611[10], _memRequest_bits_data_T_514[10]};
  wire [1:0]       memRequest_bits_data_lo_hi_18 = {_memRequest_bits_data_T_805[10], _memRequest_bits_data_T_708[10]};
  wire [3:0]       memRequest_bits_data_lo_18 = {memRequest_bits_data_lo_hi_18, memRequest_bits_data_lo_lo_18};
  wire [1:0]       memRequest_bits_data_hi_lo_18 = {_memRequest_bits_data_T_999[10], _memRequest_bits_data_T_902[10]};
  wire [1:0]       memRequest_bits_data_hi_hi_18 = {_memRequest_bits_data_T_1193[10], _memRequest_bits_data_T_1096[10]};
  wire [3:0]       memRequest_bits_data_hi_18 = {memRequest_bits_data_hi_hi_18, memRequest_bits_data_hi_lo_18};
  wire [1:0]       memRequest_bits_data_lo_lo_19 = {_memRequest_bits_data_T_611[11], _memRequest_bits_data_T_514[11]};
  wire [1:0]       memRequest_bits_data_lo_hi_19 = {_memRequest_bits_data_T_805[11], _memRequest_bits_data_T_708[11]};
  wire [3:0]       memRequest_bits_data_lo_19 = {memRequest_bits_data_lo_hi_19, memRequest_bits_data_lo_lo_19};
  wire [1:0]       memRequest_bits_data_hi_lo_19 = {_memRequest_bits_data_T_999[11], _memRequest_bits_data_T_902[11]};
  wire [1:0]       memRequest_bits_data_hi_hi_19 = {_memRequest_bits_data_T_1193[11], _memRequest_bits_data_T_1096[11]};
  wire [3:0]       memRequest_bits_data_hi_19 = {memRequest_bits_data_hi_hi_19, memRequest_bits_data_hi_lo_19};
  wire [1:0]       memRequest_bits_data_lo_lo_20 = {_memRequest_bits_data_T_611[12], _memRequest_bits_data_T_514[12]};
  wire [1:0]       memRequest_bits_data_lo_hi_20 = {_memRequest_bits_data_T_805[12], _memRequest_bits_data_T_708[12]};
  wire [3:0]       memRequest_bits_data_lo_20 = {memRequest_bits_data_lo_hi_20, memRequest_bits_data_lo_lo_20};
  wire [1:0]       memRequest_bits_data_hi_lo_20 = {_memRequest_bits_data_T_999[12], _memRequest_bits_data_T_902[12]};
  wire [1:0]       memRequest_bits_data_hi_hi_20 = {_memRequest_bits_data_T_1193[12], _memRequest_bits_data_T_1096[12]};
  wire [3:0]       memRequest_bits_data_hi_20 = {memRequest_bits_data_hi_hi_20, memRequest_bits_data_hi_lo_20};
  wire [1:0]       memRequest_bits_data_lo_lo_21 = {_memRequest_bits_data_T_611[13], _memRequest_bits_data_T_514[13]};
  wire [1:0]       memRequest_bits_data_lo_hi_21 = {_memRequest_bits_data_T_805[13], _memRequest_bits_data_T_708[13]};
  wire [3:0]       memRequest_bits_data_lo_21 = {memRequest_bits_data_lo_hi_21, memRequest_bits_data_lo_lo_21};
  wire [1:0]       memRequest_bits_data_hi_lo_21 = {_memRequest_bits_data_T_999[13], _memRequest_bits_data_T_902[13]};
  wire [1:0]       memRequest_bits_data_hi_hi_21 = {_memRequest_bits_data_T_1193[13], _memRequest_bits_data_T_1096[13]};
  wire [3:0]       memRequest_bits_data_hi_21 = {memRequest_bits_data_hi_hi_21, memRequest_bits_data_hi_lo_21};
  wire [1:0]       memRequest_bits_data_lo_lo_22 = {_memRequest_bits_data_T_611[14], _memRequest_bits_data_T_514[14]};
  wire [1:0]       memRequest_bits_data_lo_hi_22 = {_memRequest_bits_data_T_805[14], _memRequest_bits_data_T_708[14]};
  wire [3:0]       memRequest_bits_data_lo_22 = {memRequest_bits_data_lo_hi_22, memRequest_bits_data_lo_lo_22};
  wire [1:0]       memRequest_bits_data_hi_lo_22 = {_memRequest_bits_data_T_999[14], _memRequest_bits_data_T_902[14]};
  wire [1:0]       memRequest_bits_data_hi_hi_22 = {_memRequest_bits_data_T_1193[14], _memRequest_bits_data_T_1096[14]};
  wire [3:0]       memRequest_bits_data_hi_22 = {memRequest_bits_data_hi_hi_22, memRequest_bits_data_hi_lo_22};
  wire [1:0]       memRequest_bits_data_lo_lo_23 = {_memRequest_bits_data_T_611[15], _memRequest_bits_data_T_514[15]};
  wire [1:0]       memRequest_bits_data_lo_hi_23 = {_memRequest_bits_data_T_805[15], _memRequest_bits_data_T_708[15]};
  wire [3:0]       memRequest_bits_data_lo_23 = {memRequest_bits_data_lo_hi_23, memRequest_bits_data_lo_lo_23};
  wire [1:0]       memRequest_bits_data_hi_lo_23 = {_memRequest_bits_data_T_999[15], _memRequest_bits_data_T_902[15]};
  wire [1:0]       memRequest_bits_data_hi_hi_23 = {_memRequest_bits_data_T_1193[15], _memRequest_bits_data_T_1096[15]};
  wire [3:0]       memRequest_bits_data_hi_23 = {memRequest_bits_data_hi_hi_23, memRequest_bits_data_hi_lo_23};
  wire [1:0]       memRequest_bits_data_lo_lo_24 = {_memRequest_bits_data_T_611[16], _memRequest_bits_data_T_514[16]};
  wire [1:0]       memRequest_bits_data_lo_hi_24 = {_memRequest_bits_data_T_805[16], _memRequest_bits_data_T_708[16]};
  wire [3:0]       memRequest_bits_data_lo_24 = {memRequest_bits_data_lo_hi_24, memRequest_bits_data_lo_lo_24};
  wire [1:0]       memRequest_bits_data_hi_lo_24 = {_memRequest_bits_data_T_999[16], _memRequest_bits_data_T_902[16]};
  wire [1:0]       memRequest_bits_data_hi_hi_24 = {_memRequest_bits_data_T_1193[16], _memRequest_bits_data_T_1096[16]};
  wire [3:0]       memRequest_bits_data_hi_24 = {memRequest_bits_data_hi_hi_24, memRequest_bits_data_hi_lo_24};
  wire [1:0]       memRequest_bits_data_lo_lo_25 = {_memRequest_bits_data_T_611[17], _memRequest_bits_data_T_514[17]};
  wire [1:0]       memRequest_bits_data_lo_hi_25 = {_memRequest_bits_data_T_805[17], _memRequest_bits_data_T_708[17]};
  wire [3:0]       memRequest_bits_data_lo_25 = {memRequest_bits_data_lo_hi_25, memRequest_bits_data_lo_lo_25};
  wire [1:0]       memRequest_bits_data_hi_lo_25 = {_memRequest_bits_data_T_999[17], _memRequest_bits_data_T_902[17]};
  wire [1:0]       memRequest_bits_data_hi_hi_25 = {_memRequest_bits_data_T_1193[17], _memRequest_bits_data_T_1096[17]};
  wire [3:0]       memRequest_bits_data_hi_25 = {memRequest_bits_data_hi_hi_25, memRequest_bits_data_hi_lo_25};
  wire [1:0]       memRequest_bits_data_lo_lo_26 = {_memRequest_bits_data_T_611[18], _memRequest_bits_data_T_514[18]};
  wire [1:0]       memRequest_bits_data_lo_hi_26 = {_memRequest_bits_data_T_805[18], _memRequest_bits_data_T_708[18]};
  wire [3:0]       memRequest_bits_data_lo_26 = {memRequest_bits_data_lo_hi_26, memRequest_bits_data_lo_lo_26};
  wire [1:0]       memRequest_bits_data_hi_lo_26 = {_memRequest_bits_data_T_999[18], _memRequest_bits_data_T_902[18]};
  wire [1:0]       memRequest_bits_data_hi_hi_26 = {_memRequest_bits_data_T_1193[18], _memRequest_bits_data_T_1096[18]};
  wire [3:0]       memRequest_bits_data_hi_26 = {memRequest_bits_data_hi_hi_26, memRequest_bits_data_hi_lo_26};
  wire [1:0]       memRequest_bits_data_lo_lo_27 = {_memRequest_bits_data_T_611[19], _memRequest_bits_data_T_514[19]};
  wire [1:0]       memRequest_bits_data_lo_hi_27 = {_memRequest_bits_data_T_805[19], _memRequest_bits_data_T_708[19]};
  wire [3:0]       memRequest_bits_data_lo_27 = {memRequest_bits_data_lo_hi_27, memRequest_bits_data_lo_lo_27};
  wire [1:0]       memRequest_bits_data_hi_lo_27 = {_memRequest_bits_data_T_999[19], _memRequest_bits_data_T_902[19]};
  wire [1:0]       memRequest_bits_data_hi_hi_27 = {_memRequest_bits_data_T_1193[19], _memRequest_bits_data_T_1096[19]};
  wire [3:0]       memRequest_bits_data_hi_27 = {memRequest_bits_data_hi_hi_27, memRequest_bits_data_hi_lo_27};
  wire [1:0]       memRequest_bits_data_lo_lo_28 = {_memRequest_bits_data_T_611[20], _memRequest_bits_data_T_514[20]};
  wire [1:0]       memRequest_bits_data_lo_hi_28 = {_memRequest_bits_data_T_805[20], _memRequest_bits_data_T_708[20]};
  wire [3:0]       memRequest_bits_data_lo_28 = {memRequest_bits_data_lo_hi_28, memRequest_bits_data_lo_lo_28};
  wire [1:0]       memRequest_bits_data_hi_lo_28 = {_memRequest_bits_data_T_999[20], _memRequest_bits_data_T_902[20]};
  wire [1:0]       memRequest_bits_data_hi_hi_28 = {_memRequest_bits_data_T_1193[20], _memRequest_bits_data_T_1096[20]};
  wire [3:0]       memRequest_bits_data_hi_28 = {memRequest_bits_data_hi_hi_28, memRequest_bits_data_hi_lo_28};
  wire [1:0]       memRequest_bits_data_lo_lo_29 = {_memRequest_bits_data_T_611[21], _memRequest_bits_data_T_514[21]};
  wire [1:0]       memRequest_bits_data_lo_hi_29 = {_memRequest_bits_data_T_805[21], _memRequest_bits_data_T_708[21]};
  wire [3:0]       memRequest_bits_data_lo_29 = {memRequest_bits_data_lo_hi_29, memRequest_bits_data_lo_lo_29};
  wire [1:0]       memRequest_bits_data_hi_lo_29 = {_memRequest_bits_data_T_999[21], _memRequest_bits_data_T_902[21]};
  wire [1:0]       memRequest_bits_data_hi_hi_29 = {_memRequest_bits_data_T_1193[21], _memRequest_bits_data_T_1096[21]};
  wire [3:0]       memRequest_bits_data_hi_29 = {memRequest_bits_data_hi_hi_29, memRequest_bits_data_hi_lo_29};
  wire [1:0]       memRequest_bits_data_lo_lo_30 = {_memRequest_bits_data_T_611[22], _memRequest_bits_data_T_514[22]};
  wire [1:0]       memRequest_bits_data_lo_hi_30 = {_memRequest_bits_data_T_805[22], _memRequest_bits_data_T_708[22]};
  wire [3:0]       memRequest_bits_data_lo_30 = {memRequest_bits_data_lo_hi_30, memRequest_bits_data_lo_lo_30};
  wire [1:0]       memRequest_bits_data_hi_lo_30 = {_memRequest_bits_data_T_999[22], _memRequest_bits_data_T_902[22]};
  wire [1:0]       memRequest_bits_data_hi_hi_30 = {_memRequest_bits_data_T_1193[22], _memRequest_bits_data_T_1096[22]};
  wire [3:0]       memRequest_bits_data_hi_30 = {memRequest_bits_data_hi_hi_30, memRequest_bits_data_hi_lo_30};
  wire [1:0]       memRequest_bits_data_lo_lo_31 = {_memRequest_bits_data_T_611[23], _memRequest_bits_data_T_514[23]};
  wire [1:0]       memRequest_bits_data_lo_hi_31 = {_memRequest_bits_data_T_805[23], _memRequest_bits_data_T_708[23]};
  wire [3:0]       memRequest_bits_data_lo_31 = {memRequest_bits_data_lo_hi_31, memRequest_bits_data_lo_lo_31};
  wire [1:0]       memRequest_bits_data_hi_lo_31 = {_memRequest_bits_data_T_999[23], _memRequest_bits_data_T_902[23]};
  wire [1:0]       memRequest_bits_data_hi_hi_31 = {_memRequest_bits_data_T_1193[23], _memRequest_bits_data_T_1096[23]};
  wire [3:0]       memRequest_bits_data_hi_31 = {memRequest_bits_data_hi_hi_31, memRequest_bits_data_hi_lo_31};
  wire [1:0]       memRequest_bits_data_lo_lo_32 = {_memRequest_bits_data_T_611[24], _memRequest_bits_data_T_514[24]};
  wire [1:0]       memRequest_bits_data_lo_hi_32 = {_memRequest_bits_data_T_805[24], _memRequest_bits_data_T_708[24]};
  wire [3:0]       memRequest_bits_data_lo_32 = {memRequest_bits_data_lo_hi_32, memRequest_bits_data_lo_lo_32};
  wire [1:0]       memRequest_bits_data_hi_lo_32 = {_memRequest_bits_data_T_999[24], _memRequest_bits_data_T_902[24]};
  wire [1:0]       memRequest_bits_data_hi_hi_32 = {_memRequest_bits_data_T_1193[24], _memRequest_bits_data_T_1096[24]};
  wire [3:0]       memRequest_bits_data_hi_32 = {memRequest_bits_data_hi_hi_32, memRequest_bits_data_hi_lo_32};
  wire [1:0]       memRequest_bits_data_lo_lo_33 = {_memRequest_bits_data_T_611[25], _memRequest_bits_data_T_514[25]};
  wire [1:0]       memRequest_bits_data_lo_hi_33 = {_memRequest_bits_data_T_805[25], _memRequest_bits_data_T_708[25]};
  wire [3:0]       memRequest_bits_data_lo_33 = {memRequest_bits_data_lo_hi_33, memRequest_bits_data_lo_lo_33};
  wire [1:0]       memRequest_bits_data_hi_lo_33 = {_memRequest_bits_data_T_999[25], _memRequest_bits_data_T_902[25]};
  wire [1:0]       memRequest_bits_data_hi_hi_33 = {_memRequest_bits_data_T_1193[25], _memRequest_bits_data_T_1096[25]};
  wire [3:0]       memRequest_bits_data_hi_33 = {memRequest_bits_data_hi_hi_33, memRequest_bits_data_hi_lo_33};
  wire [1:0]       memRequest_bits_data_lo_lo_34 = {_memRequest_bits_data_T_611[26], _memRequest_bits_data_T_514[26]};
  wire [1:0]       memRequest_bits_data_lo_hi_34 = {_memRequest_bits_data_T_805[26], _memRequest_bits_data_T_708[26]};
  wire [3:0]       memRequest_bits_data_lo_34 = {memRequest_bits_data_lo_hi_34, memRequest_bits_data_lo_lo_34};
  wire [1:0]       memRequest_bits_data_hi_lo_34 = {_memRequest_bits_data_T_999[26], _memRequest_bits_data_T_902[26]};
  wire [1:0]       memRequest_bits_data_hi_hi_34 = {_memRequest_bits_data_T_1193[26], _memRequest_bits_data_T_1096[26]};
  wire [3:0]       memRequest_bits_data_hi_34 = {memRequest_bits_data_hi_hi_34, memRequest_bits_data_hi_lo_34};
  wire [1:0]       memRequest_bits_data_lo_lo_35 = {_memRequest_bits_data_T_611[27], _memRequest_bits_data_T_514[27]};
  wire [1:0]       memRequest_bits_data_lo_hi_35 = {_memRequest_bits_data_T_805[27], _memRequest_bits_data_T_708[27]};
  wire [3:0]       memRequest_bits_data_lo_35 = {memRequest_bits_data_lo_hi_35, memRequest_bits_data_lo_lo_35};
  wire [1:0]       memRequest_bits_data_hi_lo_35 = {_memRequest_bits_data_T_999[27], _memRequest_bits_data_T_902[27]};
  wire [1:0]       memRequest_bits_data_hi_hi_35 = {_memRequest_bits_data_T_1193[27], _memRequest_bits_data_T_1096[27]};
  wire [3:0]       memRequest_bits_data_hi_35 = {memRequest_bits_data_hi_hi_35, memRequest_bits_data_hi_lo_35};
  wire [1:0]       memRequest_bits_data_lo_lo_36 = {_memRequest_bits_data_T_611[28], _memRequest_bits_data_T_514[28]};
  wire [1:0]       memRequest_bits_data_lo_hi_36 = {_memRequest_bits_data_T_805[28], _memRequest_bits_data_T_708[28]};
  wire [3:0]       memRequest_bits_data_lo_36 = {memRequest_bits_data_lo_hi_36, memRequest_bits_data_lo_lo_36};
  wire [1:0]       memRequest_bits_data_hi_lo_36 = {_memRequest_bits_data_T_999[28], _memRequest_bits_data_T_902[28]};
  wire [1:0]       memRequest_bits_data_hi_hi_36 = {_memRequest_bits_data_T_1193[28], _memRequest_bits_data_T_1096[28]};
  wire [3:0]       memRequest_bits_data_hi_36 = {memRequest_bits_data_hi_hi_36, memRequest_bits_data_hi_lo_36};
  wire [1:0]       memRequest_bits_data_lo_lo_37 = {_memRequest_bits_data_T_611[29], _memRequest_bits_data_T_514[29]};
  wire [1:0]       memRequest_bits_data_lo_hi_37 = {_memRequest_bits_data_T_805[29], _memRequest_bits_data_T_708[29]};
  wire [3:0]       memRequest_bits_data_lo_37 = {memRequest_bits_data_lo_hi_37, memRequest_bits_data_lo_lo_37};
  wire [1:0]       memRequest_bits_data_hi_lo_37 = {_memRequest_bits_data_T_999[29], _memRequest_bits_data_T_902[29]};
  wire [1:0]       memRequest_bits_data_hi_hi_37 = {_memRequest_bits_data_T_1193[29], _memRequest_bits_data_T_1096[29]};
  wire [3:0]       memRequest_bits_data_hi_37 = {memRequest_bits_data_hi_hi_37, memRequest_bits_data_hi_lo_37};
  wire [1:0]       memRequest_bits_data_lo_lo_38 = {_memRequest_bits_data_T_611[30], _memRequest_bits_data_T_514[30]};
  wire [1:0]       memRequest_bits_data_lo_hi_38 = {_memRequest_bits_data_T_805[30], _memRequest_bits_data_T_708[30]};
  wire [3:0]       memRequest_bits_data_lo_38 = {memRequest_bits_data_lo_hi_38, memRequest_bits_data_lo_lo_38};
  wire [1:0]       memRequest_bits_data_hi_lo_38 = {_memRequest_bits_data_T_999[30], _memRequest_bits_data_T_902[30]};
  wire [1:0]       memRequest_bits_data_hi_hi_38 = {_memRequest_bits_data_T_1193[30], _memRequest_bits_data_T_1096[30]};
  wire [3:0]       memRequest_bits_data_hi_38 = {memRequest_bits_data_hi_hi_38, memRequest_bits_data_hi_lo_38};
  wire [1:0]       memRequest_bits_data_lo_lo_39 = {_memRequest_bits_data_T_611[31], _memRequest_bits_data_T_514[31]};
  wire [1:0]       memRequest_bits_data_lo_hi_39 = {_memRequest_bits_data_T_805[31], _memRequest_bits_data_T_708[31]};
  wire [3:0]       memRequest_bits_data_lo_39 = {memRequest_bits_data_lo_hi_39, memRequest_bits_data_lo_lo_39};
  wire [1:0]       memRequest_bits_data_hi_lo_39 = {_memRequest_bits_data_T_999[31], _memRequest_bits_data_T_902[31]};
  wire [1:0]       memRequest_bits_data_hi_hi_39 = {_memRequest_bits_data_T_1193[31], _memRequest_bits_data_T_1096[31]};
  wire [3:0]       memRequest_bits_data_hi_39 = {memRequest_bits_data_hi_hi_39, memRequest_bits_data_hi_lo_39};
  wire [1:0]       memRequest_bits_data_lo_lo_40 = {_memRequest_bits_data_T_611[32], _memRequest_bits_data_T_514[32]};
  wire [1:0]       memRequest_bits_data_lo_hi_40 = {_memRequest_bits_data_T_805[32], _memRequest_bits_data_T_708[32]};
  wire [3:0]       memRequest_bits_data_lo_40 = {memRequest_bits_data_lo_hi_40, memRequest_bits_data_lo_lo_40};
  wire [1:0]       memRequest_bits_data_hi_lo_40 = {_memRequest_bits_data_T_999[32], _memRequest_bits_data_T_902[32]};
  wire [1:0]       memRequest_bits_data_hi_hi_40 = {_memRequest_bits_data_T_1193[32], _memRequest_bits_data_T_1096[32]};
  wire [3:0]       memRequest_bits_data_hi_40 = {memRequest_bits_data_hi_hi_40, memRequest_bits_data_hi_lo_40};
  wire [1:0]       memRequest_bits_data_lo_lo_41 = {_memRequest_bits_data_T_611[33], _memRequest_bits_data_T_514[33]};
  wire [1:0]       memRequest_bits_data_lo_hi_41 = {_memRequest_bits_data_T_805[33], _memRequest_bits_data_T_708[33]};
  wire [3:0]       memRequest_bits_data_lo_41 = {memRequest_bits_data_lo_hi_41, memRequest_bits_data_lo_lo_41};
  wire [1:0]       memRequest_bits_data_hi_lo_41 = {_memRequest_bits_data_T_999[33], _memRequest_bits_data_T_902[33]};
  wire [1:0]       memRequest_bits_data_hi_hi_41 = {_memRequest_bits_data_T_1193[33], _memRequest_bits_data_T_1096[33]};
  wire [3:0]       memRequest_bits_data_hi_41 = {memRequest_bits_data_hi_hi_41, memRequest_bits_data_hi_lo_41};
  wire [1:0]       memRequest_bits_data_lo_lo_42 = {_memRequest_bits_data_T_611[34], _memRequest_bits_data_T_514[34]};
  wire [1:0]       memRequest_bits_data_lo_hi_42 = {_memRequest_bits_data_T_805[34], _memRequest_bits_data_T_708[34]};
  wire [3:0]       memRequest_bits_data_lo_42 = {memRequest_bits_data_lo_hi_42, memRequest_bits_data_lo_lo_42};
  wire [1:0]       memRequest_bits_data_hi_lo_42 = {_memRequest_bits_data_T_999[34], _memRequest_bits_data_T_902[34]};
  wire [1:0]       memRequest_bits_data_hi_hi_42 = {_memRequest_bits_data_T_1193[34], _memRequest_bits_data_T_1096[34]};
  wire [3:0]       memRequest_bits_data_hi_42 = {memRequest_bits_data_hi_hi_42, memRequest_bits_data_hi_lo_42};
  wire [1:0]       memRequest_bits_data_lo_lo_43 = {_memRequest_bits_data_T_611[35], _memRequest_bits_data_T_514[35]};
  wire [1:0]       memRequest_bits_data_lo_hi_43 = {_memRequest_bits_data_T_805[35], _memRequest_bits_data_T_708[35]};
  wire [3:0]       memRequest_bits_data_lo_43 = {memRequest_bits_data_lo_hi_43, memRequest_bits_data_lo_lo_43};
  wire [1:0]       memRequest_bits_data_hi_lo_43 = {_memRequest_bits_data_T_999[35], _memRequest_bits_data_T_902[35]};
  wire [1:0]       memRequest_bits_data_hi_hi_43 = {_memRequest_bits_data_T_1193[35], _memRequest_bits_data_T_1096[35]};
  wire [3:0]       memRequest_bits_data_hi_43 = {memRequest_bits_data_hi_hi_43, memRequest_bits_data_hi_lo_43};
  wire [1:0]       memRequest_bits_data_lo_lo_44 = {_memRequest_bits_data_T_611[36], _memRequest_bits_data_T_514[36]};
  wire [1:0]       memRequest_bits_data_lo_hi_44 = {_memRequest_bits_data_T_805[36], _memRequest_bits_data_T_708[36]};
  wire [3:0]       memRequest_bits_data_lo_44 = {memRequest_bits_data_lo_hi_44, memRequest_bits_data_lo_lo_44};
  wire [1:0]       memRequest_bits_data_hi_lo_44 = {_memRequest_bits_data_T_999[36], _memRequest_bits_data_T_902[36]};
  wire [1:0]       memRequest_bits_data_hi_hi_44 = {_memRequest_bits_data_T_1193[36], _memRequest_bits_data_T_1096[36]};
  wire [3:0]       memRequest_bits_data_hi_44 = {memRequest_bits_data_hi_hi_44, memRequest_bits_data_hi_lo_44};
  wire [1:0]       memRequest_bits_data_lo_lo_45 = {_memRequest_bits_data_T_611[37], _memRequest_bits_data_T_514[37]};
  wire [1:0]       memRequest_bits_data_lo_hi_45 = {_memRequest_bits_data_T_805[37], _memRequest_bits_data_T_708[37]};
  wire [3:0]       memRequest_bits_data_lo_45 = {memRequest_bits_data_lo_hi_45, memRequest_bits_data_lo_lo_45};
  wire [1:0]       memRequest_bits_data_hi_lo_45 = {_memRequest_bits_data_T_999[37], _memRequest_bits_data_T_902[37]};
  wire [1:0]       memRequest_bits_data_hi_hi_45 = {_memRequest_bits_data_T_1193[37], _memRequest_bits_data_T_1096[37]};
  wire [3:0]       memRequest_bits_data_hi_45 = {memRequest_bits_data_hi_hi_45, memRequest_bits_data_hi_lo_45};
  wire [1:0]       memRequest_bits_data_lo_lo_46 = {_memRequest_bits_data_T_611[38], _memRequest_bits_data_T_514[38]};
  wire [1:0]       memRequest_bits_data_lo_hi_46 = {_memRequest_bits_data_T_805[38], _memRequest_bits_data_T_708[38]};
  wire [3:0]       memRequest_bits_data_lo_46 = {memRequest_bits_data_lo_hi_46, memRequest_bits_data_lo_lo_46};
  wire [1:0]       memRequest_bits_data_hi_lo_46 = {_memRequest_bits_data_T_999[38], _memRequest_bits_data_T_902[38]};
  wire [1:0]       memRequest_bits_data_hi_hi_46 = {_memRequest_bits_data_T_1193[38], _memRequest_bits_data_T_1096[38]};
  wire [3:0]       memRequest_bits_data_hi_46 = {memRequest_bits_data_hi_hi_46, memRequest_bits_data_hi_lo_46};
  wire [1:0]       memRequest_bits_data_lo_lo_47 = {_memRequest_bits_data_T_611[39], _memRequest_bits_data_T_514[39]};
  wire [1:0]       memRequest_bits_data_lo_hi_47 = {_memRequest_bits_data_T_805[39], _memRequest_bits_data_T_708[39]};
  wire [3:0]       memRequest_bits_data_lo_47 = {memRequest_bits_data_lo_hi_47, memRequest_bits_data_lo_lo_47};
  wire [1:0]       memRequest_bits_data_hi_lo_47 = {_memRequest_bits_data_T_999[39], _memRequest_bits_data_T_902[39]};
  wire [1:0]       memRequest_bits_data_hi_hi_47 = {_memRequest_bits_data_T_1193[39], _memRequest_bits_data_T_1096[39]};
  wire [3:0]       memRequest_bits_data_hi_47 = {memRequest_bits_data_hi_hi_47, memRequest_bits_data_hi_lo_47};
  wire [1:0]       memRequest_bits_data_lo_lo_48 = {_memRequest_bits_data_T_611[40], _memRequest_bits_data_T_514[40]};
  wire [1:0]       memRequest_bits_data_lo_hi_48 = {_memRequest_bits_data_T_805[40], _memRequest_bits_data_T_708[40]};
  wire [3:0]       memRequest_bits_data_lo_48 = {memRequest_bits_data_lo_hi_48, memRequest_bits_data_lo_lo_48};
  wire [1:0]       memRequest_bits_data_hi_lo_48 = {_memRequest_bits_data_T_999[40], _memRequest_bits_data_T_902[40]};
  wire [1:0]       memRequest_bits_data_hi_hi_48 = {_memRequest_bits_data_T_1193[40], _memRequest_bits_data_T_1096[40]};
  wire [3:0]       memRequest_bits_data_hi_48 = {memRequest_bits_data_hi_hi_48, memRequest_bits_data_hi_lo_48};
  wire [1:0]       memRequest_bits_data_lo_lo_49 = {_memRequest_bits_data_T_611[41], _memRequest_bits_data_T_514[41]};
  wire [1:0]       memRequest_bits_data_lo_hi_49 = {_memRequest_bits_data_T_805[41], _memRequest_bits_data_T_708[41]};
  wire [3:0]       memRequest_bits_data_lo_49 = {memRequest_bits_data_lo_hi_49, memRequest_bits_data_lo_lo_49};
  wire [1:0]       memRequest_bits_data_hi_lo_49 = {_memRequest_bits_data_T_999[41], _memRequest_bits_data_T_902[41]};
  wire [1:0]       memRequest_bits_data_hi_hi_49 = {_memRequest_bits_data_T_1193[41], _memRequest_bits_data_T_1096[41]};
  wire [3:0]       memRequest_bits_data_hi_49 = {memRequest_bits_data_hi_hi_49, memRequest_bits_data_hi_lo_49};
  wire [1:0]       memRequest_bits_data_lo_lo_50 = {_memRequest_bits_data_T_611[42], _memRequest_bits_data_T_514[42]};
  wire [1:0]       memRequest_bits_data_lo_hi_50 = {_memRequest_bits_data_T_805[42], _memRequest_bits_data_T_708[42]};
  wire [3:0]       memRequest_bits_data_lo_50 = {memRequest_bits_data_lo_hi_50, memRequest_bits_data_lo_lo_50};
  wire [1:0]       memRequest_bits_data_hi_lo_50 = {_memRequest_bits_data_T_999[42], _memRequest_bits_data_T_902[42]};
  wire [1:0]       memRequest_bits_data_hi_hi_50 = {_memRequest_bits_data_T_1193[42], _memRequest_bits_data_T_1096[42]};
  wire [3:0]       memRequest_bits_data_hi_50 = {memRequest_bits_data_hi_hi_50, memRequest_bits_data_hi_lo_50};
  wire [1:0]       memRequest_bits_data_lo_lo_51 = {_memRequest_bits_data_T_611[43], _memRequest_bits_data_T_514[43]};
  wire [1:0]       memRequest_bits_data_lo_hi_51 = {_memRequest_bits_data_T_805[43], _memRequest_bits_data_T_708[43]};
  wire [3:0]       memRequest_bits_data_lo_51 = {memRequest_bits_data_lo_hi_51, memRequest_bits_data_lo_lo_51};
  wire [1:0]       memRequest_bits_data_hi_lo_51 = {_memRequest_bits_data_T_999[43], _memRequest_bits_data_T_902[43]};
  wire [1:0]       memRequest_bits_data_hi_hi_51 = {_memRequest_bits_data_T_1193[43], _memRequest_bits_data_T_1096[43]};
  wire [3:0]       memRequest_bits_data_hi_51 = {memRequest_bits_data_hi_hi_51, memRequest_bits_data_hi_lo_51};
  wire [1:0]       memRequest_bits_data_lo_lo_52 = {_memRequest_bits_data_T_611[44], _memRequest_bits_data_T_514[44]};
  wire [1:0]       memRequest_bits_data_lo_hi_52 = {_memRequest_bits_data_T_805[44], _memRequest_bits_data_T_708[44]};
  wire [3:0]       memRequest_bits_data_lo_52 = {memRequest_bits_data_lo_hi_52, memRequest_bits_data_lo_lo_52};
  wire [1:0]       memRequest_bits_data_hi_lo_52 = {_memRequest_bits_data_T_999[44], _memRequest_bits_data_T_902[44]};
  wire [1:0]       memRequest_bits_data_hi_hi_52 = {_memRequest_bits_data_T_1193[44], _memRequest_bits_data_T_1096[44]};
  wire [3:0]       memRequest_bits_data_hi_52 = {memRequest_bits_data_hi_hi_52, memRequest_bits_data_hi_lo_52};
  wire [1:0]       memRequest_bits_data_lo_lo_53 = {_memRequest_bits_data_T_611[45], _memRequest_bits_data_T_514[45]};
  wire [1:0]       memRequest_bits_data_lo_hi_53 = {_memRequest_bits_data_T_805[45], _memRequest_bits_data_T_708[45]};
  wire [3:0]       memRequest_bits_data_lo_53 = {memRequest_bits_data_lo_hi_53, memRequest_bits_data_lo_lo_53};
  wire [1:0]       memRequest_bits_data_hi_lo_53 = {_memRequest_bits_data_T_999[45], _memRequest_bits_data_T_902[45]};
  wire [1:0]       memRequest_bits_data_hi_hi_53 = {_memRequest_bits_data_T_1193[45], _memRequest_bits_data_T_1096[45]};
  wire [3:0]       memRequest_bits_data_hi_53 = {memRequest_bits_data_hi_hi_53, memRequest_bits_data_hi_lo_53};
  wire [1:0]       memRequest_bits_data_lo_lo_54 = {_memRequest_bits_data_T_611[46], _memRequest_bits_data_T_514[46]};
  wire [1:0]       memRequest_bits_data_lo_hi_54 = {_memRequest_bits_data_T_805[46], _memRequest_bits_data_T_708[46]};
  wire [3:0]       memRequest_bits_data_lo_54 = {memRequest_bits_data_lo_hi_54, memRequest_bits_data_lo_lo_54};
  wire [1:0]       memRequest_bits_data_hi_lo_54 = {_memRequest_bits_data_T_999[46], _memRequest_bits_data_T_902[46]};
  wire [1:0]       memRequest_bits_data_hi_hi_54 = {_memRequest_bits_data_T_1193[46], _memRequest_bits_data_T_1096[46]};
  wire [3:0]       memRequest_bits_data_hi_54 = {memRequest_bits_data_hi_hi_54, memRequest_bits_data_hi_lo_54};
  wire [1:0]       memRequest_bits_data_lo_lo_55 = {_memRequest_bits_data_T_611[47], _memRequest_bits_data_T_514[47]};
  wire [1:0]       memRequest_bits_data_lo_hi_55 = {_memRequest_bits_data_T_805[47], _memRequest_bits_data_T_708[47]};
  wire [3:0]       memRequest_bits_data_lo_55 = {memRequest_bits_data_lo_hi_55, memRequest_bits_data_lo_lo_55};
  wire [1:0]       memRequest_bits_data_hi_lo_55 = {_memRequest_bits_data_T_999[47], _memRequest_bits_data_T_902[47]};
  wire [1:0]       memRequest_bits_data_hi_hi_55 = {_memRequest_bits_data_T_1193[47], _memRequest_bits_data_T_1096[47]};
  wire [3:0]       memRequest_bits_data_hi_55 = {memRequest_bits_data_hi_hi_55, memRequest_bits_data_hi_lo_55};
  wire [1:0]       memRequest_bits_data_lo_lo_56 = {_memRequest_bits_data_T_611[48], _memRequest_bits_data_T_514[48]};
  wire [1:0]       memRequest_bits_data_lo_hi_56 = {_memRequest_bits_data_T_805[48], _memRequest_bits_data_T_708[48]};
  wire [3:0]       memRequest_bits_data_lo_56 = {memRequest_bits_data_lo_hi_56, memRequest_bits_data_lo_lo_56};
  wire [1:0]       memRequest_bits_data_hi_lo_56 = {_memRequest_bits_data_T_999[48], _memRequest_bits_data_T_902[48]};
  wire [1:0]       memRequest_bits_data_hi_hi_56 = {_memRequest_bits_data_T_1193[48], _memRequest_bits_data_T_1096[48]};
  wire [3:0]       memRequest_bits_data_hi_56 = {memRequest_bits_data_hi_hi_56, memRequest_bits_data_hi_lo_56};
  wire [1:0]       memRequest_bits_data_lo_lo_57 = {_memRequest_bits_data_T_611[49], _memRequest_bits_data_T_514[49]};
  wire [1:0]       memRequest_bits_data_lo_hi_57 = {_memRequest_bits_data_T_805[49], _memRequest_bits_data_T_708[49]};
  wire [3:0]       memRequest_bits_data_lo_57 = {memRequest_bits_data_lo_hi_57, memRequest_bits_data_lo_lo_57};
  wire [1:0]       memRequest_bits_data_hi_lo_57 = {_memRequest_bits_data_T_999[49], _memRequest_bits_data_T_902[49]};
  wire [1:0]       memRequest_bits_data_hi_hi_57 = {_memRequest_bits_data_T_1193[49], _memRequest_bits_data_T_1096[49]};
  wire [3:0]       memRequest_bits_data_hi_57 = {memRequest_bits_data_hi_hi_57, memRequest_bits_data_hi_lo_57};
  wire [1:0]       memRequest_bits_data_lo_lo_58 = {_memRequest_bits_data_T_611[50], _memRequest_bits_data_T_514[50]};
  wire [1:0]       memRequest_bits_data_lo_hi_58 = {_memRequest_bits_data_T_805[50], _memRequest_bits_data_T_708[50]};
  wire [3:0]       memRequest_bits_data_lo_58 = {memRequest_bits_data_lo_hi_58, memRequest_bits_data_lo_lo_58};
  wire [1:0]       memRequest_bits_data_hi_lo_58 = {_memRequest_bits_data_T_999[50], _memRequest_bits_data_T_902[50]};
  wire [1:0]       memRequest_bits_data_hi_hi_58 = {_memRequest_bits_data_T_1193[50], _memRequest_bits_data_T_1096[50]};
  wire [3:0]       memRequest_bits_data_hi_58 = {memRequest_bits_data_hi_hi_58, memRequest_bits_data_hi_lo_58};
  wire [1:0]       memRequest_bits_data_lo_lo_59 = {_memRequest_bits_data_T_611[51], _memRequest_bits_data_T_514[51]};
  wire [1:0]       memRequest_bits_data_lo_hi_59 = {_memRequest_bits_data_T_805[51], _memRequest_bits_data_T_708[51]};
  wire [3:0]       memRequest_bits_data_lo_59 = {memRequest_bits_data_lo_hi_59, memRequest_bits_data_lo_lo_59};
  wire [1:0]       memRequest_bits_data_hi_lo_59 = {_memRequest_bits_data_T_999[51], _memRequest_bits_data_T_902[51]};
  wire [1:0]       memRequest_bits_data_hi_hi_59 = {_memRequest_bits_data_T_1193[51], _memRequest_bits_data_T_1096[51]};
  wire [3:0]       memRequest_bits_data_hi_59 = {memRequest_bits_data_hi_hi_59, memRequest_bits_data_hi_lo_59};
  wire [1:0]       memRequest_bits_data_lo_lo_60 = {_memRequest_bits_data_T_611[52], _memRequest_bits_data_T_514[52]};
  wire [1:0]       memRequest_bits_data_lo_hi_60 = {_memRequest_bits_data_T_805[52], _memRequest_bits_data_T_708[52]};
  wire [3:0]       memRequest_bits_data_lo_60 = {memRequest_bits_data_lo_hi_60, memRequest_bits_data_lo_lo_60};
  wire [1:0]       memRequest_bits_data_hi_lo_60 = {_memRequest_bits_data_T_999[52], _memRequest_bits_data_T_902[52]};
  wire [1:0]       memRequest_bits_data_hi_hi_60 = {_memRequest_bits_data_T_1193[52], _memRequest_bits_data_T_1096[52]};
  wire [3:0]       memRequest_bits_data_hi_60 = {memRequest_bits_data_hi_hi_60, memRequest_bits_data_hi_lo_60};
  wire [1:0]       memRequest_bits_data_lo_lo_61 = {_memRequest_bits_data_T_611[53], _memRequest_bits_data_T_514[53]};
  wire [1:0]       memRequest_bits_data_lo_hi_61 = {_memRequest_bits_data_T_805[53], _memRequest_bits_data_T_708[53]};
  wire [3:0]       memRequest_bits_data_lo_61 = {memRequest_bits_data_lo_hi_61, memRequest_bits_data_lo_lo_61};
  wire [1:0]       memRequest_bits_data_hi_lo_61 = {_memRequest_bits_data_T_999[53], _memRequest_bits_data_T_902[53]};
  wire [1:0]       memRequest_bits_data_hi_hi_61 = {_memRequest_bits_data_T_1193[53], _memRequest_bits_data_T_1096[53]};
  wire [3:0]       memRequest_bits_data_hi_61 = {memRequest_bits_data_hi_hi_61, memRequest_bits_data_hi_lo_61};
  wire [1:0]       memRequest_bits_data_lo_lo_62 = {_memRequest_bits_data_T_611[54], _memRequest_bits_data_T_514[54]};
  wire [1:0]       memRequest_bits_data_lo_hi_62 = {_memRequest_bits_data_T_805[54], _memRequest_bits_data_T_708[54]};
  wire [3:0]       memRequest_bits_data_lo_62 = {memRequest_bits_data_lo_hi_62, memRequest_bits_data_lo_lo_62};
  wire [1:0]       memRequest_bits_data_hi_lo_62 = {_memRequest_bits_data_T_999[54], _memRequest_bits_data_T_902[54]};
  wire [1:0]       memRequest_bits_data_hi_hi_62 = {_memRequest_bits_data_T_1193[54], _memRequest_bits_data_T_1096[54]};
  wire [3:0]       memRequest_bits_data_hi_62 = {memRequest_bits_data_hi_hi_62, memRequest_bits_data_hi_lo_62};
  wire [1:0]       memRequest_bits_data_lo_lo_63 = {_memRequest_bits_data_T_611[55], _memRequest_bits_data_T_514[55]};
  wire [1:0]       memRequest_bits_data_lo_hi_63 = {_memRequest_bits_data_T_805[55], _memRequest_bits_data_T_708[55]};
  wire [3:0]       memRequest_bits_data_lo_63 = {memRequest_bits_data_lo_hi_63, memRequest_bits_data_lo_lo_63};
  wire [1:0]       memRequest_bits_data_hi_lo_63 = {_memRequest_bits_data_T_999[55], _memRequest_bits_data_T_902[55]};
  wire [1:0]       memRequest_bits_data_hi_hi_63 = {_memRequest_bits_data_T_1193[55], _memRequest_bits_data_T_1096[55]};
  wire [3:0]       memRequest_bits_data_hi_63 = {memRequest_bits_data_hi_hi_63, memRequest_bits_data_hi_lo_63};
  wire [1:0]       memRequest_bits_data_lo_lo_64 = {_memRequest_bits_data_T_611[56], _memRequest_bits_data_T_514[56]};
  wire [1:0]       memRequest_bits_data_lo_hi_64 = {_memRequest_bits_data_T_805[56], _memRequest_bits_data_T_708[56]};
  wire [3:0]       memRequest_bits_data_lo_64 = {memRequest_bits_data_lo_hi_64, memRequest_bits_data_lo_lo_64};
  wire [1:0]       memRequest_bits_data_hi_lo_64 = {_memRequest_bits_data_T_999[56], _memRequest_bits_data_T_902[56]};
  wire [1:0]       memRequest_bits_data_hi_hi_64 = {_memRequest_bits_data_T_1193[56], _memRequest_bits_data_T_1096[56]};
  wire [3:0]       memRequest_bits_data_hi_64 = {memRequest_bits_data_hi_hi_64, memRequest_bits_data_hi_lo_64};
  wire [1:0]       memRequest_bits_data_lo_lo_65 = {_memRequest_bits_data_T_611[57], _memRequest_bits_data_T_514[57]};
  wire [1:0]       memRequest_bits_data_lo_hi_65 = {_memRequest_bits_data_T_805[57], _memRequest_bits_data_T_708[57]};
  wire [3:0]       memRequest_bits_data_lo_65 = {memRequest_bits_data_lo_hi_65, memRequest_bits_data_lo_lo_65};
  wire [1:0]       memRequest_bits_data_hi_lo_65 = {_memRequest_bits_data_T_999[57], _memRequest_bits_data_T_902[57]};
  wire [1:0]       memRequest_bits_data_hi_hi_65 = {_memRequest_bits_data_T_1193[57], _memRequest_bits_data_T_1096[57]};
  wire [3:0]       memRequest_bits_data_hi_65 = {memRequest_bits_data_hi_hi_65, memRequest_bits_data_hi_lo_65};
  wire [1:0]       memRequest_bits_data_lo_lo_66 = {_memRequest_bits_data_T_611[58], _memRequest_bits_data_T_514[58]};
  wire [1:0]       memRequest_bits_data_lo_hi_66 = {_memRequest_bits_data_T_805[58], _memRequest_bits_data_T_708[58]};
  wire [3:0]       memRequest_bits_data_lo_66 = {memRequest_bits_data_lo_hi_66, memRequest_bits_data_lo_lo_66};
  wire [1:0]       memRequest_bits_data_hi_lo_66 = {_memRequest_bits_data_T_999[58], _memRequest_bits_data_T_902[58]};
  wire [1:0]       memRequest_bits_data_hi_hi_66 = {_memRequest_bits_data_T_1193[58], _memRequest_bits_data_T_1096[58]};
  wire [3:0]       memRequest_bits_data_hi_66 = {memRequest_bits_data_hi_hi_66, memRequest_bits_data_hi_lo_66};
  wire [1:0]       memRequest_bits_data_lo_lo_67 = {_memRequest_bits_data_T_611[59], _memRequest_bits_data_T_514[59]};
  wire [1:0]       memRequest_bits_data_lo_hi_67 = {_memRequest_bits_data_T_805[59], _memRequest_bits_data_T_708[59]};
  wire [3:0]       memRequest_bits_data_lo_67 = {memRequest_bits_data_lo_hi_67, memRequest_bits_data_lo_lo_67};
  wire [1:0]       memRequest_bits_data_hi_lo_67 = {_memRequest_bits_data_T_999[59], _memRequest_bits_data_T_902[59]};
  wire [1:0]       memRequest_bits_data_hi_hi_67 = {_memRequest_bits_data_T_1193[59], _memRequest_bits_data_T_1096[59]};
  wire [3:0]       memRequest_bits_data_hi_67 = {memRequest_bits_data_hi_hi_67, memRequest_bits_data_hi_lo_67};
  wire [1:0]       memRequest_bits_data_lo_lo_68 = {_memRequest_bits_data_T_611[60], _memRequest_bits_data_T_514[60]};
  wire [1:0]       memRequest_bits_data_lo_hi_68 = {_memRequest_bits_data_T_805[60], _memRequest_bits_data_T_708[60]};
  wire [3:0]       memRequest_bits_data_lo_68 = {memRequest_bits_data_lo_hi_68, memRequest_bits_data_lo_lo_68};
  wire [1:0]       memRequest_bits_data_hi_lo_68 = {_memRequest_bits_data_T_999[60], _memRequest_bits_data_T_902[60]};
  wire [1:0]       memRequest_bits_data_hi_hi_68 = {_memRequest_bits_data_T_1193[60], _memRequest_bits_data_T_1096[60]};
  wire [3:0]       memRequest_bits_data_hi_68 = {memRequest_bits_data_hi_hi_68, memRequest_bits_data_hi_lo_68};
  wire [1:0]       memRequest_bits_data_lo_lo_69 = {_memRequest_bits_data_T_611[61], _memRequest_bits_data_T_514[61]};
  wire [1:0]       memRequest_bits_data_lo_hi_69 = {_memRequest_bits_data_T_805[61], _memRequest_bits_data_T_708[61]};
  wire [3:0]       memRequest_bits_data_lo_69 = {memRequest_bits_data_lo_hi_69, memRequest_bits_data_lo_lo_69};
  wire [1:0]       memRequest_bits_data_hi_lo_69 = {_memRequest_bits_data_T_999[61], _memRequest_bits_data_T_902[61]};
  wire [1:0]       memRequest_bits_data_hi_hi_69 = {_memRequest_bits_data_T_1193[61], _memRequest_bits_data_T_1096[61]};
  wire [3:0]       memRequest_bits_data_hi_69 = {memRequest_bits_data_hi_hi_69, memRequest_bits_data_hi_lo_69};
  wire [1:0]       memRequest_bits_data_lo_lo_70 = {_memRequest_bits_data_T_611[62], _memRequest_bits_data_T_514[62]};
  wire [1:0]       memRequest_bits_data_lo_hi_70 = {_memRequest_bits_data_T_805[62], _memRequest_bits_data_T_708[62]};
  wire [3:0]       memRequest_bits_data_lo_70 = {memRequest_bits_data_lo_hi_70, memRequest_bits_data_lo_lo_70};
  wire [1:0]       memRequest_bits_data_hi_lo_70 = {_memRequest_bits_data_T_999[62], _memRequest_bits_data_T_902[62]};
  wire [1:0]       memRequest_bits_data_hi_hi_70 = {_memRequest_bits_data_T_1193[62], _memRequest_bits_data_T_1096[62]};
  wire [3:0]       memRequest_bits_data_hi_70 = {memRequest_bits_data_hi_hi_70, memRequest_bits_data_hi_lo_70};
  wire [1:0]       memRequest_bits_data_lo_lo_71 = {_memRequest_bits_data_T_611[63], _memRequest_bits_data_T_514[63]};
  wire [1:0]       memRequest_bits_data_lo_hi_71 = {_memRequest_bits_data_T_805[63], _memRequest_bits_data_T_708[63]};
  wire [3:0]       memRequest_bits_data_lo_71 = {memRequest_bits_data_lo_hi_71, memRequest_bits_data_lo_lo_71};
  wire [1:0]       memRequest_bits_data_hi_lo_71 = {_memRequest_bits_data_T_999[63], _memRequest_bits_data_T_902[63]};
  wire [1:0]       memRequest_bits_data_hi_hi_71 = {_memRequest_bits_data_T_1193[63], _memRequest_bits_data_T_1096[63]};
  wire [3:0]       memRequest_bits_data_hi_71 = {memRequest_bits_data_hi_hi_71, memRequest_bits_data_hi_lo_71};
  wire [1:0]       memRequest_bits_data_lo_lo_72 = {_memRequest_bits_data_T_611[64], _memRequest_bits_data_T_514[64]};
  wire [1:0]       memRequest_bits_data_lo_hi_72 = {_memRequest_bits_data_T_805[64], _memRequest_bits_data_T_708[64]};
  wire [3:0]       memRequest_bits_data_lo_72 = {memRequest_bits_data_lo_hi_72, memRequest_bits_data_lo_lo_72};
  wire [1:0]       memRequest_bits_data_hi_lo_72 = {_memRequest_bits_data_T_999[64], _memRequest_bits_data_T_902[64]};
  wire [1:0]       memRequest_bits_data_hi_hi_72 = {_memRequest_bits_data_T_1193[64], _memRequest_bits_data_T_1096[64]};
  wire [3:0]       memRequest_bits_data_hi_72 = {memRequest_bits_data_hi_hi_72, memRequest_bits_data_hi_lo_72};
  wire [1:0]       memRequest_bits_data_lo_lo_73 = {_memRequest_bits_data_T_611[65], _memRequest_bits_data_T_514[65]};
  wire [1:0]       memRequest_bits_data_lo_hi_73 = {_memRequest_bits_data_T_805[65], _memRequest_bits_data_T_708[65]};
  wire [3:0]       memRequest_bits_data_lo_73 = {memRequest_bits_data_lo_hi_73, memRequest_bits_data_lo_lo_73};
  wire [1:0]       memRequest_bits_data_hi_lo_73 = {_memRequest_bits_data_T_999[65], _memRequest_bits_data_T_902[65]};
  wire [1:0]       memRequest_bits_data_hi_hi_73 = {_memRequest_bits_data_T_1193[65], _memRequest_bits_data_T_1096[65]};
  wire [3:0]       memRequest_bits_data_hi_73 = {memRequest_bits_data_hi_hi_73, memRequest_bits_data_hi_lo_73};
  wire [1:0]       memRequest_bits_data_lo_lo_74 = {_memRequest_bits_data_T_611[66], _memRequest_bits_data_T_514[66]};
  wire [1:0]       memRequest_bits_data_lo_hi_74 = {_memRequest_bits_data_T_805[66], _memRequest_bits_data_T_708[66]};
  wire [3:0]       memRequest_bits_data_lo_74 = {memRequest_bits_data_lo_hi_74, memRequest_bits_data_lo_lo_74};
  wire [1:0]       memRequest_bits_data_hi_lo_74 = {_memRequest_bits_data_T_999[66], _memRequest_bits_data_T_902[66]};
  wire [1:0]       memRequest_bits_data_hi_hi_74 = {_memRequest_bits_data_T_1193[66], _memRequest_bits_data_T_1096[66]};
  wire [3:0]       memRequest_bits_data_hi_74 = {memRequest_bits_data_hi_hi_74, memRequest_bits_data_hi_lo_74};
  wire [1:0]       memRequest_bits_data_lo_lo_75 = {_memRequest_bits_data_T_611[67], _memRequest_bits_data_T_514[67]};
  wire [1:0]       memRequest_bits_data_lo_hi_75 = {_memRequest_bits_data_T_805[67], _memRequest_bits_data_T_708[67]};
  wire [3:0]       memRequest_bits_data_lo_75 = {memRequest_bits_data_lo_hi_75, memRequest_bits_data_lo_lo_75};
  wire [1:0]       memRequest_bits_data_hi_lo_75 = {_memRequest_bits_data_T_999[67], _memRequest_bits_data_T_902[67]};
  wire [1:0]       memRequest_bits_data_hi_hi_75 = {_memRequest_bits_data_T_1193[67], _memRequest_bits_data_T_1096[67]};
  wire [3:0]       memRequest_bits_data_hi_75 = {memRequest_bits_data_hi_hi_75, memRequest_bits_data_hi_lo_75};
  wire [1:0]       memRequest_bits_data_lo_lo_76 = {_memRequest_bits_data_T_611[68], _memRequest_bits_data_T_514[68]};
  wire [1:0]       memRequest_bits_data_lo_hi_76 = {_memRequest_bits_data_T_805[68], _memRequest_bits_data_T_708[68]};
  wire [3:0]       memRequest_bits_data_lo_76 = {memRequest_bits_data_lo_hi_76, memRequest_bits_data_lo_lo_76};
  wire [1:0]       memRequest_bits_data_hi_lo_76 = {_memRequest_bits_data_T_999[68], _memRequest_bits_data_T_902[68]};
  wire [1:0]       memRequest_bits_data_hi_hi_76 = {_memRequest_bits_data_T_1193[68], _memRequest_bits_data_T_1096[68]};
  wire [3:0]       memRequest_bits_data_hi_76 = {memRequest_bits_data_hi_hi_76, memRequest_bits_data_hi_lo_76};
  wire [1:0]       memRequest_bits_data_lo_lo_77 = {_memRequest_bits_data_T_611[69], _memRequest_bits_data_T_514[69]};
  wire [1:0]       memRequest_bits_data_lo_hi_77 = {_memRequest_bits_data_T_805[69], _memRequest_bits_data_T_708[69]};
  wire [3:0]       memRequest_bits_data_lo_77 = {memRequest_bits_data_lo_hi_77, memRequest_bits_data_lo_lo_77};
  wire [1:0]       memRequest_bits_data_hi_lo_77 = {_memRequest_bits_data_T_999[69], _memRequest_bits_data_T_902[69]};
  wire [1:0]       memRequest_bits_data_hi_hi_77 = {_memRequest_bits_data_T_1193[69], _memRequest_bits_data_T_1096[69]};
  wire [3:0]       memRequest_bits_data_hi_77 = {memRequest_bits_data_hi_hi_77, memRequest_bits_data_hi_lo_77};
  wire [1:0]       memRequest_bits_data_lo_lo_78 = {_memRequest_bits_data_T_611[70], _memRequest_bits_data_T_514[70]};
  wire [1:0]       memRequest_bits_data_lo_hi_78 = {_memRequest_bits_data_T_805[70], _memRequest_bits_data_T_708[70]};
  wire [3:0]       memRequest_bits_data_lo_78 = {memRequest_bits_data_lo_hi_78, memRequest_bits_data_lo_lo_78};
  wire [1:0]       memRequest_bits_data_hi_lo_78 = {_memRequest_bits_data_T_999[70], _memRequest_bits_data_T_902[70]};
  wire [1:0]       memRequest_bits_data_hi_hi_78 = {_memRequest_bits_data_T_1193[70], _memRequest_bits_data_T_1096[70]};
  wire [3:0]       memRequest_bits_data_hi_78 = {memRequest_bits_data_hi_hi_78, memRequest_bits_data_hi_lo_78};
  wire [1:0]       memRequest_bits_data_lo_lo_79 = {_memRequest_bits_data_T_611[71], _memRequest_bits_data_T_514[71]};
  wire [1:0]       memRequest_bits_data_lo_hi_79 = {_memRequest_bits_data_T_805[71], _memRequest_bits_data_T_708[71]};
  wire [3:0]       memRequest_bits_data_lo_79 = {memRequest_bits_data_lo_hi_79, memRequest_bits_data_lo_lo_79};
  wire [1:0]       memRequest_bits_data_hi_lo_79 = {_memRequest_bits_data_T_999[71], _memRequest_bits_data_T_902[71]};
  wire [1:0]       memRequest_bits_data_hi_hi_79 = {_memRequest_bits_data_T_1193[71], _memRequest_bits_data_T_1096[71]};
  wire [3:0]       memRequest_bits_data_hi_79 = {memRequest_bits_data_hi_hi_79, memRequest_bits_data_hi_lo_79};
  wire [1:0]       memRequest_bits_data_lo_lo_80 = {_memRequest_bits_data_T_611[72], _memRequest_bits_data_T_514[72]};
  wire [1:0]       memRequest_bits_data_lo_hi_80 = {_memRequest_bits_data_T_805[72], _memRequest_bits_data_T_708[72]};
  wire [3:0]       memRequest_bits_data_lo_80 = {memRequest_bits_data_lo_hi_80, memRequest_bits_data_lo_lo_80};
  wire [1:0]       memRequest_bits_data_hi_lo_80 = {_memRequest_bits_data_T_999[72], _memRequest_bits_data_T_902[72]};
  wire [1:0]       memRequest_bits_data_hi_hi_80 = {_memRequest_bits_data_T_1193[72], _memRequest_bits_data_T_1096[72]};
  wire [3:0]       memRequest_bits_data_hi_80 = {memRequest_bits_data_hi_hi_80, memRequest_bits_data_hi_lo_80};
  wire [1:0]       memRequest_bits_data_lo_lo_81 = {_memRequest_bits_data_T_611[73], _memRequest_bits_data_T_514[73]};
  wire [1:0]       memRequest_bits_data_lo_hi_81 = {_memRequest_bits_data_T_805[73], _memRequest_bits_data_T_708[73]};
  wire [3:0]       memRequest_bits_data_lo_81 = {memRequest_bits_data_lo_hi_81, memRequest_bits_data_lo_lo_81};
  wire [1:0]       memRequest_bits_data_hi_lo_81 = {_memRequest_bits_data_T_999[73], _memRequest_bits_data_T_902[73]};
  wire [1:0]       memRequest_bits_data_hi_hi_81 = {_memRequest_bits_data_T_1193[73], _memRequest_bits_data_T_1096[73]};
  wire [3:0]       memRequest_bits_data_hi_81 = {memRequest_bits_data_hi_hi_81, memRequest_bits_data_hi_lo_81};
  wire [1:0]       memRequest_bits_data_lo_lo_82 = {_memRequest_bits_data_T_611[74], _memRequest_bits_data_T_514[74]};
  wire [1:0]       memRequest_bits_data_lo_hi_82 = {_memRequest_bits_data_T_805[74], _memRequest_bits_data_T_708[74]};
  wire [3:0]       memRequest_bits_data_lo_82 = {memRequest_bits_data_lo_hi_82, memRequest_bits_data_lo_lo_82};
  wire [1:0]       memRequest_bits_data_hi_lo_82 = {_memRequest_bits_data_T_999[74], _memRequest_bits_data_T_902[74]};
  wire [1:0]       memRequest_bits_data_hi_hi_82 = {_memRequest_bits_data_T_1193[74], _memRequest_bits_data_T_1096[74]};
  wire [3:0]       memRequest_bits_data_hi_82 = {memRequest_bits_data_hi_hi_82, memRequest_bits_data_hi_lo_82};
  wire [1:0]       memRequest_bits_data_lo_lo_83 = {_memRequest_bits_data_T_611[75], _memRequest_bits_data_T_514[75]};
  wire [1:0]       memRequest_bits_data_lo_hi_83 = {_memRequest_bits_data_T_805[75], _memRequest_bits_data_T_708[75]};
  wire [3:0]       memRequest_bits_data_lo_83 = {memRequest_bits_data_lo_hi_83, memRequest_bits_data_lo_lo_83};
  wire [1:0]       memRequest_bits_data_hi_lo_83 = {_memRequest_bits_data_T_999[75], _memRequest_bits_data_T_902[75]};
  wire [1:0]       memRequest_bits_data_hi_hi_83 = {_memRequest_bits_data_T_1193[75], _memRequest_bits_data_T_1096[75]};
  wire [3:0]       memRequest_bits_data_hi_83 = {memRequest_bits_data_hi_hi_83, memRequest_bits_data_hi_lo_83};
  wire [1:0]       memRequest_bits_data_lo_lo_84 = {_memRequest_bits_data_T_611[76], _memRequest_bits_data_T_514[76]};
  wire [1:0]       memRequest_bits_data_lo_hi_84 = {_memRequest_bits_data_T_805[76], _memRequest_bits_data_T_708[76]};
  wire [3:0]       memRequest_bits_data_lo_84 = {memRequest_bits_data_lo_hi_84, memRequest_bits_data_lo_lo_84};
  wire [1:0]       memRequest_bits_data_hi_lo_84 = {_memRequest_bits_data_T_999[76], _memRequest_bits_data_T_902[76]};
  wire [1:0]       memRequest_bits_data_hi_hi_84 = {_memRequest_bits_data_T_1193[76], _memRequest_bits_data_T_1096[76]};
  wire [3:0]       memRequest_bits_data_hi_84 = {memRequest_bits_data_hi_hi_84, memRequest_bits_data_hi_lo_84};
  wire [1:0]       memRequest_bits_data_lo_lo_85 = {_memRequest_bits_data_T_611[77], _memRequest_bits_data_T_514[77]};
  wire [1:0]       memRequest_bits_data_lo_hi_85 = {_memRequest_bits_data_T_805[77], _memRequest_bits_data_T_708[77]};
  wire [3:0]       memRequest_bits_data_lo_85 = {memRequest_bits_data_lo_hi_85, memRequest_bits_data_lo_lo_85};
  wire [1:0]       memRequest_bits_data_hi_lo_85 = {_memRequest_bits_data_T_999[77], _memRequest_bits_data_T_902[77]};
  wire [1:0]       memRequest_bits_data_hi_hi_85 = {_memRequest_bits_data_T_1193[77], _memRequest_bits_data_T_1096[77]};
  wire [3:0]       memRequest_bits_data_hi_85 = {memRequest_bits_data_hi_hi_85, memRequest_bits_data_hi_lo_85};
  wire [1:0]       memRequest_bits_data_lo_lo_86 = {_memRequest_bits_data_T_611[78], _memRequest_bits_data_T_514[78]};
  wire [1:0]       memRequest_bits_data_lo_hi_86 = {_memRequest_bits_data_T_805[78], _memRequest_bits_data_T_708[78]};
  wire [3:0]       memRequest_bits_data_lo_86 = {memRequest_bits_data_lo_hi_86, memRequest_bits_data_lo_lo_86};
  wire [1:0]       memRequest_bits_data_hi_lo_86 = {_memRequest_bits_data_T_999[78], _memRequest_bits_data_T_902[78]};
  wire [1:0]       memRequest_bits_data_hi_hi_86 = {_memRequest_bits_data_T_1193[78], _memRequest_bits_data_T_1096[78]};
  wire [3:0]       memRequest_bits_data_hi_86 = {memRequest_bits_data_hi_hi_86, memRequest_bits_data_hi_lo_86};
  wire [1:0]       memRequest_bits_data_lo_lo_87 = {_memRequest_bits_data_T_611[79], _memRequest_bits_data_T_514[79]};
  wire [1:0]       memRequest_bits_data_lo_hi_87 = {_memRequest_bits_data_T_805[79], _memRequest_bits_data_T_708[79]};
  wire [3:0]       memRequest_bits_data_lo_87 = {memRequest_bits_data_lo_hi_87, memRequest_bits_data_lo_lo_87};
  wire [1:0]       memRequest_bits_data_hi_lo_87 = {_memRequest_bits_data_T_999[79], _memRequest_bits_data_T_902[79]};
  wire [1:0]       memRequest_bits_data_hi_hi_87 = {_memRequest_bits_data_T_1193[79], _memRequest_bits_data_T_1096[79]};
  wire [3:0]       memRequest_bits_data_hi_87 = {memRequest_bits_data_hi_hi_87, memRequest_bits_data_hi_lo_87};
  wire [1:0]       memRequest_bits_data_lo_lo_88 = {_memRequest_bits_data_T_611[80], _memRequest_bits_data_T_514[80]};
  wire [1:0]       memRequest_bits_data_lo_hi_88 = {_memRequest_bits_data_T_805[80], _memRequest_bits_data_T_708[80]};
  wire [3:0]       memRequest_bits_data_lo_88 = {memRequest_bits_data_lo_hi_88, memRequest_bits_data_lo_lo_88};
  wire [1:0]       memRequest_bits_data_hi_lo_88 = {_memRequest_bits_data_T_999[80], _memRequest_bits_data_T_902[80]};
  wire [1:0]       memRequest_bits_data_hi_hi_88 = {_memRequest_bits_data_T_1193[80], _memRequest_bits_data_T_1096[80]};
  wire [3:0]       memRequest_bits_data_hi_88 = {memRequest_bits_data_hi_hi_88, memRequest_bits_data_hi_lo_88};
  wire [1:0]       memRequest_bits_data_lo_lo_89 = {_memRequest_bits_data_T_611[81], _memRequest_bits_data_T_514[81]};
  wire [1:0]       memRequest_bits_data_lo_hi_89 = {_memRequest_bits_data_T_805[81], _memRequest_bits_data_T_708[81]};
  wire [3:0]       memRequest_bits_data_lo_89 = {memRequest_bits_data_lo_hi_89, memRequest_bits_data_lo_lo_89};
  wire [1:0]       memRequest_bits_data_hi_lo_89 = {_memRequest_bits_data_T_999[81], _memRequest_bits_data_T_902[81]};
  wire [1:0]       memRequest_bits_data_hi_hi_89 = {_memRequest_bits_data_T_1193[81], _memRequest_bits_data_T_1096[81]};
  wire [3:0]       memRequest_bits_data_hi_89 = {memRequest_bits_data_hi_hi_89, memRequest_bits_data_hi_lo_89};
  wire [1:0]       memRequest_bits_data_lo_lo_90 = {_memRequest_bits_data_T_611[82], _memRequest_bits_data_T_514[82]};
  wire [1:0]       memRequest_bits_data_lo_hi_90 = {_memRequest_bits_data_T_805[82], _memRequest_bits_data_T_708[82]};
  wire [3:0]       memRequest_bits_data_lo_90 = {memRequest_bits_data_lo_hi_90, memRequest_bits_data_lo_lo_90};
  wire [1:0]       memRequest_bits_data_hi_lo_90 = {_memRequest_bits_data_T_999[82], _memRequest_bits_data_T_902[82]};
  wire [1:0]       memRequest_bits_data_hi_hi_90 = {_memRequest_bits_data_T_1193[82], _memRequest_bits_data_T_1096[82]};
  wire [3:0]       memRequest_bits_data_hi_90 = {memRequest_bits_data_hi_hi_90, memRequest_bits_data_hi_lo_90};
  wire [1:0]       memRequest_bits_data_lo_lo_91 = {_memRequest_bits_data_T_611[83], _memRequest_bits_data_T_514[83]};
  wire [1:0]       memRequest_bits_data_lo_hi_91 = {_memRequest_bits_data_T_805[83], _memRequest_bits_data_T_708[83]};
  wire [3:0]       memRequest_bits_data_lo_91 = {memRequest_bits_data_lo_hi_91, memRequest_bits_data_lo_lo_91};
  wire [1:0]       memRequest_bits_data_hi_lo_91 = {_memRequest_bits_data_T_999[83], _memRequest_bits_data_T_902[83]};
  wire [1:0]       memRequest_bits_data_hi_hi_91 = {_memRequest_bits_data_T_1193[83], _memRequest_bits_data_T_1096[83]};
  wire [3:0]       memRequest_bits_data_hi_91 = {memRequest_bits_data_hi_hi_91, memRequest_bits_data_hi_lo_91};
  wire [1:0]       memRequest_bits_data_lo_lo_92 = {_memRequest_bits_data_T_611[84], _memRequest_bits_data_T_514[84]};
  wire [1:0]       memRequest_bits_data_lo_hi_92 = {_memRequest_bits_data_T_805[84], _memRequest_bits_data_T_708[84]};
  wire [3:0]       memRequest_bits_data_lo_92 = {memRequest_bits_data_lo_hi_92, memRequest_bits_data_lo_lo_92};
  wire [1:0]       memRequest_bits_data_hi_lo_92 = {_memRequest_bits_data_T_999[84], _memRequest_bits_data_T_902[84]};
  wire [1:0]       memRequest_bits_data_hi_hi_92 = {_memRequest_bits_data_T_1193[84], _memRequest_bits_data_T_1096[84]};
  wire [3:0]       memRequest_bits_data_hi_92 = {memRequest_bits_data_hi_hi_92, memRequest_bits_data_hi_lo_92};
  wire [1:0]       memRequest_bits_data_lo_lo_93 = {_memRequest_bits_data_T_611[85], _memRequest_bits_data_T_514[85]};
  wire [1:0]       memRequest_bits_data_lo_hi_93 = {_memRequest_bits_data_T_805[85], _memRequest_bits_data_T_708[85]};
  wire [3:0]       memRequest_bits_data_lo_93 = {memRequest_bits_data_lo_hi_93, memRequest_bits_data_lo_lo_93};
  wire [1:0]       memRequest_bits_data_hi_lo_93 = {_memRequest_bits_data_T_999[85], _memRequest_bits_data_T_902[85]};
  wire [1:0]       memRequest_bits_data_hi_hi_93 = {_memRequest_bits_data_T_1193[85], _memRequest_bits_data_T_1096[85]};
  wire [3:0]       memRequest_bits_data_hi_93 = {memRequest_bits_data_hi_hi_93, memRequest_bits_data_hi_lo_93};
  wire [1:0]       memRequest_bits_data_lo_lo_94 = {_memRequest_bits_data_T_611[86], _memRequest_bits_data_T_514[86]};
  wire [1:0]       memRequest_bits_data_lo_hi_94 = {_memRequest_bits_data_T_805[86], _memRequest_bits_data_T_708[86]};
  wire [3:0]       memRequest_bits_data_lo_94 = {memRequest_bits_data_lo_hi_94, memRequest_bits_data_lo_lo_94};
  wire [1:0]       memRequest_bits_data_hi_lo_94 = {_memRequest_bits_data_T_999[86], _memRequest_bits_data_T_902[86]};
  wire [1:0]       memRequest_bits_data_hi_hi_94 = {_memRequest_bits_data_T_1193[86], _memRequest_bits_data_T_1096[86]};
  wire [3:0]       memRequest_bits_data_hi_94 = {memRequest_bits_data_hi_hi_94, memRequest_bits_data_hi_lo_94};
  wire [1:0]       memRequest_bits_data_lo_lo_95 = {_memRequest_bits_data_T_611[87], _memRequest_bits_data_T_514[87]};
  wire [1:0]       memRequest_bits_data_lo_hi_95 = {_memRequest_bits_data_T_805[87], _memRequest_bits_data_T_708[87]};
  wire [3:0]       memRequest_bits_data_lo_95 = {memRequest_bits_data_lo_hi_95, memRequest_bits_data_lo_lo_95};
  wire [1:0]       memRequest_bits_data_hi_lo_95 = {_memRequest_bits_data_T_999[87], _memRequest_bits_data_T_902[87]};
  wire [1:0]       memRequest_bits_data_hi_hi_95 = {_memRequest_bits_data_T_1193[87], _memRequest_bits_data_T_1096[87]};
  wire [3:0]       memRequest_bits_data_hi_95 = {memRequest_bits_data_hi_hi_95, memRequest_bits_data_hi_lo_95};
  wire [1:0]       memRequest_bits_data_lo_lo_96 = {_memRequest_bits_data_T_611[88], _memRequest_bits_data_T_514[88]};
  wire [1:0]       memRequest_bits_data_lo_hi_96 = {_memRequest_bits_data_T_805[88], _memRequest_bits_data_T_708[88]};
  wire [3:0]       memRequest_bits_data_lo_96 = {memRequest_bits_data_lo_hi_96, memRequest_bits_data_lo_lo_96};
  wire [1:0]       memRequest_bits_data_hi_lo_96 = {_memRequest_bits_data_T_999[88], _memRequest_bits_data_T_902[88]};
  wire [1:0]       memRequest_bits_data_hi_hi_96 = {_memRequest_bits_data_T_1193[88], _memRequest_bits_data_T_1096[88]};
  wire [3:0]       memRequest_bits_data_hi_96 = {memRequest_bits_data_hi_hi_96, memRequest_bits_data_hi_lo_96};
  wire [1:0]       memRequest_bits_data_lo_lo_97 = {_memRequest_bits_data_T_611[89], _memRequest_bits_data_T_514[89]};
  wire [1:0]       memRequest_bits_data_lo_hi_97 = {_memRequest_bits_data_T_805[89], _memRequest_bits_data_T_708[89]};
  wire [3:0]       memRequest_bits_data_lo_97 = {memRequest_bits_data_lo_hi_97, memRequest_bits_data_lo_lo_97};
  wire [1:0]       memRequest_bits_data_hi_lo_97 = {_memRequest_bits_data_T_999[89], _memRequest_bits_data_T_902[89]};
  wire [1:0]       memRequest_bits_data_hi_hi_97 = {_memRequest_bits_data_T_1193[89], _memRequest_bits_data_T_1096[89]};
  wire [3:0]       memRequest_bits_data_hi_97 = {memRequest_bits_data_hi_hi_97, memRequest_bits_data_hi_lo_97};
  wire [1:0]       memRequest_bits_data_lo_lo_98 = {_memRequest_bits_data_T_611[90], _memRequest_bits_data_T_514[90]};
  wire [1:0]       memRequest_bits_data_lo_hi_98 = {_memRequest_bits_data_T_805[90], _memRequest_bits_data_T_708[90]};
  wire [3:0]       memRequest_bits_data_lo_98 = {memRequest_bits_data_lo_hi_98, memRequest_bits_data_lo_lo_98};
  wire [1:0]       memRequest_bits_data_hi_lo_98 = {_memRequest_bits_data_T_999[90], _memRequest_bits_data_T_902[90]};
  wire [1:0]       memRequest_bits_data_hi_hi_98 = {_memRequest_bits_data_T_1193[90], _memRequest_bits_data_T_1096[90]};
  wire [3:0]       memRequest_bits_data_hi_98 = {memRequest_bits_data_hi_hi_98, memRequest_bits_data_hi_lo_98};
  wire [1:0]       memRequest_bits_data_lo_lo_99 = {_memRequest_bits_data_T_611[91], _memRequest_bits_data_T_514[91]};
  wire [1:0]       memRequest_bits_data_lo_hi_99 = {_memRequest_bits_data_T_805[91], _memRequest_bits_data_T_708[91]};
  wire [3:0]       memRequest_bits_data_lo_99 = {memRequest_bits_data_lo_hi_99, memRequest_bits_data_lo_lo_99};
  wire [1:0]       memRequest_bits_data_hi_lo_99 = {_memRequest_bits_data_T_999[91], _memRequest_bits_data_T_902[91]};
  wire [1:0]       memRequest_bits_data_hi_hi_99 = {_memRequest_bits_data_T_1193[91], _memRequest_bits_data_T_1096[91]};
  wire [3:0]       memRequest_bits_data_hi_99 = {memRequest_bits_data_hi_hi_99, memRequest_bits_data_hi_lo_99};
  wire [1:0]       memRequest_bits_data_lo_lo_100 = {_memRequest_bits_data_T_611[92], _memRequest_bits_data_T_514[92]};
  wire [1:0]       memRequest_bits_data_lo_hi_100 = {_memRequest_bits_data_T_805[92], _memRequest_bits_data_T_708[92]};
  wire [3:0]       memRequest_bits_data_lo_100 = {memRequest_bits_data_lo_hi_100, memRequest_bits_data_lo_lo_100};
  wire [1:0]       memRequest_bits_data_hi_lo_100 = {_memRequest_bits_data_T_999[92], _memRequest_bits_data_T_902[92]};
  wire [1:0]       memRequest_bits_data_hi_hi_100 = {_memRequest_bits_data_T_1193[92], _memRequest_bits_data_T_1096[92]};
  wire [3:0]       memRequest_bits_data_hi_100 = {memRequest_bits_data_hi_hi_100, memRequest_bits_data_hi_lo_100};
  wire [1:0]       memRequest_bits_data_lo_lo_101 = {_memRequest_bits_data_T_611[93], _memRequest_bits_data_T_514[93]};
  wire [1:0]       memRequest_bits_data_lo_hi_101 = {_memRequest_bits_data_T_805[93], _memRequest_bits_data_T_708[93]};
  wire [3:0]       memRequest_bits_data_lo_101 = {memRequest_bits_data_lo_hi_101, memRequest_bits_data_lo_lo_101};
  wire [1:0]       memRequest_bits_data_hi_lo_101 = {_memRequest_bits_data_T_999[93], _memRequest_bits_data_T_902[93]};
  wire [1:0]       memRequest_bits_data_hi_hi_101 = {_memRequest_bits_data_T_1193[93], _memRequest_bits_data_T_1096[93]};
  wire [3:0]       memRequest_bits_data_hi_101 = {memRequest_bits_data_hi_hi_101, memRequest_bits_data_hi_lo_101};
  wire [1:0]       memRequest_bits_data_lo_lo_102 = {_memRequest_bits_data_T_611[94], _memRequest_bits_data_T_514[94]};
  wire [1:0]       memRequest_bits_data_lo_hi_102 = {_memRequest_bits_data_T_805[94], _memRequest_bits_data_T_708[94]};
  wire [3:0]       memRequest_bits_data_lo_102 = {memRequest_bits_data_lo_hi_102, memRequest_bits_data_lo_lo_102};
  wire [1:0]       memRequest_bits_data_hi_lo_102 = {_memRequest_bits_data_T_999[94], _memRequest_bits_data_T_902[94]};
  wire [1:0]       memRequest_bits_data_hi_hi_102 = {_memRequest_bits_data_T_1193[94], _memRequest_bits_data_T_1096[94]};
  wire [3:0]       memRequest_bits_data_hi_102 = {memRequest_bits_data_hi_hi_102, memRequest_bits_data_hi_lo_102};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_9, memRequest_bits_data_lo_9, memRequest_bits_data_hi_8, memRequest_bits_data_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_12, memRequest_bits_data_lo_12, memRequest_bits_data_hi_11, memRequest_bits_data_lo_11};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_10, memRequest_bits_data_lo_10};
  wire [39:0]      memRequest_bits_data_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_15, memRequest_bits_data_lo_15, memRequest_bits_data_hi_14, memRequest_bits_data_lo_14};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_13, memRequest_bits_data_lo_13};
  wire [15:0]      memRequest_bits_data_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_18, memRequest_bits_data_lo_18, memRequest_bits_data_hi_17, memRequest_bits_data_lo_17};
  wire [23:0]      memRequest_bits_data_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_16, memRequest_bits_data_lo_16};
  wire [47:0]      memRequest_bits_data_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_lo_hi_lo_8};
  wire [87:0]      memRequest_bits_data_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_21, memRequest_bits_data_lo_21, memRequest_bits_data_hi_20, memRequest_bits_data_lo_20};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_19, memRequest_bits_data_lo_19};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_24, memRequest_bits_data_lo_24, memRequest_bits_data_hi_23, memRequest_bits_data_lo_23};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_22, memRequest_bits_data_lo_22};
  wire [47:0]      memRequest_bits_data_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_8, memRequest_bits_data_lo_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_27, memRequest_bits_data_lo_27, memRequest_bits_data_hi_26, memRequest_bits_data_lo_26};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_25, memRequest_bits_data_lo_25};
  wire [15:0]      memRequest_bits_data_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_30, memRequest_bits_data_lo_30, memRequest_bits_data_hi_29, memRequest_bits_data_lo_29};
  wire [23:0]      memRequest_bits_data_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_28, memRequest_bits_data_lo_28};
  wire [47:0]      memRequest_bits_data_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_8, memRequest_bits_data_lo_lo_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_8};
  wire [183:0]     memRequest_bits_data_lo_lo_103 = {memRequest_bits_data_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_33, memRequest_bits_data_lo_33, memRequest_bits_data_hi_32, memRequest_bits_data_lo_32};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_31, memRequest_bits_data_lo_31};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_36, memRequest_bits_data_lo_36, memRequest_bits_data_hi_35, memRequest_bits_data_lo_35};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_34, memRequest_bits_data_lo_34};
  wire [47:0]      memRequest_bits_data_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_39, memRequest_bits_data_lo_39, memRequest_bits_data_hi_38, memRequest_bits_data_lo_38};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_37, memRequest_bits_data_lo_37};
  wire [15:0]      memRequest_bits_data_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_42, memRequest_bits_data_lo_42, memRequest_bits_data_hi_41, memRequest_bits_data_lo_41};
  wire [23:0]      memRequest_bits_data_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_40, memRequest_bits_data_lo_40};
  wire [47:0]      memRequest_bits_data_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_45, memRequest_bits_data_lo_45, memRequest_bits_data_hi_44, memRequest_bits_data_lo_44};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_43, memRequest_bits_data_lo_43};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_48, memRequest_bits_data_lo_48, memRequest_bits_data_hi_47, memRequest_bits_data_lo_47};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_46, memRequest_bits_data_lo_46};
  wire [47:0]      memRequest_bits_data_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_8, memRequest_bits_data_lo_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_51, memRequest_bits_data_lo_51, memRequest_bits_data_hi_50, memRequest_bits_data_lo_50};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_49, memRequest_bits_data_lo_49};
  wire [15:0]      memRequest_bits_data_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_54, memRequest_bits_data_lo_54, memRequest_bits_data_hi_53, memRequest_bits_data_lo_53};
  wire [23:0]      memRequest_bits_data_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_52, memRequest_bits_data_lo_52};
  wire [47:0]      memRequest_bits_data_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_8};
  wire [191:0]     memRequest_bits_data_lo_hi_103 = {memRequest_bits_data_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_8};
  wire [375:0]     memRequest_bits_data_lo_103 = {memRequest_bits_data_lo_hi_103, memRequest_bits_data_lo_lo_103};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_57, memRequest_bits_data_lo_57, memRequest_bits_data_hi_56, memRequest_bits_data_lo_56};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_55, memRequest_bits_data_lo_55};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_60, memRequest_bits_data_lo_60, memRequest_bits_data_hi_59, memRequest_bits_data_lo_59};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_58, memRequest_bits_data_lo_58};
  wire [47:0]      memRequest_bits_data_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_63, memRequest_bits_data_lo_63, memRequest_bits_data_hi_62, memRequest_bits_data_lo_62};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_61, memRequest_bits_data_lo_61};
  wire [15:0]      memRequest_bits_data_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_66, memRequest_bits_data_lo_66, memRequest_bits_data_hi_65, memRequest_bits_data_lo_65};
  wire [23:0]      memRequest_bits_data_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_64, memRequest_bits_data_lo_64};
  wire [47:0]      memRequest_bits_data_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_8, memRequest_bits_data_hi_lo_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_69, memRequest_bits_data_lo_69, memRequest_bits_data_hi_68, memRequest_bits_data_lo_68};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_67, memRequest_bits_data_lo_67};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_72, memRequest_bits_data_lo_72, memRequest_bits_data_hi_71, memRequest_bits_data_lo_71};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_70, memRequest_bits_data_lo_70};
  wire [47:0]      memRequest_bits_data_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_8, memRequest_bits_data_hi_lo_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_75, memRequest_bits_data_lo_75, memRequest_bits_data_hi_74, memRequest_bits_data_lo_74};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_73, memRequest_bits_data_lo_73};
  wire [15:0]      memRequest_bits_data_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_78, memRequest_bits_data_lo_78, memRequest_bits_data_hi_77, memRequest_bits_data_lo_77};
  wire [23:0]      memRequest_bits_data_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_76, memRequest_bits_data_lo_76};
  wire [47:0]      memRequest_bits_data_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_8, memRequest_bits_data_hi_lo_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_8};
  wire [191:0]     memRequest_bits_data_hi_lo_103 = {memRequest_bits_data_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_81, memRequest_bits_data_lo_81, memRequest_bits_data_hi_80, memRequest_bits_data_lo_80};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_79, memRequest_bits_data_lo_79};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_84, memRequest_bits_data_lo_84, memRequest_bits_data_hi_83, memRequest_bits_data_lo_83};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_82, memRequest_bits_data_lo_82};
  wire [47:0]      memRequest_bits_data_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_87, memRequest_bits_data_lo_87, memRequest_bits_data_hi_86, memRequest_bits_data_lo_86};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_85, memRequest_bits_data_lo_85};
  wire [15:0]      memRequest_bits_data_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_90, memRequest_bits_data_lo_90, memRequest_bits_data_hi_89, memRequest_bits_data_lo_89};
  wire [23:0]      memRequest_bits_data_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_88, memRequest_bits_data_lo_88};
  wire [47:0]      memRequest_bits_data_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_8, memRequest_bits_data_hi_hi_lo_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_93, memRequest_bits_data_lo_93, memRequest_bits_data_hi_92, memRequest_bits_data_lo_92};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_91, memRequest_bits_data_lo_91};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_96, memRequest_bits_data_lo_96, memRequest_bits_data_hi_95, memRequest_bits_data_lo_95};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_94, memRequest_bits_data_lo_94};
  wire [47:0]      memRequest_bits_data_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_hi_lo_lo_8};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_99, memRequest_bits_data_lo_99, memRequest_bits_data_hi_98, memRequest_bits_data_lo_98};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_97, memRequest_bits_data_lo_97};
  wire [15:0]      memRequest_bits_data_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_102, memRequest_bits_data_lo_102, memRequest_bits_data_hi_101, memRequest_bits_data_lo_101};
  wire [23:0]      memRequest_bits_data_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_100, memRequest_bits_data_lo_100};
  wire [47:0]      memRequest_bits_data_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_hi_lo_8};
  wire [95:0]      memRequest_bits_data_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_8};
  wire [191:0]     memRequest_bits_data_hi_hi_103 = {memRequest_bits_data_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_8};
  wire [383:0]     memRequest_bits_data_hi_103 = {memRequest_bits_data_hi_hi_103, memRequest_bits_data_hi_lo_103};
  wire [255:0]     memRequest_bits_data_0 = {memRequest_bits_data_hi_103[135:0], memRequest_bits_data_lo_103[375:256]};
  wire [31:0]      selectMaskForTail = bufferValid ? _GEN_287 : 32'h0;
  wire [94:0]      _memRequest_bits_mask_T_1 = {31'h0, selectMaskForTail, maskTemp} << _GEN_288;
  wire [31:0]      memRequest_bits_mask_0 = _memRequest_bits_mask_T_1[63:32];
  assign alignedDequeueAddress = {lsuRequestReg_rs1Data[31:5] + {20'h0, bufferBaseCacheLineIndex}, 5'h0};
  wire [31:0]      memRequest_bits_address_0 = alignedDequeueAddress;
  wire [31:0]      addressQueue_enq_bits = alignedDequeueAddress;
  assign addressQueueFree = addressQueue_enq_ready;
  wire             addressQueue_deq_valid;
  assign addressQueue_deq_valid = ~_addressQueue_fifo_empty;
  assign addressQueue_enq_ready = ~_addressQueue_fifo_full;
  wire             _status_idle_output = ~bufferValid & ~readStageValid & readQueueClear & ~bufferFull & ~addressQueue_deq_valid;
  reg              idleNext;
  wire [31:0]      addressQueue_deq_bits;
  always @(posedge clock) begin
    if (reset) begin
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 12'h0;
      csrInterfaceReg_vStart <= 12'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      requestFireNext <= 1'h0;
      dataEEW <= 2'h0;
      maskReg <= 32'h0;
      needAmend <= 1'h0;
      lastMaskAmendReg <= 31'h0;
      maskGroupCounter <= 6'h0;
      maskCounterInGroup <= 2'h0;
      isLastMaskGroup <= 1'h0;
      accessData_0 <= 256'h0;
      accessData_1 <= 256'h0;
      accessData_2 <= 256'h0;
      accessData_3 <= 256'h0;
      accessData_4 <= 256'h0;
      accessData_5 <= 256'h0;
      accessData_6 <= 256'h0;
      accessData_7 <= 256'h0;
      accessPtr <= 3'h0;
      dataGroup <= 6'h0;
      dataBuffer_0 <= 256'h0;
      dataBuffer_1 <= 256'h0;
      dataBuffer_2 <= 256'h0;
      dataBuffer_3 <= 256'h0;
      dataBuffer_4 <= 256'h0;
      dataBuffer_5 <= 256'h0;
      dataBuffer_6 <= 256'h0;
      dataBuffer_7 <= 256'h0;
      bufferBaseCacheLineIndex <= 7'h0;
      cacheLineIndexInBuffer <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      lastWriteVrfIndexReg <= 14'h0;
      lastCacheNeedPush <= 1'h0;
      cacheLineNumberReg <= 14'h0;
      lastDataGroupReg <= 10'h0;
      hazardCheck <= 1'h0;
      readStageValid_segPtr <= 3'h0;
      readStageValid_readCount <= 6'h0;
      readStageValid_stageValid <= 1'h0;
      readStageValid_readCounter <= 4'h0;
      readStageValid_segPtr_1 <= 3'h0;
      readStageValid_readCount_1 <= 6'h0;
      readStageValid_stageValid_1 <= 1'h0;
      readStageValid_readCounter_1 <= 4'h0;
      readStageValid_segPtr_2 <= 3'h0;
      readStageValid_readCount_2 <= 6'h0;
      readStageValid_stageValid_2 <= 1'h0;
      readStageValid_readCounter_2 <= 4'h0;
      readStageValid_segPtr_3 <= 3'h0;
      readStageValid_readCount_3 <= 6'h0;
      readStageValid_stageValid_3 <= 1'h0;
      readStageValid_readCounter_3 <= 4'h0;
      readStageValid_segPtr_4 <= 3'h0;
      readStageValid_readCount_4 <= 6'h0;
      readStageValid_stageValid_4 <= 1'h0;
      readStageValid_readCounter_4 <= 4'h0;
      readStageValid_segPtr_5 <= 3'h0;
      readStageValid_readCount_5 <= 6'h0;
      readStageValid_stageValid_5 <= 1'h0;
      readStageValid_readCounter_5 <= 4'h0;
      readStageValid_segPtr_6 <= 3'h0;
      readStageValid_readCount_6 <= 6'h0;
      readStageValid_stageValid_6 <= 1'h0;
      readStageValid_readCounter_6 <= 4'h0;
      readStageValid_segPtr_7 <= 3'h0;
      readStageValid_readCount_7 <= 6'h0;
      readStageValid_stageValid_7 <= 1'h0;
      readStageValid_readCounter_7 <= 4'h0;
      bufferFull <= 1'h0;
      bufferValid <= 1'h0;
      maskForBufferData_0 <= 32'h0;
      maskForBufferData_1 <= 32'h0;
      maskForBufferData_2 <= 32'h0;
      maskForBufferData_3 <= 32'h0;
      maskForBufferData_4 <= 32'h0;
      maskForBufferData_5 <= 32'h0;
      maskForBufferData_6 <= 32'h0;
      maskForBufferData_7 <= 32'h0;
      lastDataGroupInDataBuffer <= 1'h0;
      cacheLineTemp <= 256'h0;
      maskTemp <= 32'h0;
      canSendTail <= 1'h0;
      idleNext <= 1'h1;
    end
    else begin
      if (lsuRequest_valid) begin
        lsuRequestReg_instructionInformation_nf <= nfCorrection;
        lsuRequestReg_instructionInformation_mew <= ~invalidInstruction & lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataEEW <= lsuRequest_bits_instructionInformation_eew;
        needAmend <= |(csrInterface_vl[4:0]);
        lastMaskAmendReg <= lastMaskAmend;
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
        lastWriteVrfIndexReg <= lastWriteVrfIndex;
        lastCacheNeedPush <= lastCacheLineIndex == lastWriteVrfIndex;
        cacheLineNumberReg <= lastCacheLineIndex;
        lastDataGroupReg <= lastDataGroupForInstruction;
      end
      requestFireNext <= lsuRequest_valid;
      if (_maskSelect_valid_output | lsuRequest_valid) begin
        maskReg <= maskAmend;
        isLastMaskGroup <= lsuRequest_valid ? csrInterface_vl[11:5] == 7'h0 : {1'h0, _maskSelect_bits_output} == csrInterfaceReg_vl[11:5];
      end
      if (_GEN_284 & (_GEN_285 | lsuRequest_valid))
        maskGroupCounter <= _maskSelect_bits_output;
      if (_GEN_284) begin
        maskCounterInGroup <= isLastDataGroup | lsuRequest_valid ? 2'h0 : nextMaskCount;
        dataGroup <= nextDataGroup;
      end
      if (accessBufferDequeueFire | accessBufferEnqueueFire | requestFireNext) begin
        accessData_0 <= accessDataUpdate_0;
        accessData_1 <= accessDataUpdate_1;
        accessData_2 <= accessDataUpdate_2;
        accessData_3 <= accessDataUpdate_3;
        accessData_4 <= accessDataUpdate_4;
        accessData_5 <= accessDataUpdate_5;
        accessData_6 <= accessDataUpdate_6;
        accessData_7 <= accessDataUpdate_7;
        accessPtr <= accessBufferDequeueFire | lastPtr | requestFireNext ? lsuRequestReg_instructionInformation_nf - {2'h0, accessBufferEnqueueFire & ~lastPtr} : accessPtr - 3'h1;
      end
      if (accessBufferDequeueFire) begin
        automatic logic [2047:0] _GEN_289 =
          (dataEEWOH[0]
             ? (_fillBySeg_T[0] ? regroupLoadData_0_0 : 2048'h0) | (_fillBySeg_T[1] ? regroupLoadData_0_1 : 2048'h0) | (_fillBySeg_T[2] ? regroupLoadData_0_2 : 2048'h0) | (_fillBySeg_T[3] ? regroupLoadData_0_3 : 2048'h0)
               | (_fillBySeg_T[4] ? regroupLoadData_0_4 : 2048'h0) | (_fillBySeg_T[5] ? regroupLoadData_0_5 : 2048'h0) | (_fillBySeg_T[6] ? regroupLoadData_0_6 : 2048'h0) | (_fillBySeg_T[7] ? regroupLoadData_0_7 : 2048'h0)
             : 2048'h0)
          | (dataEEWOH[1]
               ? (_fillBySeg_T[0] ? regroupLoadData_1_0 : 2048'h0) | (_fillBySeg_T[1] ? regroupLoadData_1_1 : 2048'h0) | (_fillBySeg_T[2] ? regroupLoadData_1_2 : 2048'h0) | (_fillBySeg_T[3] ? regroupLoadData_1_3 : 2048'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_1_4 : 2048'h0) | (_fillBySeg_T[5] ? regroupLoadData_1_5 : 2048'h0) | (_fillBySeg_T[6] ? regroupLoadData_1_6 : 2048'h0) | (_fillBySeg_T[7] ? regroupLoadData_1_7 : 2048'h0)
               : 2048'h0)
          | (dataEEWOH[2]
               ? (_fillBySeg_T[0] ? regroupLoadData_2_0 : 2048'h0) | (_fillBySeg_T[1] ? regroupLoadData_2_1 : 2048'h0) | (_fillBySeg_T[2] ? regroupLoadData_2_2 : 2048'h0) | (_fillBySeg_T[3] ? regroupLoadData_2_3 : 2048'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_2_4 : 2048'h0) | (_fillBySeg_T[5] ? regroupLoadData_2_5 : 2048'h0) | (_fillBySeg_T[6] ? regroupLoadData_2_6 : 2048'h0) | (_fillBySeg_T[7] ? regroupLoadData_2_7 : 2048'h0)
               : 2048'h0);
        dataBuffer_0 <= _GEN_289[255:0];
        dataBuffer_1 <= _GEN_289[511:256];
        dataBuffer_2 <= _GEN_289[767:512];
        dataBuffer_3 <= _GEN_289[1023:768];
        dataBuffer_4 <= _GEN_289[1279:1024];
        dataBuffer_5 <= _GEN_289[1535:1280];
        dataBuffer_6 <= _GEN_289[1791:1536];
        dataBuffer_7 <= _GEN_289[2047:1792];
        maskForBufferData_0 <= fillBySeg[31:0];
        maskForBufferData_1 <= fillBySeg[63:32];
        maskForBufferData_2 <= fillBySeg[95:64];
        maskForBufferData_3 <= fillBySeg[127:96];
        maskForBufferData_4 <= fillBySeg[159:128];
        maskForBufferData_5 <= fillBySeg[191:160];
        maskForBufferData_6 <= fillBySeg[223:192];
        maskForBufferData_7 <= fillBySeg[255:224];
        lastDataGroupInDataBuffer <= isLastRead;
      end
      else if (alignedDequeueFire) begin
        dataBuffer_0 <= dataBuffer_1;
        dataBuffer_1 <= dataBuffer_2;
        dataBuffer_2 <= dataBuffer_3;
        dataBuffer_3 <= dataBuffer_4;
        dataBuffer_4 <= dataBuffer_5;
        dataBuffer_5 <= dataBuffer_6;
        dataBuffer_6 <= dataBuffer_7;
        dataBuffer_7 <= 256'h0;
      end
      if (lsuRequest_valid | alignedDequeueFire) begin
        bufferBaseCacheLineIndex <= lsuRequest_valid ? 7'h0 : bufferBaseCacheLineIndex + 7'h1;
        maskTemp <= lsuRequest_valid ? 32'h0 : _GEN_287;
        canSendTail <= ~lsuRequest_valid & bufferValid & isLastCacheLineInBuffer & lastDataGroupInDataBuffer;
      end
      if (accessBufferDequeueFire | alignedDequeueFire)
        cacheLineIndexInBuffer <= accessBufferDequeueFire ? 3'h0 : cacheLineIndexInBuffer + 3'h1;
      hazardCheck <= ~lsuRequest_valid;
      if (lsuRequest_valid | _readStageValid_T_11)
        readStageValid_segPtr <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_11 & readStageValid_lastReadPtr)
        readStageValid_readCount <= readStageValid_nextReadCount;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup & readStageValid_lastReadPtr & _readStageValid_T_11)
        readStageValid_stageValid <= lsuRequest_valid;
      if (_readStageValid_T_11 ^ vrfReadQueueVec_0_deq_ready & vrfReadQueueVec_0_deq_valid)
        readStageValid_readCounter <= readStageValid_readCounter + readStageValid_counterChange;
      if (lsuRequest_valid | _readStageValid_T_30)
        readStageValid_segPtr_1 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_1 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_1 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_30 & readStageValid_lastReadPtr_1)
        readStageValid_readCount_1 <= readStageValid_nextReadCount_1;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_1 & readStageValid_lastReadPtr_1 & _readStageValid_T_30)
        readStageValid_stageValid_1 <= lsuRequest_valid;
      if (_readStageValid_T_30 ^ vrfReadQueueVec_1_deq_ready & vrfReadQueueVec_1_deq_valid)
        readStageValid_readCounter_1 <= readStageValid_readCounter_1 + readStageValid_counterChange_1;
      if (lsuRequest_valid | _readStageValid_T_49)
        readStageValid_segPtr_2 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_2 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_2 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_49 & readStageValid_lastReadPtr_2)
        readStageValid_readCount_2 <= readStageValid_nextReadCount_2;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_2 & readStageValid_lastReadPtr_2 & _readStageValid_T_49)
        readStageValid_stageValid_2 <= lsuRequest_valid;
      if (_readStageValid_T_49 ^ vrfReadQueueVec_2_deq_ready & vrfReadQueueVec_2_deq_valid)
        readStageValid_readCounter_2 <= readStageValid_readCounter_2 + readStageValid_counterChange_2;
      if (lsuRequest_valid | _readStageValid_T_68)
        readStageValid_segPtr_3 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_3 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_3 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_68 & readStageValid_lastReadPtr_3)
        readStageValid_readCount_3 <= readStageValid_nextReadCount_3;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_3 & readStageValid_lastReadPtr_3 & _readStageValid_T_68)
        readStageValid_stageValid_3 <= lsuRequest_valid;
      if (_readStageValid_T_68 ^ vrfReadQueueVec_3_deq_ready & vrfReadQueueVec_3_deq_valid)
        readStageValid_readCounter_3 <= readStageValid_readCounter_3 + readStageValid_counterChange_3;
      if (lsuRequest_valid | _readStageValid_T_87)
        readStageValid_segPtr_4 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_4 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_4 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_87 & readStageValid_lastReadPtr_4)
        readStageValid_readCount_4 <= readStageValid_nextReadCount_4;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_4 & readStageValid_lastReadPtr_4 & _readStageValid_T_87)
        readStageValid_stageValid_4 <= lsuRequest_valid;
      if (_readStageValid_T_87 ^ vrfReadQueueVec_4_deq_ready & vrfReadQueueVec_4_deq_valid)
        readStageValid_readCounter_4 <= readStageValid_readCounter_4 + readStageValid_counterChange_4;
      if (lsuRequest_valid | _readStageValid_T_106)
        readStageValid_segPtr_5 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_5 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_5 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_106 & readStageValid_lastReadPtr_5)
        readStageValid_readCount_5 <= readStageValid_nextReadCount_5;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_5 & readStageValid_lastReadPtr_5 & _readStageValid_T_106)
        readStageValid_stageValid_5 <= lsuRequest_valid;
      if (_readStageValid_T_106 ^ vrfReadQueueVec_5_deq_ready & vrfReadQueueVec_5_deq_valid)
        readStageValid_readCounter_5 <= readStageValid_readCounter_5 + readStageValid_counterChange_5;
      if (lsuRequest_valid | _readStageValid_T_125)
        readStageValid_segPtr_6 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_6 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_6 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_125 & readStageValid_lastReadPtr_6)
        readStageValid_readCount_6 <= readStageValid_nextReadCount_6;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_6 & readStageValid_lastReadPtr_6 & _readStageValid_T_125)
        readStageValid_stageValid_6 <= lsuRequest_valid;
      if (_readStageValid_T_125 ^ vrfReadQueueVec_6_deq_ready & vrfReadQueueVec_6_deq_valid)
        readStageValid_readCounter_6 <= readStageValid_readCounter_6 + readStageValid_counterChange_6;
      if (lsuRequest_valid | _readStageValid_T_144)
        readStageValid_segPtr_7 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_7 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_7 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_144 & readStageValid_lastReadPtr_7)
        readStageValid_readCount_7 <= readStageValid_nextReadCount_7;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_7 & readStageValid_lastReadPtr_7 & _readStageValid_T_144)
        readStageValid_stageValid_7 <= lsuRequest_valid;
      if (_readStageValid_T_144 ^ vrfReadQueueVec_7_deq_ready & vrfReadQueueVec_7_deq_valid)
        readStageValid_readCounter_7 <= readStageValid_readCounter_7 + readStageValid_counterChange_7;
      if (lastPtrEnq ^ accessBufferDequeueFire)
        bufferFull <= lastPtrEnq;
      if (accessBufferDequeueFire ^ bufferWillClear)
        bufferValid <= accessBufferDequeueFire;
      if (alignedDequeueFire)
        cacheLineTemp <= dataBuffer_0;
      idleNext <= _status_idle_output;
    end
    invalidInstructionNext <= invalidInstruction & lsuRequest_valid;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:158];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [7:0] i = 8'h0; i < 8'h9F; i += 8'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        lsuRequestReg_instructionInformation_nf = _RANDOM[8'h0][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[8'h0][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[8'h0][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[8'h0][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[8'h0][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[8'h0][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[8'h0][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[8'h0][19];
        lsuRequestReg_rs1Data = {_RANDOM[8'h0][31:20], _RANDOM[8'h1][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[8'h1][31:20], _RANDOM[8'h2][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[8'h2][22:20];
        csrInterfaceReg_vl = {_RANDOM[8'h2][31:23], _RANDOM[8'h3][2:0]};
        csrInterfaceReg_vStart = _RANDOM[8'h3][14:3];
        csrInterfaceReg_vlmul = _RANDOM[8'h3][17:15];
        csrInterfaceReg_vSew = _RANDOM[8'h3][19:18];
        csrInterfaceReg_vxrm = _RANDOM[8'h3][21:20];
        csrInterfaceReg_vta = _RANDOM[8'h3][22];
        csrInterfaceReg_vma = _RANDOM[8'h3][23];
        requestFireNext = _RANDOM[8'h3][24];
        dataEEW = _RANDOM[8'h3][26:25];
        maskReg = {_RANDOM[8'h3][31:27], _RANDOM[8'h4][26:0]};
        needAmend = _RANDOM[8'h4][27];
        lastMaskAmendReg = {_RANDOM[8'h4][31:28], _RANDOM[8'h5][26:0]};
        maskGroupCounter = {_RANDOM[8'h5][31:27], _RANDOM[8'h6][0]};
        maskCounterInGroup = _RANDOM[8'h6][2:1];
        isLastMaskGroup = _RANDOM[8'h7][3];
        accessData_0 = {_RANDOM[8'h7][31:4], _RANDOM[8'h8], _RANDOM[8'h9], _RANDOM[8'hA], _RANDOM[8'hB], _RANDOM[8'hC], _RANDOM[8'hD], _RANDOM[8'hE], _RANDOM[8'hF][3:0]};
        accessData_1 = {_RANDOM[8'hF][31:4], _RANDOM[8'h10], _RANDOM[8'h11], _RANDOM[8'h12], _RANDOM[8'h13], _RANDOM[8'h14], _RANDOM[8'h15], _RANDOM[8'h16], _RANDOM[8'h17][3:0]};
        accessData_2 = {_RANDOM[8'h17][31:4], _RANDOM[8'h18], _RANDOM[8'h19], _RANDOM[8'h1A], _RANDOM[8'h1B], _RANDOM[8'h1C], _RANDOM[8'h1D], _RANDOM[8'h1E], _RANDOM[8'h1F][3:0]};
        accessData_3 = {_RANDOM[8'h1F][31:4], _RANDOM[8'h20], _RANDOM[8'h21], _RANDOM[8'h22], _RANDOM[8'h23], _RANDOM[8'h24], _RANDOM[8'h25], _RANDOM[8'h26], _RANDOM[8'h27][3:0]};
        accessData_4 = {_RANDOM[8'h27][31:4], _RANDOM[8'h28], _RANDOM[8'h29], _RANDOM[8'h2A], _RANDOM[8'h2B], _RANDOM[8'h2C], _RANDOM[8'h2D], _RANDOM[8'h2E], _RANDOM[8'h2F][3:0]};
        accessData_5 = {_RANDOM[8'h2F][31:4], _RANDOM[8'h30], _RANDOM[8'h31], _RANDOM[8'h32], _RANDOM[8'h33], _RANDOM[8'h34], _RANDOM[8'h35], _RANDOM[8'h36], _RANDOM[8'h37][3:0]};
        accessData_6 = {_RANDOM[8'h37][31:4], _RANDOM[8'h38], _RANDOM[8'h39], _RANDOM[8'h3A], _RANDOM[8'h3B], _RANDOM[8'h3C], _RANDOM[8'h3D], _RANDOM[8'h3E], _RANDOM[8'h3F][3:0]};
        accessData_7 = {_RANDOM[8'h3F][31:4], _RANDOM[8'h40], _RANDOM[8'h41], _RANDOM[8'h42], _RANDOM[8'h43], _RANDOM[8'h44], _RANDOM[8'h45], _RANDOM[8'h46], _RANDOM[8'h47][3:0]};
        accessPtr = _RANDOM[8'h47][6:4];
        dataGroup = _RANDOM[8'h47][20:15];
        dataBuffer_0 = {_RANDOM[8'h47][31:21], _RANDOM[8'h48], _RANDOM[8'h49], _RANDOM[8'h4A], _RANDOM[8'h4B], _RANDOM[8'h4C], _RANDOM[8'h4D], _RANDOM[8'h4E], _RANDOM[8'h4F][20:0]};
        dataBuffer_1 = {_RANDOM[8'h4F][31:21], _RANDOM[8'h50], _RANDOM[8'h51], _RANDOM[8'h52], _RANDOM[8'h53], _RANDOM[8'h54], _RANDOM[8'h55], _RANDOM[8'h56], _RANDOM[8'h57][20:0]};
        dataBuffer_2 = {_RANDOM[8'h57][31:21], _RANDOM[8'h58], _RANDOM[8'h59], _RANDOM[8'h5A], _RANDOM[8'h5B], _RANDOM[8'h5C], _RANDOM[8'h5D], _RANDOM[8'h5E], _RANDOM[8'h5F][20:0]};
        dataBuffer_3 = {_RANDOM[8'h5F][31:21], _RANDOM[8'h60], _RANDOM[8'h61], _RANDOM[8'h62], _RANDOM[8'h63], _RANDOM[8'h64], _RANDOM[8'h65], _RANDOM[8'h66], _RANDOM[8'h67][20:0]};
        dataBuffer_4 = {_RANDOM[8'h67][31:21], _RANDOM[8'h68], _RANDOM[8'h69], _RANDOM[8'h6A], _RANDOM[8'h6B], _RANDOM[8'h6C], _RANDOM[8'h6D], _RANDOM[8'h6E], _RANDOM[8'h6F][20:0]};
        dataBuffer_5 = {_RANDOM[8'h6F][31:21], _RANDOM[8'h70], _RANDOM[8'h71], _RANDOM[8'h72], _RANDOM[8'h73], _RANDOM[8'h74], _RANDOM[8'h75], _RANDOM[8'h76], _RANDOM[8'h77][20:0]};
        dataBuffer_6 = {_RANDOM[8'h77][31:21], _RANDOM[8'h78], _RANDOM[8'h79], _RANDOM[8'h7A], _RANDOM[8'h7B], _RANDOM[8'h7C], _RANDOM[8'h7D], _RANDOM[8'h7E], _RANDOM[8'h7F][20:0]};
        dataBuffer_7 = {_RANDOM[8'h7F][31:21], _RANDOM[8'h80], _RANDOM[8'h81], _RANDOM[8'h82], _RANDOM[8'h83], _RANDOM[8'h84], _RANDOM[8'h85], _RANDOM[8'h86], _RANDOM[8'h87][20:0]};
        bufferBaseCacheLineIndex = _RANDOM[8'h87][27:21];
        cacheLineIndexInBuffer = _RANDOM[8'h87][30:28];
        invalidInstructionNext = _RANDOM[8'h87][31];
        segmentInstructionIndexInterval = _RANDOM[8'h88][3:0];
        lastWriteVrfIndexReg = _RANDOM[8'h88][17:4];
        lastCacheNeedPush = _RANDOM[8'h88][18];
        cacheLineNumberReg = {_RANDOM[8'h88][31:19], _RANDOM[8'h89][0]};
        lastDataGroupReg = _RANDOM[8'h89][10:1];
        hazardCheck = _RANDOM[8'h89][11];
        readStageValid_segPtr = _RANDOM[8'h89][14:12];
        readStageValid_readCount = _RANDOM[8'h89][20:15];
        readStageValid_stageValid = _RANDOM[8'h89][21];
        readStageValid_readCounter = _RANDOM[8'h89][25:22];
        readStageValid_segPtr_1 = _RANDOM[8'h89][28:26];
        readStageValid_readCount_1 = {_RANDOM[8'h89][31:29], _RANDOM[8'h8A][2:0]};
        readStageValid_stageValid_1 = _RANDOM[8'h8A][3];
        readStageValid_readCounter_1 = _RANDOM[8'h8A][7:4];
        readStageValid_segPtr_2 = _RANDOM[8'h8A][10:8];
        readStageValid_readCount_2 = _RANDOM[8'h8A][16:11];
        readStageValid_stageValid_2 = _RANDOM[8'h8A][17];
        readStageValid_readCounter_2 = _RANDOM[8'h8A][21:18];
        readStageValid_segPtr_3 = _RANDOM[8'h8A][24:22];
        readStageValid_readCount_3 = _RANDOM[8'h8A][30:25];
        readStageValid_stageValid_3 = _RANDOM[8'h8A][31];
        readStageValid_readCounter_3 = _RANDOM[8'h8B][3:0];
        readStageValid_segPtr_4 = _RANDOM[8'h8B][6:4];
        readStageValid_readCount_4 = _RANDOM[8'h8B][12:7];
        readStageValid_stageValid_4 = _RANDOM[8'h8B][13];
        readStageValid_readCounter_4 = _RANDOM[8'h8B][17:14];
        readStageValid_segPtr_5 = _RANDOM[8'h8B][20:18];
        readStageValid_readCount_5 = _RANDOM[8'h8B][26:21];
        readStageValid_stageValid_5 = _RANDOM[8'h8B][27];
        readStageValid_readCounter_5 = _RANDOM[8'h8B][31:28];
        readStageValid_segPtr_6 = _RANDOM[8'h8C][2:0];
        readStageValid_readCount_6 = _RANDOM[8'h8C][8:3];
        readStageValid_stageValid_6 = _RANDOM[8'h8C][9];
        readStageValid_readCounter_6 = _RANDOM[8'h8C][13:10];
        readStageValid_segPtr_7 = _RANDOM[8'h8C][16:14];
        readStageValid_readCount_7 = _RANDOM[8'h8C][22:17];
        readStageValid_stageValid_7 = _RANDOM[8'h8C][23];
        readStageValid_readCounter_7 = _RANDOM[8'h8C][27:24];
        bufferFull = _RANDOM[8'h8C][28];
        bufferValid = _RANDOM[8'h8C][29];
        maskForBufferData_0 = {_RANDOM[8'h8C][31:30], _RANDOM[8'h8D][29:0]};
        maskForBufferData_1 = {_RANDOM[8'h8D][31:30], _RANDOM[8'h8E][29:0]};
        maskForBufferData_2 = {_RANDOM[8'h8E][31:30], _RANDOM[8'h8F][29:0]};
        maskForBufferData_3 = {_RANDOM[8'h8F][31:30], _RANDOM[8'h90][29:0]};
        maskForBufferData_4 = {_RANDOM[8'h90][31:30], _RANDOM[8'h91][29:0]};
        maskForBufferData_5 = {_RANDOM[8'h91][31:30], _RANDOM[8'h92][29:0]};
        maskForBufferData_6 = {_RANDOM[8'h92][31:30], _RANDOM[8'h93][29:0]};
        maskForBufferData_7 = {_RANDOM[8'h93][31:30], _RANDOM[8'h94][29:0]};
        lastDataGroupInDataBuffer = _RANDOM[8'h94][30];
        cacheLineTemp = {_RANDOM[8'h94][31], _RANDOM[8'h95], _RANDOM[8'h96], _RANDOM[8'h97], _RANDOM[8'h98], _RANDOM[8'h99], _RANDOM[8'h9A], _RANDOM[8'h9B], _RANDOM[8'h9C][30:0]};
        maskTemp = {_RANDOM[8'h9C][31], _RANDOM[8'h9D][30:0]};
        canSendTail = _RANDOM[8'h9D][31];
        idleNext = _RANDOM[8'h9E][0];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire             vrfReadQueueVec_0_empty;
  assign vrfReadQueueVec_0_empty = _vrfReadQueueVec_fifo_empty;
  wire             vrfReadQueueVec_0_full;
  assign vrfReadQueueVec_0_full = _vrfReadQueueVec_fifo_full;
  wire             vrfReadQueueVec_1_empty;
  assign vrfReadQueueVec_1_empty = _vrfReadQueueVec_fifo_1_empty;
  wire             vrfReadQueueVec_1_full;
  assign vrfReadQueueVec_1_full = _vrfReadQueueVec_fifo_1_full;
  wire             vrfReadQueueVec_2_empty;
  assign vrfReadQueueVec_2_empty = _vrfReadQueueVec_fifo_2_empty;
  wire             vrfReadQueueVec_2_full;
  assign vrfReadQueueVec_2_full = _vrfReadQueueVec_fifo_2_full;
  wire             vrfReadQueueVec_3_empty;
  assign vrfReadQueueVec_3_empty = _vrfReadQueueVec_fifo_3_empty;
  wire             vrfReadQueueVec_3_full;
  assign vrfReadQueueVec_3_full = _vrfReadQueueVec_fifo_3_full;
  wire             vrfReadQueueVec_4_empty;
  assign vrfReadQueueVec_4_empty = _vrfReadQueueVec_fifo_4_empty;
  wire             vrfReadQueueVec_4_full;
  assign vrfReadQueueVec_4_full = _vrfReadQueueVec_fifo_4_full;
  wire             vrfReadQueueVec_5_empty;
  assign vrfReadQueueVec_5_empty = _vrfReadQueueVec_fifo_5_empty;
  wire             vrfReadQueueVec_5_full;
  assign vrfReadQueueVec_5_full = _vrfReadQueueVec_fifo_5_full;
  wire             vrfReadQueueVec_6_empty;
  assign vrfReadQueueVec_6_empty = _vrfReadQueueVec_fifo_6_empty;
  wire             vrfReadQueueVec_6_full;
  assign vrfReadQueueVec_6_full = _vrfReadQueueVec_fifo_6_full;
  wire             vrfReadQueueVec_7_empty;
  assign vrfReadQueueVec_7_empty = _vrfReadQueueVec_fifo_7_empty;
  wire             vrfReadQueueVec_7_full;
  assign vrfReadQueueVec_7_full = _vrfReadQueueVec_fifo_7_full;
  wire             addressQueue_empty;
  assign addressQueue_empty = _addressQueue_fifo_empty;
  wire             addressQueue_full;
  assign addressQueue_full = _addressQueue_fifo_full;
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_0_enq_ready & vrfReadQueueVec_0_enq_valid & ~(_vrfReadQueueVec_fifo_empty & vrfReadQueueVec_0_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_0_deq_ready & ~_vrfReadQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_0_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_empty),
    .almost_empty (vrfReadQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_0_almostFull),
    .full         (_vrfReadQueueVec_fifo_full),
    .error        (_vrfReadQueueVec_fifo_error),
    .data_out     (_vrfReadQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_1_enq_ready & vrfReadQueueVec_1_enq_valid & ~(_vrfReadQueueVec_fifo_1_empty & vrfReadQueueVec_1_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_1_deq_ready & ~_vrfReadQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_1_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_1_empty),
    .almost_empty (vrfReadQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_1_almostFull),
    .full         (_vrfReadQueueVec_fifo_1_full),
    .error        (_vrfReadQueueVec_fifo_1_error),
    .data_out     (_vrfReadQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_2_enq_ready & vrfReadQueueVec_2_enq_valid & ~(_vrfReadQueueVec_fifo_2_empty & vrfReadQueueVec_2_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_2_deq_ready & ~_vrfReadQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_2_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_2_empty),
    .almost_empty (vrfReadQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_2_almostFull),
    .full         (_vrfReadQueueVec_fifo_2_full),
    .error        (_vrfReadQueueVec_fifo_2_error),
    .data_out     (_vrfReadQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_3_enq_ready & vrfReadQueueVec_3_enq_valid & ~(_vrfReadQueueVec_fifo_3_empty & vrfReadQueueVec_3_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_3_deq_ready & ~_vrfReadQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_3_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_3_empty),
    .almost_empty (vrfReadQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_3_almostFull),
    .full         (_vrfReadQueueVec_fifo_3_full),
    .error        (_vrfReadQueueVec_fifo_3_error),
    .data_out     (_vrfReadQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_4_enq_ready & vrfReadQueueVec_4_enq_valid & ~(_vrfReadQueueVec_fifo_4_empty & vrfReadQueueVec_4_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_4_deq_ready & ~_vrfReadQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_4_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_4_empty),
    .almost_empty (vrfReadQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_4_almostFull),
    .full         (_vrfReadQueueVec_fifo_4_full),
    .error        (_vrfReadQueueVec_fifo_4_error),
    .data_out     (_vrfReadQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_5_enq_ready & vrfReadQueueVec_5_enq_valid & ~(_vrfReadQueueVec_fifo_5_empty & vrfReadQueueVec_5_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_5_deq_ready & ~_vrfReadQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_5_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_5_empty),
    .almost_empty (vrfReadQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_5_almostFull),
    .full         (_vrfReadQueueVec_fifo_5_full),
    .error        (_vrfReadQueueVec_fifo_5_error),
    .data_out     (_vrfReadQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_6_enq_ready & vrfReadQueueVec_6_enq_valid & ~(_vrfReadQueueVec_fifo_6_empty & vrfReadQueueVec_6_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_6_deq_ready & ~_vrfReadQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_6_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_6_empty),
    .almost_empty (vrfReadQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_6_almostFull),
    .full         (_vrfReadQueueVec_fifo_6_full),
    .error        (_vrfReadQueueVec_fifo_6_error),
    .data_out     (_vrfReadQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_7_enq_ready & vrfReadQueueVec_7_enq_valid & ~(_vrfReadQueueVec_fifo_7_empty & vrfReadQueueVec_7_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_7_deq_ready & ~_vrfReadQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_7_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_7_empty),
    .almost_empty (vrfReadQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_7_almostFull),
    .full         (_vrfReadQueueVec_fifo_7_full),
    .error        (_vrfReadQueueVec_fifo_7_error),
    .data_out     (_vrfReadQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(32),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) addressQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(addressQueue_enq_ready & addressQueue_enq_valid)),
    .pop_req_n    (~(addressQueue_deq_ready & ~_addressQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (addressQueue_enq_bits),
    .empty        (_addressQueue_fifo_empty),
    .almost_empty (addressQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (addressQueue_almostFull),
    .full         (_addressQueue_fifo_full),
    .error        (_addressQueue_fifo_error),
    .data_out     (addressQueue_deq_bits)
  );
  assign maskSelect_valid = _maskSelect_valid_output;
  assign maskSelect_bits = _maskSelect_bits_output;
  assign memRequest_valid = memRequest_valid_0;
  assign memRequest_bits_data = memRequest_bits_data_0;
  assign memRequest_bits_mask = memRequest_bits_mask_0;
  assign memRequest_bits_index = memRequest_bits_index_0;
  assign memRequest_bits_address = memRequest_bits_address_0;
  assign status_idle = _status_idle_output;
  assign status_last = ~idleNext & _status_idle_output | invalidInstructionNext;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_changeMaskGroup = _maskSelect_valid_output & ~lsuRequest_valid;
  assign status_startAddress = addressQueue_deq_valid ? addressQueue_deq_bits : alignedDequeueAddress;
  assign status_endAddress = {lsuRequestReg_rs1Data[31:5] + {13'h0, cacheLineNumberReg}, 5'h0};
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_offset = vrfReadDataPorts_0_bits_offset_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_offset = vrfReadDataPorts_1_bits_offset_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_offset = vrfReadDataPorts_2_bits_offset_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_offset = vrfReadDataPorts_3_bits_offset_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfReadDataPorts_4_valid = vrfReadDataPorts_4_valid_0;
  assign vrfReadDataPorts_4_bits_vs = vrfReadDataPorts_4_bits_vs_0;
  assign vrfReadDataPorts_4_bits_offset = vrfReadDataPorts_4_bits_offset_0;
  assign vrfReadDataPorts_4_bits_instructionIndex = vrfReadDataPorts_4_bits_instructionIndex_0;
  assign vrfReadDataPorts_5_valid = vrfReadDataPorts_5_valid_0;
  assign vrfReadDataPorts_5_bits_vs = vrfReadDataPorts_5_bits_vs_0;
  assign vrfReadDataPorts_5_bits_offset = vrfReadDataPorts_5_bits_offset_0;
  assign vrfReadDataPorts_5_bits_instructionIndex = vrfReadDataPorts_5_bits_instructionIndex_0;
  assign vrfReadDataPorts_6_valid = vrfReadDataPorts_6_valid_0;
  assign vrfReadDataPorts_6_bits_vs = vrfReadDataPorts_6_bits_vs_0;
  assign vrfReadDataPorts_6_bits_offset = vrfReadDataPorts_6_bits_offset_0;
  assign vrfReadDataPorts_6_bits_instructionIndex = vrfReadDataPorts_6_bits_instructionIndex_0;
  assign vrfReadDataPorts_7_valid = vrfReadDataPorts_7_valid_0;
  assign vrfReadDataPorts_7_bits_vs = vrfReadDataPorts_7_bits_vs_0;
  assign vrfReadDataPorts_7_bits_offset = vrfReadDataPorts_7_bits_offset_0;
  assign vrfReadDataPorts_7_bits_instructionIndex = vrfReadDataPorts_7_bits_instructionIndex_0;
endmodule

