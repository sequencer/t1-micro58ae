module MaskExtend(
  input  [1:0]   in_eew,
  input  [2:0]   in_uop,
  input  [127:0] in_source2,
  input  [4:0]   in_groupCounter,
  output [127:0] out
);

  wire [3:0]   _eew1H_T = 4'h1 << in_eew;
  wire [2:0]   eew1H = _eew1H_T[2:0];
  wire         isMaskDestination = in_uop == 3'h0;
  wire [31:0]  sourceDataVec_0 = in_source2[31:0];
  wire [31:0]  sourceDataVec_1 = in_source2[63:32];
  wire [31:0]  sourceDataVec_2 = in_source2[95:64];
  wire [31:0]  sourceDataVec_3 = in_source2[127:96];
  wire [1:0]   maskDestinationResult_lo = sourceDataVec_0[1:0];
  wire [1:0]   maskDestinationResult_hi = sourceDataVec_0[3:2];
  wire [1:0]   maskDestinationResult_lo_1 = sourceDataVec_0[5:4];
  wire [1:0]   maskDestinationResult_hi_1 = sourceDataVec_0[7:6];
  wire [1:0]   maskDestinationResult_lo_2 = sourceDataVec_0[9:8];
  wire [1:0]   maskDestinationResult_hi_2 = sourceDataVec_0[11:10];
  wire [1:0]   maskDestinationResult_lo_3 = sourceDataVec_0[13:12];
  wire [1:0]   maskDestinationResult_hi_3 = sourceDataVec_0[15:14];
  wire [1:0]   maskDestinationResult_lo_4 = sourceDataVec_0[17:16];
  wire [1:0]   maskDestinationResult_hi_4 = sourceDataVec_0[19:18];
  wire [1:0]   maskDestinationResult_lo_5 = sourceDataVec_0[21:20];
  wire [1:0]   maskDestinationResult_hi_5 = sourceDataVec_0[23:22];
  wire [1:0]   maskDestinationResult_lo_6 = sourceDataVec_0[25:24];
  wire [1:0]   maskDestinationResult_hi_6 = sourceDataVec_0[27:26];
  wire [1:0]   maskDestinationResult_lo_7 = sourceDataVec_0[29:28];
  wire [1:0]   maskDestinationResult_hi_7 = sourceDataVec_0[31:30];
  wire [1:0]   maskDestinationResult_lo_8 = sourceDataVec_1[1:0];
  wire [1:0]   maskDestinationResult_hi_8 = sourceDataVec_1[3:2];
  wire [1:0]   maskDestinationResult_lo_9 = sourceDataVec_1[5:4];
  wire [1:0]   maskDestinationResult_hi_9 = sourceDataVec_1[7:6];
  wire [1:0]   maskDestinationResult_lo_10 = sourceDataVec_1[9:8];
  wire [1:0]   maskDestinationResult_hi_10 = sourceDataVec_1[11:10];
  wire [1:0]   maskDestinationResult_lo_11 = sourceDataVec_1[13:12];
  wire [1:0]   maskDestinationResult_hi_11 = sourceDataVec_1[15:14];
  wire [1:0]   maskDestinationResult_lo_12 = sourceDataVec_1[17:16];
  wire [1:0]   maskDestinationResult_hi_12 = sourceDataVec_1[19:18];
  wire [1:0]   maskDestinationResult_lo_13 = sourceDataVec_1[21:20];
  wire [1:0]   maskDestinationResult_hi_13 = sourceDataVec_1[23:22];
  wire [1:0]   maskDestinationResult_lo_14 = sourceDataVec_1[25:24];
  wire [1:0]   maskDestinationResult_hi_14 = sourceDataVec_1[27:26];
  wire [1:0]   maskDestinationResult_lo_15 = sourceDataVec_1[29:28];
  wire [1:0]   maskDestinationResult_hi_15 = sourceDataVec_1[31:30];
  wire [1:0]   maskDestinationResult_lo_16 = sourceDataVec_2[1:0];
  wire [1:0]   maskDestinationResult_hi_16 = sourceDataVec_2[3:2];
  wire [1:0]   maskDestinationResult_lo_17 = sourceDataVec_2[5:4];
  wire [1:0]   maskDestinationResult_hi_17 = sourceDataVec_2[7:6];
  wire [1:0]   maskDestinationResult_lo_18 = sourceDataVec_2[9:8];
  wire [1:0]   maskDestinationResult_hi_18 = sourceDataVec_2[11:10];
  wire [1:0]   maskDestinationResult_lo_19 = sourceDataVec_2[13:12];
  wire [1:0]   maskDestinationResult_hi_19 = sourceDataVec_2[15:14];
  wire [1:0]   maskDestinationResult_lo_20 = sourceDataVec_2[17:16];
  wire [1:0]   maskDestinationResult_hi_20 = sourceDataVec_2[19:18];
  wire [1:0]   maskDestinationResult_lo_21 = sourceDataVec_2[21:20];
  wire [1:0]   maskDestinationResult_hi_21 = sourceDataVec_2[23:22];
  wire [1:0]   maskDestinationResult_lo_22 = sourceDataVec_2[25:24];
  wire [1:0]   maskDestinationResult_hi_22 = sourceDataVec_2[27:26];
  wire [1:0]   maskDestinationResult_lo_23 = sourceDataVec_2[29:28];
  wire [1:0]   maskDestinationResult_hi_23 = sourceDataVec_2[31:30];
  wire [1:0]   maskDestinationResult_lo_24 = sourceDataVec_3[1:0];
  wire [1:0]   maskDestinationResult_hi_24 = sourceDataVec_3[3:2];
  wire [1:0]   maskDestinationResult_lo_25 = sourceDataVec_3[5:4];
  wire [1:0]   maskDestinationResult_hi_25 = sourceDataVec_3[7:6];
  wire [1:0]   maskDestinationResult_lo_26 = sourceDataVec_3[9:8];
  wire [1:0]   maskDestinationResult_hi_26 = sourceDataVec_3[11:10];
  wire [1:0]   maskDestinationResult_lo_27 = sourceDataVec_3[13:12];
  wire [1:0]   maskDestinationResult_hi_27 = sourceDataVec_3[15:14];
  wire [1:0]   maskDestinationResult_lo_28 = sourceDataVec_3[17:16];
  wire [1:0]   maskDestinationResult_hi_28 = sourceDataVec_3[19:18];
  wire [1:0]   maskDestinationResult_lo_29 = sourceDataVec_3[21:20];
  wire [1:0]   maskDestinationResult_hi_29 = sourceDataVec_3[23:22];
  wire [1:0]   maskDestinationResult_lo_30 = sourceDataVec_3[25:24];
  wire [1:0]   maskDestinationResult_hi_30 = sourceDataVec_3[27:26];
  wire [1:0]   maskDestinationResult_lo_31 = sourceDataVec_3[29:28];
  wire [1:0]   maskDestinationResult_hi_31 = sourceDataVec_3[31:30];
  wire [7:0]   maskDestinationResult_lo_32 = {maskDestinationResult_hi_8, maskDestinationResult_lo_8, maskDestinationResult_hi, maskDestinationResult_lo};
  wire [7:0]   maskDestinationResult_hi_32 = {maskDestinationResult_hi_24, maskDestinationResult_lo_24, maskDestinationResult_hi_16, maskDestinationResult_lo_16};
  wire [7:0]   maskDestinationResult_lo_33 = {maskDestinationResult_hi_9, maskDestinationResult_lo_9, maskDestinationResult_hi_1, maskDestinationResult_lo_1};
  wire [7:0]   maskDestinationResult_hi_33 = {maskDestinationResult_hi_25, maskDestinationResult_lo_25, maskDestinationResult_hi_17, maskDestinationResult_lo_17};
  wire [7:0]   maskDestinationResult_lo_34 = {maskDestinationResult_hi_10, maskDestinationResult_lo_10, maskDestinationResult_hi_2, maskDestinationResult_lo_2};
  wire [7:0]   maskDestinationResult_hi_34 = {maskDestinationResult_hi_26, maskDestinationResult_lo_26, maskDestinationResult_hi_18, maskDestinationResult_lo_18};
  wire [7:0]   maskDestinationResult_lo_35 = {maskDestinationResult_hi_11, maskDestinationResult_lo_11, maskDestinationResult_hi_3, maskDestinationResult_lo_3};
  wire [7:0]   maskDestinationResult_hi_35 = {maskDestinationResult_hi_27, maskDestinationResult_lo_27, maskDestinationResult_hi_19, maskDestinationResult_lo_19};
  wire [7:0]   maskDestinationResult_lo_36 = {maskDestinationResult_hi_12, maskDestinationResult_lo_12, maskDestinationResult_hi_4, maskDestinationResult_lo_4};
  wire [7:0]   maskDestinationResult_hi_36 = {maskDestinationResult_hi_28, maskDestinationResult_lo_28, maskDestinationResult_hi_20, maskDestinationResult_lo_20};
  wire [7:0]   maskDestinationResult_lo_37 = {maskDestinationResult_hi_13, maskDestinationResult_lo_13, maskDestinationResult_hi_5, maskDestinationResult_lo_5};
  wire [7:0]   maskDestinationResult_hi_37 = {maskDestinationResult_hi_29, maskDestinationResult_lo_29, maskDestinationResult_hi_21, maskDestinationResult_lo_21};
  wire [7:0]   maskDestinationResult_lo_38 = {maskDestinationResult_hi_14, maskDestinationResult_lo_14, maskDestinationResult_hi_6, maskDestinationResult_lo_6};
  wire [7:0]   maskDestinationResult_hi_38 = {maskDestinationResult_hi_30, maskDestinationResult_lo_30, maskDestinationResult_hi_22, maskDestinationResult_lo_22};
  wire [7:0]   maskDestinationResult_lo_39 = {maskDestinationResult_hi_15, maskDestinationResult_lo_15, maskDestinationResult_hi_7, maskDestinationResult_lo_7};
  wire [7:0]   maskDestinationResult_hi_39 = {maskDestinationResult_hi_31, maskDestinationResult_lo_31, maskDestinationResult_hi_23, maskDestinationResult_lo_23};
  wire [31:0]  maskDestinationResult_lo_lo = {maskDestinationResult_hi_33, maskDestinationResult_lo_33, maskDestinationResult_hi_32, maskDestinationResult_lo_32};
  wire [31:0]  maskDestinationResult_lo_hi = {maskDestinationResult_hi_35, maskDestinationResult_lo_35, maskDestinationResult_hi_34, maskDestinationResult_lo_34};
  wire [63:0]  maskDestinationResult_lo_40 = {maskDestinationResult_lo_hi, maskDestinationResult_lo_lo};
  wire [31:0]  maskDestinationResult_hi_lo = {maskDestinationResult_hi_37, maskDestinationResult_lo_37, maskDestinationResult_hi_36, maskDestinationResult_lo_36};
  wire [31:0]  maskDestinationResult_hi_hi = {maskDestinationResult_hi_39, maskDestinationResult_lo_39, maskDestinationResult_hi_38, maskDestinationResult_lo_38};
  wire [63:0]  maskDestinationResult_hi_40 = {maskDestinationResult_hi_hi, maskDestinationResult_hi_lo};
  wire [3:0]   maskDestinationResult_lo_41 = {sourceDataVec_1[1:0], sourceDataVec_0[1:0]};
  wire [3:0]   maskDestinationResult_hi_41 = {sourceDataVec_3[1:0], sourceDataVec_2[1:0]};
  wire [3:0]   maskDestinationResult_lo_42 = {sourceDataVec_1[3:2], sourceDataVec_0[3:2]};
  wire [3:0]   maskDestinationResult_hi_42 = {sourceDataVec_3[3:2], sourceDataVec_2[3:2]};
  wire [3:0]   maskDestinationResult_lo_43 = {sourceDataVec_1[5:4], sourceDataVec_0[5:4]};
  wire [3:0]   maskDestinationResult_hi_43 = {sourceDataVec_3[5:4], sourceDataVec_2[5:4]};
  wire [3:0]   maskDestinationResult_lo_44 = {sourceDataVec_1[7:6], sourceDataVec_0[7:6]};
  wire [3:0]   maskDestinationResult_hi_44 = {sourceDataVec_3[7:6], sourceDataVec_2[7:6]};
  wire [3:0]   maskDestinationResult_lo_45 = {sourceDataVec_1[9:8], sourceDataVec_0[9:8]};
  wire [3:0]   maskDestinationResult_hi_45 = {sourceDataVec_3[9:8], sourceDataVec_2[9:8]};
  wire [3:0]   maskDestinationResult_lo_46 = {sourceDataVec_1[11:10], sourceDataVec_0[11:10]};
  wire [3:0]   maskDestinationResult_hi_46 = {sourceDataVec_3[11:10], sourceDataVec_2[11:10]};
  wire [3:0]   maskDestinationResult_lo_47 = {sourceDataVec_1[13:12], sourceDataVec_0[13:12]};
  wire [3:0]   maskDestinationResult_hi_47 = {sourceDataVec_3[13:12], sourceDataVec_2[13:12]};
  wire [3:0]   maskDestinationResult_lo_48 = {sourceDataVec_1[15:14], sourceDataVec_0[15:14]};
  wire [3:0]   maskDestinationResult_hi_48 = {sourceDataVec_3[15:14], sourceDataVec_2[15:14]};
  wire [3:0]   maskDestinationResult_lo_49 = {sourceDataVec_1[17:16], sourceDataVec_0[17:16]};
  wire [3:0]   maskDestinationResult_hi_49 = {sourceDataVec_3[17:16], sourceDataVec_2[17:16]};
  wire [3:0]   maskDestinationResult_lo_50 = {sourceDataVec_1[19:18], sourceDataVec_0[19:18]};
  wire [3:0]   maskDestinationResult_hi_50 = {sourceDataVec_3[19:18], sourceDataVec_2[19:18]};
  wire [3:0]   maskDestinationResult_lo_51 = {sourceDataVec_1[21:20], sourceDataVec_0[21:20]};
  wire [3:0]   maskDestinationResult_hi_51 = {sourceDataVec_3[21:20], sourceDataVec_2[21:20]};
  wire [3:0]   maskDestinationResult_lo_52 = {sourceDataVec_1[23:22], sourceDataVec_0[23:22]};
  wire [3:0]   maskDestinationResult_hi_52 = {sourceDataVec_3[23:22], sourceDataVec_2[23:22]};
  wire [3:0]   maskDestinationResult_lo_53 = {sourceDataVec_1[25:24], sourceDataVec_0[25:24]};
  wire [3:0]   maskDestinationResult_hi_53 = {sourceDataVec_3[25:24], sourceDataVec_2[25:24]};
  wire [3:0]   maskDestinationResult_lo_54 = {sourceDataVec_1[27:26], sourceDataVec_0[27:26]};
  wire [3:0]   maskDestinationResult_hi_54 = {sourceDataVec_3[27:26], sourceDataVec_2[27:26]};
  wire [3:0]   maskDestinationResult_lo_55 = {sourceDataVec_1[29:28], sourceDataVec_0[29:28]};
  wire [3:0]   maskDestinationResult_hi_55 = {sourceDataVec_3[29:28], sourceDataVec_2[29:28]};
  wire [3:0]   maskDestinationResult_lo_56 = {sourceDataVec_1[31:30], sourceDataVec_0[31:30]};
  wire [3:0]   maskDestinationResult_hi_56 = {sourceDataVec_3[31:30], sourceDataVec_2[31:30]};
  wire [15:0]  maskDestinationResult_lo_lo_lo = {maskDestinationResult_hi_42, maskDestinationResult_lo_42, maskDestinationResult_hi_41, maskDestinationResult_lo_41};
  wire [15:0]  maskDestinationResult_lo_lo_hi = {maskDestinationResult_hi_44, maskDestinationResult_lo_44, maskDestinationResult_hi_43, maskDestinationResult_lo_43};
  wire [31:0]  maskDestinationResult_lo_lo_1 = {maskDestinationResult_lo_lo_hi, maskDestinationResult_lo_lo_lo};
  wire [15:0]  maskDestinationResult_lo_hi_lo = {maskDestinationResult_hi_46, maskDestinationResult_lo_46, maskDestinationResult_hi_45, maskDestinationResult_lo_45};
  wire [15:0]  maskDestinationResult_lo_hi_hi = {maskDestinationResult_hi_48, maskDestinationResult_lo_48, maskDestinationResult_hi_47, maskDestinationResult_lo_47};
  wire [31:0]  maskDestinationResult_lo_hi_1 = {maskDestinationResult_lo_hi_hi, maskDestinationResult_lo_hi_lo};
  wire [63:0]  maskDestinationResult_lo_57 = {maskDestinationResult_lo_hi_1, maskDestinationResult_lo_lo_1};
  wire [15:0]  maskDestinationResult_hi_lo_lo = {maskDestinationResult_hi_50, maskDestinationResult_lo_50, maskDestinationResult_hi_49, maskDestinationResult_lo_49};
  wire [15:0]  maskDestinationResult_hi_lo_hi = {maskDestinationResult_hi_52, maskDestinationResult_lo_52, maskDestinationResult_hi_51, maskDestinationResult_lo_51};
  wire [31:0]  maskDestinationResult_hi_lo_1 = {maskDestinationResult_hi_lo_hi, maskDestinationResult_hi_lo_lo};
  wire [15:0]  maskDestinationResult_hi_hi_lo = {maskDestinationResult_hi_54, maskDestinationResult_lo_54, maskDestinationResult_hi_53, maskDestinationResult_lo_53};
  wire [15:0]  maskDestinationResult_hi_hi_hi = {maskDestinationResult_hi_56, maskDestinationResult_lo_56, maskDestinationResult_hi_55, maskDestinationResult_lo_55};
  wire [31:0]  maskDestinationResult_hi_hi_1 = {maskDestinationResult_hi_hi_hi, maskDestinationResult_hi_hi_lo};
  wire [63:0]  maskDestinationResult_hi_57 = {maskDestinationResult_hi_hi_1, maskDestinationResult_hi_lo_1};
  wire [1:0]   maskDestinationResult_lo_58 = {sourceDataVec_1[0], sourceDataVec_0[0]};
  wire [1:0]   maskDestinationResult_hi_58 = {sourceDataVec_3[0], sourceDataVec_2[0]};
  wire [1:0]   maskDestinationResult_lo_59 = {sourceDataVec_1[1], sourceDataVec_0[1]};
  wire [1:0]   maskDestinationResult_hi_59 = {sourceDataVec_3[1], sourceDataVec_2[1]};
  wire [1:0]   maskDestinationResult_lo_60 = {sourceDataVec_1[2], sourceDataVec_0[2]};
  wire [1:0]   maskDestinationResult_hi_60 = {sourceDataVec_3[2], sourceDataVec_2[2]};
  wire [1:0]   maskDestinationResult_lo_61 = {sourceDataVec_1[3], sourceDataVec_0[3]};
  wire [1:0]   maskDestinationResult_hi_61 = {sourceDataVec_3[3], sourceDataVec_2[3]};
  wire [1:0]   maskDestinationResult_lo_62 = {sourceDataVec_1[4], sourceDataVec_0[4]};
  wire [1:0]   maskDestinationResult_hi_62 = {sourceDataVec_3[4], sourceDataVec_2[4]};
  wire [1:0]   maskDestinationResult_lo_63 = {sourceDataVec_1[5], sourceDataVec_0[5]};
  wire [1:0]   maskDestinationResult_hi_63 = {sourceDataVec_3[5], sourceDataVec_2[5]};
  wire [1:0]   maskDestinationResult_lo_64 = {sourceDataVec_1[6], sourceDataVec_0[6]};
  wire [1:0]   maskDestinationResult_hi_64 = {sourceDataVec_3[6], sourceDataVec_2[6]};
  wire [1:0]   maskDestinationResult_lo_65 = {sourceDataVec_1[7], sourceDataVec_0[7]};
  wire [1:0]   maskDestinationResult_hi_65 = {sourceDataVec_3[7], sourceDataVec_2[7]};
  wire [1:0]   maskDestinationResult_lo_66 = {sourceDataVec_1[8], sourceDataVec_0[8]};
  wire [1:0]   maskDestinationResult_hi_66 = {sourceDataVec_3[8], sourceDataVec_2[8]};
  wire [1:0]   maskDestinationResult_lo_67 = {sourceDataVec_1[9], sourceDataVec_0[9]};
  wire [1:0]   maskDestinationResult_hi_67 = {sourceDataVec_3[9], sourceDataVec_2[9]};
  wire [1:0]   maskDestinationResult_lo_68 = {sourceDataVec_1[10], sourceDataVec_0[10]};
  wire [1:0]   maskDestinationResult_hi_68 = {sourceDataVec_3[10], sourceDataVec_2[10]};
  wire [1:0]   maskDestinationResult_lo_69 = {sourceDataVec_1[11], sourceDataVec_0[11]};
  wire [1:0]   maskDestinationResult_hi_69 = {sourceDataVec_3[11], sourceDataVec_2[11]};
  wire [1:0]   maskDestinationResult_lo_70 = {sourceDataVec_1[12], sourceDataVec_0[12]};
  wire [1:0]   maskDestinationResult_hi_70 = {sourceDataVec_3[12], sourceDataVec_2[12]};
  wire [1:0]   maskDestinationResult_lo_71 = {sourceDataVec_1[13], sourceDataVec_0[13]};
  wire [1:0]   maskDestinationResult_hi_71 = {sourceDataVec_3[13], sourceDataVec_2[13]};
  wire [1:0]   maskDestinationResult_lo_72 = {sourceDataVec_1[14], sourceDataVec_0[14]};
  wire [1:0]   maskDestinationResult_hi_72 = {sourceDataVec_3[14], sourceDataVec_2[14]};
  wire [1:0]   maskDestinationResult_lo_73 = {sourceDataVec_1[15], sourceDataVec_0[15]};
  wire [1:0]   maskDestinationResult_hi_73 = {sourceDataVec_3[15], sourceDataVec_2[15]};
  wire [1:0]   maskDestinationResult_lo_74 = {sourceDataVec_1[16], sourceDataVec_0[16]};
  wire [1:0]   maskDestinationResult_hi_74 = {sourceDataVec_3[16], sourceDataVec_2[16]};
  wire [1:0]   maskDestinationResult_lo_75 = {sourceDataVec_1[17], sourceDataVec_0[17]};
  wire [1:0]   maskDestinationResult_hi_75 = {sourceDataVec_3[17], sourceDataVec_2[17]};
  wire [1:0]   maskDestinationResult_lo_76 = {sourceDataVec_1[18], sourceDataVec_0[18]};
  wire [1:0]   maskDestinationResult_hi_76 = {sourceDataVec_3[18], sourceDataVec_2[18]};
  wire [1:0]   maskDestinationResult_lo_77 = {sourceDataVec_1[19], sourceDataVec_0[19]};
  wire [1:0]   maskDestinationResult_hi_77 = {sourceDataVec_3[19], sourceDataVec_2[19]};
  wire [1:0]   maskDestinationResult_lo_78 = {sourceDataVec_1[20], sourceDataVec_0[20]};
  wire [1:0]   maskDestinationResult_hi_78 = {sourceDataVec_3[20], sourceDataVec_2[20]};
  wire [1:0]   maskDestinationResult_lo_79 = {sourceDataVec_1[21], sourceDataVec_0[21]};
  wire [1:0]   maskDestinationResult_hi_79 = {sourceDataVec_3[21], sourceDataVec_2[21]};
  wire [1:0]   maskDestinationResult_lo_80 = {sourceDataVec_1[22], sourceDataVec_0[22]};
  wire [1:0]   maskDestinationResult_hi_80 = {sourceDataVec_3[22], sourceDataVec_2[22]};
  wire [1:0]   maskDestinationResult_lo_81 = {sourceDataVec_1[23], sourceDataVec_0[23]};
  wire [1:0]   maskDestinationResult_hi_81 = {sourceDataVec_3[23], sourceDataVec_2[23]};
  wire [1:0]   maskDestinationResult_lo_82 = {sourceDataVec_1[24], sourceDataVec_0[24]};
  wire [1:0]   maskDestinationResult_hi_82 = {sourceDataVec_3[24], sourceDataVec_2[24]};
  wire [1:0]   maskDestinationResult_lo_83 = {sourceDataVec_1[25], sourceDataVec_0[25]};
  wire [1:0]   maskDestinationResult_hi_83 = {sourceDataVec_3[25], sourceDataVec_2[25]};
  wire [1:0]   maskDestinationResult_lo_84 = {sourceDataVec_1[26], sourceDataVec_0[26]};
  wire [1:0]   maskDestinationResult_hi_84 = {sourceDataVec_3[26], sourceDataVec_2[26]};
  wire [1:0]   maskDestinationResult_lo_85 = {sourceDataVec_1[27], sourceDataVec_0[27]};
  wire [1:0]   maskDestinationResult_hi_85 = {sourceDataVec_3[27], sourceDataVec_2[27]};
  wire [1:0]   maskDestinationResult_lo_86 = {sourceDataVec_1[28], sourceDataVec_0[28]};
  wire [1:0]   maskDestinationResult_hi_86 = {sourceDataVec_3[28], sourceDataVec_2[28]};
  wire [1:0]   maskDestinationResult_lo_87 = {sourceDataVec_1[29], sourceDataVec_0[29]};
  wire [1:0]   maskDestinationResult_hi_87 = {sourceDataVec_3[29], sourceDataVec_2[29]};
  wire [1:0]   maskDestinationResult_lo_88 = {sourceDataVec_1[30], sourceDataVec_0[30]};
  wire [1:0]   maskDestinationResult_hi_88 = {sourceDataVec_3[30], sourceDataVec_2[30]};
  wire [1:0]   maskDestinationResult_lo_89 = {sourceDataVec_1[31], sourceDataVec_0[31]};
  wire [1:0]   maskDestinationResult_hi_89 = {sourceDataVec_3[31], sourceDataVec_2[31]};
  wire [7:0]   maskDestinationResult_lo_lo_lo_lo = {maskDestinationResult_hi_59, maskDestinationResult_lo_59, maskDestinationResult_hi_58, maskDestinationResult_lo_58};
  wire [7:0]   maskDestinationResult_lo_lo_lo_hi = {maskDestinationResult_hi_61, maskDestinationResult_lo_61, maskDestinationResult_hi_60, maskDestinationResult_lo_60};
  wire [15:0]  maskDestinationResult_lo_lo_lo_1 = {maskDestinationResult_lo_lo_lo_hi, maskDestinationResult_lo_lo_lo_lo};
  wire [7:0]   maskDestinationResult_lo_lo_hi_lo = {maskDestinationResult_hi_63, maskDestinationResult_lo_63, maskDestinationResult_hi_62, maskDestinationResult_lo_62};
  wire [7:0]   maskDestinationResult_lo_lo_hi_hi = {maskDestinationResult_hi_65, maskDestinationResult_lo_65, maskDestinationResult_hi_64, maskDestinationResult_lo_64};
  wire [15:0]  maskDestinationResult_lo_lo_hi_1 = {maskDestinationResult_lo_lo_hi_hi, maskDestinationResult_lo_lo_hi_lo};
  wire [31:0]  maskDestinationResult_lo_lo_2 = {maskDestinationResult_lo_lo_hi_1, maskDestinationResult_lo_lo_lo_1};
  wire [7:0]   maskDestinationResult_lo_hi_lo_lo = {maskDestinationResult_hi_67, maskDestinationResult_lo_67, maskDestinationResult_hi_66, maskDestinationResult_lo_66};
  wire [7:0]   maskDestinationResult_lo_hi_lo_hi = {maskDestinationResult_hi_69, maskDestinationResult_lo_69, maskDestinationResult_hi_68, maskDestinationResult_lo_68};
  wire [15:0]  maskDestinationResult_lo_hi_lo_1 = {maskDestinationResult_lo_hi_lo_hi, maskDestinationResult_lo_hi_lo_lo};
  wire [7:0]   maskDestinationResult_lo_hi_hi_lo = {maskDestinationResult_hi_71, maskDestinationResult_lo_71, maskDestinationResult_hi_70, maskDestinationResult_lo_70};
  wire [7:0]   maskDestinationResult_lo_hi_hi_hi = {maskDestinationResult_hi_73, maskDestinationResult_lo_73, maskDestinationResult_hi_72, maskDestinationResult_lo_72};
  wire [15:0]  maskDestinationResult_lo_hi_hi_1 = {maskDestinationResult_lo_hi_hi_hi, maskDestinationResult_lo_hi_hi_lo};
  wire [31:0]  maskDestinationResult_lo_hi_2 = {maskDestinationResult_lo_hi_hi_1, maskDestinationResult_lo_hi_lo_1};
  wire [63:0]  maskDestinationResult_lo_90 = {maskDestinationResult_lo_hi_2, maskDestinationResult_lo_lo_2};
  wire [7:0]   maskDestinationResult_hi_lo_lo_lo = {maskDestinationResult_hi_75, maskDestinationResult_lo_75, maskDestinationResult_hi_74, maskDestinationResult_lo_74};
  wire [7:0]   maskDestinationResult_hi_lo_lo_hi = {maskDestinationResult_hi_77, maskDestinationResult_lo_77, maskDestinationResult_hi_76, maskDestinationResult_lo_76};
  wire [15:0]  maskDestinationResult_hi_lo_lo_1 = {maskDestinationResult_hi_lo_lo_hi, maskDestinationResult_hi_lo_lo_lo};
  wire [7:0]   maskDestinationResult_hi_lo_hi_lo = {maskDestinationResult_hi_79, maskDestinationResult_lo_79, maskDestinationResult_hi_78, maskDestinationResult_lo_78};
  wire [7:0]   maskDestinationResult_hi_lo_hi_hi = {maskDestinationResult_hi_81, maskDestinationResult_lo_81, maskDestinationResult_hi_80, maskDestinationResult_lo_80};
  wire [15:0]  maskDestinationResult_hi_lo_hi_1 = {maskDestinationResult_hi_lo_hi_hi, maskDestinationResult_hi_lo_hi_lo};
  wire [31:0]  maskDestinationResult_hi_lo_2 = {maskDestinationResult_hi_lo_hi_1, maskDestinationResult_hi_lo_lo_1};
  wire [7:0]   maskDestinationResult_hi_hi_lo_lo = {maskDestinationResult_hi_83, maskDestinationResult_lo_83, maskDestinationResult_hi_82, maskDestinationResult_lo_82};
  wire [7:0]   maskDestinationResult_hi_hi_lo_hi = {maskDestinationResult_hi_85, maskDestinationResult_lo_85, maskDestinationResult_hi_84, maskDestinationResult_lo_84};
  wire [15:0]  maskDestinationResult_hi_hi_lo_1 = {maskDestinationResult_hi_hi_lo_hi, maskDestinationResult_hi_hi_lo_lo};
  wire [7:0]   maskDestinationResult_hi_hi_hi_lo = {maskDestinationResult_hi_87, maskDestinationResult_lo_87, maskDestinationResult_hi_86, maskDestinationResult_lo_86};
  wire [7:0]   maskDestinationResult_hi_hi_hi_hi = {maskDestinationResult_hi_89, maskDestinationResult_lo_89, maskDestinationResult_hi_88, maskDestinationResult_lo_88};
  wire [15:0]  maskDestinationResult_hi_hi_hi_1 = {maskDestinationResult_hi_hi_hi_hi, maskDestinationResult_hi_hi_hi_lo};
  wire [31:0]  maskDestinationResult_hi_hi_2 = {maskDestinationResult_hi_hi_hi_1, maskDestinationResult_hi_hi_lo_1};
  wire [63:0]  maskDestinationResult_hi_90 = {maskDestinationResult_hi_hi_2, maskDestinationResult_hi_lo_2};
  wire [127:0] maskDestinationResult =
    (eew1H[0] ? {maskDestinationResult_hi_40, maskDestinationResult_lo_40} : 128'h0) | (eew1H[1] ? {maskDestinationResult_hi_57, maskDestinationResult_lo_57} : 128'h0)
    | (eew1H[2] ? {maskDestinationResult_hi_90, maskDestinationResult_lo_90} : 128'h0);
  wire         sign = in_uop[0];
  wire         extendRatio = in_uop[2];
  wire [3:0]   _source2_T_1 = 4'h1 << in_groupCounter[1:0];
  wire [1:0]   _source2_T_18 = 2'h1 << in_groupCounter[0];
  wire [63:0]  source2 =
    extendRatio
      ? {32'h0, (_source2_T_1[0] ? sourceDataVec_0 : 32'h0) | (_source2_T_1[1] ? sourceDataVec_1 : 32'h0) | (_source2_T_1[2] ? sourceDataVec_2 : 32'h0) | (_source2_T_1[3] ? sourceDataVec_3 : 32'h0)}
      : (_source2_T_18[0] ? in_source2[63:0] : 64'h0) | (_source2_T_18[1] ? in_source2[127:64] : 64'h0);
  wire [1:0]   _extendResult_T_129 = 2'h1 << extendRatio;
  wire [31:0]  extendResult_lo_lo = {{8{source2[15] & sign}}, source2[15:8], {8{source2[7] & sign}}, source2[7:0]};
  wire [31:0]  extendResult_lo_hi = {{8{source2[31] & sign}}, source2[31:24], {8{source2[23] & sign}}, source2[23:16]};
  wire [63:0]  extendResult_lo = {extendResult_lo_hi, extendResult_lo_lo};
  wire [31:0]  extendResult_hi_lo = {{8{source2[47] & sign}}, source2[47:40], {8{source2[39] & sign}}, source2[39:32]};
  wire [31:0]  extendResult_hi_hi = {{8{source2[63] & sign}}, source2[63:56], {8{source2[55] & sign}}, source2[55:48]};
  wire [63:0]  extendResult_hi = {extendResult_hi_hi, extendResult_hi_lo};
  wire [31:0]  extendResult_lo_lo_lo = {{12{source2[7] & sign}}, source2[7:4], {12{source2[3] & sign}}, source2[3:0]};
  wire [31:0]  extendResult_lo_lo_hi = {{12{source2[15] & sign}}, source2[15:12], {12{source2[11] & sign}}, source2[11:8]};
  wire [63:0]  extendResult_lo_lo_1 = {extendResult_lo_lo_hi, extendResult_lo_lo_lo};
  wire [31:0]  extendResult_lo_hi_lo = {{12{source2[23] & sign}}, source2[23:20], {12{source2[19] & sign}}, source2[19:16]};
  wire [31:0]  extendResult_lo_hi_hi = {{12{source2[31] & sign}}, source2[31:28], {12{source2[27] & sign}}, source2[27:24]};
  wire [63:0]  extendResult_lo_hi_1 = {extendResult_lo_hi_hi, extendResult_lo_hi_lo};
  wire [127:0] extendResult_lo_1 = {extendResult_lo_hi_1, extendResult_lo_lo_1};
  wire [31:0]  extendResult_hi_lo_lo = {{12{source2[39] & sign}}, source2[39:36], {12{source2[35] & sign}}, source2[35:32]};
  wire [31:0]  extendResult_hi_lo_hi = {{12{source2[47] & sign}}, source2[47:44], {12{source2[43] & sign}}, source2[43:40]};
  wire [63:0]  extendResult_hi_lo_1 = {extendResult_hi_lo_hi, extendResult_hi_lo_lo};
  wire [31:0]  extendResult_hi_hi_lo = {{12{source2[55] & sign}}, source2[55:52], {12{source2[51] & sign}}, source2[51:48]};
  wire [31:0]  extendResult_hi_hi_hi = {{12{source2[63] & sign}}, source2[63:60], {12{source2[59] & sign}}, source2[59:56]};
  wire [63:0]  extendResult_hi_hi_1 = {extendResult_hi_hi_hi, extendResult_hi_hi_lo};
  wire [127:0] extendResult_hi_1 = {extendResult_hi_hi_1, extendResult_hi_lo_1};
  wire [63:0]  extendResult_lo_2 = {{16{source2[31] & sign}}, source2[31:16], {16{source2[15] & sign}}, source2[15:0]};
  wire [63:0]  extendResult_hi_2 = {{16{source2[63] & sign}}, source2[63:48], {16{source2[47] & sign}}, source2[47:32]};
  wire [63:0]  extendResult_lo_lo_2 = {{24{source2[15] & sign}}, source2[15:8], {24{source2[7] & sign}}, source2[7:0]};
  wire [63:0]  extendResult_lo_hi_2 = {{24{source2[31] & sign}}, source2[31:24], {24{source2[23] & sign}}, source2[23:16]};
  wire [127:0] extendResult_lo_3 = {extendResult_lo_hi_2, extendResult_lo_lo_2};
  wire [63:0]  extendResult_hi_lo_2 = {{24{source2[47] & sign}}, source2[47:40], {24{source2[39] & sign}}, source2[39:32]};
  wire [63:0]  extendResult_hi_hi_2 = {{24{source2[63] & sign}}, source2[63:56], {24{source2[55] & sign}}, source2[55:48]};
  wire [127:0] extendResult_hi_3 = {extendResult_hi_hi_2, extendResult_hi_lo_2};
  wire [255:0] extendResult =
    (eew1H[1] ? {128'h0, _extendResult_T_129[0] ? {extendResult_hi, extendResult_lo} : 128'h0} | (_extendResult_T_129[1] ? {extendResult_hi_1, extendResult_lo_1} : 256'h0) : 256'h0)
    | (eew1H[2] ? {128'h0, _extendResult_T_129[0] ? {extendResult_hi_2, extendResult_lo_2} : 128'h0} | (_extendResult_T_129[1] ? {extendResult_hi_3, extendResult_lo_3} : 256'h0) : 256'h0);
  assign out = isMaskDestination ? maskDestinationResult : extendResult[127:0];
endmodule

