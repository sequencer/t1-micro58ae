module MaskExtend(
  input  [1:0]   in_eew,
  input  [2:0]   in_uop,
  input  [255:0] in_source2,
  input  [5:0]   in_groupCounter,
  output [255:0] out
);

  wire [3:0]   _eew1H_T = 4'h1 << in_eew;
  wire [2:0]   eew1H = _eew1H_T[2:0];
  wire         isMaskDestination = in_uop == 3'h0;
  wire [31:0]  sourceDataVec_0 = in_source2[31:0];
  wire [31:0]  sourceDataVec_1 = in_source2[63:32];
  wire [31:0]  sourceDataVec_2 = in_source2[95:64];
  wire [31:0]  sourceDataVec_3 = in_source2[127:96];
  wire [31:0]  sourceDataVec_4 = in_source2[159:128];
  wire [31:0]  sourceDataVec_5 = in_source2[191:160];
  wire [31:0]  sourceDataVec_6 = in_source2[223:192];
  wire [31:0]  sourceDataVec_7 = in_source2[255:224];
  wire [1:0]   maskDestinationResult_lo = sourceDataVec_0[1:0];
  wire [1:0]   maskDestinationResult_hi = sourceDataVec_0[3:2];
  wire [1:0]   maskDestinationResult_lo_1 = sourceDataVec_0[5:4];
  wire [1:0]   maskDestinationResult_hi_1 = sourceDataVec_0[7:6];
  wire [1:0]   maskDestinationResult_lo_2 = sourceDataVec_0[9:8];
  wire [1:0]   maskDestinationResult_hi_2 = sourceDataVec_0[11:10];
  wire [1:0]   maskDestinationResult_lo_3 = sourceDataVec_0[13:12];
  wire [1:0]   maskDestinationResult_hi_3 = sourceDataVec_0[15:14];
  wire [1:0]   maskDestinationResult_lo_4 = sourceDataVec_0[17:16];
  wire [1:0]   maskDestinationResult_hi_4 = sourceDataVec_0[19:18];
  wire [1:0]   maskDestinationResult_lo_5 = sourceDataVec_0[21:20];
  wire [1:0]   maskDestinationResult_hi_5 = sourceDataVec_0[23:22];
  wire [1:0]   maskDestinationResult_lo_6 = sourceDataVec_0[25:24];
  wire [1:0]   maskDestinationResult_hi_6 = sourceDataVec_0[27:26];
  wire [1:0]   maskDestinationResult_lo_7 = sourceDataVec_0[29:28];
  wire [1:0]   maskDestinationResult_hi_7 = sourceDataVec_0[31:30];
  wire [1:0]   maskDestinationResult_lo_8 = sourceDataVec_1[1:0];
  wire [1:0]   maskDestinationResult_hi_8 = sourceDataVec_1[3:2];
  wire [1:0]   maskDestinationResult_lo_9 = sourceDataVec_1[5:4];
  wire [1:0]   maskDestinationResult_hi_9 = sourceDataVec_1[7:6];
  wire [1:0]   maskDestinationResult_lo_10 = sourceDataVec_1[9:8];
  wire [1:0]   maskDestinationResult_hi_10 = sourceDataVec_1[11:10];
  wire [1:0]   maskDestinationResult_lo_11 = sourceDataVec_1[13:12];
  wire [1:0]   maskDestinationResult_hi_11 = sourceDataVec_1[15:14];
  wire [1:0]   maskDestinationResult_lo_12 = sourceDataVec_1[17:16];
  wire [1:0]   maskDestinationResult_hi_12 = sourceDataVec_1[19:18];
  wire [1:0]   maskDestinationResult_lo_13 = sourceDataVec_1[21:20];
  wire [1:0]   maskDestinationResult_hi_13 = sourceDataVec_1[23:22];
  wire [1:0]   maskDestinationResult_lo_14 = sourceDataVec_1[25:24];
  wire [1:0]   maskDestinationResult_hi_14 = sourceDataVec_1[27:26];
  wire [1:0]   maskDestinationResult_lo_15 = sourceDataVec_1[29:28];
  wire [1:0]   maskDestinationResult_hi_15 = sourceDataVec_1[31:30];
  wire [1:0]   maskDestinationResult_lo_16 = sourceDataVec_2[1:0];
  wire [1:0]   maskDestinationResult_hi_16 = sourceDataVec_2[3:2];
  wire [1:0]   maskDestinationResult_lo_17 = sourceDataVec_2[5:4];
  wire [1:0]   maskDestinationResult_hi_17 = sourceDataVec_2[7:6];
  wire [1:0]   maskDestinationResult_lo_18 = sourceDataVec_2[9:8];
  wire [1:0]   maskDestinationResult_hi_18 = sourceDataVec_2[11:10];
  wire [1:0]   maskDestinationResult_lo_19 = sourceDataVec_2[13:12];
  wire [1:0]   maskDestinationResult_hi_19 = sourceDataVec_2[15:14];
  wire [1:0]   maskDestinationResult_lo_20 = sourceDataVec_2[17:16];
  wire [1:0]   maskDestinationResult_hi_20 = sourceDataVec_2[19:18];
  wire [1:0]   maskDestinationResult_lo_21 = sourceDataVec_2[21:20];
  wire [1:0]   maskDestinationResult_hi_21 = sourceDataVec_2[23:22];
  wire [1:0]   maskDestinationResult_lo_22 = sourceDataVec_2[25:24];
  wire [1:0]   maskDestinationResult_hi_22 = sourceDataVec_2[27:26];
  wire [1:0]   maskDestinationResult_lo_23 = sourceDataVec_2[29:28];
  wire [1:0]   maskDestinationResult_hi_23 = sourceDataVec_2[31:30];
  wire [1:0]   maskDestinationResult_lo_24 = sourceDataVec_3[1:0];
  wire [1:0]   maskDestinationResult_hi_24 = sourceDataVec_3[3:2];
  wire [1:0]   maskDestinationResult_lo_25 = sourceDataVec_3[5:4];
  wire [1:0]   maskDestinationResult_hi_25 = sourceDataVec_3[7:6];
  wire [1:0]   maskDestinationResult_lo_26 = sourceDataVec_3[9:8];
  wire [1:0]   maskDestinationResult_hi_26 = sourceDataVec_3[11:10];
  wire [1:0]   maskDestinationResult_lo_27 = sourceDataVec_3[13:12];
  wire [1:0]   maskDestinationResult_hi_27 = sourceDataVec_3[15:14];
  wire [1:0]   maskDestinationResult_lo_28 = sourceDataVec_3[17:16];
  wire [1:0]   maskDestinationResult_hi_28 = sourceDataVec_3[19:18];
  wire [1:0]   maskDestinationResult_lo_29 = sourceDataVec_3[21:20];
  wire [1:0]   maskDestinationResult_hi_29 = sourceDataVec_3[23:22];
  wire [1:0]   maskDestinationResult_lo_30 = sourceDataVec_3[25:24];
  wire [1:0]   maskDestinationResult_hi_30 = sourceDataVec_3[27:26];
  wire [1:0]   maskDestinationResult_lo_31 = sourceDataVec_3[29:28];
  wire [1:0]   maskDestinationResult_hi_31 = sourceDataVec_3[31:30];
  wire [1:0]   maskDestinationResult_lo_32 = sourceDataVec_4[1:0];
  wire [1:0]   maskDestinationResult_hi_32 = sourceDataVec_4[3:2];
  wire [1:0]   maskDestinationResult_lo_33 = sourceDataVec_4[5:4];
  wire [1:0]   maskDestinationResult_hi_33 = sourceDataVec_4[7:6];
  wire [1:0]   maskDestinationResult_lo_34 = sourceDataVec_4[9:8];
  wire [1:0]   maskDestinationResult_hi_34 = sourceDataVec_4[11:10];
  wire [1:0]   maskDestinationResult_lo_35 = sourceDataVec_4[13:12];
  wire [1:0]   maskDestinationResult_hi_35 = sourceDataVec_4[15:14];
  wire [1:0]   maskDestinationResult_lo_36 = sourceDataVec_4[17:16];
  wire [1:0]   maskDestinationResult_hi_36 = sourceDataVec_4[19:18];
  wire [1:0]   maskDestinationResult_lo_37 = sourceDataVec_4[21:20];
  wire [1:0]   maskDestinationResult_hi_37 = sourceDataVec_4[23:22];
  wire [1:0]   maskDestinationResult_lo_38 = sourceDataVec_4[25:24];
  wire [1:0]   maskDestinationResult_hi_38 = sourceDataVec_4[27:26];
  wire [1:0]   maskDestinationResult_lo_39 = sourceDataVec_4[29:28];
  wire [1:0]   maskDestinationResult_hi_39 = sourceDataVec_4[31:30];
  wire [1:0]   maskDestinationResult_lo_40 = sourceDataVec_5[1:0];
  wire [1:0]   maskDestinationResult_hi_40 = sourceDataVec_5[3:2];
  wire [1:0]   maskDestinationResult_lo_41 = sourceDataVec_5[5:4];
  wire [1:0]   maskDestinationResult_hi_41 = sourceDataVec_5[7:6];
  wire [1:0]   maskDestinationResult_lo_42 = sourceDataVec_5[9:8];
  wire [1:0]   maskDestinationResult_hi_42 = sourceDataVec_5[11:10];
  wire [1:0]   maskDestinationResult_lo_43 = sourceDataVec_5[13:12];
  wire [1:0]   maskDestinationResult_hi_43 = sourceDataVec_5[15:14];
  wire [1:0]   maskDestinationResult_lo_44 = sourceDataVec_5[17:16];
  wire [1:0]   maskDestinationResult_hi_44 = sourceDataVec_5[19:18];
  wire [1:0]   maskDestinationResult_lo_45 = sourceDataVec_5[21:20];
  wire [1:0]   maskDestinationResult_hi_45 = sourceDataVec_5[23:22];
  wire [1:0]   maskDestinationResult_lo_46 = sourceDataVec_5[25:24];
  wire [1:0]   maskDestinationResult_hi_46 = sourceDataVec_5[27:26];
  wire [1:0]   maskDestinationResult_lo_47 = sourceDataVec_5[29:28];
  wire [1:0]   maskDestinationResult_hi_47 = sourceDataVec_5[31:30];
  wire [1:0]   maskDestinationResult_lo_48 = sourceDataVec_6[1:0];
  wire [1:0]   maskDestinationResult_hi_48 = sourceDataVec_6[3:2];
  wire [1:0]   maskDestinationResult_lo_49 = sourceDataVec_6[5:4];
  wire [1:0]   maskDestinationResult_hi_49 = sourceDataVec_6[7:6];
  wire [1:0]   maskDestinationResult_lo_50 = sourceDataVec_6[9:8];
  wire [1:0]   maskDestinationResult_hi_50 = sourceDataVec_6[11:10];
  wire [1:0]   maskDestinationResult_lo_51 = sourceDataVec_6[13:12];
  wire [1:0]   maskDestinationResult_hi_51 = sourceDataVec_6[15:14];
  wire [1:0]   maskDestinationResult_lo_52 = sourceDataVec_6[17:16];
  wire [1:0]   maskDestinationResult_hi_52 = sourceDataVec_6[19:18];
  wire [1:0]   maskDestinationResult_lo_53 = sourceDataVec_6[21:20];
  wire [1:0]   maskDestinationResult_hi_53 = sourceDataVec_6[23:22];
  wire [1:0]   maskDestinationResult_lo_54 = sourceDataVec_6[25:24];
  wire [1:0]   maskDestinationResult_hi_54 = sourceDataVec_6[27:26];
  wire [1:0]   maskDestinationResult_lo_55 = sourceDataVec_6[29:28];
  wire [1:0]   maskDestinationResult_hi_55 = sourceDataVec_6[31:30];
  wire [1:0]   maskDestinationResult_lo_56 = sourceDataVec_7[1:0];
  wire [1:0]   maskDestinationResult_hi_56 = sourceDataVec_7[3:2];
  wire [1:0]   maskDestinationResult_lo_57 = sourceDataVec_7[5:4];
  wire [1:0]   maskDestinationResult_hi_57 = sourceDataVec_7[7:6];
  wire [1:0]   maskDestinationResult_lo_58 = sourceDataVec_7[9:8];
  wire [1:0]   maskDestinationResult_hi_58 = sourceDataVec_7[11:10];
  wire [1:0]   maskDestinationResult_lo_59 = sourceDataVec_7[13:12];
  wire [1:0]   maskDestinationResult_hi_59 = sourceDataVec_7[15:14];
  wire [1:0]   maskDestinationResult_lo_60 = sourceDataVec_7[17:16];
  wire [1:0]   maskDestinationResult_hi_60 = sourceDataVec_7[19:18];
  wire [1:0]   maskDestinationResult_lo_61 = sourceDataVec_7[21:20];
  wire [1:0]   maskDestinationResult_hi_61 = sourceDataVec_7[23:22];
  wire [1:0]   maskDestinationResult_lo_62 = sourceDataVec_7[25:24];
  wire [1:0]   maskDestinationResult_hi_62 = sourceDataVec_7[27:26];
  wire [1:0]   maskDestinationResult_lo_63 = sourceDataVec_7[29:28];
  wire [1:0]   maskDestinationResult_hi_63 = sourceDataVec_7[31:30];
  wire [7:0]   maskDestinationResult_lo_lo = {maskDestinationResult_hi_8, maskDestinationResult_lo_8, maskDestinationResult_hi, maskDestinationResult_lo};
  wire [7:0]   maskDestinationResult_lo_hi = {maskDestinationResult_hi_24, maskDestinationResult_lo_24, maskDestinationResult_hi_16, maskDestinationResult_lo_16};
  wire [15:0]  maskDestinationResult_lo_64 = {maskDestinationResult_lo_hi, maskDestinationResult_lo_lo};
  wire [7:0]   maskDestinationResult_hi_lo = {maskDestinationResult_hi_40, maskDestinationResult_lo_40, maskDestinationResult_hi_32, maskDestinationResult_lo_32};
  wire [7:0]   maskDestinationResult_hi_hi = {maskDestinationResult_hi_56, maskDestinationResult_lo_56, maskDestinationResult_hi_48, maskDestinationResult_lo_48};
  wire [15:0]  maskDestinationResult_hi_64 = {maskDestinationResult_hi_hi, maskDestinationResult_hi_lo};
  wire [7:0]   maskDestinationResult_lo_lo_1 = {maskDestinationResult_hi_9, maskDestinationResult_lo_9, maskDestinationResult_hi_1, maskDestinationResult_lo_1};
  wire [7:0]   maskDestinationResult_lo_hi_1 = {maskDestinationResult_hi_25, maskDestinationResult_lo_25, maskDestinationResult_hi_17, maskDestinationResult_lo_17};
  wire [15:0]  maskDestinationResult_lo_65 = {maskDestinationResult_lo_hi_1, maskDestinationResult_lo_lo_1};
  wire [7:0]   maskDestinationResult_hi_lo_1 = {maskDestinationResult_hi_41, maskDestinationResult_lo_41, maskDestinationResult_hi_33, maskDestinationResult_lo_33};
  wire [7:0]   maskDestinationResult_hi_hi_1 = {maskDestinationResult_hi_57, maskDestinationResult_lo_57, maskDestinationResult_hi_49, maskDestinationResult_lo_49};
  wire [15:0]  maskDestinationResult_hi_65 = {maskDestinationResult_hi_hi_1, maskDestinationResult_hi_lo_1};
  wire [7:0]   maskDestinationResult_lo_lo_2 = {maskDestinationResult_hi_10, maskDestinationResult_lo_10, maskDestinationResult_hi_2, maskDestinationResult_lo_2};
  wire [7:0]   maskDestinationResult_lo_hi_2 = {maskDestinationResult_hi_26, maskDestinationResult_lo_26, maskDestinationResult_hi_18, maskDestinationResult_lo_18};
  wire [15:0]  maskDestinationResult_lo_66 = {maskDestinationResult_lo_hi_2, maskDestinationResult_lo_lo_2};
  wire [7:0]   maskDestinationResult_hi_lo_2 = {maskDestinationResult_hi_42, maskDestinationResult_lo_42, maskDestinationResult_hi_34, maskDestinationResult_lo_34};
  wire [7:0]   maskDestinationResult_hi_hi_2 = {maskDestinationResult_hi_58, maskDestinationResult_lo_58, maskDestinationResult_hi_50, maskDestinationResult_lo_50};
  wire [15:0]  maskDestinationResult_hi_66 = {maskDestinationResult_hi_hi_2, maskDestinationResult_hi_lo_2};
  wire [7:0]   maskDestinationResult_lo_lo_3 = {maskDestinationResult_hi_11, maskDestinationResult_lo_11, maskDestinationResult_hi_3, maskDestinationResult_lo_3};
  wire [7:0]   maskDestinationResult_lo_hi_3 = {maskDestinationResult_hi_27, maskDestinationResult_lo_27, maskDestinationResult_hi_19, maskDestinationResult_lo_19};
  wire [15:0]  maskDestinationResult_lo_67 = {maskDestinationResult_lo_hi_3, maskDestinationResult_lo_lo_3};
  wire [7:0]   maskDestinationResult_hi_lo_3 = {maskDestinationResult_hi_43, maskDestinationResult_lo_43, maskDestinationResult_hi_35, maskDestinationResult_lo_35};
  wire [7:0]   maskDestinationResult_hi_hi_3 = {maskDestinationResult_hi_59, maskDestinationResult_lo_59, maskDestinationResult_hi_51, maskDestinationResult_lo_51};
  wire [15:0]  maskDestinationResult_hi_67 = {maskDestinationResult_hi_hi_3, maskDestinationResult_hi_lo_3};
  wire [7:0]   maskDestinationResult_lo_lo_4 = {maskDestinationResult_hi_12, maskDestinationResult_lo_12, maskDestinationResult_hi_4, maskDestinationResult_lo_4};
  wire [7:0]   maskDestinationResult_lo_hi_4 = {maskDestinationResult_hi_28, maskDestinationResult_lo_28, maskDestinationResult_hi_20, maskDestinationResult_lo_20};
  wire [15:0]  maskDestinationResult_lo_68 = {maskDestinationResult_lo_hi_4, maskDestinationResult_lo_lo_4};
  wire [7:0]   maskDestinationResult_hi_lo_4 = {maskDestinationResult_hi_44, maskDestinationResult_lo_44, maskDestinationResult_hi_36, maskDestinationResult_lo_36};
  wire [7:0]   maskDestinationResult_hi_hi_4 = {maskDestinationResult_hi_60, maskDestinationResult_lo_60, maskDestinationResult_hi_52, maskDestinationResult_lo_52};
  wire [15:0]  maskDestinationResult_hi_68 = {maskDestinationResult_hi_hi_4, maskDestinationResult_hi_lo_4};
  wire [7:0]   maskDestinationResult_lo_lo_5 = {maskDestinationResult_hi_13, maskDestinationResult_lo_13, maskDestinationResult_hi_5, maskDestinationResult_lo_5};
  wire [7:0]   maskDestinationResult_lo_hi_5 = {maskDestinationResult_hi_29, maskDestinationResult_lo_29, maskDestinationResult_hi_21, maskDestinationResult_lo_21};
  wire [15:0]  maskDestinationResult_lo_69 = {maskDestinationResult_lo_hi_5, maskDestinationResult_lo_lo_5};
  wire [7:0]   maskDestinationResult_hi_lo_5 = {maskDestinationResult_hi_45, maskDestinationResult_lo_45, maskDestinationResult_hi_37, maskDestinationResult_lo_37};
  wire [7:0]   maskDestinationResult_hi_hi_5 = {maskDestinationResult_hi_61, maskDestinationResult_lo_61, maskDestinationResult_hi_53, maskDestinationResult_lo_53};
  wire [15:0]  maskDestinationResult_hi_69 = {maskDestinationResult_hi_hi_5, maskDestinationResult_hi_lo_5};
  wire [7:0]   maskDestinationResult_lo_lo_6 = {maskDestinationResult_hi_14, maskDestinationResult_lo_14, maskDestinationResult_hi_6, maskDestinationResult_lo_6};
  wire [7:0]   maskDestinationResult_lo_hi_6 = {maskDestinationResult_hi_30, maskDestinationResult_lo_30, maskDestinationResult_hi_22, maskDestinationResult_lo_22};
  wire [15:0]  maskDestinationResult_lo_70 = {maskDestinationResult_lo_hi_6, maskDestinationResult_lo_lo_6};
  wire [7:0]   maskDestinationResult_hi_lo_6 = {maskDestinationResult_hi_46, maskDestinationResult_lo_46, maskDestinationResult_hi_38, maskDestinationResult_lo_38};
  wire [7:0]   maskDestinationResult_hi_hi_6 = {maskDestinationResult_hi_62, maskDestinationResult_lo_62, maskDestinationResult_hi_54, maskDestinationResult_lo_54};
  wire [15:0]  maskDestinationResult_hi_70 = {maskDestinationResult_hi_hi_6, maskDestinationResult_hi_lo_6};
  wire [7:0]   maskDestinationResult_lo_lo_7 = {maskDestinationResult_hi_15, maskDestinationResult_lo_15, maskDestinationResult_hi_7, maskDestinationResult_lo_7};
  wire [7:0]   maskDestinationResult_lo_hi_7 = {maskDestinationResult_hi_31, maskDestinationResult_lo_31, maskDestinationResult_hi_23, maskDestinationResult_lo_23};
  wire [15:0]  maskDestinationResult_lo_71 = {maskDestinationResult_lo_hi_7, maskDestinationResult_lo_lo_7};
  wire [7:0]   maskDestinationResult_hi_lo_7 = {maskDestinationResult_hi_47, maskDestinationResult_lo_47, maskDestinationResult_hi_39, maskDestinationResult_lo_39};
  wire [7:0]   maskDestinationResult_hi_hi_7 = {maskDestinationResult_hi_63, maskDestinationResult_lo_63, maskDestinationResult_hi_55, maskDestinationResult_lo_55};
  wire [15:0]  maskDestinationResult_hi_71 = {maskDestinationResult_hi_hi_7, maskDestinationResult_hi_lo_7};
  wire [63:0]  maskDestinationResult_lo_lo_8 = {maskDestinationResult_hi_65, maskDestinationResult_lo_65, maskDestinationResult_hi_64, maskDestinationResult_lo_64};
  wire [63:0]  maskDestinationResult_lo_hi_8 = {maskDestinationResult_hi_67, maskDestinationResult_lo_67, maskDestinationResult_hi_66, maskDestinationResult_lo_66};
  wire [127:0] maskDestinationResult_lo_72 = {maskDestinationResult_lo_hi_8, maskDestinationResult_lo_lo_8};
  wire [63:0]  maskDestinationResult_hi_lo_8 = {maskDestinationResult_hi_69, maskDestinationResult_lo_69, maskDestinationResult_hi_68, maskDestinationResult_lo_68};
  wire [63:0]  maskDestinationResult_hi_hi_8 = {maskDestinationResult_hi_71, maskDestinationResult_lo_71, maskDestinationResult_hi_70, maskDestinationResult_lo_70};
  wire [127:0] maskDestinationResult_hi_72 = {maskDestinationResult_hi_hi_8, maskDestinationResult_hi_lo_8};
  wire [3:0]   maskDestinationResult_lo_lo_9 = {sourceDataVec_1[1:0], sourceDataVec_0[1:0]};
  wire [3:0]   maskDestinationResult_lo_hi_9 = {sourceDataVec_3[1:0], sourceDataVec_2[1:0]};
  wire [7:0]   maskDestinationResult_lo_73 = {maskDestinationResult_lo_hi_9, maskDestinationResult_lo_lo_9};
  wire [3:0]   maskDestinationResult_hi_lo_9 = {sourceDataVec_5[1:0], sourceDataVec_4[1:0]};
  wire [3:0]   maskDestinationResult_hi_hi_9 = {sourceDataVec_7[1:0], sourceDataVec_6[1:0]};
  wire [7:0]   maskDestinationResult_hi_73 = {maskDestinationResult_hi_hi_9, maskDestinationResult_hi_lo_9};
  wire [3:0]   maskDestinationResult_lo_lo_10 = {sourceDataVec_1[3:2], sourceDataVec_0[3:2]};
  wire [3:0]   maskDestinationResult_lo_hi_10 = {sourceDataVec_3[3:2], sourceDataVec_2[3:2]};
  wire [7:0]   maskDestinationResult_lo_74 = {maskDestinationResult_lo_hi_10, maskDestinationResult_lo_lo_10};
  wire [3:0]   maskDestinationResult_hi_lo_10 = {sourceDataVec_5[3:2], sourceDataVec_4[3:2]};
  wire [3:0]   maskDestinationResult_hi_hi_10 = {sourceDataVec_7[3:2], sourceDataVec_6[3:2]};
  wire [7:0]   maskDestinationResult_hi_74 = {maskDestinationResult_hi_hi_10, maskDestinationResult_hi_lo_10};
  wire [3:0]   maskDestinationResult_lo_lo_11 = {sourceDataVec_1[5:4], sourceDataVec_0[5:4]};
  wire [3:0]   maskDestinationResult_lo_hi_11 = {sourceDataVec_3[5:4], sourceDataVec_2[5:4]};
  wire [7:0]   maskDestinationResult_lo_75 = {maskDestinationResult_lo_hi_11, maskDestinationResult_lo_lo_11};
  wire [3:0]   maskDestinationResult_hi_lo_11 = {sourceDataVec_5[5:4], sourceDataVec_4[5:4]};
  wire [3:0]   maskDestinationResult_hi_hi_11 = {sourceDataVec_7[5:4], sourceDataVec_6[5:4]};
  wire [7:0]   maskDestinationResult_hi_75 = {maskDestinationResult_hi_hi_11, maskDestinationResult_hi_lo_11};
  wire [3:0]   maskDestinationResult_lo_lo_12 = {sourceDataVec_1[7:6], sourceDataVec_0[7:6]};
  wire [3:0]   maskDestinationResult_lo_hi_12 = {sourceDataVec_3[7:6], sourceDataVec_2[7:6]};
  wire [7:0]   maskDestinationResult_lo_76 = {maskDestinationResult_lo_hi_12, maskDestinationResult_lo_lo_12};
  wire [3:0]   maskDestinationResult_hi_lo_12 = {sourceDataVec_5[7:6], sourceDataVec_4[7:6]};
  wire [3:0]   maskDestinationResult_hi_hi_12 = {sourceDataVec_7[7:6], sourceDataVec_6[7:6]};
  wire [7:0]   maskDestinationResult_hi_76 = {maskDestinationResult_hi_hi_12, maskDestinationResult_hi_lo_12};
  wire [3:0]   maskDestinationResult_lo_lo_13 = {sourceDataVec_1[9:8], sourceDataVec_0[9:8]};
  wire [3:0]   maskDestinationResult_lo_hi_13 = {sourceDataVec_3[9:8], sourceDataVec_2[9:8]};
  wire [7:0]   maskDestinationResult_lo_77 = {maskDestinationResult_lo_hi_13, maskDestinationResult_lo_lo_13};
  wire [3:0]   maskDestinationResult_hi_lo_13 = {sourceDataVec_5[9:8], sourceDataVec_4[9:8]};
  wire [3:0]   maskDestinationResult_hi_hi_13 = {sourceDataVec_7[9:8], sourceDataVec_6[9:8]};
  wire [7:0]   maskDestinationResult_hi_77 = {maskDestinationResult_hi_hi_13, maskDestinationResult_hi_lo_13};
  wire [3:0]   maskDestinationResult_lo_lo_14 = {sourceDataVec_1[11:10], sourceDataVec_0[11:10]};
  wire [3:0]   maskDestinationResult_lo_hi_14 = {sourceDataVec_3[11:10], sourceDataVec_2[11:10]};
  wire [7:0]   maskDestinationResult_lo_78 = {maskDestinationResult_lo_hi_14, maskDestinationResult_lo_lo_14};
  wire [3:0]   maskDestinationResult_hi_lo_14 = {sourceDataVec_5[11:10], sourceDataVec_4[11:10]};
  wire [3:0]   maskDestinationResult_hi_hi_14 = {sourceDataVec_7[11:10], sourceDataVec_6[11:10]};
  wire [7:0]   maskDestinationResult_hi_78 = {maskDestinationResult_hi_hi_14, maskDestinationResult_hi_lo_14};
  wire [3:0]   maskDestinationResult_lo_lo_15 = {sourceDataVec_1[13:12], sourceDataVec_0[13:12]};
  wire [3:0]   maskDestinationResult_lo_hi_15 = {sourceDataVec_3[13:12], sourceDataVec_2[13:12]};
  wire [7:0]   maskDestinationResult_lo_79 = {maskDestinationResult_lo_hi_15, maskDestinationResult_lo_lo_15};
  wire [3:0]   maskDestinationResult_hi_lo_15 = {sourceDataVec_5[13:12], sourceDataVec_4[13:12]};
  wire [3:0]   maskDestinationResult_hi_hi_15 = {sourceDataVec_7[13:12], sourceDataVec_6[13:12]};
  wire [7:0]   maskDestinationResult_hi_79 = {maskDestinationResult_hi_hi_15, maskDestinationResult_hi_lo_15};
  wire [3:0]   maskDestinationResult_lo_lo_16 = {sourceDataVec_1[15:14], sourceDataVec_0[15:14]};
  wire [3:0]   maskDestinationResult_lo_hi_16 = {sourceDataVec_3[15:14], sourceDataVec_2[15:14]};
  wire [7:0]   maskDestinationResult_lo_80 = {maskDestinationResult_lo_hi_16, maskDestinationResult_lo_lo_16};
  wire [3:0]   maskDestinationResult_hi_lo_16 = {sourceDataVec_5[15:14], sourceDataVec_4[15:14]};
  wire [3:0]   maskDestinationResult_hi_hi_16 = {sourceDataVec_7[15:14], sourceDataVec_6[15:14]};
  wire [7:0]   maskDestinationResult_hi_80 = {maskDestinationResult_hi_hi_16, maskDestinationResult_hi_lo_16};
  wire [3:0]   maskDestinationResult_lo_lo_17 = {sourceDataVec_1[17:16], sourceDataVec_0[17:16]};
  wire [3:0]   maskDestinationResult_lo_hi_17 = {sourceDataVec_3[17:16], sourceDataVec_2[17:16]};
  wire [7:0]   maskDestinationResult_lo_81 = {maskDestinationResult_lo_hi_17, maskDestinationResult_lo_lo_17};
  wire [3:0]   maskDestinationResult_hi_lo_17 = {sourceDataVec_5[17:16], sourceDataVec_4[17:16]};
  wire [3:0]   maskDestinationResult_hi_hi_17 = {sourceDataVec_7[17:16], sourceDataVec_6[17:16]};
  wire [7:0]   maskDestinationResult_hi_81 = {maskDestinationResult_hi_hi_17, maskDestinationResult_hi_lo_17};
  wire [3:0]   maskDestinationResult_lo_lo_18 = {sourceDataVec_1[19:18], sourceDataVec_0[19:18]};
  wire [3:0]   maskDestinationResult_lo_hi_18 = {sourceDataVec_3[19:18], sourceDataVec_2[19:18]};
  wire [7:0]   maskDestinationResult_lo_82 = {maskDestinationResult_lo_hi_18, maskDestinationResult_lo_lo_18};
  wire [3:0]   maskDestinationResult_hi_lo_18 = {sourceDataVec_5[19:18], sourceDataVec_4[19:18]};
  wire [3:0]   maskDestinationResult_hi_hi_18 = {sourceDataVec_7[19:18], sourceDataVec_6[19:18]};
  wire [7:0]   maskDestinationResult_hi_82 = {maskDestinationResult_hi_hi_18, maskDestinationResult_hi_lo_18};
  wire [3:0]   maskDestinationResult_lo_lo_19 = {sourceDataVec_1[21:20], sourceDataVec_0[21:20]};
  wire [3:0]   maskDestinationResult_lo_hi_19 = {sourceDataVec_3[21:20], sourceDataVec_2[21:20]};
  wire [7:0]   maskDestinationResult_lo_83 = {maskDestinationResult_lo_hi_19, maskDestinationResult_lo_lo_19};
  wire [3:0]   maskDestinationResult_hi_lo_19 = {sourceDataVec_5[21:20], sourceDataVec_4[21:20]};
  wire [3:0]   maskDestinationResult_hi_hi_19 = {sourceDataVec_7[21:20], sourceDataVec_6[21:20]};
  wire [7:0]   maskDestinationResult_hi_83 = {maskDestinationResult_hi_hi_19, maskDestinationResult_hi_lo_19};
  wire [3:0]   maskDestinationResult_lo_lo_20 = {sourceDataVec_1[23:22], sourceDataVec_0[23:22]};
  wire [3:0]   maskDestinationResult_lo_hi_20 = {sourceDataVec_3[23:22], sourceDataVec_2[23:22]};
  wire [7:0]   maskDestinationResult_lo_84 = {maskDestinationResult_lo_hi_20, maskDestinationResult_lo_lo_20};
  wire [3:0]   maskDestinationResult_hi_lo_20 = {sourceDataVec_5[23:22], sourceDataVec_4[23:22]};
  wire [3:0]   maskDestinationResult_hi_hi_20 = {sourceDataVec_7[23:22], sourceDataVec_6[23:22]};
  wire [7:0]   maskDestinationResult_hi_84 = {maskDestinationResult_hi_hi_20, maskDestinationResult_hi_lo_20};
  wire [3:0]   maskDestinationResult_lo_lo_21 = {sourceDataVec_1[25:24], sourceDataVec_0[25:24]};
  wire [3:0]   maskDestinationResult_lo_hi_21 = {sourceDataVec_3[25:24], sourceDataVec_2[25:24]};
  wire [7:0]   maskDestinationResult_lo_85 = {maskDestinationResult_lo_hi_21, maskDestinationResult_lo_lo_21};
  wire [3:0]   maskDestinationResult_hi_lo_21 = {sourceDataVec_5[25:24], sourceDataVec_4[25:24]};
  wire [3:0]   maskDestinationResult_hi_hi_21 = {sourceDataVec_7[25:24], sourceDataVec_6[25:24]};
  wire [7:0]   maskDestinationResult_hi_85 = {maskDestinationResult_hi_hi_21, maskDestinationResult_hi_lo_21};
  wire [3:0]   maskDestinationResult_lo_lo_22 = {sourceDataVec_1[27:26], sourceDataVec_0[27:26]};
  wire [3:0]   maskDestinationResult_lo_hi_22 = {sourceDataVec_3[27:26], sourceDataVec_2[27:26]};
  wire [7:0]   maskDestinationResult_lo_86 = {maskDestinationResult_lo_hi_22, maskDestinationResult_lo_lo_22};
  wire [3:0]   maskDestinationResult_hi_lo_22 = {sourceDataVec_5[27:26], sourceDataVec_4[27:26]};
  wire [3:0]   maskDestinationResult_hi_hi_22 = {sourceDataVec_7[27:26], sourceDataVec_6[27:26]};
  wire [7:0]   maskDestinationResult_hi_86 = {maskDestinationResult_hi_hi_22, maskDestinationResult_hi_lo_22};
  wire [3:0]   maskDestinationResult_lo_lo_23 = {sourceDataVec_1[29:28], sourceDataVec_0[29:28]};
  wire [3:0]   maskDestinationResult_lo_hi_23 = {sourceDataVec_3[29:28], sourceDataVec_2[29:28]};
  wire [7:0]   maskDestinationResult_lo_87 = {maskDestinationResult_lo_hi_23, maskDestinationResult_lo_lo_23};
  wire [3:0]   maskDestinationResult_hi_lo_23 = {sourceDataVec_5[29:28], sourceDataVec_4[29:28]};
  wire [3:0]   maskDestinationResult_hi_hi_23 = {sourceDataVec_7[29:28], sourceDataVec_6[29:28]};
  wire [7:0]   maskDestinationResult_hi_87 = {maskDestinationResult_hi_hi_23, maskDestinationResult_hi_lo_23};
  wire [3:0]   maskDestinationResult_lo_lo_24 = {sourceDataVec_1[31:30], sourceDataVec_0[31:30]};
  wire [3:0]   maskDestinationResult_lo_hi_24 = {sourceDataVec_3[31:30], sourceDataVec_2[31:30]};
  wire [7:0]   maskDestinationResult_lo_88 = {maskDestinationResult_lo_hi_24, maskDestinationResult_lo_lo_24};
  wire [3:0]   maskDestinationResult_hi_lo_24 = {sourceDataVec_5[31:30], sourceDataVec_4[31:30]};
  wire [3:0]   maskDestinationResult_hi_hi_24 = {sourceDataVec_7[31:30], sourceDataVec_6[31:30]};
  wire [7:0]   maskDestinationResult_hi_88 = {maskDestinationResult_hi_hi_24, maskDestinationResult_hi_lo_24};
  wire [31:0]  maskDestinationResult_lo_lo_lo = {maskDestinationResult_hi_74, maskDestinationResult_lo_74, maskDestinationResult_hi_73, maskDestinationResult_lo_73};
  wire [31:0]  maskDestinationResult_lo_lo_hi = {maskDestinationResult_hi_76, maskDestinationResult_lo_76, maskDestinationResult_hi_75, maskDestinationResult_lo_75};
  wire [63:0]  maskDestinationResult_lo_lo_25 = {maskDestinationResult_lo_lo_hi, maskDestinationResult_lo_lo_lo};
  wire [31:0]  maskDestinationResult_lo_hi_lo = {maskDestinationResult_hi_78, maskDestinationResult_lo_78, maskDestinationResult_hi_77, maskDestinationResult_lo_77};
  wire [31:0]  maskDestinationResult_lo_hi_hi = {maskDestinationResult_hi_80, maskDestinationResult_lo_80, maskDestinationResult_hi_79, maskDestinationResult_lo_79};
  wire [63:0]  maskDestinationResult_lo_hi_25 = {maskDestinationResult_lo_hi_hi, maskDestinationResult_lo_hi_lo};
  wire [127:0] maskDestinationResult_lo_89 = {maskDestinationResult_lo_hi_25, maskDestinationResult_lo_lo_25};
  wire [31:0]  maskDestinationResult_hi_lo_lo = {maskDestinationResult_hi_82, maskDestinationResult_lo_82, maskDestinationResult_hi_81, maskDestinationResult_lo_81};
  wire [31:0]  maskDestinationResult_hi_lo_hi = {maskDestinationResult_hi_84, maskDestinationResult_lo_84, maskDestinationResult_hi_83, maskDestinationResult_lo_83};
  wire [63:0]  maskDestinationResult_hi_lo_25 = {maskDestinationResult_hi_lo_hi, maskDestinationResult_hi_lo_lo};
  wire [31:0]  maskDestinationResult_hi_hi_lo = {maskDestinationResult_hi_86, maskDestinationResult_lo_86, maskDestinationResult_hi_85, maskDestinationResult_lo_85};
  wire [31:0]  maskDestinationResult_hi_hi_hi = {maskDestinationResult_hi_88, maskDestinationResult_lo_88, maskDestinationResult_hi_87, maskDestinationResult_lo_87};
  wire [63:0]  maskDestinationResult_hi_hi_25 = {maskDestinationResult_hi_hi_hi, maskDestinationResult_hi_hi_lo};
  wire [127:0] maskDestinationResult_hi_89 = {maskDestinationResult_hi_hi_25, maskDestinationResult_hi_lo_25};
  wire [1:0]   maskDestinationResult_lo_lo_26 = {sourceDataVec_1[0], sourceDataVec_0[0]};
  wire [1:0]   maskDestinationResult_lo_hi_26 = {sourceDataVec_3[0], sourceDataVec_2[0]};
  wire [3:0]   maskDestinationResult_lo_90 = {maskDestinationResult_lo_hi_26, maskDestinationResult_lo_lo_26};
  wire [1:0]   maskDestinationResult_hi_lo_26 = {sourceDataVec_5[0], sourceDataVec_4[0]};
  wire [1:0]   maskDestinationResult_hi_hi_26 = {sourceDataVec_7[0], sourceDataVec_6[0]};
  wire [3:0]   maskDestinationResult_hi_90 = {maskDestinationResult_hi_hi_26, maskDestinationResult_hi_lo_26};
  wire [1:0]   maskDestinationResult_lo_lo_27 = {sourceDataVec_1[1], sourceDataVec_0[1]};
  wire [1:0]   maskDestinationResult_lo_hi_27 = {sourceDataVec_3[1], sourceDataVec_2[1]};
  wire [3:0]   maskDestinationResult_lo_91 = {maskDestinationResult_lo_hi_27, maskDestinationResult_lo_lo_27};
  wire [1:0]   maskDestinationResult_hi_lo_27 = {sourceDataVec_5[1], sourceDataVec_4[1]};
  wire [1:0]   maskDestinationResult_hi_hi_27 = {sourceDataVec_7[1], sourceDataVec_6[1]};
  wire [3:0]   maskDestinationResult_hi_91 = {maskDestinationResult_hi_hi_27, maskDestinationResult_hi_lo_27};
  wire [1:0]   maskDestinationResult_lo_lo_28 = {sourceDataVec_1[2], sourceDataVec_0[2]};
  wire [1:0]   maskDestinationResult_lo_hi_28 = {sourceDataVec_3[2], sourceDataVec_2[2]};
  wire [3:0]   maskDestinationResult_lo_92 = {maskDestinationResult_lo_hi_28, maskDestinationResult_lo_lo_28};
  wire [1:0]   maskDestinationResult_hi_lo_28 = {sourceDataVec_5[2], sourceDataVec_4[2]};
  wire [1:0]   maskDestinationResult_hi_hi_28 = {sourceDataVec_7[2], sourceDataVec_6[2]};
  wire [3:0]   maskDestinationResult_hi_92 = {maskDestinationResult_hi_hi_28, maskDestinationResult_hi_lo_28};
  wire [1:0]   maskDestinationResult_lo_lo_29 = {sourceDataVec_1[3], sourceDataVec_0[3]};
  wire [1:0]   maskDestinationResult_lo_hi_29 = {sourceDataVec_3[3], sourceDataVec_2[3]};
  wire [3:0]   maskDestinationResult_lo_93 = {maskDestinationResult_lo_hi_29, maskDestinationResult_lo_lo_29};
  wire [1:0]   maskDestinationResult_hi_lo_29 = {sourceDataVec_5[3], sourceDataVec_4[3]};
  wire [1:0]   maskDestinationResult_hi_hi_29 = {sourceDataVec_7[3], sourceDataVec_6[3]};
  wire [3:0]   maskDestinationResult_hi_93 = {maskDestinationResult_hi_hi_29, maskDestinationResult_hi_lo_29};
  wire [1:0]   maskDestinationResult_lo_lo_30 = {sourceDataVec_1[4], sourceDataVec_0[4]};
  wire [1:0]   maskDestinationResult_lo_hi_30 = {sourceDataVec_3[4], sourceDataVec_2[4]};
  wire [3:0]   maskDestinationResult_lo_94 = {maskDestinationResult_lo_hi_30, maskDestinationResult_lo_lo_30};
  wire [1:0]   maskDestinationResult_hi_lo_30 = {sourceDataVec_5[4], sourceDataVec_4[4]};
  wire [1:0]   maskDestinationResult_hi_hi_30 = {sourceDataVec_7[4], sourceDataVec_6[4]};
  wire [3:0]   maskDestinationResult_hi_94 = {maskDestinationResult_hi_hi_30, maskDestinationResult_hi_lo_30};
  wire [1:0]   maskDestinationResult_lo_lo_31 = {sourceDataVec_1[5], sourceDataVec_0[5]};
  wire [1:0]   maskDestinationResult_lo_hi_31 = {sourceDataVec_3[5], sourceDataVec_2[5]};
  wire [3:0]   maskDestinationResult_lo_95 = {maskDestinationResult_lo_hi_31, maskDestinationResult_lo_lo_31};
  wire [1:0]   maskDestinationResult_hi_lo_31 = {sourceDataVec_5[5], sourceDataVec_4[5]};
  wire [1:0]   maskDestinationResult_hi_hi_31 = {sourceDataVec_7[5], sourceDataVec_6[5]};
  wire [3:0]   maskDestinationResult_hi_95 = {maskDestinationResult_hi_hi_31, maskDestinationResult_hi_lo_31};
  wire [1:0]   maskDestinationResult_lo_lo_32 = {sourceDataVec_1[6], sourceDataVec_0[6]};
  wire [1:0]   maskDestinationResult_lo_hi_32 = {sourceDataVec_3[6], sourceDataVec_2[6]};
  wire [3:0]   maskDestinationResult_lo_96 = {maskDestinationResult_lo_hi_32, maskDestinationResult_lo_lo_32};
  wire [1:0]   maskDestinationResult_hi_lo_32 = {sourceDataVec_5[6], sourceDataVec_4[6]};
  wire [1:0]   maskDestinationResult_hi_hi_32 = {sourceDataVec_7[6], sourceDataVec_6[6]};
  wire [3:0]   maskDestinationResult_hi_96 = {maskDestinationResult_hi_hi_32, maskDestinationResult_hi_lo_32};
  wire [1:0]   maskDestinationResult_lo_lo_33 = {sourceDataVec_1[7], sourceDataVec_0[7]};
  wire [1:0]   maskDestinationResult_lo_hi_33 = {sourceDataVec_3[7], sourceDataVec_2[7]};
  wire [3:0]   maskDestinationResult_lo_97 = {maskDestinationResult_lo_hi_33, maskDestinationResult_lo_lo_33};
  wire [1:0]   maskDestinationResult_hi_lo_33 = {sourceDataVec_5[7], sourceDataVec_4[7]};
  wire [1:0]   maskDestinationResult_hi_hi_33 = {sourceDataVec_7[7], sourceDataVec_6[7]};
  wire [3:0]   maskDestinationResult_hi_97 = {maskDestinationResult_hi_hi_33, maskDestinationResult_hi_lo_33};
  wire [1:0]   maskDestinationResult_lo_lo_34 = {sourceDataVec_1[8], sourceDataVec_0[8]};
  wire [1:0]   maskDestinationResult_lo_hi_34 = {sourceDataVec_3[8], sourceDataVec_2[8]};
  wire [3:0]   maskDestinationResult_lo_98 = {maskDestinationResult_lo_hi_34, maskDestinationResult_lo_lo_34};
  wire [1:0]   maskDestinationResult_hi_lo_34 = {sourceDataVec_5[8], sourceDataVec_4[8]};
  wire [1:0]   maskDestinationResult_hi_hi_34 = {sourceDataVec_7[8], sourceDataVec_6[8]};
  wire [3:0]   maskDestinationResult_hi_98 = {maskDestinationResult_hi_hi_34, maskDestinationResult_hi_lo_34};
  wire [1:0]   maskDestinationResult_lo_lo_35 = {sourceDataVec_1[9], sourceDataVec_0[9]};
  wire [1:0]   maskDestinationResult_lo_hi_35 = {sourceDataVec_3[9], sourceDataVec_2[9]};
  wire [3:0]   maskDestinationResult_lo_99 = {maskDestinationResult_lo_hi_35, maskDestinationResult_lo_lo_35};
  wire [1:0]   maskDestinationResult_hi_lo_35 = {sourceDataVec_5[9], sourceDataVec_4[9]};
  wire [1:0]   maskDestinationResult_hi_hi_35 = {sourceDataVec_7[9], sourceDataVec_6[9]};
  wire [3:0]   maskDestinationResult_hi_99 = {maskDestinationResult_hi_hi_35, maskDestinationResult_hi_lo_35};
  wire [1:0]   maskDestinationResult_lo_lo_36 = {sourceDataVec_1[10], sourceDataVec_0[10]};
  wire [1:0]   maskDestinationResult_lo_hi_36 = {sourceDataVec_3[10], sourceDataVec_2[10]};
  wire [3:0]   maskDestinationResult_lo_100 = {maskDestinationResult_lo_hi_36, maskDestinationResult_lo_lo_36};
  wire [1:0]   maskDestinationResult_hi_lo_36 = {sourceDataVec_5[10], sourceDataVec_4[10]};
  wire [1:0]   maskDestinationResult_hi_hi_36 = {sourceDataVec_7[10], sourceDataVec_6[10]};
  wire [3:0]   maskDestinationResult_hi_100 = {maskDestinationResult_hi_hi_36, maskDestinationResult_hi_lo_36};
  wire [1:0]   maskDestinationResult_lo_lo_37 = {sourceDataVec_1[11], sourceDataVec_0[11]};
  wire [1:0]   maskDestinationResult_lo_hi_37 = {sourceDataVec_3[11], sourceDataVec_2[11]};
  wire [3:0]   maskDestinationResult_lo_101 = {maskDestinationResult_lo_hi_37, maskDestinationResult_lo_lo_37};
  wire [1:0]   maskDestinationResult_hi_lo_37 = {sourceDataVec_5[11], sourceDataVec_4[11]};
  wire [1:0]   maskDestinationResult_hi_hi_37 = {sourceDataVec_7[11], sourceDataVec_6[11]};
  wire [3:0]   maskDestinationResult_hi_101 = {maskDestinationResult_hi_hi_37, maskDestinationResult_hi_lo_37};
  wire [1:0]   maskDestinationResult_lo_lo_38 = {sourceDataVec_1[12], sourceDataVec_0[12]};
  wire [1:0]   maskDestinationResult_lo_hi_38 = {sourceDataVec_3[12], sourceDataVec_2[12]};
  wire [3:0]   maskDestinationResult_lo_102 = {maskDestinationResult_lo_hi_38, maskDestinationResult_lo_lo_38};
  wire [1:0]   maskDestinationResult_hi_lo_38 = {sourceDataVec_5[12], sourceDataVec_4[12]};
  wire [1:0]   maskDestinationResult_hi_hi_38 = {sourceDataVec_7[12], sourceDataVec_6[12]};
  wire [3:0]   maskDestinationResult_hi_102 = {maskDestinationResult_hi_hi_38, maskDestinationResult_hi_lo_38};
  wire [1:0]   maskDestinationResult_lo_lo_39 = {sourceDataVec_1[13], sourceDataVec_0[13]};
  wire [1:0]   maskDestinationResult_lo_hi_39 = {sourceDataVec_3[13], sourceDataVec_2[13]};
  wire [3:0]   maskDestinationResult_lo_103 = {maskDestinationResult_lo_hi_39, maskDestinationResult_lo_lo_39};
  wire [1:0]   maskDestinationResult_hi_lo_39 = {sourceDataVec_5[13], sourceDataVec_4[13]};
  wire [1:0]   maskDestinationResult_hi_hi_39 = {sourceDataVec_7[13], sourceDataVec_6[13]};
  wire [3:0]   maskDestinationResult_hi_103 = {maskDestinationResult_hi_hi_39, maskDestinationResult_hi_lo_39};
  wire [1:0]   maskDestinationResult_lo_lo_40 = {sourceDataVec_1[14], sourceDataVec_0[14]};
  wire [1:0]   maskDestinationResult_lo_hi_40 = {sourceDataVec_3[14], sourceDataVec_2[14]};
  wire [3:0]   maskDestinationResult_lo_104 = {maskDestinationResult_lo_hi_40, maskDestinationResult_lo_lo_40};
  wire [1:0]   maskDestinationResult_hi_lo_40 = {sourceDataVec_5[14], sourceDataVec_4[14]};
  wire [1:0]   maskDestinationResult_hi_hi_40 = {sourceDataVec_7[14], sourceDataVec_6[14]};
  wire [3:0]   maskDestinationResult_hi_104 = {maskDestinationResult_hi_hi_40, maskDestinationResult_hi_lo_40};
  wire [1:0]   maskDestinationResult_lo_lo_41 = {sourceDataVec_1[15], sourceDataVec_0[15]};
  wire [1:0]   maskDestinationResult_lo_hi_41 = {sourceDataVec_3[15], sourceDataVec_2[15]};
  wire [3:0]   maskDestinationResult_lo_105 = {maskDestinationResult_lo_hi_41, maskDestinationResult_lo_lo_41};
  wire [1:0]   maskDestinationResult_hi_lo_41 = {sourceDataVec_5[15], sourceDataVec_4[15]};
  wire [1:0]   maskDestinationResult_hi_hi_41 = {sourceDataVec_7[15], sourceDataVec_6[15]};
  wire [3:0]   maskDestinationResult_hi_105 = {maskDestinationResult_hi_hi_41, maskDestinationResult_hi_lo_41};
  wire [1:0]   maskDestinationResult_lo_lo_42 = {sourceDataVec_1[16], sourceDataVec_0[16]};
  wire [1:0]   maskDestinationResult_lo_hi_42 = {sourceDataVec_3[16], sourceDataVec_2[16]};
  wire [3:0]   maskDestinationResult_lo_106 = {maskDestinationResult_lo_hi_42, maskDestinationResult_lo_lo_42};
  wire [1:0]   maskDestinationResult_hi_lo_42 = {sourceDataVec_5[16], sourceDataVec_4[16]};
  wire [1:0]   maskDestinationResult_hi_hi_42 = {sourceDataVec_7[16], sourceDataVec_6[16]};
  wire [3:0]   maskDestinationResult_hi_106 = {maskDestinationResult_hi_hi_42, maskDestinationResult_hi_lo_42};
  wire [1:0]   maskDestinationResult_lo_lo_43 = {sourceDataVec_1[17], sourceDataVec_0[17]};
  wire [1:0]   maskDestinationResult_lo_hi_43 = {sourceDataVec_3[17], sourceDataVec_2[17]};
  wire [3:0]   maskDestinationResult_lo_107 = {maskDestinationResult_lo_hi_43, maskDestinationResult_lo_lo_43};
  wire [1:0]   maskDestinationResult_hi_lo_43 = {sourceDataVec_5[17], sourceDataVec_4[17]};
  wire [1:0]   maskDestinationResult_hi_hi_43 = {sourceDataVec_7[17], sourceDataVec_6[17]};
  wire [3:0]   maskDestinationResult_hi_107 = {maskDestinationResult_hi_hi_43, maskDestinationResult_hi_lo_43};
  wire [1:0]   maskDestinationResult_lo_lo_44 = {sourceDataVec_1[18], sourceDataVec_0[18]};
  wire [1:0]   maskDestinationResult_lo_hi_44 = {sourceDataVec_3[18], sourceDataVec_2[18]};
  wire [3:0]   maskDestinationResult_lo_108 = {maskDestinationResult_lo_hi_44, maskDestinationResult_lo_lo_44};
  wire [1:0]   maskDestinationResult_hi_lo_44 = {sourceDataVec_5[18], sourceDataVec_4[18]};
  wire [1:0]   maskDestinationResult_hi_hi_44 = {sourceDataVec_7[18], sourceDataVec_6[18]};
  wire [3:0]   maskDestinationResult_hi_108 = {maskDestinationResult_hi_hi_44, maskDestinationResult_hi_lo_44};
  wire [1:0]   maskDestinationResult_lo_lo_45 = {sourceDataVec_1[19], sourceDataVec_0[19]};
  wire [1:0]   maskDestinationResult_lo_hi_45 = {sourceDataVec_3[19], sourceDataVec_2[19]};
  wire [3:0]   maskDestinationResult_lo_109 = {maskDestinationResult_lo_hi_45, maskDestinationResult_lo_lo_45};
  wire [1:0]   maskDestinationResult_hi_lo_45 = {sourceDataVec_5[19], sourceDataVec_4[19]};
  wire [1:0]   maskDestinationResult_hi_hi_45 = {sourceDataVec_7[19], sourceDataVec_6[19]};
  wire [3:0]   maskDestinationResult_hi_109 = {maskDestinationResult_hi_hi_45, maskDestinationResult_hi_lo_45};
  wire [1:0]   maskDestinationResult_lo_lo_46 = {sourceDataVec_1[20], sourceDataVec_0[20]};
  wire [1:0]   maskDestinationResult_lo_hi_46 = {sourceDataVec_3[20], sourceDataVec_2[20]};
  wire [3:0]   maskDestinationResult_lo_110 = {maskDestinationResult_lo_hi_46, maskDestinationResult_lo_lo_46};
  wire [1:0]   maskDestinationResult_hi_lo_46 = {sourceDataVec_5[20], sourceDataVec_4[20]};
  wire [1:0]   maskDestinationResult_hi_hi_46 = {sourceDataVec_7[20], sourceDataVec_6[20]};
  wire [3:0]   maskDestinationResult_hi_110 = {maskDestinationResult_hi_hi_46, maskDestinationResult_hi_lo_46};
  wire [1:0]   maskDestinationResult_lo_lo_47 = {sourceDataVec_1[21], sourceDataVec_0[21]};
  wire [1:0]   maskDestinationResult_lo_hi_47 = {sourceDataVec_3[21], sourceDataVec_2[21]};
  wire [3:0]   maskDestinationResult_lo_111 = {maskDestinationResult_lo_hi_47, maskDestinationResult_lo_lo_47};
  wire [1:0]   maskDestinationResult_hi_lo_47 = {sourceDataVec_5[21], sourceDataVec_4[21]};
  wire [1:0]   maskDestinationResult_hi_hi_47 = {sourceDataVec_7[21], sourceDataVec_6[21]};
  wire [3:0]   maskDestinationResult_hi_111 = {maskDestinationResult_hi_hi_47, maskDestinationResult_hi_lo_47};
  wire [1:0]   maskDestinationResult_lo_lo_48 = {sourceDataVec_1[22], sourceDataVec_0[22]};
  wire [1:0]   maskDestinationResult_lo_hi_48 = {sourceDataVec_3[22], sourceDataVec_2[22]};
  wire [3:0]   maskDestinationResult_lo_112 = {maskDestinationResult_lo_hi_48, maskDestinationResult_lo_lo_48};
  wire [1:0]   maskDestinationResult_hi_lo_48 = {sourceDataVec_5[22], sourceDataVec_4[22]};
  wire [1:0]   maskDestinationResult_hi_hi_48 = {sourceDataVec_7[22], sourceDataVec_6[22]};
  wire [3:0]   maskDestinationResult_hi_112 = {maskDestinationResult_hi_hi_48, maskDestinationResult_hi_lo_48};
  wire [1:0]   maskDestinationResult_lo_lo_49 = {sourceDataVec_1[23], sourceDataVec_0[23]};
  wire [1:0]   maskDestinationResult_lo_hi_49 = {sourceDataVec_3[23], sourceDataVec_2[23]};
  wire [3:0]   maskDestinationResult_lo_113 = {maskDestinationResult_lo_hi_49, maskDestinationResult_lo_lo_49};
  wire [1:0]   maskDestinationResult_hi_lo_49 = {sourceDataVec_5[23], sourceDataVec_4[23]};
  wire [1:0]   maskDestinationResult_hi_hi_49 = {sourceDataVec_7[23], sourceDataVec_6[23]};
  wire [3:0]   maskDestinationResult_hi_113 = {maskDestinationResult_hi_hi_49, maskDestinationResult_hi_lo_49};
  wire [1:0]   maskDestinationResult_lo_lo_50 = {sourceDataVec_1[24], sourceDataVec_0[24]};
  wire [1:0]   maskDestinationResult_lo_hi_50 = {sourceDataVec_3[24], sourceDataVec_2[24]};
  wire [3:0]   maskDestinationResult_lo_114 = {maskDestinationResult_lo_hi_50, maskDestinationResult_lo_lo_50};
  wire [1:0]   maskDestinationResult_hi_lo_50 = {sourceDataVec_5[24], sourceDataVec_4[24]};
  wire [1:0]   maskDestinationResult_hi_hi_50 = {sourceDataVec_7[24], sourceDataVec_6[24]};
  wire [3:0]   maskDestinationResult_hi_114 = {maskDestinationResult_hi_hi_50, maskDestinationResult_hi_lo_50};
  wire [1:0]   maskDestinationResult_lo_lo_51 = {sourceDataVec_1[25], sourceDataVec_0[25]};
  wire [1:0]   maskDestinationResult_lo_hi_51 = {sourceDataVec_3[25], sourceDataVec_2[25]};
  wire [3:0]   maskDestinationResult_lo_115 = {maskDestinationResult_lo_hi_51, maskDestinationResult_lo_lo_51};
  wire [1:0]   maskDestinationResult_hi_lo_51 = {sourceDataVec_5[25], sourceDataVec_4[25]};
  wire [1:0]   maskDestinationResult_hi_hi_51 = {sourceDataVec_7[25], sourceDataVec_6[25]};
  wire [3:0]   maskDestinationResult_hi_115 = {maskDestinationResult_hi_hi_51, maskDestinationResult_hi_lo_51};
  wire [1:0]   maskDestinationResult_lo_lo_52 = {sourceDataVec_1[26], sourceDataVec_0[26]};
  wire [1:0]   maskDestinationResult_lo_hi_52 = {sourceDataVec_3[26], sourceDataVec_2[26]};
  wire [3:0]   maskDestinationResult_lo_116 = {maskDestinationResult_lo_hi_52, maskDestinationResult_lo_lo_52};
  wire [1:0]   maskDestinationResult_hi_lo_52 = {sourceDataVec_5[26], sourceDataVec_4[26]};
  wire [1:0]   maskDestinationResult_hi_hi_52 = {sourceDataVec_7[26], sourceDataVec_6[26]};
  wire [3:0]   maskDestinationResult_hi_116 = {maskDestinationResult_hi_hi_52, maskDestinationResult_hi_lo_52};
  wire [1:0]   maskDestinationResult_lo_lo_53 = {sourceDataVec_1[27], sourceDataVec_0[27]};
  wire [1:0]   maskDestinationResult_lo_hi_53 = {sourceDataVec_3[27], sourceDataVec_2[27]};
  wire [3:0]   maskDestinationResult_lo_117 = {maskDestinationResult_lo_hi_53, maskDestinationResult_lo_lo_53};
  wire [1:0]   maskDestinationResult_hi_lo_53 = {sourceDataVec_5[27], sourceDataVec_4[27]};
  wire [1:0]   maskDestinationResult_hi_hi_53 = {sourceDataVec_7[27], sourceDataVec_6[27]};
  wire [3:0]   maskDestinationResult_hi_117 = {maskDestinationResult_hi_hi_53, maskDestinationResult_hi_lo_53};
  wire [1:0]   maskDestinationResult_lo_lo_54 = {sourceDataVec_1[28], sourceDataVec_0[28]};
  wire [1:0]   maskDestinationResult_lo_hi_54 = {sourceDataVec_3[28], sourceDataVec_2[28]};
  wire [3:0]   maskDestinationResult_lo_118 = {maskDestinationResult_lo_hi_54, maskDestinationResult_lo_lo_54};
  wire [1:0]   maskDestinationResult_hi_lo_54 = {sourceDataVec_5[28], sourceDataVec_4[28]};
  wire [1:0]   maskDestinationResult_hi_hi_54 = {sourceDataVec_7[28], sourceDataVec_6[28]};
  wire [3:0]   maskDestinationResult_hi_118 = {maskDestinationResult_hi_hi_54, maskDestinationResult_hi_lo_54};
  wire [1:0]   maskDestinationResult_lo_lo_55 = {sourceDataVec_1[29], sourceDataVec_0[29]};
  wire [1:0]   maskDestinationResult_lo_hi_55 = {sourceDataVec_3[29], sourceDataVec_2[29]};
  wire [3:0]   maskDestinationResult_lo_119 = {maskDestinationResult_lo_hi_55, maskDestinationResult_lo_lo_55};
  wire [1:0]   maskDestinationResult_hi_lo_55 = {sourceDataVec_5[29], sourceDataVec_4[29]};
  wire [1:0]   maskDestinationResult_hi_hi_55 = {sourceDataVec_7[29], sourceDataVec_6[29]};
  wire [3:0]   maskDestinationResult_hi_119 = {maskDestinationResult_hi_hi_55, maskDestinationResult_hi_lo_55};
  wire [1:0]   maskDestinationResult_lo_lo_56 = {sourceDataVec_1[30], sourceDataVec_0[30]};
  wire [1:0]   maskDestinationResult_lo_hi_56 = {sourceDataVec_3[30], sourceDataVec_2[30]};
  wire [3:0]   maskDestinationResult_lo_120 = {maskDestinationResult_lo_hi_56, maskDestinationResult_lo_lo_56};
  wire [1:0]   maskDestinationResult_hi_lo_56 = {sourceDataVec_5[30], sourceDataVec_4[30]};
  wire [1:0]   maskDestinationResult_hi_hi_56 = {sourceDataVec_7[30], sourceDataVec_6[30]};
  wire [3:0]   maskDestinationResult_hi_120 = {maskDestinationResult_hi_hi_56, maskDestinationResult_hi_lo_56};
  wire [1:0]   maskDestinationResult_lo_lo_57 = {sourceDataVec_1[31], sourceDataVec_0[31]};
  wire [1:0]   maskDestinationResult_lo_hi_57 = {sourceDataVec_3[31], sourceDataVec_2[31]};
  wire [3:0]   maskDestinationResult_lo_121 = {maskDestinationResult_lo_hi_57, maskDestinationResult_lo_lo_57};
  wire [1:0]   maskDestinationResult_hi_lo_57 = {sourceDataVec_5[31], sourceDataVec_4[31]};
  wire [1:0]   maskDestinationResult_hi_hi_57 = {sourceDataVec_7[31], sourceDataVec_6[31]};
  wire [3:0]   maskDestinationResult_hi_121 = {maskDestinationResult_hi_hi_57, maskDestinationResult_hi_lo_57};
  wire [15:0]  maskDestinationResult_lo_lo_lo_lo = {maskDestinationResult_hi_91, maskDestinationResult_lo_91, maskDestinationResult_hi_90, maskDestinationResult_lo_90};
  wire [15:0]  maskDestinationResult_lo_lo_lo_hi = {maskDestinationResult_hi_93, maskDestinationResult_lo_93, maskDestinationResult_hi_92, maskDestinationResult_lo_92};
  wire [31:0]  maskDestinationResult_lo_lo_lo_1 = {maskDestinationResult_lo_lo_lo_hi, maskDestinationResult_lo_lo_lo_lo};
  wire [15:0]  maskDestinationResult_lo_lo_hi_lo = {maskDestinationResult_hi_95, maskDestinationResult_lo_95, maskDestinationResult_hi_94, maskDestinationResult_lo_94};
  wire [15:0]  maskDestinationResult_lo_lo_hi_hi = {maskDestinationResult_hi_97, maskDestinationResult_lo_97, maskDestinationResult_hi_96, maskDestinationResult_lo_96};
  wire [31:0]  maskDestinationResult_lo_lo_hi_1 = {maskDestinationResult_lo_lo_hi_hi, maskDestinationResult_lo_lo_hi_lo};
  wire [63:0]  maskDestinationResult_lo_lo_58 = {maskDestinationResult_lo_lo_hi_1, maskDestinationResult_lo_lo_lo_1};
  wire [15:0]  maskDestinationResult_lo_hi_lo_lo = {maskDestinationResult_hi_99, maskDestinationResult_lo_99, maskDestinationResult_hi_98, maskDestinationResult_lo_98};
  wire [15:0]  maskDestinationResult_lo_hi_lo_hi = {maskDestinationResult_hi_101, maskDestinationResult_lo_101, maskDestinationResult_hi_100, maskDestinationResult_lo_100};
  wire [31:0]  maskDestinationResult_lo_hi_lo_1 = {maskDestinationResult_lo_hi_lo_hi, maskDestinationResult_lo_hi_lo_lo};
  wire [15:0]  maskDestinationResult_lo_hi_hi_lo = {maskDestinationResult_hi_103, maskDestinationResult_lo_103, maskDestinationResult_hi_102, maskDestinationResult_lo_102};
  wire [15:0]  maskDestinationResult_lo_hi_hi_hi = {maskDestinationResult_hi_105, maskDestinationResult_lo_105, maskDestinationResult_hi_104, maskDestinationResult_lo_104};
  wire [31:0]  maskDestinationResult_lo_hi_hi_1 = {maskDestinationResult_lo_hi_hi_hi, maskDestinationResult_lo_hi_hi_lo};
  wire [63:0]  maskDestinationResult_lo_hi_58 = {maskDestinationResult_lo_hi_hi_1, maskDestinationResult_lo_hi_lo_1};
  wire [127:0] maskDestinationResult_lo_122 = {maskDestinationResult_lo_hi_58, maskDestinationResult_lo_lo_58};
  wire [15:0]  maskDestinationResult_hi_lo_lo_lo = {maskDestinationResult_hi_107, maskDestinationResult_lo_107, maskDestinationResult_hi_106, maskDestinationResult_lo_106};
  wire [15:0]  maskDestinationResult_hi_lo_lo_hi = {maskDestinationResult_hi_109, maskDestinationResult_lo_109, maskDestinationResult_hi_108, maskDestinationResult_lo_108};
  wire [31:0]  maskDestinationResult_hi_lo_lo_1 = {maskDestinationResult_hi_lo_lo_hi, maskDestinationResult_hi_lo_lo_lo};
  wire [15:0]  maskDestinationResult_hi_lo_hi_lo = {maskDestinationResult_hi_111, maskDestinationResult_lo_111, maskDestinationResult_hi_110, maskDestinationResult_lo_110};
  wire [15:0]  maskDestinationResult_hi_lo_hi_hi = {maskDestinationResult_hi_113, maskDestinationResult_lo_113, maskDestinationResult_hi_112, maskDestinationResult_lo_112};
  wire [31:0]  maskDestinationResult_hi_lo_hi_1 = {maskDestinationResult_hi_lo_hi_hi, maskDestinationResult_hi_lo_hi_lo};
  wire [63:0]  maskDestinationResult_hi_lo_58 = {maskDestinationResult_hi_lo_hi_1, maskDestinationResult_hi_lo_lo_1};
  wire [15:0]  maskDestinationResult_hi_hi_lo_lo = {maskDestinationResult_hi_115, maskDestinationResult_lo_115, maskDestinationResult_hi_114, maskDestinationResult_lo_114};
  wire [15:0]  maskDestinationResult_hi_hi_lo_hi = {maskDestinationResult_hi_117, maskDestinationResult_lo_117, maskDestinationResult_hi_116, maskDestinationResult_lo_116};
  wire [31:0]  maskDestinationResult_hi_hi_lo_1 = {maskDestinationResult_hi_hi_lo_hi, maskDestinationResult_hi_hi_lo_lo};
  wire [15:0]  maskDestinationResult_hi_hi_hi_lo = {maskDestinationResult_hi_119, maskDestinationResult_lo_119, maskDestinationResult_hi_118, maskDestinationResult_lo_118};
  wire [15:0]  maskDestinationResult_hi_hi_hi_hi = {maskDestinationResult_hi_121, maskDestinationResult_lo_121, maskDestinationResult_hi_120, maskDestinationResult_lo_120};
  wire [31:0]  maskDestinationResult_hi_hi_hi_1 = {maskDestinationResult_hi_hi_hi_hi, maskDestinationResult_hi_hi_hi_lo};
  wire [63:0]  maskDestinationResult_hi_hi_58 = {maskDestinationResult_hi_hi_hi_1, maskDestinationResult_hi_hi_lo_1};
  wire [127:0] maskDestinationResult_hi_122 = {maskDestinationResult_hi_hi_58, maskDestinationResult_hi_lo_58};
  wire [255:0] maskDestinationResult =
    (eew1H[0] ? {maskDestinationResult_hi_72, maskDestinationResult_lo_72} : 256'h0) | (eew1H[1] ? {maskDestinationResult_hi_89, maskDestinationResult_lo_89} : 256'h0)
    | (eew1H[2] ? {maskDestinationResult_hi_122, maskDestinationResult_lo_122} : 256'h0);
  wire         sign = in_uop[0];
  wire         extendRatio = in_uop[2];
  wire [3:0]   _source2_T_1 = 4'h1 << in_groupCounter[1:0];
  wire [1:0]   _source2_T_18 = 2'h1 << in_groupCounter[0];
  wire [127:0] source2 =
    extendRatio
      ? {64'h0, (_source2_T_1[0] ? in_source2[63:0] : 64'h0) | (_source2_T_1[1] ? in_source2[127:64] : 64'h0) | (_source2_T_1[2] ? in_source2[191:128] : 64'h0) | (_source2_T_1[3] ? in_source2[255:192] : 64'h0)}
      : (_source2_T_18[0] ? in_source2[127:0] : 128'h0) | (_source2_T_18[1] ? in_source2[255:128] : 128'h0);
  wire [1:0]   _extendResult_T_249 = 2'h1 << extendRatio;
  wire [31:0]  extendResult_lo_lo_lo = {{8{source2[15] & sign}}, source2[15:8], {8{source2[7] & sign}}, source2[7:0]};
  wire [31:0]  extendResult_lo_lo_hi = {{8{source2[31] & sign}}, source2[31:24], {8{source2[23] & sign}}, source2[23:16]};
  wire [63:0]  extendResult_lo_lo = {extendResult_lo_lo_hi, extendResult_lo_lo_lo};
  wire [31:0]  extendResult_lo_hi_lo = {{8{source2[47] & sign}}, source2[47:40], {8{source2[39] & sign}}, source2[39:32]};
  wire [31:0]  extendResult_lo_hi_hi = {{8{source2[63] & sign}}, source2[63:56], {8{source2[55] & sign}}, source2[55:48]};
  wire [63:0]  extendResult_lo_hi = {extendResult_lo_hi_hi, extendResult_lo_hi_lo};
  wire [127:0] extendResult_lo = {extendResult_lo_hi, extendResult_lo_lo};
  wire [31:0]  extendResult_hi_lo_lo = {{8{source2[79] & sign}}, source2[79:72], {8{source2[71] & sign}}, source2[71:64]};
  wire [31:0]  extendResult_hi_lo_hi = {{8{source2[95] & sign}}, source2[95:88], {8{source2[87] & sign}}, source2[87:80]};
  wire [63:0]  extendResult_hi_lo = {extendResult_hi_lo_hi, extendResult_hi_lo_lo};
  wire [31:0]  extendResult_hi_hi_lo = {{8{source2[111] & sign}}, source2[111:104], {8{source2[103] & sign}}, source2[103:96]};
  wire [31:0]  extendResult_hi_hi_hi = {{8{source2[127] & sign}}, source2[127:120], {8{source2[119] & sign}}, source2[119:112]};
  wire [63:0]  extendResult_hi_hi = {extendResult_hi_hi_hi, extendResult_hi_hi_lo};
  wire [127:0] extendResult_hi = {extendResult_hi_hi, extendResult_hi_lo};
  wire [31:0]  extendResult_lo_lo_lo_lo = {{12{source2[7] & sign}}, source2[7:4], {12{source2[3] & sign}}, source2[3:0]};
  wire [31:0]  extendResult_lo_lo_lo_hi = {{12{source2[15] & sign}}, source2[15:12], {12{source2[11] & sign}}, source2[11:8]};
  wire [63:0]  extendResult_lo_lo_lo_1 = {extendResult_lo_lo_lo_hi, extendResult_lo_lo_lo_lo};
  wire [31:0]  extendResult_lo_lo_hi_lo = {{12{source2[23] & sign}}, source2[23:20], {12{source2[19] & sign}}, source2[19:16]};
  wire [31:0]  extendResult_lo_lo_hi_hi = {{12{source2[31] & sign}}, source2[31:28], {12{source2[27] & sign}}, source2[27:24]};
  wire [63:0]  extendResult_lo_lo_hi_1 = {extendResult_lo_lo_hi_hi, extendResult_lo_lo_hi_lo};
  wire [127:0] extendResult_lo_lo_1 = {extendResult_lo_lo_hi_1, extendResult_lo_lo_lo_1};
  wire [31:0]  extendResult_lo_hi_lo_lo = {{12{source2[39] & sign}}, source2[39:36], {12{source2[35] & sign}}, source2[35:32]};
  wire [31:0]  extendResult_lo_hi_lo_hi = {{12{source2[47] & sign}}, source2[47:44], {12{source2[43] & sign}}, source2[43:40]};
  wire [63:0]  extendResult_lo_hi_lo_1 = {extendResult_lo_hi_lo_hi, extendResult_lo_hi_lo_lo};
  wire [31:0]  extendResult_lo_hi_hi_lo = {{12{source2[55] & sign}}, source2[55:52], {12{source2[51] & sign}}, source2[51:48]};
  wire [31:0]  extendResult_lo_hi_hi_hi = {{12{source2[63] & sign}}, source2[63:60], {12{source2[59] & sign}}, source2[59:56]};
  wire [63:0]  extendResult_lo_hi_hi_1 = {extendResult_lo_hi_hi_hi, extendResult_lo_hi_hi_lo};
  wire [127:0] extendResult_lo_hi_1 = {extendResult_lo_hi_hi_1, extendResult_lo_hi_lo_1};
  wire [255:0] extendResult_lo_1 = {extendResult_lo_hi_1, extendResult_lo_lo_1};
  wire [31:0]  extendResult_hi_lo_lo_lo = {{12{source2[71] & sign}}, source2[71:68], {12{source2[67] & sign}}, source2[67:64]};
  wire [31:0]  extendResult_hi_lo_lo_hi = {{12{source2[79] & sign}}, source2[79:76], {12{source2[75] & sign}}, source2[75:72]};
  wire [63:0]  extendResult_hi_lo_lo_1 = {extendResult_hi_lo_lo_hi, extendResult_hi_lo_lo_lo};
  wire [31:0]  extendResult_hi_lo_hi_lo = {{12{source2[87] & sign}}, source2[87:84], {12{source2[83] & sign}}, source2[83:80]};
  wire [31:0]  extendResult_hi_lo_hi_hi = {{12{source2[95] & sign}}, source2[95:92], {12{source2[91] & sign}}, source2[91:88]};
  wire [63:0]  extendResult_hi_lo_hi_1 = {extendResult_hi_lo_hi_hi, extendResult_hi_lo_hi_lo};
  wire [127:0] extendResult_hi_lo_1 = {extendResult_hi_lo_hi_1, extendResult_hi_lo_lo_1};
  wire [31:0]  extendResult_hi_hi_lo_lo = {{12{source2[103] & sign}}, source2[103:100], {12{source2[99] & sign}}, source2[99:96]};
  wire [31:0]  extendResult_hi_hi_lo_hi = {{12{source2[111] & sign}}, source2[111:108], {12{source2[107] & sign}}, source2[107:104]};
  wire [63:0]  extendResult_hi_hi_lo_1 = {extendResult_hi_hi_lo_hi, extendResult_hi_hi_lo_lo};
  wire [31:0]  extendResult_hi_hi_hi_lo = {{12{source2[119] & sign}}, source2[119:116], {12{source2[115] & sign}}, source2[115:112]};
  wire [31:0]  extendResult_hi_hi_hi_hi = {{12{source2[127] & sign}}, source2[127:124], {12{source2[123] & sign}}, source2[123:120]};
  wire [63:0]  extendResult_hi_hi_hi_1 = {extendResult_hi_hi_hi_hi, extendResult_hi_hi_hi_lo};
  wire [127:0] extendResult_hi_hi_1 = {extendResult_hi_hi_hi_1, extendResult_hi_hi_lo_1};
  wire [255:0] extendResult_hi_1 = {extendResult_hi_hi_1, extendResult_hi_lo_1};
  wire [63:0]  extendResult_lo_lo_2 = {{16{source2[31] & sign}}, source2[31:16], {16{source2[15] & sign}}, source2[15:0]};
  wire [63:0]  extendResult_lo_hi_2 = {{16{source2[63] & sign}}, source2[63:48], {16{source2[47] & sign}}, source2[47:32]};
  wire [127:0] extendResult_lo_2 = {extendResult_lo_hi_2, extendResult_lo_lo_2};
  wire [63:0]  extendResult_hi_lo_2 = {{16{source2[95] & sign}}, source2[95:80], {16{source2[79] & sign}}, source2[79:64]};
  wire [63:0]  extendResult_hi_hi_2 = {{16{source2[127] & sign}}, source2[127:112], {16{source2[111] & sign}}, source2[111:96]};
  wire [127:0] extendResult_hi_2 = {extendResult_hi_hi_2, extendResult_hi_lo_2};
  wire [63:0]  extendResult_lo_lo_lo_2 = {{24{source2[15] & sign}}, source2[15:8], {24{source2[7] & sign}}, source2[7:0]};
  wire [63:0]  extendResult_lo_lo_hi_2 = {{24{source2[31] & sign}}, source2[31:24], {24{source2[23] & sign}}, source2[23:16]};
  wire [127:0] extendResult_lo_lo_3 = {extendResult_lo_lo_hi_2, extendResult_lo_lo_lo_2};
  wire [63:0]  extendResult_lo_hi_lo_2 = {{24{source2[47] & sign}}, source2[47:40], {24{source2[39] & sign}}, source2[39:32]};
  wire [63:0]  extendResult_lo_hi_hi_2 = {{24{source2[63] & sign}}, source2[63:56], {24{source2[55] & sign}}, source2[55:48]};
  wire [127:0] extendResult_lo_hi_3 = {extendResult_lo_hi_hi_2, extendResult_lo_hi_lo_2};
  wire [255:0] extendResult_lo_3 = {extendResult_lo_hi_3, extendResult_lo_lo_3};
  wire [63:0]  extendResult_hi_lo_lo_2 = {{24{source2[79] & sign}}, source2[79:72], {24{source2[71] & sign}}, source2[71:64]};
  wire [63:0]  extendResult_hi_lo_hi_2 = {{24{source2[95] & sign}}, source2[95:88], {24{source2[87] & sign}}, source2[87:80]};
  wire [127:0] extendResult_hi_lo_3 = {extendResult_hi_lo_hi_2, extendResult_hi_lo_lo_2};
  wire [63:0]  extendResult_hi_hi_lo_2 = {{24{source2[111] & sign}}, source2[111:104], {24{source2[103] & sign}}, source2[103:96]};
  wire [63:0]  extendResult_hi_hi_hi_2 = {{24{source2[127] & sign}}, source2[127:120], {24{source2[119] & sign}}, source2[119:112]};
  wire [127:0] extendResult_hi_hi_3 = {extendResult_hi_hi_hi_2, extendResult_hi_hi_lo_2};
  wire [255:0] extendResult_hi_3 = {extendResult_hi_hi_3, extendResult_hi_lo_3};
  wire [511:0] extendResult =
    (eew1H[1] ? {256'h0, _extendResult_T_249[0] ? {extendResult_hi, extendResult_lo} : 256'h0} | (_extendResult_T_249[1] ? {extendResult_hi_1, extendResult_lo_1} : 512'h0) : 512'h0)
    | (eew1H[2] ? {256'h0, _extendResult_T_249[0] ? {extendResult_hi_2, extendResult_lo_2} : 256'h0} | (_extendResult_T_249[1] ? {extendResult_hi_3, extendResult_lo_3} : 512'h0) : 512'h0);
  assign out = isMaskDestination ? maskDestinationResult : extendResult[255:0];
endmodule

