
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module SlideIndexGen(
  input         clock,
                reset,
                newInstruction,
  input  [4:0]  instructionReq_decodeResult_topUop,
  input  [31:0] instructionReq_readFromScala,
  input  [1:0]  instructionReq_sew,
  input  [2:0]  instructionReq_vlmul,
  input         instructionReq_maskType,
  input  [11:0] instructionReq_vl,
  input         indexDeq_ready,
  output        indexDeq_valid,
  output [31:0] indexDeq_bits_needRead,
                indexDeq_bits_elementValid,
                indexDeq_bits_replaceVs1,
                indexDeq_bits_readOffset,
  output [4:0]  indexDeq_bits_accessLane_0,
                indexDeq_bits_accessLane_1,
                indexDeq_bits_accessLane_2,
                indexDeq_bits_accessLane_3,
                indexDeq_bits_accessLane_4,
                indexDeq_bits_accessLane_5,
                indexDeq_bits_accessLane_6,
                indexDeq_bits_accessLane_7,
                indexDeq_bits_accessLane_8,
                indexDeq_bits_accessLane_9,
                indexDeq_bits_accessLane_10,
                indexDeq_bits_accessLane_11,
                indexDeq_bits_accessLane_12,
                indexDeq_bits_accessLane_13,
                indexDeq_bits_accessLane_14,
                indexDeq_bits_accessLane_15,
                indexDeq_bits_accessLane_16,
                indexDeq_bits_accessLane_17,
                indexDeq_bits_accessLane_18,
                indexDeq_bits_accessLane_19,
                indexDeq_bits_accessLane_20,
                indexDeq_bits_accessLane_21,
                indexDeq_bits_accessLane_22,
                indexDeq_bits_accessLane_23,
                indexDeq_bits_accessLane_24,
                indexDeq_bits_accessLane_25,
                indexDeq_bits_accessLane_26,
                indexDeq_bits_accessLane_27,
                indexDeq_bits_accessLane_28,
                indexDeq_bits_accessLane_29,
                indexDeq_bits_accessLane_30,
                indexDeq_bits_accessLane_31,
  output [2:0]  indexDeq_bits_vsGrowth_0,
                indexDeq_bits_vsGrowth_1,
                indexDeq_bits_vsGrowth_2,
                indexDeq_bits_vsGrowth_3,
                indexDeq_bits_vsGrowth_4,
                indexDeq_bits_vsGrowth_5,
                indexDeq_bits_vsGrowth_6,
                indexDeq_bits_vsGrowth_7,
                indexDeq_bits_vsGrowth_8,
                indexDeq_bits_vsGrowth_9,
                indexDeq_bits_vsGrowth_10,
                indexDeq_bits_vsGrowth_11,
                indexDeq_bits_vsGrowth_12,
                indexDeq_bits_vsGrowth_13,
                indexDeq_bits_vsGrowth_14,
                indexDeq_bits_vsGrowth_15,
                indexDeq_bits_vsGrowth_16,
                indexDeq_bits_vsGrowth_17,
                indexDeq_bits_vsGrowth_18,
                indexDeq_bits_vsGrowth_19,
                indexDeq_bits_vsGrowth_20,
                indexDeq_bits_vsGrowth_21,
                indexDeq_bits_vsGrowth_22,
                indexDeq_bits_vsGrowth_23,
                indexDeq_bits_vsGrowth_24,
                indexDeq_bits_vsGrowth_25,
                indexDeq_bits_vsGrowth_26,
                indexDeq_bits_vsGrowth_27,
                indexDeq_bits_vsGrowth_28,
                indexDeq_bits_vsGrowth_29,
                indexDeq_bits_vsGrowth_30,
                indexDeq_bits_vsGrowth_31,
  output [6:0]  indexDeq_bits_executeGroup,
  output [63:0] indexDeq_bits_readDataOffset,
  output        indexDeq_bits_last,
  output [6:0]  slideGroupOut,
  input  [31:0] slideMaskInput
);

  wire        indexDeq_ready_0 = indexDeq_ready;
  wire [1:0]  indexVec_checkResult_2_0 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_1 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_2 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_3 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_4 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_5 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_6 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_7 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_8 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_9 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_10 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_11 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_12 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_13 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_14 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_15 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_16 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_17 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_18 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_19 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_20 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_21 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_22 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_23 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_24 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_25 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_26 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_27 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_28 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_29 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_30 = 2'h0;
  wire [1:0]  indexVec_checkResult_2_0_31 = 2'h0;
  wire [31:0] indexDeq_bits_groupReadState = 32'h0;
  wire [31:0] replaceWithVs1;
  wire [4:0]  indexVec_0_1;
  wire [4:0]  indexVec_1_1;
  wire [4:0]  indexVec_2_1;
  wire [4:0]  indexVec_3_1;
  wire [4:0]  indexVec_4_1;
  wire [4:0]  indexVec_5_1;
  wire [4:0]  indexVec_6_1;
  wire [4:0]  indexVec_7_1;
  wire [4:0]  indexVec_8_1;
  wire [4:0]  indexVec_9_1;
  wire [4:0]  indexVec_10_1;
  wire [4:0]  indexVec_11_1;
  wire [4:0]  indexVec_12_1;
  wire [4:0]  indexVec_13_1;
  wire [4:0]  indexVec_14_1;
  wire [4:0]  indexVec_15_1;
  wire [4:0]  indexVec_16_1;
  wire [4:0]  indexVec_17_1;
  wire [4:0]  indexVec_18_1;
  wire [4:0]  indexVec_19_1;
  wire [4:0]  indexVec_20_1;
  wire [4:0]  indexVec_21_1;
  wire [4:0]  indexVec_22_1;
  wire [4:0]  indexVec_23_1;
  wire [4:0]  indexVec_24_1;
  wire [4:0]  indexVec_25_1;
  wire [4:0]  indexVec_26_1;
  wire [4:0]  indexVec_27_1;
  wire [4:0]  indexVec_28_1;
  wire [4:0]  indexVec_29_1;
  wire [4:0]  indexVec_30_1;
  wire [4:0]  indexVec_31_1;
  wire [2:0]  indexVec_0_3;
  wire [2:0]  indexVec_1_3;
  wire [2:0]  indexVec_2_3;
  wire [2:0]  indexVec_3_3;
  wire [2:0]  indexVec_4_3;
  wire [2:0]  indexVec_5_3;
  wire [2:0]  indexVec_6_3;
  wire [2:0]  indexVec_7_3;
  wire [2:0]  indexVec_8_3;
  wire [2:0]  indexVec_9_3;
  wire [2:0]  indexVec_10_3;
  wire [2:0]  indexVec_11_3;
  wire [2:0]  indexVec_12_3;
  wire [2:0]  indexVec_13_3;
  wire [2:0]  indexVec_14_3;
  wire [2:0]  indexVec_15_3;
  wire [2:0]  indexVec_16_3;
  wire [2:0]  indexVec_17_3;
  wire [2:0]  indexVec_18_3;
  wire [2:0]  indexVec_19_3;
  wire [2:0]  indexVec_20_3;
  wire [2:0]  indexVec_21_3;
  wire [2:0]  indexVec_22_3;
  wire [2:0]  indexVec_23_3;
  wire [2:0]  indexVec_24_3;
  wire [2:0]  indexVec_25_3;
  wire [2:0]  indexVec_26_3;
  wire [2:0]  indexVec_27_3;
  wire [2:0]  indexVec_28_3;
  wire [2:0]  indexVec_29_3;
  wire [2:0]  indexVec_30_3;
  wire [2:0]  indexVec_31_3;
  reg         InstructionValid;
  wire        isSlide = instructionReq_decodeResult_topUop[4:2] == 3'h0;
  wire        slideUp = instructionReq_decodeResult_topUop[0];
  wire        slide1 = instructionReq_decodeResult_topUop[1];
  reg  [6:0]  slideGroup;
  wire [6:0]  indexDeq_bits_executeGroup_0 = slideGroup;
  wire [4:0]  vlTail = instructionReq_vl[4:0];
  wire [6:0]  lastSlideGroup = instructionReq_vl[11:5] - {6'h0, vlTail == 5'h0};
  wire [31:0] _lastValidVec_T = 32'h1 << vlTail;
  wire [31:0] _lastValidVec_T_3 = _lastValidVec_T | {_lastValidVec_T[30:0], 1'h0};
  wire [31:0] _lastValidVec_T_6 = _lastValidVec_T_3 | {_lastValidVec_T_3[29:0], 2'h0};
  wire [31:0] _lastValidVec_T_9 = _lastValidVec_T_6 | {_lastValidVec_T_6[27:0], 4'h0};
  wire [31:0] _lastValidVec_T_12 = _lastValidVec_T_9 | {_lastValidVec_T_9[23:0], 8'h0};
  wire [31:0] lastValidVec = ~(_lastValidVec_T_12 | {_lastValidVec_T_12[15:0], 16'h0});
  wire        indexDeq_bits_last_0 = slideGroup == lastSlideGroup;
  wire [31:0] groupVlValid = indexDeq_bits_last_0 & (|vlTail) ? lastValidVec : 32'hFFFFFFFF;
  wire [31:0] groupMaskValid = instructionReq_maskType ? slideMaskInput : 32'hFFFFFFFF;
  wire [31:0] validVec = groupVlValid & groupMaskValid;
  wire [31:0] lastElementValid = ({1'h0, groupVlValid[31:1]} ^ groupVlValid) & groupMaskValid;
  assign replaceWithVs1 = (slideGroup == 7'h0 & slide1 & slideUp ? {31'h0, groupMaskValid[0]} : 32'h0) | (indexDeq_bits_last_0 & slide1 & ~slideUp ? lastElementValid : 32'h0);
  wire        indexDeq_valid_0;
  wire [31:0] indexDeq_bits_replaceVs1_0 = replaceWithVs1;
  wire        _lastFire_T_1 = indexDeq_ready_0 & indexDeq_valid_0;
  wire        lastFire = indexDeq_bits_last_0 & _lastFire_T_1;
  wire [31:0] slideValue = slide1 ? 32'h1 : instructionReq_readFromScala;
  wire [31:0] PNSelect = {32{slideUp}} ^ slideValue;
  wire [31:0] baseIndex = {20'h0, slideGroup, 5'h0} + PNSelect + {31'h0, slideUp};
  wire [31:0] indexVec_readIndex = baseIndex;
  wire        lagerThanVL = |(slideValue[31:12]);
  wire [3:0]  _sew1H_T = 4'h1 << instructionReq_sew;
  wire [2:0]  sew1H = _sew1H_T[2:0];
  wire [31:0] indexVec_checkResult_allDataPosition = indexVec_readIndex;
  wire [3:0]  _GEN = 4'h1 << instructionReq_vlmul[1:0];
  wire [3:0]  indexVec_checkResult_intLMULInput;
  assign indexVec_checkResult_intLMULInput = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_1;
  assign indexVec_checkResult_intLMULInput_1 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_2;
  assign indexVec_checkResult_intLMULInput_2 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_3;
  assign indexVec_checkResult_intLMULInput_3 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_4;
  assign indexVec_checkResult_intLMULInput_4 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_5;
  assign indexVec_checkResult_intLMULInput_5 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_6;
  assign indexVec_checkResult_intLMULInput_6 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_7;
  assign indexVec_checkResult_intLMULInput_7 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_8;
  assign indexVec_checkResult_intLMULInput_8 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_9;
  assign indexVec_checkResult_intLMULInput_9 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_10;
  assign indexVec_checkResult_intLMULInput_10 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_11;
  assign indexVec_checkResult_intLMULInput_11 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_12;
  assign indexVec_checkResult_intLMULInput_12 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_13;
  assign indexVec_checkResult_intLMULInput_13 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_14;
  assign indexVec_checkResult_intLMULInput_14 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_15;
  assign indexVec_checkResult_intLMULInput_15 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_16;
  assign indexVec_checkResult_intLMULInput_16 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_17;
  assign indexVec_checkResult_intLMULInput_17 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_18;
  assign indexVec_checkResult_intLMULInput_18 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_19;
  assign indexVec_checkResult_intLMULInput_19 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_20;
  assign indexVec_checkResult_intLMULInput_20 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_21;
  assign indexVec_checkResult_intLMULInput_21 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_22;
  assign indexVec_checkResult_intLMULInput_22 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_23;
  assign indexVec_checkResult_intLMULInput_23 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_24;
  assign indexVec_checkResult_intLMULInput_24 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_25;
  assign indexVec_checkResult_intLMULInput_25 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_26;
  assign indexVec_checkResult_intLMULInput_26 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_27;
  assign indexVec_checkResult_intLMULInput_27 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_28;
  assign indexVec_checkResult_intLMULInput_28 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_29;
  assign indexVec_checkResult_intLMULInput_29 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_30;
  assign indexVec_checkResult_intLMULInput_30 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_31;
  assign indexVec_checkResult_intLMULInput_31 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_32;
  assign indexVec_checkResult_intLMULInput_32 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_33;
  assign indexVec_checkResult_intLMULInput_33 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_34;
  assign indexVec_checkResult_intLMULInput_34 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_35;
  assign indexVec_checkResult_intLMULInput_35 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_36;
  assign indexVec_checkResult_intLMULInput_36 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_37;
  assign indexVec_checkResult_intLMULInput_37 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_38;
  assign indexVec_checkResult_intLMULInput_38 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_39;
  assign indexVec_checkResult_intLMULInput_39 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_40;
  assign indexVec_checkResult_intLMULInput_40 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_41;
  assign indexVec_checkResult_intLMULInput_41 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_42;
  assign indexVec_checkResult_intLMULInput_42 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_43;
  assign indexVec_checkResult_intLMULInput_43 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_44;
  assign indexVec_checkResult_intLMULInput_44 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_45;
  assign indexVec_checkResult_intLMULInput_45 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_46;
  assign indexVec_checkResult_intLMULInput_46 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_47;
  assign indexVec_checkResult_intLMULInput_47 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_48;
  assign indexVec_checkResult_intLMULInput_48 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_49;
  assign indexVec_checkResult_intLMULInput_49 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_50;
  assign indexVec_checkResult_intLMULInput_50 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_51;
  assign indexVec_checkResult_intLMULInput_51 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_52;
  assign indexVec_checkResult_intLMULInput_52 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_53;
  assign indexVec_checkResult_intLMULInput_53 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_54;
  assign indexVec_checkResult_intLMULInput_54 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_55;
  assign indexVec_checkResult_intLMULInput_55 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_56;
  assign indexVec_checkResult_intLMULInput_56 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_57;
  assign indexVec_checkResult_intLMULInput_57 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_58;
  assign indexVec_checkResult_intLMULInput_58 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_59;
  assign indexVec_checkResult_intLMULInput_59 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_60;
  assign indexVec_checkResult_intLMULInput_60 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_61;
  assign indexVec_checkResult_intLMULInput_61 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_62;
  assign indexVec_checkResult_intLMULInput_62 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_63;
  assign indexVec_checkResult_intLMULInput_63 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_64;
  assign indexVec_checkResult_intLMULInput_64 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_65;
  assign indexVec_checkResult_intLMULInput_65 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_66;
  assign indexVec_checkResult_intLMULInput_66 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_67;
  assign indexVec_checkResult_intLMULInput_67 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_68;
  assign indexVec_checkResult_intLMULInput_68 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_69;
  assign indexVec_checkResult_intLMULInput_69 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_70;
  assign indexVec_checkResult_intLMULInput_70 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_71;
  assign indexVec_checkResult_intLMULInput_71 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_72;
  assign indexVec_checkResult_intLMULInput_72 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_73;
  assign indexVec_checkResult_intLMULInput_73 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_74;
  assign indexVec_checkResult_intLMULInput_74 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_75;
  assign indexVec_checkResult_intLMULInput_75 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_76;
  assign indexVec_checkResult_intLMULInput_76 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_77;
  assign indexVec_checkResult_intLMULInput_77 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_78;
  assign indexVec_checkResult_intLMULInput_78 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_79;
  assign indexVec_checkResult_intLMULInput_79 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_80;
  assign indexVec_checkResult_intLMULInput_80 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_81;
  assign indexVec_checkResult_intLMULInput_81 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_82;
  assign indexVec_checkResult_intLMULInput_82 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_83;
  assign indexVec_checkResult_intLMULInput_83 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_84;
  assign indexVec_checkResult_intLMULInput_84 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_85;
  assign indexVec_checkResult_intLMULInput_85 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_86;
  assign indexVec_checkResult_intLMULInput_86 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_87;
  assign indexVec_checkResult_intLMULInput_87 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_88;
  assign indexVec_checkResult_intLMULInput_88 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_89;
  assign indexVec_checkResult_intLMULInput_89 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_90;
  assign indexVec_checkResult_intLMULInput_90 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_91;
  assign indexVec_checkResult_intLMULInput_91 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_92;
  assign indexVec_checkResult_intLMULInput_92 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_93;
  assign indexVec_checkResult_intLMULInput_93 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_94;
  assign indexVec_checkResult_intLMULInput_94 = _GEN;
  wire [3:0]  indexVec_checkResult_intLMULInput_95;
  assign indexVec_checkResult_intLMULInput_95 = _GEN;
  wire [10:0] indexVec_checkResult_dataPosition = indexVec_checkResult_allDataPosition[10:0];
  wire [1:0]  indexVec_checkResult_0_0 = indexVec_checkResult_dataPosition[1:0];
  wire [4:0]  indexVec_checkResult_0_1 = indexVec_checkResult_dataPosition[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup = indexVec_checkResult_dataPosition[10:7];
  wire        indexVec_checkResult_0_2 = indexVec_checkResult_dataGroup[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth = indexVec_checkResult_dataGroup[3:1];
  wire [2:0]  indexVec_checkResult_0_3 = indexVec_checkResult_accessRegGrowth;
  wire [5:0]  indexVec_checkResult_decimalProportion = {indexVec_checkResult_0_2, indexVec_checkResult_0_1};
  wire [2:0]  indexVec_checkResult_decimal = indexVec_checkResult_decimalProportion[5:3];
  wire        indexVec_checkResult_overlap =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal >= indexVec_checkResult_intLMULInput[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth} >= indexVec_checkResult_intLMULInput,
      indexVec_checkResult_allDataPosition[31:11]};
  wire        indexVec_checkResult_unChange = slideUp & (indexVec_readIndex[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5 = validVec[0] & ~indexVec_checkResult_unChange;
  wire        indexVec_checkResult_0_4 = indexVec_checkResult_overlap | ~indexVec_checkResult_0_5 | lagerThanVL | indexVec_checkResult_unChange;
  wire [32:0] indexVec_checkResult_allDataPosition_1 = {indexVec_readIndex, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_1 = indexVec_checkResult_allDataPosition_1[10:0];
  wire [1:0]  indexVec_checkResult_1_0 = {indexVec_checkResult_dataPosition_1[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1 = indexVec_checkResult_dataPosition_1[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_1 = indexVec_checkResult_dataPosition_1[10:7];
  wire        indexVec_checkResult_1_2 = indexVec_checkResult_dataGroup_1[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_1 = indexVec_checkResult_dataGroup_1[3:1];
  wire [2:0]  indexVec_checkResult_1_3 = indexVec_checkResult_accessRegGrowth_1;
  wire [5:0]  indexVec_checkResult_decimalProportion_1 = {indexVec_checkResult_1_2, indexVec_checkResult_1_1};
  wire [2:0]  indexVec_checkResult_decimal_1 = indexVec_checkResult_decimalProportion_1[5:3];
  wire        indexVec_checkResult_overlap_1 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_1 >= indexVec_checkResult_intLMULInput_1[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_1} >= indexVec_checkResult_intLMULInput_1,
      indexVec_checkResult_allDataPosition_1[32:11]};
  wire        indexVec_checkResult_unChange_1 = slideUp & (indexVec_readIndex[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5 = validVec[0] & ~indexVec_checkResult_unChange_1;
  wire        indexVec_checkResult_1_4 = indexVec_checkResult_overlap_1 | ~indexVec_checkResult_1_5 | lagerThanVL | indexVec_checkResult_unChange_1;
  wire [33:0] indexVec_checkResult_allDataPosition_2 = {indexVec_readIndex, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_2 = indexVec_checkResult_allDataPosition_2[10:0];
  wire [4:0]  indexVec_checkResult_2_1 = indexVec_checkResult_dataPosition_2[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_2 = indexVec_checkResult_dataPosition_2[10:7];
  wire        indexVec_checkResult_2_2 = indexVec_checkResult_dataGroup_2[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_2 = indexVec_checkResult_dataGroup_2[3:1];
  wire [2:0]  indexVec_checkResult_2_3 = indexVec_checkResult_accessRegGrowth_2;
  wire [5:0]  indexVec_checkResult_decimalProportion_2 = {indexVec_checkResult_2_2, indexVec_checkResult_2_1};
  wire [2:0]  indexVec_checkResult_decimal_2 = indexVec_checkResult_decimalProportion_2[5:3];
  wire        indexVec_checkResult_overlap_2 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_2 >= indexVec_checkResult_intLMULInput_2[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_2} >= indexVec_checkResult_intLMULInput_2,
      indexVec_checkResult_allDataPosition_2[33:11]};
  wire        indexVec_checkResult_unChange_2 = slideUp & (indexVec_readIndex[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5 = validVec[0] & ~indexVec_checkResult_unChange_2;
  wire        indexVec_checkResult_2_4 = indexVec_checkResult_overlap_2 | ~indexVec_checkResult_2_5 | lagerThanVL | indexVec_checkResult_unChange_2;
  wire [1:0]  indexVec_0_0 = (sew1H[0] ? indexVec_checkResult_0_0 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0 : 2'h0);
  assign indexVec_0_1 = (sew1H[0] ? indexVec_checkResult_0_1 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_0_0 = indexVec_0_1;
  wire        indexVec_0_2 = sew1H[0] & indexVec_checkResult_0_2 | sew1H[1] & indexVec_checkResult_1_2 | sew1H[2] & indexVec_checkResult_2_2;
  assign indexVec_0_3 = (sew1H[0] ? indexVec_checkResult_0_3 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_0_0 = indexVec_0_3;
  wire        indexVec_0_4 = sew1H[0] & indexVec_checkResult_0_4 | sew1H[1] & indexVec_checkResult_1_4 | sew1H[2] & indexVec_checkResult_2_4;
  wire        indexVec_0_5 = sew1H[0] & indexVec_checkResult_0_5 | sew1H[1] & indexVec_checkResult_1_5 | sew1H[2] & indexVec_checkResult_2_5;
  wire [31:0] indexVec_readIndex_1 = baseIndex + 32'h1;
  wire [31:0] indexVec_checkResult_allDataPosition_3 = indexVec_readIndex_1;
  wire [10:0] indexVec_checkResult_dataPosition_3 = indexVec_checkResult_allDataPosition_3[10:0];
  wire [1:0]  indexVec_checkResult_0_0_1 = indexVec_checkResult_dataPosition_3[1:0];
  wire [4:0]  indexVec_checkResult_0_1_1 = indexVec_checkResult_dataPosition_3[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_3 = indexVec_checkResult_dataPosition_3[10:7];
  wire        indexVec_checkResult_0_2_1 = indexVec_checkResult_dataGroup_3[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_3 = indexVec_checkResult_dataGroup_3[3:1];
  wire [2:0]  indexVec_checkResult_0_3_1 = indexVec_checkResult_accessRegGrowth_3;
  wire [5:0]  indexVec_checkResult_decimalProportion_3 = {indexVec_checkResult_0_2_1, indexVec_checkResult_0_1_1};
  wire [2:0]  indexVec_checkResult_decimal_3 = indexVec_checkResult_decimalProportion_3[5:3];
  wire        indexVec_checkResult_overlap_3 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_3 >= indexVec_checkResult_intLMULInput_3[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_3} >= indexVec_checkResult_intLMULInput_3,
      indexVec_checkResult_allDataPosition_3[31:11]};
  wire        indexVec_checkResult_unChange_3 = slideUp & (indexVec_readIndex_1[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_1 = validVec[1] & ~indexVec_checkResult_unChange_3;
  wire        indexVec_checkResult_0_4_1 = indexVec_checkResult_overlap_3 | ~indexVec_checkResult_0_5_1 | lagerThanVL | indexVec_checkResult_unChange_3;
  wire [32:0] indexVec_checkResult_allDataPosition_4 = {indexVec_readIndex_1, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_4 = indexVec_checkResult_allDataPosition_4[10:0];
  wire [1:0]  indexVec_checkResult_1_0_1 = {indexVec_checkResult_dataPosition_4[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_1 = indexVec_checkResult_dataPosition_4[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_4 = indexVec_checkResult_dataPosition_4[10:7];
  wire        indexVec_checkResult_1_2_1 = indexVec_checkResult_dataGroup_4[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_4 = indexVec_checkResult_dataGroup_4[3:1];
  wire [2:0]  indexVec_checkResult_1_3_1 = indexVec_checkResult_accessRegGrowth_4;
  wire [5:0]  indexVec_checkResult_decimalProportion_4 = {indexVec_checkResult_1_2_1, indexVec_checkResult_1_1_1};
  wire [2:0]  indexVec_checkResult_decimal_4 = indexVec_checkResult_decimalProportion_4[5:3];
  wire        indexVec_checkResult_overlap_4 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_4 >= indexVec_checkResult_intLMULInput_4[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_4} >= indexVec_checkResult_intLMULInput_4,
      indexVec_checkResult_allDataPosition_4[32:11]};
  wire        indexVec_checkResult_unChange_4 = slideUp & (indexVec_readIndex_1[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_1 = validVec[1] & ~indexVec_checkResult_unChange_4;
  wire        indexVec_checkResult_1_4_1 = indexVec_checkResult_overlap_4 | ~indexVec_checkResult_1_5_1 | lagerThanVL | indexVec_checkResult_unChange_4;
  wire [33:0] indexVec_checkResult_allDataPosition_5 = {indexVec_readIndex_1, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_5 = indexVec_checkResult_allDataPosition_5[10:0];
  wire [4:0]  indexVec_checkResult_2_1_1 = indexVec_checkResult_dataPosition_5[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_5 = indexVec_checkResult_dataPosition_5[10:7];
  wire        indexVec_checkResult_2_2_1 = indexVec_checkResult_dataGroup_5[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_5 = indexVec_checkResult_dataGroup_5[3:1];
  wire [2:0]  indexVec_checkResult_2_3_1 = indexVec_checkResult_accessRegGrowth_5;
  wire [5:0]  indexVec_checkResult_decimalProportion_5 = {indexVec_checkResult_2_2_1, indexVec_checkResult_2_1_1};
  wire [2:0]  indexVec_checkResult_decimal_5 = indexVec_checkResult_decimalProportion_5[5:3];
  wire        indexVec_checkResult_overlap_5 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_5 >= indexVec_checkResult_intLMULInput_5[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_5} >= indexVec_checkResult_intLMULInput_5,
      indexVec_checkResult_allDataPosition_5[33:11]};
  wire        indexVec_checkResult_unChange_5 = slideUp & (indexVec_readIndex_1[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_1 = validVec[1] & ~indexVec_checkResult_unChange_5;
  wire        indexVec_checkResult_2_4_1 = indexVec_checkResult_overlap_5 | ~indexVec_checkResult_2_5_1 | lagerThanVL | indexVec_checkResult_unChange_5;
  wire [1:0]  indexVec_1_0 = (sew1H[0] ? indexVec_checkResult_0_0_1 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_1 : 2'h0);
  assign indexVec_1_1 = (sew1H[0] ? indexVec_checkResult_0_1_1 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_1 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_1 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_1_0 = indexVec_1_1;
  wire        indexVec_1_2 = sew1H[0] & indexVec_checkResult_0_2_1 | sew1H[1] & indexVec_checkResult_1_2_1 | sew1H[2] & indexVec_checkResult_2_2_1;
  assign indexVec_1_3 = (sew1H[0] ? indexVec_checkResult_0_3_1 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_1 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_1 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_1_0 = indexVec_1_3;
  wire        indexVec_1_4 = sew1H[0] & indexVec_checkResult_0_4_1 | sew1H[1] & indexVec_checkResult_1_4_1 | sew1H[2] & indexVec_checkResult_2_4_1;
  wire        indexVec_1_5 = sew1H[0] & indexVec_checkResult_0_5_1 | sew1H[1] & indexVec_checkResult_1_5_1 | sew1H[2] & indexVec_checkResult_2_5_1;
  wire [31:0] indexVec_readIndex_2 = baseIndex + 32'h2;
  wire [31:0] indexVec_checkResult_allDataPosition_6 = indexVec_readIndex_2;
  wire [10:0] indexVec_checkResult_dataPosition_6 = indexVec_checkResult_allDataPosition_6[10:0];
  wire [1:0]  indexVec_checkResult_0_0_2 = indexVec_checkResult_dataPosition_6[1:0];
  wire [4:0]  indexVec_checkResult_0_1_2 = indexVec_checkResult_dataPosition_6[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_6 = indexVec_checkResult_dataPosition_6[10:7];
  wire        indexVec_checkResult_0_2_2 = indexVec_checkResult_dataGroup_6[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_6 = indexVec_checkResult_dataGroup_6[3:1];
  wire [2:0]  indexVec_checkResult_0_3_2 = indexVec_checkResult_accessRegGrowth_6;
  wire [5:0]  indexVec_checkResult_decimalProportion_6 = {indexVec_checkResult_0_2_2, indexVec_checkResult_0_1_2};
  wire [2:0]  indexVec_checkResult_decimal_6 = indexVec_checkResult_decimalProportion_6[5:3];
  wire        indexVec_checkResult_overlap_6 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_6 >= indexVec_checkResult_intLMULInput_6[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_6} >= indexVec_checkResult_intLMULInput_6,
      indexVec_checkResult_allDataPosition_6[31:11]};
  wire        indexVec_checkResult_unChange_6 = slideUp & (indexVec_readIndex_2[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_2 = validVec[2] & ~indexVec_checkResult_unChange_6;
  wire        indexVec_checkResult_0_4_2 = indexVec_checkResult_overlap_6 | ~indexVec_checkResult_0_5_2 | lagerThanVL | indexVec_checkResult_unChange_6;
  wire [32:0] indexVec_checkResult_allDataPosition_7 = {indexVec_readIndex_2, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_7 = indexVec_checkResult_allDataPosition_7[10:0];
  wire [1:0]  indexVec_checkResult_1_0_2 = {indexVec_checkResult_dataPosition_7[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_2 = indexVec_checkResult_dataPosition_7[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_7 = indexVec_checkResult_dataPosition_7[10:7];
  wire        indexVec_checkResult_1_2_2 = indexVec_checkResult_dataGroup_7[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_7 = indexVec_checkResult_dataGroup_7[3:1];
  wire [2:0]  indexVec_checkResult_1_3_2 = indexVec_checkResult_accessRegGrowth_7;
  wire [5:0]  indexVec_checkResult_decimalProportion_7 = {indexVec_checkResult_1_2_2, indexVec_checkResult_1_1_2};
  wire [2:0]  indexVec_checkResult_decimal_7 = indexVec_checkResult_decimalProportion_7[5:3];
  wire        indexVec_checkResult_overlap_7 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_7 >= indexVec_checkResult_intLMULInput_7[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_7} >= indexVec_checkResult_intLMULInput_7,
      indexVec_checkResult_allDataPosition_7[32:11]};
  wire        indexVec_checkResult_unChange_7 = slideUp & (indexVec_readIndex_2[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_2 = validVec[2] & ~indexVec_checkResult_unChange_7;
  wire        indexVec_checkResult_1_4_2 = indexVec_checkResult_overlap_7 | ~indexVec_checkResult_1_5_2 | lagerThanVL | indexVec_checkResult_unChange_7;
  wire [33:0] indexVec_checkResult_allDataPosition_8 = {indexVec_readIndex_2, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_8 = indexVec_checkResult_allDataPosition_8[10:0];
  wire [4:0]  indexVec_checkResult_2_1_2 = indexVec_checkResult_dataPosition_8[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_8 = indexVec_checkResult_dataPosition_8[10:7];
  wire        indexVec_checkResult_2_2_2 = indexVec_checkResult_dataGroup_8[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_8 = indexVec_checkResult_dataGroup_8[3:1];
  wire [2:0]  indexVec_checkResult_2_3_2 = indexVec_checkResult_accessRegGrowth_8;
  wire [5:0]  indexVec_checkResult_decimalProportion_8 = {indexVec_checkResult_2_2_2, indexVec_checkResult_2_1_2};
  wire [2:0]  indexVec_checkResult_decimal_8 = indexVec_checkResult_decimalProportion_8[5:3];
  wire        indexVec_checkResult_overlap_8 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_8 >= indexVec_checkResult_intLMULInput_8[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_8} >= indexVec_checkResult_intLMULInput_8,
      indexVec_checkResult_allDataPosition_8[33:11]};
  wire        indexVec_checkResult_unChange_8 = slideUp & (indexVec_readIndex_2[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_2 = validVec[2] & ~indexVec_checkResult_unChange_8;
  wire        indexVec_checkResult_2_4_2 = indexVec_checkResult_overlap_8 | ~indexVec_checkResult_2_5_2 | lagerThanVL | indexVec_checkResult_unChange_8;
  wire [1:0]  indexVec_2_0 = (sew1H[0] ? indexVec_checkResult_0_0_2 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_2 : 2'h0);
  assign indexVec_2_1 = (sew1H[0] ? indexVec_checkResult_0_1_2 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_2 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_2 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_2_0 = indexVec_2_1;
  wire        indexVec_2_2 = sew1H[0] & indexVec_checkResult_0_2_2 | sew1H[1] & indexVec_checkResult_1_2_2 | sew1H[2] & indexVec_checkResult_2_2_2;
  assign indexVec_2_3 = (sew1H[0] ? indexVec_checkResult_0_3_2 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_2 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_2 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_2_0 = indexVec_2_3;
  wire        indexVec_2_4 = sew1H[0] & indexVec_checkResult_0_4_2 | sew1H[1] & indexVec_checkResult_1_4_2 | sew1H[2] & indexVec_checkResult_2_4_2;
  wire        indexVec_2_5 = sew1H[0] & indexVec_checkResult_0_5_2 | sew1H[1] & indexVec_checkResult_1_5_2 | sew1H[2] & indexVec_checkResult_2_5_2;
  wire [31:0] indexVec_readIndex_3 = baseIndex + 32'h3;
  wire [31:0] indexVec_checkResult_allDataPosition_9 = indexVec_readIndex_3;
  wire [10:0] indexVec_checkResult_dataPosition_9 = indexVec_checkResult_allDataPosition_9[10:0];
  wire [1:0]  indexVec_checkResult_0_0_3 = indexVec_checkResult_dataPosition_9[1:0];
  wire [4:0]  indexVec_checkResult_0_1_3 = indexVec_checkResult_dataPosition_9[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_9 = indexVec_checkResult_dataPosition_9[10:7];
  wire        indexVec_checkResult_0_2_3 = indexVec_checkResult_dataGroup_9[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_9 = indexVec_checkResult_dataGroup_9[3:1];
  wire [2:0]  indexVec_checkResult_0_3_3 = indexVec_checkResult_accessRegGrowth_9;
  wire [5:0]  indexVec_checkResult_decimalProportion_9 = {indexVec_checkResult_0_2_3, indexVec_checkResult_0_1_3};
  wire [2:0]  indexVec_checkResult_decimal_9 = indexVec_checkResult_decimalProportion_9[5:3];
  wire        indexVec_checkResult_overlap_9 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_9 >= indexVec_checkResult_intLMULInput_9[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_9} >= indexVec_checkResult_intLMULInput_9,
      indexVec_checkResult_allDataPosition_9[31:11]};
  wire        indexVec_checkResult_unChange_9 = slideUp & (indexVec_readIndex_3[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_3 = validVec[3] & ~indexVec_checkResult_unChange_9;
  wire        indexVec_checkResult_0_4_3 = indexVec_checkResult_overlap_9 | ~indexVec_checkResult_0_5_3 | lagerThanVL | indexVec_checkResult_unChange_9;
  wire [32:0] indexVec_checkResult_allDataPosition_10 = {indexVec_readIndex_3, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_10 = indexVec_checkResult_allDataPosition_10[10:0];
  wire [1:0]  indexVec_checkResult_1_0_3 = {indexVec_checkResult_dataPosition_10[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_3 = indexVec_checkResult_dataPosition_10[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_10 = indexVec_checkResult_dataPosition_10[10:7];
  wire        indexVec_checkResult_1_2_3 = indexVec_checkResult_dataGroup_10[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_10 = indexVec_checkResult_dataGroup_10[3:1];
  wire [2:0]  indexVec_checkResult_1_3_3 = indexVec_checkResult_accessRegGrowth_10;
  wire [5:0]  indexVec_checkResult_decimalProportion_10 = {indexVec_checkResult_1_2_3, indexVec_checkResult_1_1_3};
  wire [2:0]  indexVec_checkResult_decimal_10 = indexVec_checkResult_decimalProportion_10[5:3];
  wire        indexVec_checkResult_overlap_10 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_10 >= indexVec_checkResult_intLMULInput_10[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_10} >= indexVec_checkResult_intLMULInput_10,
      indexVec_checkResult_allDataPosition_10[32:11]};
  wire        indexVec_checkResult_unChange_10 = slideUp & (indexVec_readIndex_3[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_3 = validVec[3] & ~indexVec_checkResult_unChange_10;
  wire        indexVec_checkResult_1_4_3 = indexVec_checkResult_overlap_10 | ~indexVec_checkResult_1_5_3 | lagerThanVL | indexVec_checkResult_unChange_10;
  wire [33:0] indexVec_checkResult_allDataPosition_11 = {indexVec_readIndex_3, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_11 = indexVec_checkResult_allDataPosition_11[10:0];
  wire [4:0]  indexVec_checkResult_2_1_3 = indexVec_checkResult_dataPosition_11[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_11 = indexVec_checkResult_dataPosition_11[10:7];
  wire        indexVec_checkResult_2_2_3 = indexVec_checkResult_dataGroup_11[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_11 = indexVec_checkResult_dataGroup_11[3:1];
  wire [2:0]  indexVec_checkResult_2_3_3 = indexVec_checkResult_accessRegGrowth_11;
  wire [5:0]  indexVec_checkResult_decimalProportion_11 = {indexVec_checkResult_2_2_3, indexVec_checkResult_2_1_3};
  wire [2:0]  indexVec_checkResult_decimal_11 = indexVec_checkResult_decimalProportion_11[5:3];
  wire        indexVec_checkResult_overlap_11 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_11 >= indexVec_checkResult_intLMULInput_11[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_11} >= indexVec_checkResult_intLMULInput_11,
      indexVec_checkResult_allDataPosition_11[33:11]};
  wire        indexVec_checkResult_unChange_11 = slideUp & (indexVec_readIndex_3[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_3 = validVec[3] & ~indexVec_checkResult_unChange_11;
  wire        indexVec_checkResult_2_4_3 = indexVec_checkResult_overlap_11 | ~indexVec_checkResult_2_5_3 | lagerThanVL | indexVec_checkResult_unChange_11;
  wire [1:0]  indexVec_3_0 = (sew1H[0] ? indexVec_checkResult_0_0_3 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_3 : 2'h0);
  assign indexVec_3_1 = (sew1H[0] ? indexVec_checkResult_0_1_3 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_3 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_3 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_3_0 = indexVec_3_1;
  wire        indexVec_3_2 = sew1H[0] & indexVec_checkResult_0_2_3 | sew1H[1] & indexVec_checkResult_1_2_3 | sew1H[2] & indexVec_checkResult_2_2_3;
  assign indexVec_3_3 = (sew1H[0] ? indexVec_checkResult_0_3_3 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_3 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_3 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_3_0 = indexVec_3_3;
  wire        indexVec_3_4 = sew1H[0] & indexVec_checkResult_0_4_3 | sew1H[1] & indexVec_checkResult_1_4_3 | sew1H[2] & indexVec_checkResult_2_4_3;
  wire        indexVec_3_5 = sew1H[0] & indexVec_checkResult_0_5_3 | sew1H[1] & indexVec_checkResult_1_5_3 | sew1H[2] & indexVec_checkResult_2_5_3;
  wire [31:0] indexVec_readIndex_4 = baseIndex + 32'h4;
  wire [31:0] indexVec_checkResult_allDataPosition_12 = indexVec_readIndex_4;
  wire [10:0] indexVec_checkResult_dataPosition_12 = indexVec_checkResult_allDataPosition_12[10:0];
  wire [1:0]  indexVec_checkResult_0_0_4 = indexVec_checkResult_dataPosition_12[1:0];
  wire [4:0]  indexVec_checkResult_0_1_4 = indexVec_checkResult_dataPosition_12[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_12 = indexVec_checkResult_dataPosition_12[10:7];
  wire        indexVec_checkResult_0_2_4 = indexVec_checkResult_dataGroup_12[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_12 = indexVec_checkResult_dataGroup_12[3:1];
  wire [2:0]  indexVec_checkResult_0_3_4 = indexVec_checkResult_accessRegGrowth_12;
  wire [5:0]  indexVec_checkResult_decimalProportion_12 = {indexVec_checkResult_0_2_4, indexVec_checkResult_0_1_4};
  wire [2:0]  indexVec_checkResult_decimal_12 = indexVec_checkResult_decimalProportion_12[5:3];
  wire        indexVec_checkResult_overlap_12 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_12 >= indexVec_checkResult_intLMULInput_12[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_12} >= indexVec_checkResult_intLMULInput_12,
      indexVec_checkResult_allDataPosition_12[31:11]};
  wire        indexVec_checkResult_unChange_12 = slideUp & (indexVec_readIndex_4[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_4 = validVec[4] & ~indexVec_checkResult_unChange_12;
  wire        indexVec_checkResult_0_4_4 = indexVec_checkResult_overlap_12 | ~indexVec_checkResult_0_5_4 | lagerThanVL | indexVec_checkResult_unChange_12;
  wire [32:0] indexVec_checkResult_allDataPosition_13 = {indexVec_readIndex_4, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_13 = indexVec_checkResult_allDataPosition_13[10:0];
  wire [1:0]  indexVec_checkResult_1_0_4 = {indexVec_checkResult_dataPosition_13[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_4 = indexVec_checkResult_dataPosition_13[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_13 = indexVec_checkResult_dataPosition_13[10:7];
  wire        indexVec_checkResult_1_2_4 = indexVec_checkResult_dataGroup_13[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_13 = indexVec_checkResult_dataGroup_13[3:1];
  wire [2:0]  indexVec_checkResult_1_3_4 = indexVec_checkResult_accessRegGrowth_13;
  wire [5:0]  indexVec_checkResult_decimalProportion_13 = {indexVec_checkResult_1_2_4, indexVec_checkResult_1_1_4};
  wire [2:0]  indexVec_checkResult_decimal_13 = indexVec_checkResult_decimalProportion_13[5:3];
  wire        indexVec_checkResult_overlap_13 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_13 >= indexVec_checkResult_intLMULInput_13[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_13} >= indexVec_checkResult_intLMULInput_13,
      indexVec_checkResult_allDataPosition_13[32:11]};
  wire        indexVec_checkResult_unChange_13 = slideUp & (indexVec_readIndex_4[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_4 = validVec[4] & ~indexVec_checkResult_unChange_13;
  wire        indexVec_checkResult_1_4_4 = indexVec_checkResult_overlap_13 | ~indexVec_checkResult_1_5_4 | lagerThanVL | indexVec_checkResult_unChange_13;
  wire [33:0] indexVec_checkResult_allDataPosition_14 = {indexVec_readIndex_4, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_14 = indexVec_checkResult_allDataPosition_14[10:0];
  wire [4:0]  indexVec_checkResult_2_1_4 = indexVec_checkResult_dataPosition_14[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_14 = indexVec_checkResult_dataPosition_14[10:7];
  wire        indexVec_checkResult_2_2_4 = indexVec_checkResult_dataGroup_14[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_14 = indexVec_checkResult_dataGroup_14[3:1];
  wire [2:0]  indexVec_checkResult_2_3_4 = indexVec_checkResult_accessRegGrowth_14;
  wire [5:0]  indexVec_checkResult_decimalProportion_14 = {indexVec_checkResult_2_2_4, indexVec_checkResult_2_1_4};
  wire [2:0]  indexVec_checkResult_decimal_14 = indexVec_checkResult_decimalProportion_14[5:3];
  wire        indexVec_checkResult_overlap_14 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_14 >= indexVec_checkResult_intLMULInput_14[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_14} >= indexVec_checkResult_intLMULInput_14,
      indexVec_checkResult_allDataPosition_14[33:11]};
  wire        indexVec_checkResult_unChange_14 = slideUp & (indexVec_readIndex_4[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_4 = validVec[4] & ~indexVec_checkResult_unChange_14;
  wire        indexVec_checkResult_2_4_4 = indexVec_checkResult_overlap_14 | ~indexVec_checkResult_2_5_4 | lagerThanVL | indexVec_checkResult_unChange_14;
  wire [1:0]  indexVec_4_0 = (sew1H[0] ? indexVec_checkResult_0_0_4 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_4 : 2'h0);
  assign indexVec_4_1 = (sew1H[0] ? indexVec_checkResult_0_1_4 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_4 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_4 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_4_0 = indexVec_4_1;
  wire        indexVec_4_2 = sew1H[0] & indexVec_checkResult_0_2_4 | sew1H[1] & indexVec_checkResult_1_2_4 | sew1H[2] & indexVec_checkResult_2_2_4;
  assign indexVec_4_3 = (sew1H[0] ? indexVec_checkResult_0_3_4 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_4 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_4 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_4_0 = indexVec_4_3;
  wire        indexVec_4_4 = sew1H[0] & indexVec_checkResult_0_4_4 | sew1H[1] & indexVec_checkResult_1_4_4 | sew1H[2] & indexVec_checkResult_2_4_4;
  wire        indexVec_4_5 = sew1H[0] & indexVec_checkResult_0_5_4 | sew1H[1] & indexVec_checkResult_1_5_4 | sew1H[2] & indexVec_checkResult_2_5_4;
  wire [31:0] indexVec_readIndex_5 = baseIndex + 32'h5;
  wire [31:0] indexVec_checkResult_allDataPosition_15 = indexVec_readIndex_5;
  wire [10:0] indexVec_checkResult_dataPosition_15 = indexVec_checkResult_allDataPosition_15[10:0];
  wire [1:0]  indexVec_checkResult_0_0_5 = indexVec_checkResult_dataPosition_15[1:0];
  wire [4:0]  indexVec_checkResult_0_1_5 = indexVec_checkResult_dataPosition_15[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_15 = indexVec_checkResult_dataPosition_15[10:7];
  wire        indexVec_checkResult_0_2_5 = indexVec_checkResult_dataGroup_15[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_15 = indexVec_checkResult_dataGroup_15[3:1];
  wire [2:0]  indexVec_checkResult_0_3_5 = indexVec_checkResult_accessRegGrowth_15;
  wire [5:0]  indexVec_checkResult_decimalProportion_15 = {indexVec_checkResult_0_2_5, indexVec_checkResult_0_1_5};
  wire [2:0]  indexVec_checkResult_decimal_15 = indexVec_checkResult_decimalProportion_15[5:3];
  wire        indexVec_checkResult_overlap_15 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_15 >= indexVec_checkResult_intLMULInput_15[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_15} >= indexVec_checkResult_intLMULInput_15,
      indexVec_checkResult_allDataPosition_15[31:11]};
  wire        indexVec_checkResult_unChange_15 = slideUp & (indexVec_readIndex_5[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_5 = validVec[5] & ~indexVec_checkResult_unChange_15;
  wire        indexVec_checkResult_0_4_5 = indexVec_checkResult_overlap_15 | ~indexVec_checkResult_0_5_5 | lagerThanVL | indexVec_checkResult_unChange_15;
  wire [32:0] indexVec_checkResult_allDataPosition_16 = {indexVec_readIndex_5, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_16 = indexVec_checkResult_allDataPosition_16[10:0];
  wire [1:0]  indexVec_checkResult_1_0_5 = {indexVec_checkResult_dataPosition_16[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_5 = indexVec_checkResult_dataPosition_16[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_16 = indexVec_checkResult_dataPosition_16[10:7];
  wire        indexVec_checkResult_1_2_5 = indexVec_checkResult_dataGroup_16[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_16 = indexVec_checkResult_dataGroup_16[3:1];
  wire [2:0]  indexVec_checkResult_1_3_5 = indexVec_checkResult_accessRegGrowth_16;
  wire [5:0]  indexVec_checkResult_decimalProportion_16 = {indexVec_checkResult_1_2_5, indexVec_checkResult_1_1_5};
  wire [2:0]  indexVec_checkResult_decimal_16 = indexVec_checkResult_decimalProportion_16[5:3];
  wire        indexVec_checkResult_overlap_16 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_16 >= indexVec_checkResult_intLMULInput_16[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_16} >= indexVec_checkResult_intLMULInput_16,
      indexVec_checkResult_allDataPosition_16[32:11]};
  wire        indexVec_checkResult_unChange_16 = slideUp & (indexVec_readIndex_5[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_5 = validVec[5] & ~indexVec_checkResult_unChange_16;
  wire        indexVec_checkResult_1_4_5 = indexVec_checkResult_overlap_16 | ~indexVec_checkResult_1_5_5 | lagerThanVL | indexVec_checkResult_unChange_16;
  wire [33:0] indexVec_checkResult_allDataPosition_17 = {indexVec_readIndex_5, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_17 = indexVec_checkResult_allDataPosition_17[10:0];
  wire [4:0]  indexVec_checkResult_2_1_5 = indexVec_checkResult_dataPosition_17[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_17 = indexVec_checkResult_dataPosition_17[10:7];
  wire        indexVec_checkResult_2_2_5 = indexVec_checkResult_dataGroup_17[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_17 = indexVec_checkResult_dataGroup_17[3:1];
  wire [2:0]  indexVec_checkResult_2_3_5 = indexVec_checkResult_accessRegGrowth_17;
  wire [5:0]  indexVec_checkResult_decimalProportion_17 = {indexVec_checkResult_2_2_5, indexVec_checkResult_2_1_5};
  wire [2:0]  indexVec_checkResult_decimal_17 = indexVec_checkResult_decimalProportion_17[5:3];
  wire        indexVec_checkResult_overlap_17 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_17 >= indexVec_checkResult_intLMULInput_17[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_17} >= indexVec_checkResult_intLMULInput_17,
      indexVec_checkResult_allDataPosition_17[33:11]};
  wire        indexVec_checkResult_unChange_17 = slideUp & (indexVec_readIndex_5[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_5 = validVec[5] & ~indexVec_checkResult_unChange_17;
  wire        indexVec_checkResult_2_4_5 = indexVec_checkResult_overlap_17 | ~indexVec_checkResult_2_5_5 | lagerThanVL | indexVec_checkResult_unChange_17;
  wire [1:0]  indexVec_5_0 = (sew1H[0] ? indexVec_checkResult_0_0_5 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_5 : 2'h0);
  assign indexVec_5_1 = (sew1H[0] ? indexVec_checkResult_0_1_5 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_5 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_5 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_5_0 = indexVec_5_1;
  wire        indexVec_5_2 = sew1H[0] & indexVec_checkResult_0_2_5 | sew1H[1] & indexVec_checkResult_1_2_5 | sew1H[2] & indexVec_checkResult_2_2_5;
  assign indexVec_5_3 = (sew1H[0] ? indexVec_checkResult_0_3_5 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_5 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_5 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_5_0 = indexVec_5_3;
  wire        indexVec_5_4 = sew1H[0] & indexVec_checkResult_0_4_5 | sew1H[1] & indexVec_checkResult_1_4_5 | sew1H[2] & indexVec_checkResult_2_4_5;
  wire        indexVec_5_5 = sew1H[0] & indexVec_checkResult_0_5_5 | sew1H[1] & indexVec_checkResult_1_5_5 | sew1H[2] & indexVec_checkResult_2_5_5;
  wire [31:0] indexVec_readIndex_6 = baseIndex + 32'h6;
  wire [31:0] indexVec_checkResult_allDataPosition_18 = indexVec_readIndex_6;
  wire [10:0] indexVec_checkResult_dataPosition_18 = indexVec_checkResult_allDataPosition_18[10:0];
  wire [1:0]  indexVec_checkResult_0_0_6 = indexVec_checkResult_dataPosition_18[1:0];
  wire [4:0]  indexVec_checkResult_0_1_6 = indexVec_checkResult_dataPosition_18[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_18 = indexVec_checkResult_dataPosition_18[10:7];
  wire        indexVec_checkResult_0_2_6 = indexVec_checkResult_dataGroup_18[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_18 = indexVec_checkResult_dataGroup_18[3:1];
  wire [2:0]  indexVec_checkResult_0_3_6 = indexVec_checkResult_accessRegGrowth_18;
  wire [5:0]  indexVec_checkResult_decimalProportion_18 = {indexVec_checkResult_0_2_6, indexVec_checkResult_0_1_6};
  wire [2:0]  indexVec_checkResult_decimal_18 = indexVec_checkResult_decimalProportion_18[5:3];
  wire        indexVec_checkResult_overlap_18 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_18 >= indexVec_checkResult_intLMULInput_18[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_18} >= indexVec_checkResult_intLMULInput_18,
      indexVec_checkResult_allDataPosition_18[31:11]};
  wire        indexVec_checkResult_unChange_18 = slideUp & (indexVec_readIndex_6[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_6 = validVec[6] & ~indexVec_checkResult_unChange_18;
  wire        indexVec_checkResult_0_4_6 = indexVec_checkResult_overlap_18 | ~indexVec_checkResult_0_5_6 | lagerThanVL | indexVec_checkResult_unChange_18;
  wire [32:0] indexVec_checkResult_allDataPosition_19 = {indexVec_readIndex_6, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_19 = indexVec_checkResult_allDataPosition_19[10:0];
  wire [1:0]  indexVec_checkResult_1_0_6 = {indexVec_checkResult_dataPosition_19[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_6 = indexVec_checkResult_dataPosition_19[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_19 = indexVec_checkResult_dataPosition_19[10:7];
  wire        indexVec_checkResult_1_2_6 = indexVec_checkResult_dataGroup_19[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_19 = indexVec_checkResult_dataGroup_19[3:1];
  wire [2:0]  indexVec_checkResult_1_3_6 = indexVec_checkResult_accessRegGrowth_19;
  wire [5:0]  indexVec_checkResult_decimalProportion_19 = {indexVec_checkResult_1_2_6, indexVec_checkResult_1_1_6};
  wire [2:0]  indexVec_checkResult_decimal_19 = indexVec_checkResult_decimalProportion_19[5:3];
  wire        indexVec_checkResult_overlap_19 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_19 >= indexVec_checkResult_intLMULInput_19[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_19} >= indexVec_checkResult_intLMULInput_19,
      indexVec_checkResult_allDataPosition_19[32:11]};
  wire        indexVec_checkResult_unChange_19 = slideUp & (indexVec_readIndex_6[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_6 = validVec[6] & ~indexVec_checkResult_unChange_19;
  wire        indexVec_checkResult_1_4_6 = indexVec_checkResult_overlap_19 | ~indexVec_checkResult_1_5_6 | lagerThanVL | indexVec_checkResult_unChange_19;
  wire [33:0] indexVec_checkResult_allDataPosition_20 = {indexVec_readIndex_6, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_20 = indexVec_checkResult_allDataPosition_20[10:0];
  wire [4:0]  indexVec_checkResult_2_1_6 = indexVec_checkResult_dataPosition_20[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_20 = indexVec_checkResult_dataPosition_20[10:7];
  wire        indexVec_checkResult_2_2_6 = indexVec_checkResult_dataGroup_20[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_20 = indexVec_checkResult_dataGroup_20[3:1];
  wire [2:0]  indexVec_checkResult_2_3_6 = indexVec_checkResult_accessRegGrowth_20;
  wire [5:0]  indexVec_checkResult_decimalProportion_20 = {indexVec_checkResult_2_2_6, indexVec_checkResult_2_1_6};
  wire [2:0]  indexVec_checkResult_decimal_20 = indexVec_checkResult_decimalProportion_20[5:3];
  wire        indexVec_checkResult_overlap_20 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_20 >= indexVec_checkResult_intLMULInput_20[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_20} >= indexVec_checkResult_intLMULInput_20,
      indexVec_checkResult_allDataPosition_20[33:11]};
  wire        indexVec_checkResult_unChange_20 = slideUp & (indexVec_readIndex_6[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_6 = validVec[6] & ~indexVec_checkResult_unChange_20;
  wire        indexVec_checkResult_2_4_6 = indexVec_checkResult_overlap_20 | ~indexVec_checkResult_2_5_6 | lagerThanVL | indexVec_checkResult_unChange_20;
  wire [1:0]  indexVec_6_0 = (sew1H[0] ? indexVec_checkResult_0_0_6 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_6 : 2'h0);
  assign indexVec_6_1 = (sew1H[0] ? indexVec_checkResult_0_1_6 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_6 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_6 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_6_0 = indexVec_6_1;
  wire        indexVec_6_2 = sew1H[0] & indexVec_checkResult_0_2_6 | sew1H[1] & indexVec_checkResult_1_2_6 | sew1H[2] & indexVec_checkResult_2_2_6;
  assign indexVec_6_3 = (sew1H[0] ? indexVec_checkResult_0_3_6 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_6 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_6 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_6_0 = indexVec_6_3;
  wire        indexVec_6_4 = sew1H[0] & indexVec_checkResult_0_4_6 | sew1H[1] & indexVec_checkResult_1_4_6 | sew1H[2] & indexVec_checkResult_2_4_6;
  wire        indexVec_6_5 = sew1H[0] & indexVec_checkResult_0_5_6 | sew1H[1] & indexVec_checkResult_1_5_6 | sew1H[2] & indexVec_checkResult_2_5_6;
  wire [31:0] indexVec_readIndex_7 = baseIndex + 32'h7;
  wire [31:0] indexVec_checkResult_allDataPosition_21 = indexVec_readIndex_7;
  wire [10:0] indexVec_checkResult_dataPosition_21 = indexVec_checkResult_allDataPosition_21[10:0];
  wire [1:0]  indexVec_checkResult_0_0_7 = indexVec_checkResult_dataPosition_21[1:0];
  wire [4:0]  indexVec_checkResult_0_1_7 = indexVec_checkResult_dataPosition_21[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_21 = indexVec_checkResult_dataPosition_21[10:7];
  wire        indexVec_checkResult_0_2_7 = indexVec_checkResult_dataGroup_21[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_21 = indexVec_checkResult_dataGroup_21[3:1];
  wire [2:0]  indexVec_checkResult_0_3_7 = indexVec_checkResult_accessRegGrowth_21;
  wire [5:0]  indexVec_checkResult_decimalProportion_21 = {indexVec_checkResult_0_2_7, indexVec_checkResult_0_1_7};
  wire [2:0]  indexVec_checkResult_decimal_21 = indexVec_checkResult_decimalProportion_21[5:3];
  wire        indexVec_checkResult_overlap_21 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_21 >= indexVec_checkResult_intLMULInput_21[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_21} >= indexVec_checkResult_intLMULInput_21,
      indexVec_checkResult_allDataPosition_21[31:11]};
  wire        indexVec_checkResult_unChange_21 = slideUp & (indexVec_readIndex_7[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_7 = validVec[7] & ~indexVec_checkResult_unChange_21;
  wire        indexVec_checkResult_0_4_7 = indexVec_checkResult_overlap_21 | ~indexVec_checkResult_0_5_7 | lagerThanVL | indexVec_checkResult_unChange_21;
  wire [32:0] indexVec_checkResult_allDataPosition_22 = {indexVec_readIndex_7, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_22 = indexVec_checkResult_allDataPosition_22[10:0];
  wire [1:0]  indexVec_checkResult_1_0_7 = {indexVec_checkResult_dataPosition_22[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_7 = indexVec_checkResult_dataPosition_22[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_22 = indexVec_checkResult_dataPosition_22[10:7];
  wire        indexVec_checkResult_1_2_7 = indexVec_checkResult_dataGroup_22[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_22 = indexVec_checkResult_dataGroup_22[3:1];
  wire [2:0]  indexVec_checkResult_1_3_7 = indexVec_checkResult_accessRegGrowth_22;
  wire [5:0]  indexVec_checkResult_decimalProportion_22 = {indexVec_checkResult_1_2_7, indexVec_checkResult_1_1_7};
  wire [2:0]  indexVec_checkResult_decimal_22 = indexVec_checkResult_decimalProportion_22[5:3];
  wire        indexVec_checkResult_overlap_22 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_22 >= indexVec_checkResult_intLMULInput_22[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_22} >= indexVec_checkResult_intLMULInput_22,
      indexVec_checkResult_allDataPosition_22[32:11]};
  wire        indexVec_checkResult_unChange_22 = slideUp & (indexVec_readIndex_7[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_7 = validVec[7] & ~indexVec_checkResult_unChange_22;
  wire        indexVec_checkResult_1_4_7 = indexVec_checkResult_overlap_22 | ~indexVec_checkResult_1_5_7 | lagerThanVL | indexVec_checkResult_unChange_22;
  wire [33:0] indexVec_checkResult_allDataPosition_23 = {indexVec_readIndex_7, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_23 = indexVec_checkResult_allDataPosition_23[10:0];
  wire [4:0]  indexVec_checkResult_2_1_7 = indexVec_checkResult_dataPosition_23[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_23 = indexVec_checkResult_dataPosition_23[10:7];
  wire        indexVec_checkResult_2_2_7 = indexVec_checkResult_dataGroup_23[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_23 = indexVec_checkResult_dataGroup_23[3:1];
  wire [2:0]  indexVec_checkResult_2_3_7 = indexVec_checkResult_accessRegGrowth_23;
  wire [5:0]  indexVec_checkResult_decimalProportion_23 = {indexVec_checkResult_2_2_7, indexVec_checkResult_2_1_7};
  wire [2:0]  indexVec_checkResult_decimal_23 = indexVec_checkResult_decimalProportion_23[5:3];
  wire        indexVec_checkResult_overlap_23 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_23 >= indexVec_checkResult_intLMULInput_23[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_23} >= indexVec_checkResult_intLMULInput_23,
      indexVec_checkResult_allDataPosition_23[33:11]};
  wire        indexVec_checkResult_unChange_23 = slideUp & (indexVec_readIndex_7[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_7 = validVec[7] & ~indexVec_checkResult_unChange_23;
  wire        indexVec_checkResult_2_4_7 = indexVec_checkResult_overlap_23 | ~indexVec_checkResult_2_5_7 | lagerThanVL | indexVec_checkResult_unChange_23;
  wire [1:0]  indexVec_7_0 = (sew1H[0] ? indexVec_checkResult_0_0_7 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_7 : 2'h0);
  assign indexVec_7_1 = (sew1H[0] ? indexVec_checkResult_0_1_7 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_7 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_7 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_7_0 = indexVec_7_1;
  wire        indexVec_7_2 = sew1H[0] & indexVec_checkResult_0_2_7 | sew1H[1] & indexVec_checkResult_1_2_7 | sew1H[2] & indexVec_checkResult_2_2_7;
  assign indexVec_7_3 = (sew1H[0] ? indexVec_checkResult_0_3_7 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_7 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_7 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_7_0 = indexVec_7_3;
  wire        indexVec_7_4 = sew1H[0] & indexVec_checkResult_0_4_7 | sew1H[1] & indexVec_checkResult_1_4_7 | sew1H[2] & indexVec_checkResult_2_4_7;
  wire        indexVec_7_5 = sew1H[0] & indexVec_checkResult_0_5_7 | sew1H[1] & indexVec_checkResult_1_5_7 | sew1H[2] & indexVec_checkResult_2_5_7;
  wire [31:0] indexVec_readIndex_8 = baseIndex + 32'h8;
  wire [31:0] indexVec_checkResult_allDataPosition_24 = indexVec_readIndex_8;
  wire [10:0] indexVec_checkResult_dataPosition_24 = indexVec_checkResult_allDataPosition_24[10:0];
  wire [1:0]  indexVec_checkResult_0_0_8 = indexVec_checkResult_dataPosition_24[1:0];
  wire [4:0]  indexVec_checkResult_0_1_8 = indexVec_checkResult_dataPosition_24[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_24 = indexVec_checkResult_dataPosition_24[10:7];
  wire        indexVec_checkResult_0_2_8 = indexVec_checkResult_dataGroup_24[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_24 = indexVec_checkResult_dataGroup_24[3:1];
  wire [2:0]  indexVec_checkResult_0_3_8 = indexVec_checkResult_accessRegGrowth_24;
  wire [5:0]  indexVec_checkResult_decimalProportion_24 = {indexVec_checkResult_0_2_8, indexVec_checkResult_0_1_8};
  wire [2:0]  indexVec_checkResult_decimal_24 = indexVec_checkResult_decimalProportion_24[5:3];
  wire        indexVec_checkResult_overlap_24 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_24 >= indexVec_checkResult_intLMULInput_24[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_24} >= indexVec_checkResult_intLMULInput_24,
      indexVec_checkResult_allDataPosition_24[31:11]};
  wire        indexVec_checkResult_unChange_24 = slideUp & (indexVec_readIndex_8[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_8 = validVec[8] & ~indexVec_checkResult_unChange_24;
  wire        indexVec_checkResult_0_4_8 = indexVec_checkResult_overlap_24 | ~indexVec_checkResult_0_5_8 | lagerThanVL | indexVec_checkResult_unChange_24;
  wire [32:0] indexVec_checkResult_allDataPosition_25 = {indexVec_readIndex_8, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_25 = indexVec_checkResult_allDataPosition_25[10:0];
  wire [1:0]  indexVec_checkResult_1_0_8 = {indexVec_checkResult_dataPosition_25[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_8 = indexVec_checkResult_dataPosition_25[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_25 = indexVec_checkResult_dataPosition_25[10:7];
  wire        indexVec_checkResult_1_2_8 = indexVec_checkResult_dataGroup_25[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_25 = indexVec_checkResult_dataGroup_25[3:1];
  wire [2:0]  indexVec_checkResult_1_3_8 = indexVec_checkResult_accessRegGrowth_25;
  wire [5:0]  indexVec_checkResult_decimalProportion_25 = {indexVec_checkResult_1_2_8, indexVec_checkResult_1_1_8};
  wire [2:0]  indexVec_checkResult_decimal_25 = indexVec_checkResult_decimalProportion_25[5:3];
  wire        indexVec_checkResult_overlap_25 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_25 >= indexVec_checkResult_intLMULInput_25[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_25} >= indexVec_checkResult_intLMULInput_25,
      indexVec_checkResult_allDataPosition_25[32:11]};
  wire        indexVec_checkResult_unChange_25 = slideUp & (indexVec_readIndex_8[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_8 = validVec[8] & ~indexVec_checkResult_unChange_25;
  wire        indexVec_checkResult_1_4_8 = indexVec_checkResult_overlap_25 | ~indexVec_checkResult_1_5_8 | lagerThanVL | indexVec_checkResult_unChange_25;
  wire [33:0] indexVec_checkResult_allDataPosition_26 = {indexVec_readIndex_8, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_26 = indexVec_checkResult_allDataPosition_26[10:0];
  wire [4:0]  indexVec_checkResult_2_1_8 = indexVec_checkResult_dataPosition_26[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_26 = indexVec_checkResult_dataPosition_26[10:7];
  wire        indexVec_checkResult_2_2_8 = indexVec_checkResult_dataGroup_26[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_26 = indexVec_checkResult_dataGroup_26[3:1];
  wire [2:0]  indexVec_checkResult_2_3_8 = indexVec_checkResult_accessRegGrowth_26;
  wire [5:0]  indexVec_checkResult_decimalProportion_26 = {indexVec_checkResult_2_2_8, indexVec_checkResult_2_1_8};
  wire [2:0]  indexVec_checkResult_decimal_26 = indexVec_checkResult_decimalProportion_26[5:3];
  wire        indexVec_checkResult_overlap_26 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_26 >= indexVec_checkResult_intLMULInput_26[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_26} >= indexVec_checkResult_intLMULInput_26,
      indexVec_checkResult_allDataPosition_26[33:11]};
  wire        indexVec_checkResult_unChange_26 = slideUp & (indexVec_readIndex_8[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_8 = validVec[8] & ~indexVec_checkResult_unChange_26;
  wire        indexVec_checkResult_2_4_8 = indexVec_checkResult_overlap_26 | ~indexVec_checkResult_2_5_8 | lagerThanVL | indexVec_checkResult_unChange_26;
  wire [1:0]  indexVec_8_0 = (sew1H[0] ? indexVec_checkResult_0_0_8 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_8 : 2'h0);
  assign indexVec_8_1 = (sew1H[0] ? indexVec_checkResult_0_1_8 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_8 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_8 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_8_0 = indexVec_8_1;
  wire        indexVec_8_2 = sew1H[0] & indexVec_checkResult_0_2_8 | sew1H[1] & indexVec_checkResult_1_2_8 | sew1H[2] & indexVec_checkResult_2_2_8;
  assign indexVec_8_3 = (sew1H[0] ? indexVec_checkResult_0_3_8 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_8 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_8 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_8_0 = indexVec_8_3;
  wire        indexVec_8_4 = sew1H[0] & indexVec_checkResult_0_4_8 | sew1H[1] & indexVec_checkResult_1_4_8 | sew1H[2] & indexVec_checkResult_2_4_8;
  wire        indexVec_8_5 = sew1H[0] & indexVec_checkResult_0_5_8 | sew1H[1] & indexVec_checkResult_1_5_8 | sew1H[2] & indexVec_checkResult_2_5_8;
  wire [31:0] indexVec_readIndex_9 = baseIndex + 32'h9;
  wire [31:0] indexVec_checkResult_allDataPosition_27 = indexVec_readIndex_9;
  wire [10:0] indexVec_checkResult_dataPosition_27 = indexVec_checkResult_allDataPosition_27[10:0];
  wire [1:0]  indexVec_checkResult_0_0_9 = indexVec_checkResult_dataPosition_27[1:0];
  wire [4:0]  indexVec_checkResult_0_1_9 = indexVec_checkResult_dataPosition_27[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_27 = indexVec_checkResult_dataPosition_27[10:7];
  wire        indexVec_checkResult_0_2_9 = indexVec_checkResult_dataGroup_27[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_27 = indexVec_checkResult_dataGroup_27[3:1];
  wire [2:0]  indexVec_checkResult_0_3_9 = indexVec_checkResult_accessRegGrowth_27;
  wire [5:0]  indexVec_checkResult_decimalProportion_27 = {indexVec_checkResult_0_2_9, indexVec_checkResult_0_1_9};
  wire [2:0]  indexVec_checkResult_decimal_27 = indexVec_checkResult_decimalProportion_27[5:3];
  wire        indexVec_checkResult_overlap_27 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_27 >= indexVec_checkResult_intLMULInput_27[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_27} >= indexVec_checkResult_intLMULInput_27,
      indexVec_checkResult_allDataPosition_27[31:11]};
  wire        indexVec_checkResult_unChange_27 = slideUp & (indexVec_readIndex_9[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_9 = validVec[9] & ~indexVec_checkResult_unChange_27;
  wire        indexVec_checkResult_0_4_9 = indexVec_checkResult_overlap_27 | ~indexVec_checkResult_0_5_9 | lagerThanVL | indexVec_checkResult_unChange_27;
  wire [32:0] indexVec_checkResult_allDataPosition_28 = {indexVec_readIndex_9, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_28 = indexVec_checkResult_allDataPosition_28[10:0];
  wire [1:0]  indexVec_checkResult_1_0_9 = {indexVec_checkResult_dataPosition_28[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_9 = indexVec_checkResult_dataPosition_28[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_28 = indexVec_checkResult_dataPosition_28[10:7];
  wire        indexVec_checkResult_1_2_9 = indexVec_checkResult_dataGroup_28[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_28 = indexVec_checkResult_dataGroup_28[3:1];
  wire [2:0]  indexVec_checkResult_1_3_9 = indexVec_checkResult_accessRegGrowth_28;
  wire [5:0]  indexVec_checkResult_decimalProportion_28 = {indexVec_checkResult_1_2_9, indexVec_checkResult_1_1_9};
  wire [2:0]  indexVec_checkResult_decimal_28 = indexVec_checkResult_decimalProportion_28[5:3];
  wire        indexVec_checkResult_overlap_28 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_28 >= indexVec_checkResult_intLMULInput_28[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_28} >= indexVec_checkResult_intLMULInput_28,
      indexVec_checkResult_allDataPosition_28[32:11]};
  wire        indexVec_checkResult_unChange_28 = slideUp & (indexVec_readIndex_9[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_9 = validVec[9] & ~indexVec_checkResult_unChange_28;
  wire        indexVec_checkResult_1_4_9 = indexVec_checkResult_overlap_28 | ~indexVec_checkResult_1_5_9 | lagerThanVL | indexVec_checkResult_unChange_28;
  wire [33:0] indexVec_checkResult_allDataPosition_29 = {indexVec_readIndex_9, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_29 = indexVec_checkResult_allDataPosition_29[10:0];
  wire [4:0]  indexVec_checkResult_2_1_9 = indexVec_checkResult_dataPosition_29[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_29 = indexVec_checkResult_dataPosition_29[10:7];
  wire        indexVec_checkResult_2_2_9 = indexVec_checkResult_dataGroup_29[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_29 = indexVec_checkResult_dataGroup_29[3:1];
  wire [2:0]  indexVec_checkResult_2_3_9 = indexVec_checkResult_accessRegGrowth_29;
  wire [5:0]  indexVec_checkResult_decimalProportion_29 = {indexVec_checkResult_2_2_9, indexVec_checkResult_2_1_9};
  wire [2:0]  indexVec_checkResult_decimal_29 = indexVec_checkResult_decimalProportion_29[5:3];
  wire        indexVec_checkResult_overlap_29 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_29 >= indexVec_checkResult_intLMULInput_29[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_29} >= indexVec_checkResult_intLMULInput_29,
      indexVec_checkResult_allDataPosition_29[33:11]};
  wire        indexVec_checkResult_unChange_29 = slideUp & (indexVec_readIndex_9[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_9 = validVec[9] & ~indexVec_checkResult_unChange_29;
  wire        indexVec_checkResult_2_4_9 = indexVec_checkResult_overlap_29 | ~indexVec_checkResult_2_5_9 | lagerThanVL | indexVec_checkResult_unChange_29;
  wire [1:0]  indexVec_9_0 = (sew1H[0] ? indexVec_checkResult_0_0_9 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_9 : 2'h0);
  assign indexVec_9_1 = (sew1H[0] ? indexVec_checkResult_0_1_9 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_9 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_9 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_9_0 = indexVec_9_1;
  wire        indexVec_9_2 = sew1H[0] & indexVec_checkResult_0_2_9 | sew1H[1] & indexVec_checkResult_1_2_9 | sew1H[2] & indexVec_checkResult_2_2_9;
  assign indexVec_9_3 = (sew1H[0] ? indexVec_checkResult_0_3_9 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_9 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_9 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_9_0 = indexVec_9_3;
  wire        indexVec_9_4 = sew1H[0] & indexVec_checkResult_0_4_9 | sew1H[1] & indexVec_checkResult_1_4_9 | sew1H[2] & indexVec_checkResult_2_4_9;
  wire        indexVec_9_5 = sew1H[0] & indexVec_checkResult_0_5_9 | sew1H[1] & indexVec_checkResult_1_5_9 | sew1H[2] & indexVec_checkResult_2_5_9;
  wire [31:0] indexVec_readIndex_10 = baseIndex + 32'hA;
  wire [31:0] indexVec_checkResult_allDataPosition_30 = indexVec_readIndex_10;
  wire [10:0] indexVec_checkResult_dataPosition_30 = indexVec_checkResult_allDataPosition_30[10:0];
  wire [1:0]  indexVec_checkResult_0_0_10 = indexVec_checkResult_dataPosition_30[1:0];
  wire [4:0]  indexVec_checkResult_0_1_10 = indexVec_checkResult_dataPosition_30[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_30 = indexVec_checkResult_dataPosition_30[10:7];
  wire        indexVec_checkResult_0_2_10 = indexVec_checkResult_dataGroup_30[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_30 = indexVec_checkResult_dataGroup_30[3:1];
  wire [2:0]  indexVec_checkResult_0_3_10 = indexVec_checkResult_accessRegGrowth_30;
  wire [5:0]  indexVec_checkResult_decimalProportion_30 = {indexVec_checkResult_0_2_10, indexVec_checkResult_0_1_10};
  wire [2:0]  indexVec_checkResult_decimal_30 = indexVec_checkResult_decimalProportion_30[5:3];
  wire        indexVec_checkResult_overlap_30 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_30 >= indexVec_checkResult_intLMULInput_30[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_30} >= indexVec_checkResult_intLMULInput_30,
      indexVec_checkResult_allDataPosition_30[31:11]};
  wire        indexVec_checkResult_unChange_30 = slideUp & (indexVec_readIndex_10[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_10 = validVec[10] & ~indexVec_checkResult_unChange_30;
  wire        indexVec_checkResult_0_4_10 = indexVec_checkResult_overlap_30 | ~indexVec_checkResult_0_5_10 | lagerThanVL | indexVec_checkResult_unChange_30;
  wire [32:0] indexVec_checkResult_allDataPosition_31 = {indexVec_readIndex_10, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_31 = indexVec_checkResult_allDataPosition_31[10:0];
  wire [1:0]  indexVec_checkResult_1_0_10 = {indexVec_checkResult_dataPosition_31[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_10 = indexVec_checkResult_dataPosition_31[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_31 = indexVec_checkResult_dataPosition_31[10:7];
  wire        indexVec_checkResult_1_2_10 = indexVec_checkResult_dataGroup_31[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_31 = indexVec_checkResult_dataGroup_31[3:1];
  wire [2:0]  indexVec_checkResult_1_3_10 = indexVec_checkResult_accessRegGrowth_31;
  wire [5:0]  indexVec_checkResult_decimalProportion_31 = {indexVec_checkResult_1_2_10, indexVec_checkResult_1_1_10};
  wire [2:0]  indexVec_checkResult_decimal_31 = indexVec_checkResult_decimalProportion_31[5:3];
  wire        indexVec_checkResult_overlap_31 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_31 >= indexVec_checkResult_intLMULInput_31[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_31} >= indexVec_checkResult_intLMULInput_31,
      indexVec_checkResult_allDataPosition_31[32:11]};
  wire        indexVec_checkResult_unChange_31 = slideUp & (indexVec_readIndex_10[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_10 = validVec[10] & ~indexVec_checkResult_unChange_31;
  wire        indexVec_checkResult_1_4_10 = indexVec_checkResult_overlap_31 | ~indexVec_checkResult_1_5_10 | lagerThanVL | indexVec_checkResult_unChange_31;
  wire [33:0] indexVec_checkResult_allDataPosition_32 = {indexVec_readIndex_10, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_32 = indexVec_checkResult_allDataPosition_32[10:0];
  wire [4:0]  indexVec_checkResult_2_1_10 = indexVec_checkResult_dataPosition_32[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_32 = indexVec_checkResult_dataPosition_32[10:7];
  wire        indexVec_checkResult_2_2_10 = indexVec_checkResult_dataGroup_32[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_32 = indexVec_checkResult_dataGroup_32[3:1];
  wire [2:0]  indexVec_checkResult_2_3_10 = indexVec_checkResult_accessRegGrowth_32;
  wire [5:0]  indexVec_checkResult_decimalProportion_32 = {indexVec_checkResult_2_2_10, indexVec_checkResult_2_1_10};
  wire [2:0]  indexVec_checkResult_decimal_32 = indexVec_checkResult_decimalProportion_32[5:3];
  wire        indexVec_checkResult_overlap_32 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_32 >= indexVec_checkResult_intLMULInput_32[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_32} >= indexVec_checkResult_intLMULInput_32,
      indexVec_checkResult_allDataPosition_32[33:11]};
  wire        indexVec_checkResult_unChange_32 = slideUp & (indexVec_readIndex_10[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_10 = validVec[10] & ~indexVec_checkResult_unChange_32;
  wire        indexVec_checkResult_2_4_10 = indexVec_checkResult_overlap_32 | ~indexVec_checkResult_2_5_10 | lagerThanVL | indexVec_checkResult_unChange_32;
  wire [1:0]  indexVec_10_0 = (sew1H[0] ? indexVec_checkResult_0_0_10 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_10 : 2'h0);
  assign indexVec_10_1 = (sew1H[0] ? indexVec_checkResult_0_1_10 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_10 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_10 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_10_0 = indexVec_10_1;
  wire        indexVec_10_2 = sew1H[0] & indexVec_checkResult_0_2_10 | sew1H[1] & indexVec_checkResult_1_2_10 | sew1H[2] & indexVec_checkResult_2_2_10;
  assign indexVec_10_3 = (sew1H[0] ? indexVec_checkResult_0_3_10 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_10 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_10 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_10_0 = indexVec_10_3;
  wire        indexVec_10_4 = sew1H[0] & indexVec_checkResult_0_4_10 | sew1H[1] & indexVec_checkResult_1_4_10 | sew1H[2] & indexVec_checkResult_2_4_10;
  wire        indexVec_10_5 = sew1H[0] & indexVec_checkResult_0_5_10 | sew1H[1] & indexVec_checkResult_1_5_10 | sew1H[2] & indexVec_checkResult_2_5_10;
  wire [31:0] indexVec_readIndex_11 = baseIndex + 32'hB;
  wire [31:0] indexVec_checkResult_allDataPosition_33 = indexVec_readIndex_11;
  wire [10:0] indexVec_checkResult_dataPosition_33 = indexVec_checkResult_allDataPosition_33[10:0];
  wire [1:0]  indexVec_checkResult_0_0_11 = indexVec_checkResult_dataPosition_33[1:0];
  wire [4:0]  indexVec_checkResult_0_1_11 = indexVec_checkResult_dataPosition_33[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_33 = indexVec_checkResult_dataPosition_33[10:7];
  wire        indexVec_checkResult_0_2_11 = indexVec_checkResult_dataGroup_33[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_33 = indexVec_checkResult_dataGroup_33[3:1];
  wire [2:0]  indexVec_checkResult_0_3_11 = indexVec_checkResult_accessRegGrowth_33;
  wire [5:0]  indexVec_checkResult_decimalProportion_33 = {indexVec_checkResult_0_2_11, indexVec_checkResult_0_1_11};
  wire [2:0]  indexVec_checkResult_decimal_33 = indexVec_checkResult_decimalProportion_33[5:3];
  wire        indexVec_checkResult_overlap_33 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_33 >= indexVec_checkResult_intLMULInput_33[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_33} >= indexVec_checkResult_intLMULInput_33,
      indexVec_checkResult_allDataPosition_33[31:11]};
  wire        indexVec_checkResult_unChange_33 = slideUp & (indexVec_readIndex_11[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_11 = validVec[11] & ~indexVec_checkResult_unChange_33;
  wire        indexVec_checkResult_0_4_11 = indexVec_checkResult_overlap_33 | ~indexVec_checkResult_0_5_11 | lagerThanVL | indexVec_checkResult_unChange_33;
  wire [32:0] indexVec_checkResult_allDataPosition_34 = {indexVec_readIndex_11, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_34 = indexVec_checkResult_allDataPosition_34[10:0];
  wire [1:0]  indexVec_checkResult_1_0_11 = {indexVec_checkResult_dataPosition_34[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_11 = indexVec_checkResult_dataPosition_34[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_34 = indexVec_checkResult_dataPosition_34[10:7];
  wire        indexVec_checkResult_1_2_11 = indexVec_checkResult_dataGroup_34[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_34 = indexVec_checkResult_dataGroup_34[3:1];
  wire [2:0]  indexVec_checkResult_1_3_11 = indexVec_checkResult_accessRegGrowth_34;
  wire [5:0]  indexVec_checkResult_decimalProportion_34 = {indexVec_checkResult_1_2_11, indexVec_checkResult_1_1_11};
  wire [2:0]  indexVec_checkResult_decimal_34 = indexVec_checkResult_decimalProportion_34[5:3];
  wire        indexVec_checkResult_overlap_34 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_34 >= indexVec_checkResult_intLMULInput_34[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_34} >= indexVec_checkResult_intLMULInput_34,
      indexVec_checkResult_allDataPosition_34[32:11]};
  wire        indexVec_checkResult_unChange_34 = slideUp & (indexVec_readIndex_11[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_11 = validVec[11] & ~indexVec_checkResult_unChange_34;
  wire        indexVec_checkResult_1_4_11 = indexVec_checkResult_overlap_34 | ~indexVec_checkResult_1_5_11 | lagerThanVL | indexVec_checkResult_unChange_34;
  wire [33:0] indexVec_checkResult_allDataPosition_35 = {indexVec_readIndex_11, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_35 = indexVec_checkResult_allDataPosition_35[10:0];
  wire [4:0]  indexVec_checkResult_2_1_11 = indexVec_checkResult_dataPosition_35[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_35 = indexVec_checkResult_dataPosition_35[10:7];
  wire        indexVec_checkResult_2_2_11 = indexVec_checkResult_dataGroup_35[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_35 = indexVec_checkResult_dataGroup_35[3:1];
  wire [2:0]  indexVec_checkResult_2_3_11 = indexVec_checkResult_accessRegGrowth_35;
  wire [5:0]  indexVec_checkResult_decimalProportion_35 = {indexVec_checkResult_2_2_11, indexVec_checkResult_2_1_11};
  wire [2:0]  indexVec_checkResult_decimal_35 = indexVec_checkResult_decimalProportion_35[5:3];
  wire        indexVec_checkResult_overlap_35 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_35 >= indexVec_checkResult_intLMULInput_35[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_35} >= indexVec_checkResult_intLMULInput_35,
      indexVec_checkResult_allDataPosition_35[33:11]};
  wire        indexVec_checkResult_unChange_35 = slideUp & (indexVec_readIndex_11[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_11 = validVec[11] & ~indexVec_checkResult_unChange_35;
  wire        indexVec_checkResult_2_4_11 = indexVec_checkResult_overlap_35 | ~indexVec_checkResult_2_5_11 | lagerThanVL | indexVec_checkResult_unChange_35;
  wire [1:0]  indexVec_11_0 = (sew1H[0] ? indexVec_checkResult_0_0_11 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_11 : 2'h0);
  assign indexVec_11_1 = (sew1H[0] ? indexVec_checkResult_0_1_11 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_11 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_11 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_11_0 = indexVec_11_1;
  wire        indexVec_11_2 = sew1H[0] & indexVec_checkResult_0_2_11 | sew1H[1] & indexVec_checkResult_1_2_11 | sew1H[2] & indexVec_checkResult_2_2_11;
  assign indexVec_11_3 = (sew1H[0] ? indexVec_checkResult_0_3_11 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_11 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_11 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_11_0 = indexVec_11_3;
  wire        indexVec_11_4 = sew1H[0] & indexVec_checkResult_0_4_11 | sew1H[1] & indexVec_checkResult_1_4_11 | sew1H[2] & indexVec_checkResult_2_4_11;
  wire        indexVec_11_5 = sew1H[0] & indexVec_checkResult_0_5_11 | sew1H[1] & indexVec_checkResult_1_5_11 | sew1H[2] & indexVec_checkResult_2_5_11;
  wire [31:0] indexVec_readIndex_12 = baseIndex + 32'hC;
  wire [31:0] indexVec_checkResult_allDataPosition_36 = indexVec_readIndex_12;
  wire [10:0] indexVec_checkResult_dataPosition_36 = indexVec_checkResult_allDataPosition_36[10:0];
  wire [1:0]  indexVec_checkResult_0_0_12 = indexVec_checkResult_dataPosition_36[1:0];
  wire [4:0]  indexVec_checkResult_0_1_12 = indexVec_checkResult_dataPosition_36[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_36 = indexVec_checkResult_dataPosition_36[10:7];
  wire        indexVec_checkResult_0_2_12 = indexVec_checkResult_dataGroup_36[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_36 = indexVec_checkResult_dataGroup_36[3:1];
  wire [2:0]  indexVec_checkResult_0_3_12 = indexVec_checkResult_accessRegGrowth_36;
  wire [5:0]  indexVec_checkResult_decimalProportion_36 = {indexVec_checkResult_0_2_12, indexVec_checkResult_0_1_12};
  wire [2:0]  indexVec_checkResult_decimal_36 = indexVec_checkResult_decimalProportion_36[5:3];
  wire        indexVec_checkResult_overlap_36 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_36 >= indexVec_checkResult_intLMULInput_36[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_36} >= indexVec_checkResult_intLMULInput_36,
      indexVec_checkResult_allDataPosition_36[31:11]};
  wire        indexVec_checkResult_unChange_36 = slideUp & (indexVec_readIndex_12[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_12 = validVec[12] & ~indexVec_checkResult_unChange_36;
  wire        indexVec_checkResult_0_4_12 = indexVec_checkResult_overlap_36 | ~indexVec_checkResult_0_5_12 | lagerThanVL | indexVec_checkResult_unChange_36;
  wire [32:0] indexVec_checkResult_allDataPosition_37 = {indexVec_readIndex_12, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_37 = indexVec_checkResult_allDataPosition_37[10:0];
  wire [1:0]  indexVec_checkResult_1_0_12 = {indexVec_checkResult_dataPosition_37[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_12 = indexVec_checkResult_dataPosition_37[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_37 = indexVec_checkResult_dataPosition_37[10:7];
  wire        indexVec_checkResult_1_2_12 = indexVec_checkResult_dataGroup_37[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_37 = indexVec_checkResult_dataGroup_37[3:1];
  wire [2:0]  indexVec_checkResult_1_3_12 = indexVec_checkResult_accessRegGrowth_37;
  wire [5:0]  indexVec_checkResult_decimalProportion_37 = {indexVec_checkResult_1_2_12, indexVec_checkResult_1_1_12};
  wire [2:0]  indexVec_checkResult_decimal_37 = indexVec_checkResult_decimalProportion_37[5:3];
  wire        indexVec_checkResult_overlap_37 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_37 >= indexVec_checkResult_intLMULInput_37[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_37} >= indexVec_checkResult_intLMULInput_37,
      indexVec_checkResult_allDataPosition_37[32:11]};
  wire        indexVec_checkResult_unChange_37 = slideUp & (indexVec_readIndex_12[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_12 = validVec[12] & ~indexVec_checkResult_unChange_37;
  wire        indexVec_checkResult_1_4_12 = indexVec_checkResult_overlap_37 | ~indexVec_checkResult_1_5_12 | lagerThanVL | indexVec_checkResult_unChange_37;
  wire [33:0] indexVec_checkResult_allDataPosition_38 = {indexVec_readIndex_12, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_38 = indexVec_checkResult_allDataPosition_38[10:0];
  wire [4:0]  indexVec_checkResult_2_1_12 = indexVec_checkResult_dataPosition_38[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_38 = indexVec_checkResult_dataPosition_38[10:7];
  wire        indexVec_checkResult_2_2_12 = indexVec_checkResult_dataGroup_38[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_38 = indexVec_checkResult_dataGroup_38[3:1];
  wire [2:0]  indexVec_checkResult_2_3_12 = indexVec_checkResult_accessRegGrowth_38;
  wire [5:0]  indexVec_checkResult_decimalProportion_38 = {indexVec_checkResult_2_2_12, indexVec_checkResult_2_1_12};
  wire [2:0]  indexVec_checkResult_decimal_38 = indexVec_checkResult_decimalProportion_38[5:3];
  wire        indexVec_checkResult_overlap_38 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_38 >= indexVec_checkResult_intLMULInput_38[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_38} >= indexVec_checkResult_intLMULInput_38,
      indexVec_checkResult_allDataPosition_38[33:11]};
  wire        indexVec_checkResult_unChange_38 = slideUp & (indexVec_readIndex_12[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_12 = validVec[12] & ~indexVec_checkResult_unChange_38;
  wire        indexVec_checkResult_2_4_12 = indexVec_checkResult_overlap_38 | ~indexVec_checkResult_2_5_12 | lagerThanVL | indexVec_checkResult_unChange_38;
  wire [1:0]  indexVec_12_0 = (sew1H[0] ? indexVec_checkResult_0_0_12 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_12 : 2'h0);
  assign indexVec_12_1 = (sew1H[0] ? indexVec_checkResult_0_1_12 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_12 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_12 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_12_0 = indexVec_12_1;
  wire        indexVec_12_2 = sew1H[0] & indexVec_checkResult_0_2_12 | sew1H[1] & indexVec_checkResult_1_2_12 | sew1H[2] & indexVec_checkResult_2_2_12;
  assign indexVec_12_3 = (sew1H[0] ? indexVec_checkResult_0_3_12 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_12 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_12 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_12_0 = indexVec_12_3;
  wire        indexVec_12_4 = sew1H[0] & indexVec_checkResult_0_4_12 | sew1H[1] & indexVec_checkResult_1_4_12 | sew1H[2] & indexVec_checkResult_2_4_12;
  wire        indexVec_12_5 = sew1H[0] & indexVec_checkResult_0_5_12 | sew1H[1] & indexVec_checkResult_1_5_12 | sew1H[2] & indexVec_checkResult_2_5_12;
  wire [31:0] indexVec_readIndex_13 = baseIndex + 32'hD;
  wire [31:0] indexVec_checkResult_allDataPosition_39 = indexVec_readIndex_13;
  wire [10:0] indexVec_checkResult_dataPosition_39 = indexVec_checkResult_allDataPosition_39[10:0];
  wire [1:0]  indexVec_checkResult_0_0_13 = indexVec_checkResult_dataPosition_39[1:0];
  wire [4:0]  indexVec_checkResult_0_1_13 = indexVec_checkResult_dataPosition_39[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_39 = indexVec_checkResult_dataPosition_39[10:7];
  wire        indexVec_checkResult_0_2_13 = indexVec_checkResult_dataGroup_39[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_39 = indexVec_checkResult_dataGroup_39[3:1];
  wire [2:0]  indexVec_checkResult_0_3_13 = indexVec_checkResult_accessRegGrowth_39;
  wire [5:0]  indexVec_checkResult_decimalProportion_39 = {indexVec_checkResult_0_2_13, indexVec_checkResult_0_1_13};
  wire [2:0]  indexVec_checkResult_decimal_39 = indexVec_checkResult_decimalProportion_39[5:3];
  wire        indexVec_checkResult_overlap_39 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_39 >= indexVec_checkResult_intLMULInput_39[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_39} >= indexVec_checkResult_intLMULInput_39,
      indexVec_checkResult_allDataPosition_39[31:11]};
  wire        indexVec_checkResult_unChange_39 = slideUp & (indexVec_readIndex_13[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_13 = validVec[13] & ~indexVec_checkResult_unChange_39;
  wire        indexVec_checkResult_0_4_13 = indexVec_checkResult_overlap_39 | ~indexVec_checkResult_0_5_13 | lagerThanVL | indexVec_checkResult_unChange_39;
  wire [32:0] indexVec_checkResult_allDataPosition_40 = {indexVec_readIndex_13, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_40 = indexVec_checkResult_allDataPosition_40[10:0];
  wire [1:0]  indexVec_checkResult_1_0_13 = {indexVec_checkResult_dataPosition_40[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_13 = indexVec_checkResult_dataPosition_40[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_40 = indexVec_checkResult_dataPosition_40[10:7];
  wire        indexVec_checkResult_1_2_13 = indexVec_checkResult_dataGroup_40[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_40 = indexVec_checkResult_dataGroup_40[3:1];
  wire [2:0]  indexVec_checkResult_1_3_13 = indexVec_checkResult_accessRegGrowth_40;
  wire [5:0]  indexVec_checkResult_decimalProportion_40 = {indexVec_checkResult_1_2_13, indexVec_checkResult_1_1_13};
  wire [2:0]  indexVec_checkResult_decimal_40 = indexVec_checkResult_decimalProportion_40[5:3];
  wire        indexVec_checkResult_overlap_40 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_40 >= indexVec_checkResult_intLMULInput_40[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_40} >= indexVec_checkResult_intLMULInput_40,
      indexVec_checkResult_allDataPosition_40[32:11]};
  wire        indexVec_checkResult_unChange_40 = slideUp & (indexVec_readIndex_13[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_13 = validVec[13] & ~indexVec_checkResult_unChange_40;
  wire        indexVec_checkResult_1_4_13 = indexVec_checkResult_overlap_40 | ~indexVec_checkResult_1_5_13 | lagerThanVL | indexVec_checkResult_unChange_40;
  wire [33:0] indexVec_checkResult_allDataPosition_41 = {indexVec_readIndex_13, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_41 = indexVec_checkResult_allDataPosition_41[10:0];
  wire [4:0]  indexVec_checkResult_2_1_13 = indexVec_checkResult_dataPosition_41[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_41 = indexVec_checkResult_dataPosition_41[10:7];
  wire        indexVec_checkResult_2_2_13 = indexVec_checkResult_dataGroup_41[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_41 = indexVec_checkResult_dataGroup_41[3:1];
  wire [2:0]  indexVec_checkResult_2_3_13 = indexVec_checkResult_accessRegGrowth_41;
  wire [5:0]  indexVec_checkResult_decimalProportion_41 = {indexVec_checkResult_2_2_13, indexVec_checkResult_2_1_13};
  wire [2:0]  indexVec_checkResult_decimal_41 = indexVec_checkResult_decimalProportion_41[5:3];
  wire        indexVec_checkResult_overlap_41 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_41 >= indexVec_checkResult_intLMULInput_41[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_41} >= indexVec_checkResult_intLMULInput_41,
      indexVec_checkResult_allDataPosition_41[33:11]};
  wire        indexVec_checkResult_unChange_41 = slideUp & (indexVec_readIndex_13[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_13 = validVec[13] & ~indexVec_checkResult_unChange_41;
  wire        indexVec_checkResult_2_4_13 = indexVec_checkResult_overlap_41 | ~indexVec_checkResult_2_5_13 | lagerThanVL | indexVec_checkResult_unChange_41;
  wire [1:0]  indexVec_13_0 = (sew1H[0] ? indexVec_checkResult_0_0_13 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_13 : 2'h0);
  assign indexVec_13_1 = (sew1H[0] ? indexVec_checkResult_0_1_13 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_13 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_13 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_13_0 = indexVec_13_1;
  wire        indexVec_13_2 = sew1H[0] & indexVec_checkResult_0_2_13 | sew1H[1] & indexVec_checkResult_1_2_13 | sew1H[2] & indexVec_checkResult_2_2_13;
  assign indexVec_13_3 = (sew1H[0] ? indexVec_checkResult_0_3_13 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_13 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_13 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_13_0 = indexVec_13_3;
  wire        indexVec_13_4 = sew1H[0] & indexVec_checkResult_0_4_13 | sew1H[1] & indexVec_checkResult_1_4_13 | sew1H[2] & indexVec_checkResult_2_4_13;
  wire        indexVec_13_5 = sew1H[0] & indexVec_checkResult_0_5_13 | sew1H[1] & indexVec_checkResult_1_5_13 | sew1H[2] & indexVec_checkResult_2_5_13;
  wire [31:0] indexVec_readIndex_14 = baseIndex + 32'hE;
  wire [31:0] indexVec_checkResult_allDataPosition_42 = indexVec_readIndex_14;
  wire [10:0] indexVec_checkResult_dataPosition_42 = indexVec_checkResult_allDataPosition_42[10:0];
  wire [1:0]  indexVec_checkResult_0_0_14 = indexVec_checkResult_dataPosition_42[1:0];
  wire [4:0]  indexVec_checkResult_0_1_14 = indexVec_checkResult_dataPosition_42[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_42 = indexVec_checkResult_dataPosition_42[10:7];
  wire        indexVec_checkResult_0_2_14 = indexVec_checkResult_dataGroup_42[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_42 = indexVec_checkResult_dataGroup_42[3:1];
  wire [2:0]  indexVec_checkResult_0_3_14 = indexVec_checkResult_accessRegGrowth_42;
  wire [5:0]  indexVec_checkResult_decimalProportion_42 = {indexVec_checkResult_0_2_14, indexVec_checkResult_0_1_14};
  wire [2:0]  indexVec_checkResult_decimal_42 = indexVec_checkResult_decimalProportion_42[5:3];
  wire        indexVec_checkResult_overlap_42 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_42 >= indexVec_checkResult_intLMULInput_42[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_42} >= indexVec_checkResult_intLMULInput_42,
      indexVec_checkResult_allDataPosition_42[31:11]};
  wire        indexVec_checkResult_unChange_42 = slideUp & (indexVec_readIndex_14[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_14 = validVec[14] & ~indexVec_checkResult_unChange_42;
  wire        indexVec_checkResult_0_4_14 = indexVec_checkResult_overlap_42 | ~indexVec_checkResult_0_5_14 | lagerThanVL | indexVec_checkResult_unChange_42;
  wire [32:0] indexVec_checkResult_allDataPosition_43 = {indexVec_readIndex_14, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_43 = indexVec_checkResult_allDataPosition_43[10:0];
  wire [1:0]  indexVec_checkResult_1_0_14 = {indexVec_checkResult_dataPosition_43[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_14 = indexVec_checkResult_dataPosition_43[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_43 = indexVec_checkResult_dataPosition_43[10:7];
  wire        indexVec_checkResult_1_2_14 = indexVec_checkResult_dataGroup_43[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_43 = indexVec_checkResult_dataGroup_43[3:1];
  wire [2:0]  indexVec_checkResult_1_3_14 = indexVec_checkResult_accessRegGrowth_43;
  wire [5:0]  indexVec_checkResult_decimalProportion_43 = {indexVec_checkResult_1_2_14, indexVec_checkResult_1_1_14};
  wire [2:0]  indexVec_checkResult_decimal_43 = indexVec_checkResult_decimalProportion_43[5:3];
  wire        indexVec_checkResult_overlap_43 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_43 >= indexVec_checkResult_intLMULInput_43[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_43} >= indexVec_checkResult_intLMULInput_43,
      indexVec_checkResult_allDataPosition_43[32:11]};
  wire        indexVec_checkResult_unChange_43 = slideUp & (indexVec_readIndex_14[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_14 = validVec[14] & ~indexVec_checkResult_unChange_43;
  wire        indexVec_checkResult_1_4_14 = indexVec_checkResult_overlap_43 | ~indexVec_checkResult_1_5_14 | lagerThanVL | indexVec_checkResult_unChange_43;
  wire [33:0] indexVec_checkResult_allDataPosition_44 = {indexVec_readIndex_14, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_44 = indexVec_checkResult_allDataPosition_44[10:0];
  wire [4:0]  indexVec_checkResult_2_1_14 = indexVec_checkResult_dataPosition_44[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_44 = indexVec_checkResult_dataPosition_44[10:7];
  wire        indexVec_checkResult_2_2_14 = indexVec_checkResult_dataGroup_44[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_44 = indexVec_checkResult_dataGroup_44[3:1];
  wire [2:0]  indexVec_checkResult_2_3_14 = indexVec_checkResult_accessRegGrowth_44;
  wire [5:0]  indexVec_checkResult_decimalProportion_44 = {indexVec_checkResult_2_2_14, indexVec_checkResult_2_1_14};
  wire [2:0]  indexVec_checkResult_decimal_44 = indexVec_checkResult_decimalProportion_44[5:3];
  wire        indexVec_checkResult_overlap_44 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_44 >= indexVec_checkResult_intLMULInput_44[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_44} >= indexVec_checkResult_intLMULInput_44,
      indexVec_checkResult_allDataPosition_44[33:11]};
  wire        indexVec_checkResult_unChange_44 = slideUp & (indexVec_readIndex_14[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_14 = validVec[14] & ~indexVec_checkResult_unChange_44;
  wire        indexVec_checkResult_2_4_14 = indexVec_checkResult_overlap_44 | ~indexVec_checkResult_2_5_14 | lagerThanVL | indexVec_checkResult_unChange_44;
  wire [1:0]  indexVec_14_0 = (sew1H[0] ? indexVec_checkResult_0_0_14 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_14 : 2'h0);
  assign indexVec_14_1 = (sew1H[0] ? indexVec_checkResult_0_1_14 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_14 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_14 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_14_0 = indexVec_14_1;
  wire        indexVec_14_2 = sew1H[0] & indexVec_checkResult_0_2_14 | sew1H[1] & indexVec_checkResult_1_2_14 | sew1H[2] & indexVec_checkResult_2_2_14;
  assign indexVec_14_3 = (sew1H[0] ? indexVec_checkResult_0_3_14 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_14 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_14 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_14_0 = indexVec_14_3;
  wire        indexVec_14_4 = sew1H[0] & indexVec_checkResult_0_4_14 | sew1H[1] & indexVec_checkResult_1_4_14 | sew1H[2] & indexVec_checkResult_2_4_14;
  wire        indexVec_14_5 = sew1H[0] & indexVec_checkResult_0_5_14 | sew1H[1] & indexVec_checkResult_1_5_14 | sew1H[2] & indexVec_checkResult_2_5_14;
  wire [31:0] indexVec_readIndex_15 = baseIndex + 32'hF;
  wire [31:0] indexVec_checkResult_allDataPosition_45 = indexVec_readIndex_15;
  wire [10:0] indexVec_checkResult_dataPosition_45 = indexVec_checkResult_allDataPosition_45[10:0];
  wire [1:0]  indexVec_checkResult_0_0_15 = indexVec_checkResult_dataPosition_45[1:0];
  wire [4:0]  indexVec_checkResult_0_1_15 = indexVec_checkResult_dataPosition_45[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_45 = indexVec_checkResult_dataPosition_45[10:7];
  wire        indexVec_checkResult_0_2_15 = indexVec_checkResult_dataGroup_45[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_45 = indexVec_checkResult_dataGroup_45[3:1];
  wire [2:0]  indexVec_checkResult_0_3_15 = indexVec_checkResult_accessRegGrowth_45;
  wire [5:0]  indexVec_checkResult_decimalProportion_45 = {indexVec_checkResult_0_2_15, indexVec_checkResult_0_1_15};
  wire [2:0]  indexVec_checkResult_decimal_45 = indexVec_checkResult_decimalProportion_45[5:3];
  wire        indexVec_checkResult_overlap_45 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_45 >= indexVec_checkResult_intLMULInput_45[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_45} >= indexVec_checkResult_intLMULInput_45,
      indexVec_checkResult_allDataPosition_45[31:11]};
  wire        indexVec_checkResult_unChange_45 = slideUp & (indexVec_readIndex_15[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_15 = validVec[15] & ~indexVec_checkResult_unChange_45;
  wire        indexVec_checkResult_0_4_15 = indexVec_checkResult_overlap_45 | ~indexVec_checkResult_0_5_15 | lagerThanVL | indexVec_checkResult_unChange_45;
  wire [32:0] indexVec_checkResult_allDataPosition_46 = {indexVec_readIndex_15, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_46 = indexVec_checkResult_allDataPosition_46[10:0];
  wire [1:0]  indexVec_checkResult_1_0_15 = {indexVec_checkResult_dataPosition_46[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_15 = indexVec_checkResult_dataPosition_46[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_46 = indexVec_checkResult_dataPosition_46[10:7];
  wire        indexVec_checkResult_1_2_15 = indexVec_checkResult_dataGroup_46[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_46 = indexVec_checkResult_dataGroup_46[3:1];
  wire [2:0]  indexVec_checkResult_1_3_15 = indexVec_checkResult_accessRegGrowth_46;
  wire [5:0]  indexVec_checkResult_decimalProportion_46 = {indexVec_checkResult_1_2_15, indexVec_checkResult_1_1_15};
  wire [2:0]  indexVec_checkResult_decimal_46 = indexVec_checkResult_decimalProportion_46[5:3];
  wire        indexVec_checkResult_overlap_46 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_46 >= indexVec_checkResult_intLMULInput_46[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_46} >= indexVec_checkResult_intLMULInput_46,
      indexVec_checkResult_allDataPosition_46[32:11]};
  wire        indexVec_checkResult_unChange_46 = slideUp & (indexVec_readIndex_15[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_15 = validVec[15] & ~indexVec_checkResult_unChange_46;
  wire        indexVec_checkResult_1_4_15 = indexVec_checkResult_overlap_46 | ~indexVec_checkResult_1_5_15 | lagerThanVL | indexVec_checkResult_unChange_46;
  wire [33:0] indexVec_checkResult_allDataPosition_47 = {indexVec_readIndex_15, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_47 = indexVec_checkResult_allDataPosition_47[10:0];
  wire [4:0]  indexVec_checkResult_2_1_15 = indexVec_checkResult_dataPosition_47[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_47 = indexVec_checkResult_dataPosition_47[10:7];
  wire        indexVec_checkResult_2_2_15 = indexVec_checkResult_dataGroup_47[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_47 = indexVec_checkResult_dataGroup_47[3:1];
  wire [2:0]  indexVec_checkResult_2_3_15 = indexVec_checkResult_accessRegGrowth_47;
  wire [5:0]  indexVec_checkResult_decimalProportion_47 = {indexVec_checkResult_2_2_15, indexVec_checkResult_2_1_15};
  wire [2:0]  indexVec_checkResult_decimal_47 = indexVec_checkResult_decimalProportion_47[5:3];
  wire        indexVec_checkResult_overlap_47 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_47 >= indexVec_checkResult_intLMULInput_47[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_47} >= indexVec_checkResult_intLMULInput_47,
      indexVec_checkResult_allDataPosition_47[33:11]};
  wire        indexVec_checkResult_unChange_47 = slideUp & (indexVec_readIndex_15[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_15 = validVec[15] & ~indexVec_checkResult_unChange_47;
  wire        indexVec_checkResult_2_4_15 = indexVec_checkResult_overlap_47 | ~indexVec_checkResult_2_5_15 | lagerThanVL | indexVec_checkResult_unChange_47;
  wire [1:0]  indexVec_15_0 = (sew1H[0] ? indexVec_checkResult_0_0_15 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_15 : 2'h0);
  assign indexVec_15_1 = (sew1H[0] ? indexVec_checkResult_0_1_15 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_15 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_15 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_15_0 = indexVec_15_1;
  wire        indexVec_15_2 = sew1H[0] & indexVec_checkResult_0_2_15 | sew1H[1] & indexVec_checkResult_1_2_15 | sew1H[2] & indexVec_checkResult_2_2_15;
  assign indexVec_15_3 = (sew1H[0] ? indexVec_checkResult_0_3_15 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_15 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_15 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_15_0 = indexVec_15_3;
  wire        indexVec_15_4 = sew1H[0] & indexVec_checkResult_0_4_15 | sew1H[1] & indexVec_checkResult_1_4_15 | sew1H[2] & indexVec_checkResult_2_4_15;
  wire        indexVec_15_5 = sew1H[0] & indexVec_checkResult_0_5_15 | sew1H[1] & indexVec_checkResult_1_5_15 | sew1H[2] & indexVec_checkResult_2_5_15;
  wire [31:0] indexVec_readIndex_16 = baseIndex + 32'h10;
  wire [31:0] indexVec_checkResult_allDataPosition_48 = indexVec_readIndex_16;
  wire [10:0] indexVec_checkResult_dataPosition_48 = indexVec_checkResult_allDataPosition_48[10:0];
  wire [1:0]  indexVec_checkResult_0_0_16 = indexVec_checkResult_dataPosition_48[1:0];
  wire [4:0]  indexVec_checkResult_0_1_16 = indexVec_checkResult_dataPosition_48[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_48 = indexVec_checkResult_dataPosition_48[10:7];
  wire        indexVec_checkResult_0_2_16 = indexVec_checkResult_dataGroup_48[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_48 = indexVec_checkResult_dataGroup_48[3:1];
  wire [2:0]  indexVec_checkResult_0_3_16 = indexVec_checkResult_accessRegGrowth_48;
  wire [5:0]  indexVec_checkResult_decimalProportion_48 = {indexVec_checkResult_0_2_16, indexVec_checkResult_0_1_16};
  wire [2:0]  indexVec_checkResult_decimal_48 = indexVec_checkResult_decimalProportion_48[5:3];
  wire        indexVec_checkResult_overlap_48 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_48 >= indexVec_checkResult_intLMULInput_48[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_48} >= indexVec_checkResult_intLMULInput_48,
      indexVec_checkResult_allDataPosition_48[31:11]};
  wire        indexVec_checkResult_unChange_48 = slideUp & (indexVec_readIndex_16[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_16 = validVec[16] & ~indexVec_checkResult_unChange_48;
  wire        indexVec_checkResult_0_4_16 = indexVec_checkResult_overlap_48 | ~indexVec_checkResult_0_5_16 | lagerThanVL | indexVec_checkResult_unChange_48;
  wire [32:0] indexVec_checkResult_allDataPosition_49 = {indexVec_readIndex_16, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_49 = indexVec_checkResult_allDataPosition_49[10:0];
  wire [1:0]  indexVec_checkResult_1_0_16 = {indexVec_checkResult_dataPosition_49[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_16 = indexVec_checkResult_dataPosition_49[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_49 = indexVec_checkResult_dataPosition_49[10:7];
  wire        indexVec_checkResult_1_2_16 = indexVec_checkResult_dataGroup_49[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_49 = indexVec_checkResult_dataGroup_49[3:1];
  wire [2:0]  indexVec_checkResult_1_3_16 = indexVec_checkResult_accessRegGrowth_49;
  wire [5:0]  indexVec_checkResult_decimalProportion_49 = {indexVec_checkResult_1_2_16, indexVec_checkResult_1_1_16};
  wire [2:0]  indexVec_checkResult_decimal_49 = indexVec_checkResult_decimalProportion_49[5:3];
  wire        indexVec_checkResult_overlap_49 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_49 >= indexVec_checkResult_intLMULInput_49[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_49} >= indexVec_checkResult_intLMULInput_49,
      indexVec_checkResult_allDataPosition_49[32:11]};
  wire        indexVec_checkResult_unChange_49 = slideUp & (indexVec_readIndex_16[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_16 = validVec[16] & ~indexVec_checkResult_unChange_49;
  wire        indexVec_checkResult_1_4_16 = indexVec_checkResult_overlap_49 | ~indexVec_checkResult_1_5_16 | lagerThanVL | indexVec_checkResult_unChange_49;
  wire [33:0] indexVec_checkResult_allDataPosition_50 = {indexVec_readIndex_16, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_50 = indexVec_checkResult_allDataPosition_50[10:0];
  wire [4:0]  indexVec_checkResult_2_1_16 = indexVec_checkResult_dataPosition_50[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_50 = indexVec_checkResult_dataPosition_50[10:7];
  wire        indexVec_checkResult_2_2_16 = indexVec_checkResult_dataGroup_50[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_50 = indexVec_checkResult_dataGroup_50[3:1];
  wire [2:0]  indexVec_checkResult_2_3_16 = indexVec_checkResult_accessRegGrowth_50;
  wire [5:0]  indexVec_checkResult_decimalProportion_50 = {indexVec_checkResult_2_2_16, indexVec_checkResult_2_1_16};
  wire [2:0]  indexVec_checkResult_decimal_50 = indexVec_checkResult_decimalProportion_50[5:3];
  wire        indexVec_checkResult_overlap_50 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_50 >= indexVec_checkResult_intLMULInput_50[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_50} >= indexVec_checkResult_intLMULInput_50,
      indexVec_checkResult_allDataPosition_50[33:11]};
  wire        indexVec_checkResult_unChange_50 = slideUp & (indexVec_readIndex_16[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_16 = validVec[16] & ~indexVec_checkResult_unChange_50;
  wire        indexVec_checkResult_2_4_16 = indexVec_checkResult_overlap_50 | ~indexVec_checkResult_2_5_16 | lagerThanVL | indexVec_checkResult_unChange_50;
  wire [1:0]  indexVec_16_0 = (sew1H[0] ? indexVec_checkResult_0_0_16 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_16 : 2'h0);
  assign indexVec_16_1 = (sew1H[0] ? indexVec_checkResult_0_1_16 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_16 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_16 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_16_0 = indexVec_16_1;
  wire        indexVec_16_2 = sew1H[0] & indexVec_checkResult_0_2_16 | sew1H[1] & indexVec_checkResult_1_2_16 | sew1H[2] & indexVec_checkResult_2_2_16;
  assign indexVec_16_3 = (sew1H[0] ? indexVec_checkResult_0_3_16 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_16 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_16 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_16_0 = indexVec_16_3;
  wire        indexVec_16_4 = sew1H[0] & indexVec_checkResult_0_4_16 | sew1H[1] & indexVec_checkResult_1_4_16 | sew1H[2] & indexVec_checkResult_2_4_16;
  wire        indexVec_16_5 = sew1H[0] & indexVec_checkResult_0_5_16 | sew1H[1] & indexVec_checkResult_1_5_16 | sew1H[2] & indexVec_checkResult_2_5_16;
  wire [31:0] indexVec_readIndex_17 = baseIndex + 32'h11;
  wire [31:0] indexVec_checkResult_allDataPosition_51 = indexVec_readIndex_17;
  wire [10:0] indexVec_checkResult_dataPosition_51 = indexVec_checkResult_allDataPosition_51[10:0];
  wire [1:0]  indexVec_checkResult_0_0_17 = indexVec_checkResult_dataPosition_51[1:0];
  wire [4:0]  indexVec_checkResult_0_1_17 = indexVec_checkResult_dataPosition_51[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_51 = indexVec_checkResult_dataPosition_51[10:7];
  wire        indexVec_checkResult_0_2_17 = indexVec_checkResult_dataGroup_51[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_51 = indexVec_checkResult_dataGroup_51[3:1];
  wire [2:0]  indexVec_checkResult_0_3_17 = indexVec_checkResult_accessRegGrowth_51;
  wire [5:0]  indexVec_checkResult_decimalProportion_51 = {indexVec_checkResult_0_2_17, indexVec_checkResult_0_1_17};
  wire [2:0]  indexVec_checkResult_decimal_51 = indexVec_checkResult_decimalProportion_51[5:3];
  wire        indexVec_checkResult_overlap_51 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_51 >= indexVec_checkResult_intLMULInput_51[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_51} >= indexVec_checkResult_intLMULInput_51,
      indexVec_checkResult_allDataPosition_51[31:11]};
  wire        indexVec_checkResult_unChange_51 = slideUp & (indexVec_readIndex_17[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_17 = validVec[17] & ~indexVec_checkResult_unChange_51;
  wire        indexVec_checkResult_0_4_17 = indexVec_checkResult_overlap_51 | ~indexVec_checkResult_0_5_17 | lagerThanVL | indexVec_checkResult_unChange_51;
  wire [32:0] indexVec_checkResult_allDataPosition_52 = {indexVec_readIndex_17, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_52 = indexVec_checkResult_allDataPosition_52[10:0];
  wire [1:0]  indexVec_checkResult_1_0_17 = {indexVec_checkResult_dataPosition_52[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_17 = indexVec_checkResult_dataPosition_52[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_52 = indexVec_checkResult_dataPosition_52[10:7];
  wire        indexVec_checkResult_1_2_17 = indexVec_checkResult_dataGroup_52[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_52 = indexVec_checkResult_dataGroup_52[3:1];
  wire [2:0]  indexVec_checkResult_1_3_17 = indexVec_checkResult_accessRegGrowth_52;
  wire [5:0]  indexVec_checkResult_decimalProportion_52 = {indexVec_checkResult_1_2_17, indexVec_checkResult_1_1_17};
  wire [2:0]  indexVec_checkResult_decimal_52 = indexVec_checkResult_decimalProportion_52[5:3];
  wire        indexVec_checkResult_overlap_52 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_52 >= indexVec_checkResult_intLMULInput_52[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_52} >= indexVec_checkResult_intLMULInput_52,
      indexVec_checkResult_allDataPosition_52[32:11]};
  wire        indexVec_checkResult_unChange_52 = slideUp & (indexVec_readIndex_17[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_17 = validVec[17] & ~indexVec_checkResult_unChange_52;
  wire        indexVec_checkResult_1_4_17 = indexVec_checkResult_overlap_52 | ~indexVec_checkResult_1_5_17 | lagerThanVL | indexVec_checkResult_unChange_52;
  wire [33:0] indexVec_checkResult_allDataPosition_53 = {indexVec_readIndex_17, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_53 = indexVec_checkResult_allDataPosition_53[10:0];
  wire [4:0]  indexVec_checkResult_2_1_17 = indexVec_checkResult_dataPosition_53[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_53 = indexVec_checkResult_dataPosition_53[10:7];
  wire        indexVec_checkResult_2_2_17 = indexVec_checkResult_dataGroup_53[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_53 = indexVec_checkResult_dataGroup_53[3:1];
  wire [2:0]  indexVec_checkResult_2_3_17 = indexVec_checkResult_accessRegGrowth_53;
  wire [5:0]  indexVec_checkResult_decimalProportion_53 = {indexVec_checkResult_2_2_17, indexVec_checkResult_2_1_17};
  wire [2:0]  indexVec_checkResult_decimal_53 = indexVec_checkResult_decimalProportion_53[5:3];
  wire        indexVec_checkResult_overlap_53 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_53 >= indexVec_checkResult_intLMULInput_53[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_53} >= indexVec_checkResult_intLMULInput_53,
      indexVec_checkResult_allDataPosition_53[33:11]};
  wire        indexVec_checkResult_unChange_53 = slideUp & (indexVec_readIndex_17[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_17 = validVec[17] & ~indexVec_checkResult_unChange_53;
  wire        indexVec_checkResult_2_4_17 = indexVec_checkResult_overlap_53 | ~indexVec_checkResult_2_5_17 | lagerThanVL | indexVec_checkResult_unChange_53;
  wire [1:0]  indexVec_17_0 = (sew1H[0] ? indexVec_checkResult_0_0_17 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_17 : 2'h0);
  assign indexVec_17_1 = (sew1H[0] ? indexVec_checkResult_0_1_17 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_17 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_17 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_17_0 = indexVec_17_1;
  wire        indexVec_17_2 = sew1H[0] & indexVec_checkResult_0_2_17 | sew1H[1] & indexVec_checkResult_1_2_17 | sew1H[2] & indexVec_checkResult_2_2_17;
  assign indexVec_17_3 = (sew1H[0] ? indexVec_checkResult_0_3_17 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_17 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_17 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_17_0 = indexVec_17_3;
  wire        indexVec_17_4 = sew1H[0] & indexVec_checkResult_0_4_17 | sew1H[1] & indexVec_checkResult_1_4_17 | sew1H[2] & indexVec_checkResult_2_4_17;
  wire        indexVec_17_5 = sew1H[0] & indexVec_checkResult_0_5_17 | sew1H[1] & indexVec_checkResult_1_5_17 | sew1H[2] & indexVec_checkResult_2_5_17;
  wire [31:0] indexVec_readIndex_18 = baseIndex + 32'h12;
  wire [31:0] indexVec_checkResult_allDataPosition_54 = indexVec_readIndex_18;
  wire [10:0] indexVec_checkResult_dataPosition_54 = indexVec_checkResult_allDataPosition_54[10:0];
  wire [1:0]  indexVec_checkResult_0_0_18 = indexVec_checkResult_dataPosition_54[1:0];
  wire [4:0]  indexVec_checkResult_0_1_18 = indexVec_checkResult_dataPosition_54[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_54 = indexVec_checkResult_dataPosition_54[10:7];
  wire        indexVec_checkResult_0_2_18 = indexVec_checkResult_dataGroup_54[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_54 = indexVec_checkResult_dataGroup_54[3:1];
  wire [2:0]  indexVec_checkResult_0_3_18 = indexVec_checkResult_accessRegGrowth_54;
  wire [5:0]  indexVec_checkResult_decimalProportion_54 = {indexVec_checkResult_0_2_18, indexVec_checkResult_0_1_18};
  wire [2:0]  indexVec_checkResult_decimal_54 = indexVec_checkResult_decimalProportion_54[5:3];
  wire        indexVec_checkResult_overlap_54 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_54 >= indexVec_checkResult_intLMULInput_54[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_54} >= indexVec_checkResult_intLMULInput_54,
      indexVec_checkResult_allDataPosition_54[31:11]};
  wire        indexVec_checkResult_unChange_54 = slideUp & (indexVec_readIndex_18[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_18 = validVec[18] & ~indexVec_checkResult_unChange_54;
  wire        indexVec_checkResult_0_4_18 = indexVec_checkResult_overlap_54 | ~indexVec_checkResult_0_5_18 | lagerThanVL | indexVec_checkResult_unChange_54;
  wire [32:0] indexVec_checkResult_allDataPosition_55 = {indexVec_readIndex_18, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_55 = indexVec_checkResult_allDataPosition_55[10:0];
  wire [1:0]  indexVec_checkResult_1_0_18 = {indexVec_checkResult_dataPosition_55[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_18 = indexVec_checkResult_dataPosition_55[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_55 = indexVec_checkResult_dataPosition_55[10:7];
  wire        indexVec_checkResult_1_2_18 = indexVec_checkResult_dataGroup_55[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_55 = indexVec_checkResult_dataGroup_55[3:1];
  wire [2:0]  indexVec_checkResult_1_3_18 = indexVec_checkResult_accessRegGrowth_55;
  wire [5:0]  indexVec_checkResult_decimalProportion_55 = {indexVec_checkResult_1_2_18, indexVec_checkResult_1_1_18};
  wire [2:0]  indexVec_checkResult_decimal_55 = indexVec_checkResult_decimalProportion_55[5:3];
  wire        indexVec_checkResult_overlap_55 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_55 >= indexVec_checkResult_intLMULInput_55[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_55} >= indexVec_checkResult_intLMULInput_55,
      indexVec_checkResult_allDataPosition_55[32:11]};
  wire        indexVec_checkResult_unChange_55 = slideUp & (indexVec_readIndex_18[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_18 = validVec[18] & ~indexVec_checkResult_unChange_55;
  wire        indexVec_checkResult_1_4_18 = indexVec_checkResult_overlap_55 | ~indexVec_checkResult_1_5_18 | lagerThanVL | indexVec_checkResult_unChange_55;
  wire [33:0] indexVec_checkResult_allDataPosition_56 = {indexVec_readIndex_18, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_56 = indexVec_checkResult_allDataPosition_56[10:0];
  wire [4:0]  indexVec_checkResult_2_1_18 = indexVec_checkResult_dataPosition_56[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_56 = indexVec_checkResult_dataPosition_56[10:7];
  wire        indexVec_checkResult_2_2_18 = indexVec_checkResult_dataGroup_56[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_56 = indexVec_checkResult_dataGroup_56[3:1];
  wire [2:0]  indexVec_checkResult_2_3_18 = indexVec_checkResult_accessRegGrowth_56;
  wire [5:0]  indexVec_checkResult_decimalProportion_56 = {indexVec_checkResult_2_2_18, indexVec_checkResult_2_1_18};
  wire [2:0]  indexVec_checkResult_decimal_56 = indexVec_checkResult_decimalProportion_56[5:3];
  wire        indexVec_checkResult_overlap_56 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_56 >= indexVec_checkResult_intLMULInput_56[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_56} >= indexVec_checkResult_intLMULInput_56,
      indexVec_checkResult_allDataPosition_56[33:11]};
  wire        indexVec_checkResult_unChange_56 = slideUp & (indexVec_readIndex_18[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_18 = validVec[18] & ~indexVec_checkResult_unChange_56;
  wire        indexVec_checkResult_2_4_18 = indexVec_checkResult_overlap_56 | ~indexVec_checkResult_2_5_18 | lagerThanVL | indexVec_checkResult_unChange_56;
  wire [1:0]  indexVec_18_0 = (sew1H[0] ? indexVec_checkResult_0_0_18 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_18 : 2'h0);
  assign indexVec_18_1 = (sew1H[0] ? indexVec_checkResult_0_1_18 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_18 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_18 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_18_0 = indexVec_18_1;
  wire        indexVec_18_2 = sew1H[0] & indexVec_checkResult_0_2_18 | sew1H[1] & indexVec_checkResult_1_2_18 | sew1H[2] & indexVec_checkResult_2_2_18;
  assign indexVec_18_3 = (sew1H[0] ? indexVec_checkResult_0_3_18 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_18 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_18 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_18_0 = indexVec_18_3;
  wire        indexVec_18_4 = sew1H[0] & indexVec_checkResult_0_4_18 | sew1H[1] & indexVec_checkResult_1_4_18 | sew1H[2] & indexVec_checkResult_2_4_18;
  wire        indexVec_18_5 = sew1H[0] & indexVec_checkResult_0_5_18 | sew1H[1] & indexVec_checkResult_1_5_18 | sew1H[2] & indexVec_checkResult_2_5_18;
  wire [31:0] indexVec_readIndex_19 = baseIndex + 32'h13;
  wire [31:0] indexVec_checkResult_allDataPosition_57 = indexVec_readIndex_19;
  wire [10:0] indexVec_checkResult_dataPosition_57 = indexVec_checkResult_allDataPosition_57[10:0];
  wire [1:0]  indexVec_checkResult_0_0_19 = indexVec_checkResult_dataPosition_57[1:0];
  wire [4:0]  indexVec_checkResult_0_1_19 = indexVec_checkResult_dataPosition_57[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_57 = indexVec_checkResult_dataPosition_57[10:7];
  wire        indexVec_checkResult_0_2_19 = indexVec_checkResult_dataGroup_57[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_57 = indexVec_checkResult_dataGroup_57[3:1];
  wire [2:0]  indexVec_checkResult_0_3_19 = indexVec_checkResult_accessRegGrowth_57;
  wire [5:0]  indexVec_checkResult_decimalProportion_57 = {indexVec_checkResult_0_2_19, indexVec_checkResult_0_1_19};
  wire [2:0]  indexVec_checkResult_decimal_57 = indexVec_checkResult_decimalProportion_57[5:3];
  wire        indexVec_checkResult_overlap_57 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_57 >= indexVec_checkResult_intLMULInput_57[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_57} >= indexVec_checkResult_intLMULInput_57,
      indexVec_checkResult_allDataPosition_57[31:11]};
  wire        indexVec_checkResult_unChange_57 = slideUp & (indexVec_readIndex_19[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_19 = validVec[19] & ~indexVec_checkResult_unChange_57;
  wire        indexVec_checkResult_0_4_19 = indexVec_checkResult_overlap_57 | ~indexVec_checkResult_0_5_19 | lagerThanVL | indexVec_checkResult_unChange_57;
  wire [32:0] indexVec_checkResult_allDataPosition_58 = {indexVec_readIndex_19, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_58 = indexVec_checkResult_allDataPosition_58[10:0];
  wire [1:0]  indexVec_checkResult_1_0_19 = {indexVec_checkResult_dataPosition_58[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_19 = indexVec_checkResult_dataPosition_58[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_58 = indexVec_checkResult_dataPosition_58[10:7];
  wire        indexVec_checkResult_1_2_19 = indexVec_checkResult_dataGroup_58[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_58 = indexVec_checkResult_dataGroup_58[3:1];
  wire [2:0]  indexVec_checkResult_1_3_19 = indexVec_checkResult_accessRegGrowth_58;
  wire [5:0]  indexVec_checkResult_decimalProportion_58 = {indexVec_checkResult_1_2_19, indexVec_checkResult_1_1_19};
  wire [2:0]  indexVec_checkResult_decimal_58 = indexVec_checkResult_decimalProportion_58[5:3];
  wire        indexVec_checkResult_overlap_58 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_58 >= indexVec_checkResult_intLMULInput_58[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_58} >= indexVec_checkResult_intLMULInput_58,
      indexVec_checkResult_allDataPosition_58[32:11]};
  wire        indexVec_checkResult_unChange_58 = slideUp & (indexVec_readIndex_19[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_19 = validVec[19] & ~indexVec_checkResult_unChange_58;
  wire        indexVec_checkResult_1_4_19 = indexVec_checkResult_overlap_58 | ~indexVec_checkResult_1_5_19 | lagerThanVL | indexVec_checkResult_unChange_58;
  wire [33:0] indexVec_checkResult_allDataPosition_59 = {indexVec_readIndex_19, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_59 = indexVec_checkResult_allDataPosition_59[10:0];
  wire [4:0]  indexVec_checkResult_2_1_19 = indexVec_checkResult_dataPosition_59[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_59 = indexVec_checkResult_dataPosition_59[10:7];
  wire        indexVec_checkResult_2_2_19 = indexVec_checkResult_dataGroup_59[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_59 = indexVec_checkResult_dataGroup_59[3:1];
  wire [2:0]  indexVec_checkResult_2_3_19 = indexVec_checkResult_accessRegGrowth_59;
  wire [5:0]  indexVec_checkResult_decimalProportion_59 = {indexVec_checkResult_2_2_19, indexVec_checkResult_2_1_19};
  wire [2:0]  indexVec_checkResult_decimal_59 = indexVec_checkResult_decimalProportion_59[5:3];
  wire        indexVec_checkResult_overlap_59 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_59 >= indexVec_checkResult_intLMULInput_59[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_59} >= indexVec_checkResult_intLMULInput_59,
      indexVec_checkResult_allDataPosition_59[33:11]};
  wire        indexVec_checkResult_unChange_59 = slideUp & (indexVec_readIndex_19[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_19 = validVec[19] & ~indexVec_checkResult_unChange_59;
  wire        indexVec_checkResult_2_4_19 = indexVec_checkResult_overlap_59 | ~indexVec_checkResult_2_5_19 | lagerThanVL | indexVec_checkResult_unChange_59;
  wire [1:0]  indexVec_19_0 = (sew1H[0] ? indexVec_checkResult_0_0_19 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_19 : 2'h0);
  assign indexVec_19_1 = (sew1H[0] ? indexVec_checkResult_0_1_19 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_19 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_19 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_19_0 = indexVec_19_1;
  wire        indexVec_19_2 = sew1H[0] & indexVec_checkResult_0_2_19 | sew1H[1] & indexVec_checkResult_1_2_19 | sew1H[2] & indexVec_checkResult_2_2_19;
  assign indexVec_19_3 = (sew1H[0] ? indexVec_checkResult_0_3_19 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_19 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_19 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_19_0 = indexVec_19_3;
  wire        indexVec_19_4 = sew1H[0] & indexVec_checkResult_0_4_19 | sew1H[1] & indexVec_checkResult_1_4_19 | sew1H[2] & indexVec_checkResult_2_4_19;
  wire        indexVec_19_5 = sew1H[0] & indexVec_checkResult_0_5_19 | sew1H[1] & indexVec_checkResult_1_5_19 | sew1H[2] & indexVec_checkResult_2_5_19;
  wire [31:0] indexVec_readIndex_20 = baseIndex + 32'h14;
  wire [31:0] indexVec_checkResult_allDataPosition_60 = indexVec_readIndex_20;
  wire [10:0] indexVec_checkResult_dataPosition_60 = indexVec_checkResult_allDataPosition_60[10:0];
  wire [1:0]  indexVec_checkResult_0_0_20 = indexVec_checkResult_dataPosition_60[1:0];
  wire [4:0]  indexVec_checkResult_0_1_20 = indexVec_checkResult_dataPosition_60[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_60 = indexVec_checkResult_dataPosition_60[10:7];
  wire        indexVec_checkResult_0_2_20 = indexVec_checkResult_dataGroup_60[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_60 = indexVec_checkResult_dataGroup_60[3:1];
  wire [2:0]  indexVec_checkResult_0_3_20 = indexVec_checkResult_accessRegGrowth_60;
  wire [5:0]  indexVec_checkResult_decimalProportion_60 = {indexVec_checkResult_0_2_20, indexVec_checkResult_0_1_20};
  wire [2:0]  indexVec_checkResult_decimal_60 = indexVec_checkResult_decimalProportion_60[5:3];
  wire        indexVec_checkResult_overlap_60 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_60 >= indexVec_checkResult_intLMULInput_60[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_60} >= indexVec_checkResult_intLMULInput_60,
      indexVec_checkResult_allDataPosition_60[31:11]};
  wire        indexVec_checkResult_unChange_60 = slideUp & (indexVec_readIndex_20[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_20 = validVec[20] & ~indexVec_checkResult_unChange_60;
  wire        indexVec_checkResult_0_4_20 = indexVec_checkResult_overlap_60 | ~indexVec_checkResult_0_5_20 | lagerThanVL | indexVec_checkResult_unChange_60;
  wire [32:0] indexVec_checkResult_allDataPosition_61 = {indexVec_readIndex_20, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_61 = indexVec_checkResult_allDataPosition_61[10:0];
  wire [1:0]  indexVec_checkResult_1_0_20 = {indexVec_checkResult_dataPosition_61[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_20 = indexVec_checkResult_dataPosition_61[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_61 = indexVec_checkResult_dataPosition_61[10:7];
  wire        indexVec_checkResult_1_2_20 = indexVec_checkResult_dataGroup_61[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_61 = indexVec_checkResult_dataGroup_61[3:1];
  wire [2:0]  indexVec_checkResult_1_3_20 = indexVec_checkResult_accessRegGrowth_61;
  wire [5:0]  indexVec_checkResult_decimalProportion_61 = {indexVec_checkResult_1_2_20, indexVec_checkResult_1_1_20};
  wire [2:0]  indexVec_checkResult_decimal_61 = indexVec_checkResult_decimalProportion_61[5:3];
  wire        indexVec_checkResult_overlap_61 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_61 >= indexVec_checkResult_intLMULInput_61[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_61} >= indexVec_checkResult_intLMULInput_61,
      indexVec_checkResult_allDataPosition_61[32:11]};
  wire        indexVec_checkResult_unChange_61 = slideUp & (indexVec_readIndex_20[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_20 = validVec[20] & ~indexVec_checkResult_unChange_61;
  wire        indexVec_checkResult_1_4_20 = indexVec_checkResult_overlap_61 | ~indexVec_checkResult_1_5_20 | lagerThanVL | indexVec_checkResult_unChange_61;
  wire [33:0] indexVec_checkResult_allDataPosition_62 = {indexVec_readIndex_20, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_62 = indexVec_checkResult_allDataPosition_62[10:0];
  wire [4:0]  indexVec_checkResult_2_1_20 = indexVec_checkResult_dataPosition_62[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_62 = indexVec_checkResult_dataPosition_62[10:7];
  wire        indexVec_checkResult_2_2_20 = indexVec_checkResult_dataGroup_62[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_62 = indexVec_checkResult_dataGroup_62[3:1];
  wire [2:0]  indexVec_checkResult_2_3_20 = indexVec_checkResult_accessRegGrowth_62;
  wire [5:0]  indexVec_checkResult_decimalProportion_62 = {indexVec_checkResult_2_2_20, indexVec_checkResult_2_1_20};
  wire [2:0]  indexVec_checkResult_decimal_62 = indexVec_checkResult_decimalProportion_62[5:3];
  wire        indexVec_checkResult_overlap_62 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_62 >= indexVec_checkResult_intLMULInput_62[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_62} >= indexVec_checkResult_intLMULInput_62,
      indexVec_checkResult_allDataPosition_62[33:11]};
  wire        indexVec_checkResult_unChange_62 = slideUp & (indexVec_readIndex_20[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_20 = validVec[20] & ~indexVec_checkResult_unChange_62;
  wire        indexVec_checkResult_2_4_20 = indexVec_checkResult_overlap_62 | ~indexVec_checkResult_2_5_20 | lagerThanVL | indexVec_checkResult_unChange_62;
  wire [1:0]  indexVec_20_0 = (sew1H[0] ? indexVec_checkResult_0_0_20 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_20 : 2'h0);
  assign indexVec_20_1 = (sew1H[0] ? indexVec_checkResult_0_1_20 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_20 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_20 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_20_0 = indexVec_20_1;
  wire        indexVec_20_2 = sew1H[0] & indexVec_checkResult_0_2_20 | sew1H[1] & indexVec_checkResult_1_2_20 | sew1H[2] & indexVec_checkResult_2_2_20;
  assign indexVec_20_3 = (sew1H[0] ? indexVec_checkResult_0_3_20 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_20 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_20 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_20_0 = indexVec_20_3;
  wire        indexVec_20_4 = sew1H[0] & indexVec_checkResult_0_4_20 | sew1H[1] & indexVec_checkResult_1_4_20 | sew1H[2] & indexVec_checkResult_2_4_20;
  wire        indexVec_20_5 = sew1H[0] & indexVec_checkResult_0_5_20 | sew1H[1] & indexVec_checkResult_1_5_20 | sew1H[2] & indexVec_checkResult_2_5_20;
  wire [31:0] indexVec_readIndex_21 = baseIndex + 32'h15;
  wire [31:0] indexVec_checkResult_allDataPosition_63 = indexVec_readIndex_21;
  wire [10:0] indexVec_checkResult_dataPosition_63 = indexVec_checkResult_allDataPosition_63[10:0];
  wire [1:0]  indexVec_checkResult_0_0_21 = indexVec_checkResult_dataPosition_63[1:0];
  wire [4:0]  indexVec_checkResult_0_1_21 = indexVec_checkResult_dataPosition_63[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_63 = indexVec_checkResult_dataPosition_63[10:7];
  wire        indexVec_checkResult_0_2_21 = indexVec_checkResult_dataGroup_63[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_63 = indexVec_checkResult_dataGroup_63[3:1];
  wire [2:0]  indexVec_checkResult_0_3_21 = indexVec_checkResult_accessRegGrowth_63;
  wire [5:0]  indexVec_checkResult_decimalProportion_63 = {indexVec_checkResult_0_2_21, indexVec_checkResult_0_1_21};
  wire [2:0]  indexVec_checkResult_decimal_63 = indexVec_checkResult_decimalProportion_63[5:3];
  wire        indexVec_checkResult_overlap_63 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_63 >= indexVec_checkResult_intLMULInput_63[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_63} >= indexVec_checkResult_intLMULInput_63,
      indexVec_checkResult_allDataPosition_63[31:11]};
  wire        indexVec_checkResult_unChange_63 = slideUp & (indexVec_readIndex_21[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_21 = validVec[21] & ~indexVec_checkResult_unChange_63;
  wire        indexVec_checkResult_0_4_21 = indexVec_checkResult_overlap_63 | ~indexVec_checkResult_0_5_21 | lagerThanVL | indexVec_checkResult_unChange_63;
  wire [32:0] indexVec_checkResult_allDataPosition_64 = {indexVec_readIndex_21, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_64 = indexVec_checkResult_allDataPosition_64[10:0];
  wire [1:0]  indexVec_checkResult_1_0_21 = {indexVec_checkResult_dataPosition_64[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_21 = indexVec_checkResult_dataPosition_64[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_64 = indexVec_checkResult_dataPosition_64[10:7];
  wire        indexVec_checkResult_1_2_21 = indexVec_checkResult_dataGroup_64[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_64 = indexVec_checkResult_dataGroup_64[3:1];
  wire [2:0]  indexVec_checkResult_1_3_21 = indexVec_checkResult_accessRegGrowth_64;
  wire [5:0]  indexVec_checkResult_decimalProportion_64 = {indexVec_checkResult_1_2_21, indexVec_checkResult_1_1_21};
  wire [2:0]  indexVec_checkResult_decimal_64 = indexVec_checkResult_decimalProportion_64[5:3];
  wire        indexVec_checkResult_overlap_64 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_64 >= indexVec_checkResult_intLMULInput_64[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_64} >= indexVec_checkResult_intLMULInput_64,
      indexVec_checkResult_allDataPosition_64[32:11]};
  wire        indexVec_checkResult_unChange_64 = slideUp & (indexVec_readIndex_21[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_21 = validVec[21] & ~indexVec_checkResult_unChange_64;
  wire        indexVec_checkResult_1_4_21 = indexVec_checkResult_overlap_64 | ~indexVec_checkResult_1_5_21 | lagerThanVL | indexVec_checkResult_unChange_64;
  wire [33:0] indexVec_checkResult_allDataPosition_65 = {indexVec_readIndex_21, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_65 = indexVec_checkResult_allDataPosition_65[10:0];
  wire [4:0]  indexVec_checkResult_2_1_21 = indexVec_checkResult_dataPosition_65[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_65 = indexVec_checkResult_dataPosition_65[10:7];
  wire        indexVec_checkResult_2_2_21 = indexVec_checkResult_dataGroup_65[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_65 = indexVec_checkResult_dataGroup_65[3:1];
  wire [2:0]  indexVec_checkResult_2_3_21 = indexVec_checkResult_accessRegGrowth_65;
  wire [5:0]  indexVec_checkResult_decimalProportion_65 = {indexVec_checkResult_2_2_21, indexVec_checkResult_2_1_21};
  wire [2:0]  indexVec_checkResult_decimal_65 = indexVec_checkResult_decimalProportion_65[5:3];
  wire        indexVec_checkResult_overlap_65 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_65 >= indexVec_checkResult_intLMULInput_65[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_65} >= indexVec_checkResult_intLMULInput_65,
      indexVec_checkResult_allDataPosition_65[33:11]};
  wire        indexVec_checkResult_unChange_65 = slideUp & (indexVec_readIndex_21[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_21 = validVec[21] & ~indexVec_checkResult_unChange_65;
  wire        indexVec_checkResult_2_4_21 = indexVec_checkResult_overlap_65 | ~indexVec_checkResult_2_5_21 | lagerThanVL | indexVec_checkResult_unChange_65;
  wire [1:0]  indexVec_21_0 = (sew1H[0] ? indexVec_checkResult_0_0_21 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_21 : 2'h0);
  assign indexVec_21_1 = (sew1H[0] ? indexVec_checkResult_0_1_21 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_21 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_21 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_21_0 = indexVec_21_1;
  wire        indexVec_21_2 = sew1H[0] & indexVec_checkResult_0_2_21 | sew1H[1] & indexVec_checkResult_1_2_21 | sew1H[2] & indexVec_checkResult_2_2_21;
  assign indexVec_21_3 = (sew1H[0] ? indexVec_checkResult_0_3_21 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_21 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_21 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_21_0 = indexVec_21_3;
  wire        indexVec_21_4 = sew1H[0] & indexVec_checkResult_0_4_21 | sew1H[1] & indexVec_checkResult_1_4_21 | sew1H[2] & indexVec_checkResult_2_4_21;
  wire        indexVec_21_5 = sew1H[0] & indexVec_checkResult_0_5_21 | sew1H[1] & indexVec_checkResult_1_5_21 | sew1H[2] & indexVec_checkResult_2_5_21;
  wire [31:0] indexVec_readIndex_22 = baseIndex + 32'h16;
  wire [31:0] indexVec_checkResult_allDataPosition_66 = indexVec_readIndex_22;
  wire [10:0] indexVec_checkResult_dataPosition_66 = indexVec_checkResult_allDataPosition_66[10:0];
  wire [1:0]  indexVec_checkResult_0_0_22 = indexVec_checkResult_dataPosition_66[1:0];
  wire [4:0]  indexVec_checkResult_0_1_22 = indexVec_checkResult_dataPosition_66[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_66 = indexVec_checkResult_dataPosition_66[10:7];
  wire        indexVec_checkResult_0_2_22 = indexVec_checkResult_dataGroup_66[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_66 = indexVec_checkResult_dataGroup_66[3:1];
  wire [2:0]  indexVec_checkResult_0_3_22 = indexVec_checkResult_accessRegGrowth_66;
  wire [5:0]  indexVec_checkResult_decimalProportion_66 = {indexVec_checkResult_0_2_22, indexVec_checkResult_0_1_22};
  wire [2:0]  indexVec_checkResult_decimal_66 = indexVec_checkResult_decimalProportion_66[5:3];
  wire        indexVec_checkResult_overlap_66 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_66 >= indexVec_checkResult_intLMULInput_66[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_66} >= indexVec_checkResult_intLMULInput_66,
      indexVec_checkResult_allDataPosition_66[31:11]};
  wire        indexVec_checkResult_unChange_66 = slideUp & (indexVec_readIndex_22[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_22 = validVec[22] & ~indexVec_checkResult_unChange_66;
  wire        indexVec_checkResult_0_4_22 = indexVec_checkResult_overlap_66 | ~indexVec_checkResult_0_5_22 | lagerThanVL | indexVec_checkResult_unChange_66;
  wire [32:0] indexVec_checkResult_allDataPosition_67 = {indexVec_readIndex_22, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_67 = indexVec_checkResult_allDataPosition_67[10:0];
  wire [1:0]  indexVec_checkResult_1_0_22 = {indexVec_checkResult_dataPosition_67[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_22 = indexVec_checkResult_dataPosition_67[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_67 = indexVec_checkResult_dataPosition_67[10:7];
  wire        indexVec_checkResult_1_2_22 = indexVec_checkResult_dataGroup_67[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_67 = indexVec_checkResult_dataGroup_67[3:1];
  wire [2:0]  indexVec_checkResult_1_3_22 = indexVec_checkResult_accessRegGrowth_67;
  wire [5:0]  indexVec_checkResult_decimalProportion_67 = {indexVec_checkResult_1_2_22, indexVec_checkResult_1_1_22};
  wire [2:0]  indexVec_checkResult_decimal_67 = indexVec_checkResult_decimalProportion_67[5:3];
  wire        indexVec_checkResult_overlap_67 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_67 >= indexVec_checkResult_intLMULInput_67[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_67} >= indexVec_checkResult_intLMULInput_67,
      indexVec_checkResult_allDataPosition_67[32:11]};
  wire        indexVec_checkResult_unChange_67 = slideUp & (indexVec_readIndex_22[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_22 = validVec[22] & ~indexVec_checkResult_unChange_67;
  wire        indexVec_checkResult_1_4_22 = indexVec_checkResult_overlap_67 | ~indexVec_checkResult_1_5_22 | lagerThanVL | indexVec_checkResult_unChange_67;
  wire [33:0] indexVec_checkResult_allDataPosition_68 = {indexVec_readIndex_22, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_68 = indexVec_checkResult_allDataPosition_68[10:0];
  wire [4:0]  indexVec_checkResult_2_1_22 = indexVec_checkResult_dataPosition_68[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_68 = indexVec_checkResult_dataPosition_68[10:7];
  wire        indexVec_checkResult_2_2_22 = indexVec_checkResult_dataGroup_68[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_68 = indexVec_checkResult_dataGroup_68[3:1];
  wire [2:0]  indexVec_checkResult_2_3_22 = indexVec_checkResult_accessRegGrowth_68;
  wire [5:0]  indexVec_checkResult_decimalProportion_68 = {indexVec_checkResult_2_2_22, indexVec_checkResult_2_1_22};
  wire [2:0]  indexVec_checkResult_decimal_68 = indexVec_checkResult_decimalProportion_68[5:3];
  wire        indexVec_checkResult_overlap_68 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_68 >= indexVec_checkResult_intLMULInput_68[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_68} >= indexVec_checkResult_intLMULInput_68,
      indexVec_checkResult_allDataPosition_68[33:11]};
  wire        indexVec_checkResult_unChange_68 = slideUp & (indexVec_readIndex_22[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_22 = validVec[22] & ~indexVec_checkResult_unChange_68;
  wire        indexVec_checkResult_2_4_22 = indexVec_checkResult_overlap_68 | ~indexVec_checkResult_2_5_22 | lagerThanVL | indexVec_checkResult_unChange_68;
  wire [1:0]  indexVec_22_0 = (sew1H[0] ? indexVec_checkResult_0_0_22 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_22 : 2'h0);
  assign indexVec_22_1 = (sew1H[0] ? indexVec_checkResult_0_1_22 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_22 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_22 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_22_0 = indexVec_22_1;
  wire        indexVec_22_2 = sew1H[0] & indexVec_checkResult_0_2_22 | sew1H[1] & indexVec_checkResult_1_2_22 | sew1H[2] & indexVec_checkResult_2_2_22;
  assign indexVec_22_3 = (sew1H[0] ? indexVec_checkResult_0_3_22 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_22 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_22 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_22_0 = indexVec_22_3;
  wire        indexVec_22_4 = sew1H[0] & indexVec_checkResult_0_4_22 | sew1H[1] & indexVec_checkResult_1_4_22 | sew1H[2] & indexVec_checkResult_2_4_22;
  wire        indexVec_22_5 = sew1H[0] & indexVec_checkResult_0_5_22 | sew1H[1] & indexVec_checkResult_1_5_22 | sew1H[2] & indexVec_checkResult_2_5_22;
  wire [31:0] indexVec_readIndex_23 = baseIndex + 32'h17;
  wire [31:0] indexVec_checkResult_allDataPosition_69 = indexVec_readIndex_23;
  wire [10:0] indexVec_checkResult_dataPosition_69 = indexVec_checkResult_allDataPosition_69[10:0];
  wire [1:0]  indexVec_checkResult_0_0_23 = indexVec_checkResult_dataPosition_69[1:0];
  wire [4:0]  indexVec_checkResult_0_1_23 = indexVec_checkResult_dataPosition_69[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_69 = indexVec_checkResult_dataPosition_69[10:7];
  wire        indexVec_checkResult_0_2_23 = indexVec_checkResult_dataGroup_69[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_69 = indexVec_checkResult_dataGroup_69[3:1];
  wire [2:0]  indexVec_checkResult_0_3_23 = indexVec_checkResult_accessRegGrowth_69;
  wire [5:0]  indexVec_checkResult_decimalProportion_69 = {indexVec_checkResult_0_2_23, indexVec_checkResult_0_1_23};
  wire [2:0]  indexVec_checkResult_decimal_69 = indexVec_checkResult_decimalProportion_69[5:3];
  wire        indexVec_checkResult_overlap_69 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_69 >= indexVec_checkResult_intLMULInput_69[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_69} >= indexVec_checkResult_intLMULInput_69,
      indexVec_checkResult_allDataPosition_69[31:11]};
  wire        indexVec_checkResult_unChange_69 = slideUp & (indexVec_readIndex_23[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_23 = validVec[23] & ~indexVec_checkResult_unChange_69;
  wire        indexVec_checkResult_0_4_23 = indexVec_checkResult_overlap_69 | ~indexVec_checkResult_0_5_23 | lagerThanVL | indexVec_checkResult_unChange_69;
  wire [32:0] indexVec_checkResult_allDataPosition_70 = {indexVec_readIndex_23, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_70 = indexVec_checkResult_allDataPosition_70[10:0];
  wire [1:0]  indexVec_checkResult_1_0_23 = {indexVec_checkResult_dataPosition_70[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_23 = indexVec_checkResult_dataPosition_70[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_70 = indexVec_checkResult_dataPosition_70[10:7];
  wire        indexVec_checkResult_1_2_23 = indexVec_checkResult_dataGroup_70[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_70 = indexVec_checkResult_dataGroup_70[3:1];
  wire [2:0]  indexVec_checkResult_1_3_23 = indexVec_checkResult_accessRegGrowth_70;
  wire [5:0]  indexVec_checkResult_decimalProportion_70 = {indexVec_checkResult_1_2_23, indexVec_checkResult_1_1_23};
  wire [2:0]  indexVec_checkResult_decimal_70 = indexVec_checkResult_decimalProportion_70[5:3];
  wire        indexVec_checkResult_overlap_70 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_70 >= indexVec_checkResult_intLMULInput_70[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_70} >= indexVec_checkResult_intLMULInput_70,
      indexVec_checkResult_allDataPosition_70[32:11]};
  wire        indexVec_checkResult_unChange_70 = slideUp & (indexVec_readIndex_23[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_23 = validVec[23] & ~indexVec_checkResult_unChange_70;
  wire        indexVec_checkResult_1_4_23 = indexVec_checkResult_overlap_70 | ~indexVec_checkResult_1_5_23 | lagerThanVL | indexVec_checkResult_unChange_70;
  wire [33:0] indexVec_checkResult_allDataPosition_71 = {indexVec_readIndex_23, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_71 = indexVec_checkResult_allDataPosition_71[10:0];
  wire [4:0]  indexVec_checkResult_2_1_23 = indexVec_checkResult_dataPosition_71[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_71 = indexVec_checkResult_dataPosition_71[10:7];
  wire        indexVec_checkResult_2_2_23 = indexVec_checkResult_dataGroup_71[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_71 = indexVec_checkResult_dataGroup_71[3:1];
  wire [2:0]  indexVec_checkResult_2_3_23 = indexVec_checkResult_accessRegGrowth_71;
  wire [5:0]  indexVec_checkResult_decimalProportion_71 = {indexVec_checkResult_2_2_23, indexVec_checkResult_2_1_23};
  wire [2:0]  indexVec_checkResult_decimal_71 = indexVec_checkResult_decimalProportion_71[5:3];
  wire        indexVec_checkResult_overlap_71 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_71 >= indexVec_checkResult_intLMULInput_71[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_71} >= indexVec_checkResult_intLMULInput_71,
      indexVec_checkResult_allDataPosition_71[33:11]};
  wire        indexVec_checkResult_unChange_71 = slideUp & (indexVec_readIndex_23[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_23 = validVec[23] & ~indexVec_checkResult_unChange_71;
  wire        indexVec_checkResult_2_4_23 = indexVec_checkResult_overlap_71 | ~indexVec_checkResult_2_5_23 | lagerThanVL | indexVec_checkResult_unChange_71;
  wire [1:0]  indexVec_23_0 = (sew1H[0] ? indexVec_checkResult_0_0_23 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_23 : 2'h0);
  assign indexVec_23_1 = (sew1H[0] ? indexVec_checkResult_0_1_23 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_23 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_23 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_23_0 = indexVec_23_1;
  wire        indexVec_23_2 = sew1H[0] & indexVec_checkResult_0_2_23 | sew1H[1] & indexVec_checkResult_1_2_23 | sew1H[2] & indexVec_checkResult_2_2_23;
  assign indexVec_23_3 = (sew1H[0] ? indexVec_checkResult_0_3_23 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_23 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_23 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_23_0 = indexVec_23_3;
  wire        indexVec_23_4 = sew1H[0] & indexVec_checkResult_0_4_23 | sew1H[1] & indexVec_checkResult_1_4_23 | sew1H[2] & indexVec_checkResult_2_4_23;
  wire        indexVec_23_5 = sew1H[0] & indexVec_checkResult_0_5_23 | sew1H[1] & indexVec_checkResult_1_5_23 | sew1H[2] & indexVec_checkResult_2_5_23;
  wire [31:0] indexVec_readIndex_24 = baseIndex + 32'h18;
  wire [31:0] indexVec_checkResult_allDataPosition_72 = indexVec_readIndex_24;
  wire [10:0] indexVec_checkResult_dataPosition_72 = indexVec_checkResult_allDataPosition_72[10:0];
  wire [1:0]  indexVec_checkResult_0_0_24 = indexVec_checkResult_dataPosition_72[1:0];
  wire [4:0]  indexVec_checkResult_0_1_24 = indexVec_checkResult_dataPosition_72[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_72 = indexVec_checkResult_dataPosition_72[10:7];
  wire        indexVec_checkResult_0_2_24 = indexVec_checkResult_dataGroup_72[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_72 = indexVec_checkResult_dataGroup_72[3:1];
  wire [2:0]  indexVec_checkResult_0_3_24 = indexVec_checkResult_accessRegGrowth_72;
  wire [5:0]  indexVec_checkResult_decimalProportion_72 = {indexVec_checkResult_0_2_24, indexVec_checkResult_0_1_24};
  wire [2:0]  indexVec_checkResult_decimal_72 = indexVec_checkResult_decimalProportion_72[5:3];
  wire        indexVec_checkResult_overlap_72 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_72 >= indexVec_checkResult_intLMULInput_72[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_72} >= indexVec_checkResult_intLMULInput_72,
      indexVec_checkResult_allDataPosition_72[31:11]};
  wire        indexVec_checkResult_unChange_72 = slideUp & (indexVec_readIndex_24[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_24 = validVec[24] & ~indexVec_checkResult_unChange_72;
  wire        indexVec_checkResult_0_4_24 = indexVec_checkResult_overlap_72 | ~indexVec_checkResult_0_5_24 | lagerThanVL | indexVec_checkResult_unChange_72;
  wire [32:0] indexVec_checkResult_allDataPosition_73 = {indexVec_readIndex_24, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_73 = indexVec_checkResult_allDataPosition_73[10:0];
  wire [1:0]  indexVec_checkResult_1_0_24 = {indexVec_checkResult_dataPosition_73[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_24 = indexVec_checkResult_dataPosition_73[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_73 = indexVec_checkResult_dataPosition_73[10:7];
  wire        indexVec_checkResult_1_2_24 = indexVec_checkResult_dataGroup_73[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_73 = indexVec_checkResult_dataGroup_73[3:1];
  wire [2:0]  indexVec_checkResult_1_3_24 = indexVec_checkResult_accessRegGrowth_73;
  wire [5:0]  indexVec_checkResult_decimalProportion_73 = {indexVec_checkResult_1_2_24, indexVec_checkResult_1_1_24};
  wire [2:0]  indexVec_checkResult_decimal_73 = indexVec_checkResult_decimalProportion_73[5:3];
  wire        indexVec_checkResult_overlap_73 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_73 >= indexVec_checkResult_intLMULInput_73[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_73} >= indexVec_checkResult_intLMULInput_73,
      indexVec_checkResult_allDataPosition_73[32:11]};
  wire        indexVec_checkResult_unChange_73 = slideUp & (indexVec_readIndex_24[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_24 = validVec[24] & ~indexVec_checkResult_unChange_73;
  wire        indexVec_checkResult_1_4_24 = indexVec_checkResult_overlap_73 | ~indexVec_checkResult_1_5_24 | lagerThanVL | indexVec_checkResult_unChange_73;
  wire [33:0] indexVec_checkResult_allDataPosition_74 = {indexVec_readIndex_24, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_74 = indexVec_checkResult_allDataPosition_74[10:0];
  wire [4:0]  indexVec_checkResult_2_1_24 = indexVec_checkResult_dataPosition_74[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_74 = indexVec_checkResult_dataPosition_74[10:7];
  wire        indexVec_checkResult_2_2_24 = indexVec_checkResult_dataGroup_74[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_74 = indexVec_checkResult_dataGroup_74[3:1];
  wire [2:0]  indexVec_checkResult_2_3_24 = indexVec_checkResult_accessRegGrowth_74;
  wire [5:0]  indexVec_checkResult_decimalProportion_74 = {indexVec_checkResult_2_2_24, indexVec_checkResult_2_1_24};
  wire [2:0]  indexVec_checkResult_decimal_74 = indexVec_checkResult_decimalProportion_74[5:3];
  wire        indexVec_checkResult_overlap_74 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_74 >= indexVec_checkResult_intLMULInput_74[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_74} >= indexVec_checkResult_intLMULInput_74,
      indexVec_checkResult_allDataPosition_74[33:11]};
  wire        indexVec_checkResult_unChange_74 = slideUp & (indexVec_readIndex_24[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_24 = validVec[24] & ~indexVec_checkResult_unChange_74;
  wire        indexVec_checkResult_2_4_24 = indexVec_checkResult_overlap_74 | ~indexVec_checkResult_2_5_24 | lagerThanVL | indexVec_checkResult_unChange_74;
  wire [1:0]  indexVec_24_0 = (sew1H[0] ? indexVec_checkResult_0_0_24 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_24 : 2'h0);
  assign indexVec_24_1 = (sew1H[0] ? indexVec_checkResult_0_1_24 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_24 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_24 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_24_0 = indexVec_24_1;
  wire        indexVec_24_2 = sew1H[0] & indexVec_checkResult_0_2_24 | sew1H[1] & indexVec_checkResult_1_2_24 | sew1H[2] & indexVec_checkResult_2_2_24;
  assign indexVec_24_3 = (sew1H[0] ? indexVec_checkResult_0_3_24 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_24 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_24 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_24_0 = indexVec_24_3;
  wire        indexVec_24_4 = sew1H[0] & indexVec_checkResult_0_4_24 | sew1H[1] & indexVec_checkResult_1_4_24 | sew1H[2] & indexVec_checkResult_2_4_24;
  wire        indexVec_24_5 = sew1H[0] & indexVec_checkResult_0_5_24 | sew1H[1] & indexVec_checkResult_1_5_24 | sew1H[2] & indexVec_checkResult_2_5_24;
  wire [31:0] indexVec_readIndex_25 = baseIndex + 32'h19;
  wire [31:0] indexVec_checkResult_allDataPosition_75 = indexVec_readIndex_25;
  wire [10:0] indexVec_checkResult_dataPosition_75 = indexVec_checkResult_allDataPosition_75[10:0];
  wire [1:0]  indexVec_checkResult_0_0_25 = indexVec_checkResult_dataPosition_75[1:0];
  wire [4:0]  indexVec_checkResult_0_1_25 = indexVec_checkResult_dataPosition_75[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_75 = indexVec_checkResult_dataPosition_75[10:7];
  wire        indexVec_checkResult_0_2_25 = indexVec_checkResult_dataGroup_75[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_75 = indexVec_checkResult_dataGroup_75[3:1];
  wire [2:0]  indexVec_checkResult_0_3_25 = indexVec_checkResult_accessRegGrowth_75;
  wire [5:0]  indexVec_checkResult_decimalProportion_75 = {indexVec_checkResult_0_2_25, indexVec_checkResult_0_1_25};
  wire [2:0]  indexVec_checkResult_decimal_75 = indexVec_checkResult_decimalProportion_75[5:3];
  wire        indexVec_checkResult_overlap_75 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_75 >= indexVec_checkResult_intLMULInput_75[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_75} >= indexVec_checkResult_intLMULInput_75,
      indexVec_checkResult_allDataPosition_75[31:11]};
  wire        indexVec_checkResult_unChange_75 = slideUp & (indexVec_readIndex_25[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_25 = validVec[25] & ~indexVec_checkResult_unChange_75;
  wire        indexVec_checkResult_0_4_25 = indexVec_checkResult_overlap_75 | ~indexVec_checkResult_0_5_25 | lagerThanVL | indexVec_checkResult_unChange_75;
  wire [32:0] indexVec_checkResult_allDataPosition_76 = {indexVec_readIndex_25, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_76 = indexVec_checkResult_allDataPosition_76[10:0];
  wire [1:0]  indexVec_checkResult_1_0_25 = {indexVec_checkResult_dataPosition_76[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_25 = indexVec_checkResult_dataPosition_76[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_76 = indexVec_checkResult_dataPosition_76[10:7];
  wire        indexVec_checkResult_1_2_25 = indexVec_checkResult_dataGroup_76[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_76 = indexVec_checkResult_dataGroup_76[3:1];
  wire [2:0]  indexVec_checkResult_1_3_25 = indexVec_checkResult_accessRegGrowth_76;
  wire [5:0]  indexVec_checkResult_decimalProportion_76 = {indexVec_checkResult_1_2_25, indexVec_checkResult_1_1_25};
  wire [2:0]  indexVec_checkResult_decimal_76 = indexVec_checkResult_decimalProportion_76[5:3];
  wire        indexVec_checkResult_overlap_76 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_76 >= indexVec_checkResult_intLMULInput_76[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_76} >= indexVec_checkResult_intLMULInput_76,
      indexVec_checkResult_allDataPosition_76[32:11]};
  wire        indexVec_checkResult_unChange_76 = slideUp & (indexVec_readIndex_25[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_25 = validVec[25] & ~indexVec_checkResult_unChange_76;
  wire        indexVec_checkResult_1_4_25 = indexVec_checkResult_overlap_76 | ~indexVec_checkResult_1_5_25 | lagerThanVL | indexVec_checkResult_unChange_76;
  wire [33:0] indexVec_checkResult_allDataPosition_77 = {indexVec_readIndex_25, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_77 = indexVec_checkResult_allDataPosition_77[10:0];
  wire [4:0]  indexVec_checkResult_2_1_25 = indexVec_checkResult_dataPosition_77[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_77 = indexVec_checkResult_dataPosition_77[10:7];
  wire        indexVec_checkResult_2_2_25 = indexVec_checkResult_dataGroup_77[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_77 = indexVec_checkResult_dataGroup_77[3:1];
  wire [2:0]  indexVec_checkResult_2_3_25 = indexVec_checkResult_accessRegGrowth_77;
  wire [5:0]  indexVec_checkResult_decimalProportion_77 = {indexVec_checkResult_2_2_25, indexVec_checkResult_2_1_25};
  wire [2:0]  indexVec_checkResult_decimal_77 = indexVec_checkResult_decimalProportion_77[5:3];
  wire        indexVec_checkResult_overlap_77 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_77 >= indexVec_checkResult_intLMULInput_77[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_77} >= indexVec_checkResult_intLMULInput_77,
      indexVec_checkResult_allDataPosition_77[33:11]};
  wire        indexVec_checkResult_unChange_77 = slideUp & (indexVec_readIndex_25[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_25 = validVec[25] & ~indexVec_checkResult_unChange_77;
  wire        indexVec_checkResult_2_4_25 = indexVec_checkResult_overlap_77 | ~indexVec_checkResult_2_5_25 | lagerThanVL | indexVec_checkResult_unChange_77;
  wire [1:0]  indexVec_25_0 = (sew1H[0] ? indexVec_checkResult_0_0_25 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_25 : 2'h0);
  assign indexVec_25_1 = (sew1H[0] ? indexVec_checkResult_0_1_25 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_25 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_25 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_25_0 = indexVec_25_1;
  wire        indexVec_25_2 = sew1H[0] & indexVec_checkResult_0_2_25 | sew1H[1] & indexVec_checkResult_1_2_25 | sew1H[2] & indexVec_checkResult_2_2_25;
  assign indexVec_25_3 = (sew1H[0] ? indexVec_checkResult_0_3_25 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_25 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_25 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_25_0 = indexVec_25_3;
  wire        indexVec_25_4 = sew1H[0] & indexVec_checkResult_0_4_25 | sew1H[1] & indexVec_checkResult_1_4_25 | sew1H[2] & indexVec_checkResult_2_4_25;
  wire        indexVec_25_5 = sew1H[0] & indexVec_checkResult_0_5_25 | sew1H[1] & indexVec_checkResult_1_5_25 | sew1H[2] & indexVec_checkResult_2_5_25;
  wire [31:0] indexVec_readIndex_26 = baseIndex + 32'h1A;
  wire [31:0] indexVec_checkResult_allDataPosition_78 = indexVec_readIndex_26;
  wire [10:0] indexVec_checkResult_dataPosition_78 = indexVec_checkResult_allDataPosition_78[10:0];
  wire [1:0]  indexVec_checkResult_0_0_26 = indexVec_checkResult_dataPosition_78[1:0];
  wire [4:0]  indexVec_checkResult_0_1_26 = indexVec_checkResult_dataPosition_78[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_78 = indexVec_checkResult_dataPosition_78[10:7];
  wire        indexVec_checkResult_0_2_26 = indexVec_checkResult_dataGroup_78[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_78 = indexVec_checkResult_dataGroup_78[3:1];
  wire [2:0]  indexVec_checkResult_0_3_26 = indexVec_checkResult_accessRegGrowth_78;
  wire [5:0]  indexVec_checkResult_decimalProportion_78 = {indexVec_checkResult_0_2_26, indexVec_checkResult_0_1_26};
  wire [2:0]  indexVec_checkResult_decimal_78 = indexVec_checkResult_decimalProportion_78[5:3];
  wire        indexVec_checkResult_overlap_78 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_78 >= indexVec_checkResult_intLMULInput_78[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_78} >= indexVec_checkResult_intLMULInput_78,
      indexVec_checkResult_allDataPosition_78[31:11]};
  wire        indexVec_checkResult_unChange_78 = slideUp & (indexVec_readIndex_26[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_26 = validVec[26] & ~indexVec_checkResult_unChange_78;
  wire        indexVec_checkResult_0_4_26 = indexVec_checkResult_overlap_78 | ~indexVec_checkResult_0_5_26 | lagerThanVL | indexVec_checkResult_unChange_78;
  wire [32:0] indexVec_checkResult_allDataPosition_79 = {indexVec_readIndex_26, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_79 = indexVec_checkResult_allDataPosition_79[10:0];
  wire [1:0]  indexVec_checkResult_1_0_26 = {indexVec_checkResult_dataPosition_79[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_26 = indexVec_checkResult_dataPosition_79[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_79 = indexVec_checkResult_dataPosition_79[10:7];
  wire        indexVec_checkResult_1_2_26 = indexVec_checkResult_dataGroup_79[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_79 = indexVec_checkResult_dataGroup_79[3:1];
  wire [2:0]  indexVec_checkResult_1_3_26 = indexVec_checkResult_accessRegGrowth_79;
  wire [5:0]  indexVec_checkResult_decimalProportion_79 = {indexVec_checkResult_1_2_26, indexVec_checkResult_1_1_26};
  wire [2:0]  indexVec_checkResult_decimal_79 = indexVec_checkResult_decimalProportion_79[5:3];
  wire        indexVec_checkResult_overlap_79 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_79 >= indexVec_checkResult_intLMULInput_79[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_79} >= indexVec_checkResult_intLMULInput_79,
      indexVec_checkResult_allDataPosition_79[32:11]};
  wire        indexVec_checkResult_unChange_79 = slideUp & (indexVec_readIndex_26[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_26 = validVec[26] & ~indexVec_checkResult_unChange_79;
  wire        indexVec_checkResult_1_4_26 = indexVec_checkResult_overlap_79 | ~indexVec_checkResult_1_5_26 | lagerThanVL | indexVec_checkResult_unChange_79;
  wire [33:0] indexVec_checkResult_allDataPosition_80 = {indexVec_readIndex_26, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_80 = indexVec_checkResult_allDataPosition_80[10:0];
  wire [4:0]  indexVec_checkResult_2_1_26 = indexVec_checkResult_dataPosition_80[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_80 = indexVec_checkResult_dataPosition_80[10:7];
  wire        indexVec_checkResult_2_2_26 = indexVec_checkResult_dataGroup_80[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_80 = indexVec_checkResult_dataGroup_80[3:1];
  wire [2:0]  indexVec_checkResult_2_3_26 = indexVec_checkResult_accessRegGrowth_80;
  wire [5:0]  indexVec_checkResult_decimalProportion_80 = {indexVec_checkResult_2_2_26, indexVec_checkResult_2_1_26};
  wire [2:0]  indexVec_checkResult_decimal_80 = indexVec_checkResult_decimalProportion_80[5:3];
  wire        indexVec_checkResult_overlap_80 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_80 >= indexVec_checkResult_intLMULInput_80[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_80} >= indexVec_checkResult_intLMULInput_80,
      indexVec_checkResult_allDataPosition_80[33:11]};
  wire        indexVec_checkResult_unChange_80 = slideUp & (indexVec_readIndex_26[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_26 = validVec[26] & ~indexVec_checkResult_unChange_80;
  wire        indexVec_checkResult_2_4_26 = indexVec_checkResult_overlap_80 | ~indexVec_checkResult_2_5_26 | lagerThanVL | indexVec_checkResult_unChange_80;
  wire [1:0]  indexVec_26_0 = (sew1H[0] ? indexVec_checkResult_0_0_26 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_26 : 2'h0);
  assign indexVec_26_1 = (sew1H[0] ? indexVec_checkResult_0_1_26 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_26 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_26 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_26_0 = indexVec_26_1;
  wire        indexVec_26_2 = sew1H[0] & indexVec_checkResult_0_2_26 | sew1H[1] & indexVec_checkResult_1_2_26 | sew1H[2] & indexVec_checkResult_2_2_26;
  assign indexVec_26_3 = (sew1H[0] ? indexVec_checkResult_0_3_26 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_26 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_26 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_26_0 = indexVec_26_3;
  wire        indexVec_26_4 = sew1H[0] & indexVec_checkResult_0_4_26 | sew1H[1] & indexVec_checkResult_1_4_26 | sew1H[2] & indexVec_checkResult_2_4_26;
  wire        indexVec_26_5 = sew1H[0] & indexVec_checkResult_0_5_26 | sew1H[1] & indexVec_checkResult_1_5_26 | sew1H[2] & indexVec_checkResult_2_5_26;
  wire [31:0] indexVec_readIndex_27 = baseIndex + 32'h1B;
  wire [31:0] indexVec_checkResult_allDataPosition_81 = indexVec_readIndex_27;
  wire [10:0] indexVec_checkResult_dataPosition_81 = indexVec_checkResult_allDataPosition_81[10:0];
  wire [1:0]  indexVec_checkResult_0_0_27 = indexVec_checkResult_dataPosition_81[1:0];
  wire [4:0]  indexVec_checkResult_0_1_27 = indexVec_checkResult_dataPosition_81[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_81 = indexVec_checkResult_dataPosition_81[10:7];
  wire        indexVec_checkResult_0_2_27 = indexVec_checkResult_dataGroup_81[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_81 = indexVec_checkResult_dataGroup_81[3:1];
  wire [2:0]  indexVec_checkResult_0_3_27 = indexVec_checkResult_accessRegGrowth_81;
  wire [5:0]  indexVec_checkResult_decimalProportion_81 = {indexVec_checkResult_0_2_27, indexVec_checkResult_0_1_27};
  wire [2:0]  indexVec_checkResult_decimal_81 = indexVec_checkResult_decimalProportion_81[5:3];
  wire        indexVec_checkResult_overlap_81 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_81 >= indexVec_checkResult_intLMULInput_81[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_81} >= indexVec_checkResult_intLMULInput_81,
      indexVec_checkResult_allDataPosition_81[31:11]};
  wire        indexVec_checkResult_unChange_81 = slideUp & (indexVec_readIndex_27[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_27 = validVec[27] & ~indexVec_checkResult_unChange_81;
  wire        indexVec_checkResult_0_4_27 = indexVec_checkResult_overlap_81 | ~indexVec_checkResult_0_5_27 | lagerThanVL | indexVec_checkResult_unChange_81;
  wire [32:0] indexVec_checkResult_allDataPosition_82 = {indexVec_readIndex_27, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_82 = indexVec_checkResult_allDataPosition_82[10:0];
  wire [1:0]  indexVec_checkResult_1_0_27 = {indexVec_checkResult_dataPosition_82[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_27 = indexVec_checkResult_dataPosition_82[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_82 = indexVec_checkResult_dataPosition_82[10:7];
  wire        indexVec_checkResult_1_2_27 = indexVec_checkResult_dataGroup_82[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_82 = indexVec_checkResult_dataGroup_82[3:1];
  wire [2:0]  indexVec_checkResult_1_3_27 = indexVec_checkResult_accessRegGrowth_82;
  wire [5:0]  indexVec_checkResult_decimalProportion_82 = {indexVec_checkResult_1_2_27, indexVec_checkResult_1_1_27};
  wire [2:0]  indexVec_checkResult_decimal_82 = indexVec_checkResult_decimalProportion_82[5:3];
  wire        indexVec_checkResult_overlap_82 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_82 >= indexVec_checkResult_intLMULInput_82[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_82} >= indexVec_checkResult_intLMULInput_82,
      indexVec_checkResult_allDataPosition_82[32:11]};
  wire        indexVec_checkResult_unChange_82 = slideUp & (indexVec_readIndex_27[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_27 = validVec[27] & ~indexVec_checkResult_unChange_82;
  wire        indexVec_checkResult_1_4_27 = indexVec_checkResult_overlap_82 | ~indexVec_checkResult_1_5_27 | lagerThanVL | indexVec_checkResult_unChange_82;
  wire [33:0] indexVec_checkResult_allDataPosition_83 = {indexVec_readIndex_27, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_83 = indexVec_checkResult_allDataPosition_83[10:0];
  wire [4:0]  indexVec_checkResult_2_1_27 = indexVec_checkResult_dataPosition_83[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_83 = indexVec_checkResult_dataPosition_83[10:7];
  wire        indexVec_checkResult_2_2_27 = indexVec_checkResult_dataGroup_83[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_83 = indexVec_checkResult_dataGroup_83[3:1];
  wire [2:0]  indexVec_checkResult_2_3_27 = indexVec_checkResult_accessRegGrowth_83;
  wire [5:0]  indexVec_checkResult_decimalProportion_83 = {indexVec_checkResult_2_2_27, indexVec_checkResult_2_1_27};
  wire [2:0]  indexVec_checkResult_decimal_83 = indexVec_checkResult_decimalProportion_83[5:3];
  wire        indexVec_checkResult_overlap_83 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_83 >= indexVec_checkResult_intLMULInput_83[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_83} >= indexVec_checkResult_intLMULInput_83,
      indexVec_checkResult_allDataPosition_83[33:11]};
  wire        indexVec_checkResult_unChange_83 = slideUp & (indexVec_readIndex_27[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_27 = validVec[27] & ~indexVec_checkResult_unChange_83;
  wire        indexVec_checkResult_2_4_27 = indexVec_checkResult_overlap_83 | ~indexVec_checkResult_2_5_27 | lagerThanVL | indexVec_checkResult_unChange_83;
  wire [1:0]  indexVec_27_0 = (sew1H[0] ? indexVec_checkResult_0_0_27 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_27 : 2'h0);
  assign indexVec_27_1 = (sew1H[0] ? indexVec_checkResult_0_1_27 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_27 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_27 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_27_0 = indexVec_27_1;
  wire        indexVec_27_2 = sew1H[0] & indexVec_checkResult_0_2_27 | sew1H[1] & indexVec_checkResult_1_2_27 | sew1H[2] & indexVec_checkResult_2_2_27;
  assign indexVec_27_3 = (sew1H[0] ? indexVec_checkResult_0_3_27 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_27 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_27 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_27_0 = indexVec_27_3;
  wire        indexVec_27_4 = sew1H[0] & indexVec_checkResult_0_4_27 | sew1H[1] & indexVec_checkResult_1_4_27 | sew1H[2] & indexVec_checkResult_2_4_27;
  wire        indexVec_27_5 = sew1H[0] & indexVec_checkResult_0_5_27 | sew1H[1] & indexVec_checkResult_1_5_27 | sew1H[2] & indexVec_checkResult_2_5_27;
  wire [31:0] indexVec_readIndex_28 = baseIndex + 32'h1C;
  wire [31:0] indexVec_checkResult_allDataPosition_84 = indexVec_readIndex_28;
  wire [10:0] indexVec_checkResult_dataPosition_84 = indexVec_checkResult_allDataPosition_84[10:0];
  wire [1:0]  indexVec_checkResult_0_0_28 = indexVec_checkResult_dataPosition_84[1:0];
  wire [4:0]  indexVec_checkResult_0_1_28 = indexVec_checkResult_dataPosition_84[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_84 = indexVec_checkResult_dataPosition_84[10:7];
  wire        indexVec_checkResult_0_2_28 = indexVec_checkResult_dataGroup_84[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_84 = indexVec_checkResult_dataGroup_84[3:1];
  wire [2:0]  indexVec_checkResult_0_3_28 = indexVec_checkResult_accessRegGrowth_84;
  wire [5:0]  indexVec_checkResult_decimalProportion_84 = {indexVec_checkResult_0_2_28, indexVec_checkResult_0_1_28};
  wire [2:0]  indexVec_checkResult_decimal_84 = indexVec_checkResult_decimalProportion_84[5:3];
  wire        indexVec_checkResult_overlap_84 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_84 >= indexVec_checkResult_intLMULInput_84[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_84} >= indexVec_checkResult_intLMULInput_84,
      indexVec_checkResult_allDataPosition_84[31:11]};
  wire        indexVec_checkResult_unChange_84 = slideUp & (indexVec_readIndex_28[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_28 = validVec[28] & ~indexVec_checkResult_unChange_84;
  wire        indexVec_checkResult_0_4_28 = indexVec_checkResult_overlap_84 | ~indexVec_checkResult_0_5_28 | lagerThanVL | indexVec_checkResult_unChange_84;
  wire [32:0] indexVec_checkResult_allDataPosition_85 = {indexVec_readIndex_28, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_85 = indexVec_checkResult_allDataPosition_85[10:0];
  wire [1:0]  indexVec_checkResult_1_0_28 = {indexVec_checkResult_dataPosition_85[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_28 = indexVec_checkResult_dataPosition_85[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_85 = indexVec_checkResult_dataPosition_85[10:7];
  wire        indexVec_checkResult_1_2_28 = indexVec_checkResult_dataGroup_85[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_85 = indexVec_checkResult_dataGroup_85[3:1];
  wire [2:0]  indexVec_checkResult_1_3_28 = indexVec_checkResult_accessRegGrowth_85;
  wire [5:0]  indexVec_checkResult_decimalProportion_85 = {indexVec_checkResult_1_2_28, indexVec_checkResult_1_1_28};
  wire [2:0]  indexVec_checkResult_decimal_85 = indexVec_checkResult_decimalProportion_85[5:3];
  wire        indexVec_checkResult_overlap_85 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_85 >= indexVec_checkResult_intLMULInput_85[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_85} >= indexVec_checkResult_intLMULInput_85,
      indexVec_checkResult_allDataPosition_85[32:11]};
  wire        indexVec_checkResult_unChange_85 = slideUp & (indexVec_readIndex_28[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_28 = validVec[28] & ~indexVec_checkResult_unChange_85;
  wire        indexVec_checkResult_1_4_28 = indexVec_checkResult_overlap_85 | ~indexVec_checkResult_1_5_28 | lagerThanVL | indexVec_checkResult_unChange_85;
  wire [33:0] indexVec_checkResult_allDataPosition_86 = {indexVec_readIndex_28, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_86 = indexVec_checkResult_allDataPosition_86[10:0];
  wire [4:0]  indexVec_checkResult_2_1_28 = indexVec_checkResult_dataPosition_86[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_86 = indexVec_checkResult_dataPosition_86[10:7];
  wire        indexVec_checkResult_2_2_28 = indexVec_checkResult_dataGroup_86[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_86 = indexVec_checkResult_dataGroup_86[3:1];
  wire [2:0]  indexVec_checkResult_2_3_28 = indexVec_checkResult_accessRegGrowth_86;
  wire [5:0]  indexVec_checkResult_decimalProportion_86 = {indexVec_checkResult_2_2_28, indexVec_checkResult_2_1_28};
  wire [2:0]  indexVec_checkResult_decimal_86 = indexVec_checkResult_decimalProportion_86[5:3];
  wire        indexVec_checkResult_overlap_86 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_86 >= indexVec_checkResult_intLMULInput_86[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_86} >= indexVec_checkResult_intLMULInput_86,
      indexVec_checkResult_allDataPosition_86[33:11]};
  wire        indexVec_checkResult_unChange_86 = slideUp & (indexVec_readIndex_28[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_28 = validVec[28] & ~indexVec_checkResult_unChange_86;
  wire        indexVec_checkResult_2_4_28 = indexVec_checkResult_overlap_86 | ~indexVec_checkResult_2_5_28 | lagerThanVL | indexVec_checkResult_unChange_86;
  wire [1:0]  indexVec_28_0 = (sew1H[0] ? indexVec_checkResult_0_0_28 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_28 : 2'h0);
  assign indexVec_28_1 = (sew1H[0] ? indexVec_checkResult_0_1_28 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_28 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_28 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_28_0 = indexVec_28_1;
  wire        indexVec_28_2 = sew1H[0] & indexVec_checkResult_0_2_28 | sew1H[1] & indexVec_checkResult_1_2_28 | sew1H[2] & indexVec_checkResult_2_2_28;
  assign indexVec_28_3 = (sew1H[0] ? indexVec_checkResult_0_3_28 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_28 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_28 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_28_0 = indexVec_28_3;
  wire        indexVec_28_4 = sew1H[0] & indexVec_checkResult_0_4_28 | sew1H[1] & indexVec_checkResult_1_4_28 | sew1H[2] & indexVec_checkResult_2_4_28;
  wire        indexVec_28_5 = sew1H[0] & indexVec_checkResult_0_5_28 | sew1H[1] & indexVec_checkResult_1_5_28 | sew1H[2] & indexVec_checkResult_2_5_28;
  wire [31:0] indexVec_readIndex_29 = baseIndex + 32'h1D;
  wire [31:0] indexVec_checkResult_allDataPosition_87 = indexVec_readIndex_29;
  wire [10:0] indexVec_checkResult_dataPosition_87 = indexVec_checkResult_allDataPosition_87[10:0];
  wire [1:0]  indexVec_checkResult_0_0_29 = indexVec_checkResult_dataPosition_87[1:0];
  wire [4:0]  indexVec_checkResult_0_1_29 = indexVec_checkResult_dataPosition_87[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_87 = indexVec_checkResult_dataPosition_87[10:7];
  wire        indexVec_checkResult_0_2_29 = indexVec_checkResult_dataGroup_87[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_87 = indexVec_checkResult_dataGroup_87[3:1];
  wire [2:0]  indexVec_checkResult_0_3_29 = indexVec_checkResult_accessRegGrowth_87;
  wire [5:0]  indexVec_checkResult_decimalProportion_87 = {indexVec_checkResult_0_2_29, indexVec_checkResult_0_1_29};
  wire [2:0]  indexVec_checkResult_decimal_87 = indexVec_checkResult_decimalProportion_87[5:3];
  wire        indexVec_checkResult_overlap_87 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_87 >= indexVec_checkResult_intLMULInput_87[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_87} >= indexVec_checkResult_intLMULInput_87,
      indexVec_checkResult_allDataPosition_87[31:11]};
  wire        indexVec_checkResult_unChange_87 = slideUp & (indexVec_readIndex_29[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_29 = validVec[29] & ~indexVec_checkResult_unChange_87;
  wire        indexVec_checkResult_0_4_29 = indexVec_checkResult_overlap_87 | ~indexVec_checkResult_0_5_29 | lagerThanVL | indexVec_checkResult_unChange_87;
  wire [32:0] indexVec_checkResult_allDataPosition_88 = {indexVec_readIndex_29, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_88 = indexVec_checkResult_allDataPosition_88[10:0];
  wire [1:0]  indexVec_checkResult_1_0_29 = {indexVec_checkResult_dataPosition_88[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_29 = indexVec_checkResult_dataPosition_88[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_88 = indexVec_checkResult_dataPosition_88[10:7];
  wire        indexVec_checkResult_1_2_29 = indexVec_checkResult_dataGroup_88[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_88 = indexVec_checkResult_dataGroup_88[3:1];
  wire [2:0]  indexVec_checkResult_1_3_29 = indexVec_checkResult_accessRegGrowth_88;
  wire [5:0]  indexVec_checkResult_decimalProportion_88 = {indexVec_checkResult_1_2_29, indexVec_checkResult_1_1_29};
  wire [2:0]  indexVec_checkResult_decimal_88 = indexVec_checkResult_decimalProportion_88[5:3];
  wire        indexVec_checkResult_overlap_88 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_88 >= indexVec_checkResult_intLMULInput_88[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_88} >= indexVec_checkResult_intLMULInput_88,
      indexVec_checkResult_allDataPosition_88[32:11]};
  wire        indexVec_checkResult_unChange_88 = slideUp & (indexVec_readIndex_29[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_29 = validVec[29] & ~indexVec_checkResult_unChange_88;
  wire        indexVec_checkResult_1_4_29 = indexVec_checkResult_overlap_88 | ~indexVec_checkResult_1_5_29 | lagerThanVL | indexVec_checkResult_unChange_88;
  wire [33:0] indexVec_checkResult_allDataPosition_89 = {indexVec_readIndex_29, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_89 = indexVec_checkResult_allDataPosition_89[10:0];
  wire [4:0]  indexVec_checkResult_2_1_29 = indexVec_checkResult_dataPosition_89[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_89 = indexVec_checkResult_dataPosition_89[10:7];
  wire        indexVec_checkResult_2_2_29 = indexVec_checkResult_dataGroup_89[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_89 = indexVec_checkResult_dataGroup_89[3:1];
  wire [2:0]  indexVec_checkResult_2_3_29 = indexVec_checkResult_accessRegGrowth_89;
  wire [5:0]  indexVec_checkResult_decimalProportion_89 = {indexVec_checkResult_2_2_29, indexVec_checkResult_2_1_29};
  wire [2:0]  indexVec_checkResult_decimal_89 = indexVec_checkResult_decimalProportion_89[5:3];
  wire        indexVec_checkResult_overlap_89 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_89 >= indexVec_checkResult_intLMULInput_89[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_89} >= indexVec_checkResult_intLMULInput_89,
      indexVec_checkResult_allDataPosition_89[33:11]};
  wire        indexVec_checkResult_unChange_89 = slideUp & (indexVec_readIndex_29[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_29 = validVec[29] & ~indexVec_checkResult_unChange_89;
  wire        indexVec_checkResult_2_4_29 = indexVec_checkResult_overlap_89 | ~indexVec_checkResult_2_5_29 | lagerThanVL | indexVec_checkResult_unChange_89;
  wire [1:0]  indexVec_29_0 = (sew1H[0] ? indexVec_checkResult_0_0_29 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_29 : 2'h0);
  assign indexVec_29_1 = (sew1H[0] ? indexVec_checkResult_0_1_29 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_29 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_29 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_29_0 = indexVec_29_1;
  wire        indexVec_29_2 = sew1H[0] & indexVec_checkResult_0_2_29 | sew1H[1] & indexVec_checkResult_1_2_29 | sew1H[2] & indexVec_checkResult_2_2_29;
  assign indexVec_29_3 = (sew1H[0] ? indexVec_checkResult_0_3_29 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_29 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_29 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_29_0 = indexVec_29_3;
  wire        indexVec_29_4 = sew1H[0] & indexVec_checkResult_0_4_29 | sew1H[1] & indexVec_checkResult_1_4_29 | sew1H[2] & indexVec_checkResult_2_4_29;
  wire        indexVec_29_5 = sew1H[0] & indexVec_checkResult_0_5_29 | sew1H[1] & indexVec_checkResult_1_5_29 | sew1H[2] & indexVec_checkResult_2_5_29;
  wire [31:0] indexVec_readIndex_30 = baseIndex + 32'h1E;
  wire [31:0] indexVec_checkResult_allDataPosition_90 = indexVec_readIndex_30;
  wire [10:0] indexVec_checkResult_dataPosition_90 = indexVec_checkResult_allDataPosition_90[10:0];
  wire [1:0]  indexVec_checkResult_0_0_30 = indexVec_checkResult_dataPosition_90[1:0];
  wire [4:0]  indexVec_checkResult_0_1_30 = indexVec_checkResult_dataPosition_90[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_90 = indexVec_checkResult_dataPosition_90[10:7];
  wire        indexVec_checkResult_0_2_30 = indexVec_checkResult_dataGroup_90[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_90 = indexVec_checkResult_dataGroup_90[3:1];
  wire [2:0]  indexVec_checkResult_0_3_30 = indexVec_checkResult_accessRegGrowth_90;
  wire [5:0]  indexVec_checkResult_decimalProportion_90 = {indexVec_checkResult_0_2_30, indexVec_checkResult_0_1_30};
  wire [2:0]  indexVec_checkResult_decimal_90 = indexVec_checkResult_decimalProportion_90[5:3];
  wire        indexVec_checkResult_overlap_90 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_90 >= indexVec_checkResult_intLMULInput_90[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_90} >= indexVec_checkResult_intLMULInput_90,
      indexVec_checkResult_allDataPosition_90[31:11]};
  wire        indexVec_checkResult_unChange_90 = slideUp & (indexVec_readIndex_30[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_30 = validVec[30] & ~indexVec_checkResult_unChange_90;
  wire        indexVec_checkResult_0_4_30 = indexVec_checkResult_overlap_90 | ~indexVec_checkResult_0_5_30 | lagerThanVL | indexVec_checkResult_unChange_90;
  wire [32:0] indexVec_checkResult_allDataPosition_91 = {indexVec_readIndex_30, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_91 = indexVec_checkResult_allDataPosition_91[10:0];
  wire [1:0]  indexVec_checkResult_1_0_30 = {indexVec_checkResult_dataPosition_91[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_30 = indexVec_checkResult_dataPosition_91[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_91 = indexVec_checkResult_dataPosition_91[10:7];
  wire        indexVec_checkResult_1_2_30 = indexVec_checkResult_dataGroup_91[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_91 = indexVec_checkResult_dataGroup_91[3:1];
  wire [2:0]  indexVec_checkResult_1_3_30 = indexVec_checkResult_accessRegGrowth_91;
  wire [5:0]  indexVec_checkResult_decimalProportion_91 = {indexVec_checkResult_1_2_30, indexVec_checkResult_1_1_30};
  wire [2:0]  indexVec_checkResult_decimal_91 = indexVec_checkResult_decimalProportion_91[5:3];
  wire        indexVec_checkResult_overlap_91 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_91 >= indexVec_checkResult_intLMULInput_91[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_91} >= indexVec_checkResult_intLMULInput_91,
      indexVec_checkResult_allDataPosition_91[32:11]};
  wire        indexVec_checkResult_unChange_91 = slideUp & (indexVec_readIndex_30[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_30 = validVec[30] & ~indexVec_checkResult_unChange_91;
  wire        indexVec_checkResult_1_4_30 = indexVec_checkResult_overlap_91 | ~indexVec_checkResult_1_5_30 | lagerThanVL | indexVec_checkResult_unChange_91;
  wire [33:0] indexVec_checkResult_allDataPosition_92 = {indexVec_readIndex_30, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_92 = indexVec_checkResult_allDataPosition_92[10:0];
  wire [4:0]  indexVec_checkResult_2_1_30 = indexVec_checkResult_dataPosition_92[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_92 = indexVec_checkResult_dataPosition_92[10:7];
  wire        indexVec_checkResult_2_2_30 = indexVec_checkResult_dataGroup_92[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_92 = indexVec_checkResult_dataGroup_92[3:1];
  wire [2:0]  indexVec_checkResult_2_3_30 = indexVec_checkResult_accessRegGrowth_92;
  wire [5:0]  indexVec_checkResult_decimalProportion_92 = {indexVec_checkResult_2_2_30, indexVec_checkResult_2_1_30};
  wire [2:0]  indexVec_checkResult_decimal_92 = indexVec_checkResult_decimalProportion_92[5:3];
  wire        indexVec_checkResult_overlap_92 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_92 >= indexVec_checkResult_intLMULInput_92[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_92} >= indexVec_checkResult_intLMULInput_92,
      indexVec_checkResult_allDataPosition_92[33:11]};
  wire        indexVec_checkResult_unChange_92 = slideUp & (indexVec_readIndex_30[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_30 = validVec[30] & ~indexVec_checkResult_unChange_92;
  wire        indexVec_checkResult_2_4_30 = indexVec_checkResult_overlap_92 | ~indexVec_checkResult_2_5_30 | lagerThanVL | indexVec_checkResult_unChange_92;
  wire [1:0]  indexVec_30_0 = (sew1H[0] ? indexVec_checkResult_0_0_30 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_30 : 2'h0);
  assign indexVec_30_1 = (sew1H[0] ? indexVec_checkResult_0_1_30 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_30 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_30 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_30_0 = indexVec_30_1;
  wire        indexVec_30_2 = sew1H[0] & indexVec_checkResult_0_2_30 | sew1H[1] & indexVec_checkResult_1_2_30 | sew1H[2] & indexVec_checkResult_2_2_30;
  assign indexVec_30_3 = (sew1H[0] ? indexVec_checkResult_0_3_30 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_30 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_30 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_30_0 = indexVec_30_3;
  wire        indexVec_30_4 = sew1H[0] & indexVec_checkResult_0_4_30 | sew1H[1] & indexVec_checkResult_1_4_30 | sew1H[2] & indexVec_checkResult_2_4_30;
  wire        indexVec_30_5 = sew1H[0] & indexVec_checkResult_0_5_30 | sew1H[1] & indexVec_checkResult_1_5_30 | sew1H[2] & indexVec_checkResult_2_5_30;
  wire [31:0] indexVec_readIndex_31 = baseIndex + 32'h1F;
  wire [31:0] indexVec_checkResult_allDataPosition_93 = indexVec_readIndex_31;
  wire [10:0] indexVec_checkResult_dataPosition_93 = indexVec_checkResult_allDataPosition_93[10:0];
  wire [1:0]  indexVec_checkResult_0_0_31 = indexVec_checkResult_dataPosition_93[1:0];
  wire [4:0]  indexVec_checkResult_0_1_31 = indexVec_checkResult_dataPosition_93[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_93 = indexVec_checkResult_dataPosition_93[10:7];
  wire        indexVec_checkResult_0_2_31 = indexVec_checkResult_dataGroup_93[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_93 = indexVec_checkResult_dataGroup_93[3:1];
  wire [2:0]  indexVec_checkResult_0_3_31 = indexVec_checkResult_accessRegGrowth_93;
  wire [5:0]  indexVec_checkResult_decimalProportion_93 = {indexVec_checkResult_0_2_31, indexVec_checkResult_0_1_31};
  wire [2:0]  indexVec_checkResult_decimal_93 = indexVec_checkResult_decimalProportion_93[5:3];
  wire        indexVec_checkResult_overlap_93 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_93 >= indexVec_checkResult_intLMULInput_93[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_93} >= indexVec_checkResult_intLMULInput_93,
      indexVec_checkResult_allDataPosition_93[31:11]};
  wire        indexVec_checkResult_unChange_93 = slideUp & (indexVec_readIndex_31[31] | lagerThanVL);
  wire        indexVec_checkResult_0_5_31 = validVec[31] & ~indexVec_checkResult_unChange_93;
  wire        indexVec_checkResult_0_4_31 = indexVec_checkResult_overlap_93 | ~indexVec_checkResult_0_5_31 | lagerThanVL | indexVec_checkResult_unChange_93;
  wire [32:0] indexVec_checkResult_allDataPosition_94 = {indexVec_readIndex_31, 1'h0};
  wire [10:0] indexVec_checkResult_dataPosition_94 = indexVec_checkResult_allDataPosition_94[10:0];
  wire [1:0]  indexVec_checkResult_1_0_31 = {indexVec_checkResult_dataPosition_94[1], 1'h0};
  wire [4:0]  indexVec_checkResult_1_1_31 = indexVec_checkResult_dataPosition_94[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_94 = indexVec_checkResult_dataPosition_94[10:7];
  wire        indexVec_checkResult_1_2_31 = indexVec_checkResult_dataGroup_94[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_94 = indexVec_checkResult_dataGroup_94[3:1];
  wire [2:0]  indexVec_checkResult_1_3_31 = indexVec_checkResult_accessRegGrowth_94;
  wire [5:0]  indexVec_checkResult_decimalProportion_94 = {indexVec_checkResult_1_2_31, indexVec_checkResult_1_1_31};
  wire [2:0]  indexVec_checkResult_decimal_94 = indexVec_checkResult_decimalProportion_94[5:3];
  wire        indexVec_checkResult_overlap_94 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_94 >= indexVec_checkResult_intLMULInput_94[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_94} >= indexVec_checkResult_intLMULInput_94,
      indexVec_checkResult_allDataPosition_94[32:11]};
  wire        indexVec_checkResult_unChange_94 = slideUp & (indexVec_readIndex_31[31] | lagerThanVL);
  wire        indexVec_checkResult_1_5_31 = validVec[31] & ~indexVec_checkResult_unChange_94;
  wire        indexVec_checkResult_1_4_31 = indexVec_checkResult_overlap_94 | ~indexVec_checkResult_1_5_31 | lagerThanVL | indexVec_checkResult_unChange_94;
  wire [33:0] indexVec_checkResult_allDataPosition_95 = {indexVec_readIndex_31, 2'h0};
  wire [10:0] indexVec_checkResult_dataPosition_95 = indexVec_checkResult_allDataPosition_95[10:0];
  wire [4:0]  indexVec_checkResult_2_1_31 = indexVec_checkResult_dataPosition_95[6:2];
  wire [3:0]  indexVec_checkResult_dataGroup_95 = indexVec_checkResult_dataPosition_95[10:7];
  wire        indexVec_checkResult_2_2_31 = indexVec_checkResult_dataGroup_95[0];
  wire [2:0]  indexVec_checkResult_accessRegGrowth_95 = indexVec_checkResult_dataGroup_95[3:1];
  wire [2:0]  indexVec_checkResult_2_3_31 = indexVec_checkResult_accessRegGrowth_95;
  wire [5:0]  indexVec_checkResult_decimalProportion_95 = {indexVec_checkResult_2_2_31, indexVec_checkResult_2_1_31};
  wire [2:0]  indexVec_checkResult_decimal_95 = indexVec_checkResult_decimalProportion_95[5:3];
  wire        indexVec_checkResult_overlap_95 =
    |{instructionReq_vlmul[2] & indexVec_checkResult_decimal_95 >= indexVec_checkResult_intLMULInput_95[3:1] | ~(instructionReq_vlmul[2]) & {1'h0, indexVec_checkResult_accessRegGrowth_95} >= indexVec_checkResult_intLMULInput_95,
      indexVec_checkResult_allDataPosition_95[33:11]};
  wire        indexVec_checkResult_unChange_95 = slideUp & (indexVec_readIndex_31[31] | lagerThanVL);
  wire        indexVec_checkResult_2_5_31 = validVec[31] & ~indexVec_checkResult_unChange_95;
  wire        indexVec_checkResult_2_4_31 = indexVec_checkResult_overlap_95 | ~indexVec_checkResult_2_5_31 | lagerThanVL | indexVec_checkResult_unChange_95;
  wire [1:0]  indexVec_31_0 = (sew1H[0] ? indexVec_checkResult_0_0_31 : 2'h0) | (sew1H[1] ? indexVec_checkResult_1_0_31 : 2'h0);
  assign indexVec_31_1 = (sew1H[0] ? indexVec_checkResult_0_1_31 : 5'h0) | (sew1H[1] ? indexVec_checkResult_1_1_31 : 5'h0) | (sew1H[2] ? indexVec_checkResult_2_1_31 : 5'h0);
  wire [4:0]  indexDeq_bits_accessLane_31_0 = indexVec_31_1;
  wire        indexVec_31_2 = sew1H[0] & indexVec_checkResult_0_2_31 | sew1H[1] & indexVec_checkResult_1_2_31 | sew1H[2] & indexVec_checkResult_2_2_31;
  assign indexVec_31_3 = (sew1H[0] ? indexVec_checkResult_0_3_31 : 3'h0) | (sew1H[1] ? indexVec_checkResult_1_3_31 : 3'h0) | (sew1H[2] ? indexVec_checkResult_2_3_31 : 3'h0);
  wire [2:0]  indexDeq_bits_vsGrowth_31_0 = indexVec_31_3;
  wire        indexVec_31_4 = sew1H[0] & indexVec_checkResult_0_4_31 | sew1H[1] & indexVec_checkResult_1_4_31 | sew1H[2] & indexVec_checkResult_2_4_31;
  wire        indexVec_31_5 = sew1H[0] & indexVec_checkResult_0_5_31 | sew1H[1] & indexVec_checkResult_1_5_31 | sew1H[2] & indexVec_checkResult_2_5_31;
  assign indexDeq_valid_0 = InstructionValid & isSlide;
  wire [1:0]  indexDeq_bits_needRead_lo_lo_lo_lo = {~indexVec_1_4, ~indexVec_0_4};
  wire [1:0]  indexDeq_bits_needRead_lo_lo_lo_hi = {~indexVec_3_4, ~indexVec_2_4};
  wire [3:0]  indexDeq_bits_needRead_lo_lo_lo = {indexDeq_bits_needRead_lo_lo_lo_hi, indexDeq_bits_needRead_lo_lo_lo_lo};
  wire [1:0]  indexDeq_bits_needRead_lo_lo_hi_lo = {~indexVec_5_4, ~indexVec_4_4};
  wire [1:0]  indexDeq_bits_needRead_lo_lo_hi_hi = {~indexVec_7_4, ~indexVec_6_4};
  wire [3:0]  indexDeq_bits_needRead_lo_lo_hi = {indexDeq_bits_needRead_lo_lo_hi_hi, indexDeq_bits_needRead_lo_lo_hi_lo};
  wire [7:0]  indexDeq_bits_needRead_lo_lo = {indexDeq_bits_needRead_lo_lo_hi, indexDeq_bits_needRead_lo_lo_lo};
  wire [1:0]  indexDeq_bits_needRead_lo_hi_lo_lo = {~indexVec_9_4, ~indexVec_8_4};
  wire [1:0]  indexDeq_bits_needRead_lo_hi_lo_hi = {~indexVec_11_4, ~indexVec_10_4};
  wire [3:0]  indexDeq_bits_needRead_lo_hi_lo = {indexDeq_bits_needRead_lo_hi_lo_hi, indexDeq_bits_needRead_lo_hi_lo_lo};
  wire [1:0]  indexDeq_bits_needRead_lo_hi_hi_lo = {~indexVec_13_4, ~indexVec_12_4};
  wire [1:0]  indexDeq_bits_needRead_lo_hi_hi_hi = {~indexVec_15_4, ~indexVec_14_4};
  wire [3:0]  indexDeq_bits_needRead_lo_hi_hi = {indexDeq_bits_needRead_lo_hi_hi_hi, indexDeq_bits_needRead_lo_hi_hi_lo};
  wire [7:0]  indexDeq_bits_needRead_lo_hi = {indexDeq_bits_needRead_lo_hi_hi, indexDeq_bits_needRead_lo_hi_lo};
  wire [15:0] indexDeq_bits_needRead_lo = {indexDeq_bits_needRead_lo_hi, indexDeq_bits_needRead_lo_lo};
  wire [1:0]  indexDeq_bits_needRead_hi_lo_lo_lo = {~indexVec_17_4, ~indexVec_16_4};
  wire [1:0]  indexDeq_bits_needRead_hi_lo_lo_hi = {~indexVec_19_4, ~indexVec_18_4};
  wire [3:0]  indexDeq_bits_needRead_hi_lo_lo = {indexDeq_bits_needRead_hi_lo_lo_hi, indexDeq_bits_needRead_hi_lo_lo_lo};
  wire [1:0]  indexDeq_bits_needRead_hi_lo_hi_lo = {~indexVec_21_4, ~indexVec_20_4};
  wire [1:0]  indexDeq_bits_needRead_hi_lo_hi_hi = {~indexVec_23_4, ~indexVec_22_4};
  wire [3:0]  indexDeq_bits_needRead_hi_lo_hi = {indexDeq_bits_needRead_hi_lo_hi_hi, indexDeq_bits_needRead_hi_lo_hi_lo};
  wire [7:0]  indexDeq_bits_needRead_hi_lo = {indexDeq_bits_needRead_hi_lo_hi, indexDeq_bits_needRead_hi_lo_lo};
  wire [1:0]  indexDeq_bits_needRead_hi_hi_lo_lo = {~indexVec_25_4, ~indexVec_24_4};
  wire [1:0]  indexDeq_bits_needRead_hi_hi_lo_hi = {~indexVec_27_4, ~indexVec_26_4};
  wire [3:0]  indexDeq_bits_needRead_hi_hi_lo = {indexDeq_bits_needRead_hi_hi_lo_hi, indexDeq_bits_needRead_hi_hi_lo_lo};
  wire [1:0]  indexDeq_bits_needRead_hi_hi_hi_lo = {~indexVec_29_4, ~indexVec_28_4};
  wire [1:0]  indexDeq_bits_needRead_hi_hi_hi_hi = {~indexVec_31_4, ~indexVec_30_4};
  wire [3:0]  indexDeq_bits_needRead_hi_hi_hi = {indexDeq_bits_needRead_hi_hi_hi_hi, indexDeq_bits_needRead_hi_hi_hi_lo};
  wire [7:0]  indexDeq_bits_needRead_hi_hi = {indexDeq_bits_needRead_hi_hi_hi, indexDeq_bits_needRead_hi_hi_lo};
  wire [15:0] indexDeq_bits_needRead_hi = {indexDeq_bits_needRead_hi_hi, indexDeq_bits_needRead_hi_lo};
  wire [31:0] indexDeq_bits_needRead_0 = {indexDeq_bits_needRead_hi, indexDeq_bits_needRead_lo} & ~replaceWithVs1;
  wire [1:0]  indexDeq_bits_elementValid_lo_lo_lo_lo = {indexVec_1_5, indexVec_0_5};
  wire [1:0]  indexDeq_bits_elementValid_lo_lo_lo_hi = {indexVec_3_5, indexVec_2_5};
  wire [3:0]  indexDeq_bits_elementValid_lo_lo_lo = {indexDeq_bits_elementValid_lo_lo_lo_hi, indexDeq_bits_elementValid_lo_lo_lo_lo};
  wire [1:0]  indexDeq_bits_elementValid_lo_lo_hi_lo = {indexVec_5_5, indexVec_4_5};
  wire [1:0]  indexDeq_bits_elementValid_lo_lo_hi_hi = {indexVec_7_5, indexVec_6_5};
  wire [3:0]  indexDeq_bits_elementValid_lo_lo_hi = {indexDeq_bits_elementValid_lo_lo_hi_hi, indexDeq_bits_elementValid_lo_lo_hi_lo};
  wire [7:0]  indexDeq_bits_elementValid_lo_lo = {indexDeq_bits_elementValid_lo_lo_hi, indexDeq_bits_elementValid_lo_lo_lo};
  wire [1:0]  indexDeq_bits_elementValid_lo_hi_lo_lo = {indexVec_9_5, indexVec_8_5};
  wire [1:0]  indexDeq_bits_elementValid_lo_hi_lo_hi = {indexVec_11_5, indexVec_10_5};
  wire [3:0]  indexDeq_bits_elementValid_lo_hi_lo = {indexDeq_bits_elementValid_lo_hi_lo_hi, indexDeq_bits_elementValid_lo_hi_lo_lo};
  wire [1:0]  indexDeq_bits_elementValid_lo_hi_hi_lo = {indexVec_13_5, indexVec_12_5};
  wire [1:0]  indexDeq_bits_elementValid_lo_hi_hi_hi = {indexVec_15_5, indexVec_14_5};
  wire [3:0]  indexDeq_bits_elementValid_lo_hi_hi = {indexDeq_bits_elementValid_lo_hi_hi_hi, indexDeq_bits_elementValid_lo_hi_hi_lo};
  wire [7:0]  indexDeq_bits_elementValid_lo_hi = {indexDeq_bits_elementValid_lo_hi_hi, indexDeq_bits_elementValid_lo_hi_lo};
  wire [15:0] indexDeq_bits_elementValid_lo = {indexDeq_bits_elementValid_lo_hi, indexDeq_bits_elementValid_lo_lo};
  wire [1:0]  indexDeq_bits_elementValid_hi_lo_lo_lo = {indexVec_17_5, indexVec_16_5};
  wire [1:0]  indexDeq_bits_elementValid_hi_lo_lo_hi = {indexVec_19_5, indexVec_18_5};
  wire [3:0]  indexDeq_bits_elementValid_hi_lo_lo = {indexDeq_bits_elementValid_hi_lo_lo_hi, indexDeq_bits_elementValid_hi_lo_lo_lo};
  wire [1:0]  indexDeq_bits_elementValid_hi_lo_hi_lo = {indexVec_21_5, indexVec_20_5};
  wire [1:0]  indexDeq_bits_elementValid_hi_lo_hi_hi = {indexVec_23_5, indexVec_22_5};
  wire [3:0]  indexDeq_bits_elementValid_hi_lo_hi = {indexDeq_bits_elementValid_hi_lo_hi_hi, indexDeq_bits_elementValid_hi_lo_hi_lo};
  wire [7:0]  indexDeq_bits_elementValid_hi_lo = {indexDeq_bits_elementValid_hi_lo_hi, indexDeq_bits_elementValid_hi_lo_lo};
  wire [1:0]  indexDeq_bits_elementValid_hi_hi_lo_lo = {indexVec_25_5, indexVec_24_5};
  wire [1:0]  indexDeq_bits_elementValid_hi_hi_lo_hi = {indexVec_27_5, indexVec_26_5};
  wire [3:0]  indexDeq_bits_elementValid_hi_hi_lo = {indexDeq_bits_elementValid_hi_hi_lo_hi, indexDeq_bits_elementValid_hi_hi_lo_lo};
  wire [1:0]  indexDeq_bits_elementValid_hi_hi_hi_lo = {indexVec_29_5, indexVec_28_5};
  wire [1:0]  indexDeq_bits_elementValid_hi_hi_hi_hi = {indexVec_31_5, indexVec_30_5};
  wire [3:0]  indexDeq_bits_elementValid_hi_hi_hi = {indexDeq_bits_elementValid_hi_hi_hi_hi, indexDeq_bits_elementValid_hi_hi_hi_lo};
  wire [7:0]  indexDeq_bits_elementValid_hi_hi = {indexDeq_bits_elementValid_hi_hi_hi, indexDeq_bits_elementValid_hi_hi_lo};
  wire [15:0] indexDeq_bits_elementValid_hi = {indexDeq_bits_elementValid_hi_hi, indexDeq_bits_elementValid_hi_lo};
  wire [31:0] indexDeq_bits_elementValid_0 = {indexDeq_bits_elementValid_hi, indexDeq_bits_elementValid_lo} | replaceWithVs1;
  wire [1:0]  indexDeq_bits_readOffset_lo_lo_lo_lo = {indexVec_1_2, indexVec_0_2};
  wire [1:0]  indexDeq_bits_readOffset_lo_lo_lo_hi = {indexVec_3_2, indexVec_2_2};
  wire [3:0]  indexDeq_bits_readOffset_lo_lo_lo = {indexDeq_bits_readOffset_lo_lo_lo_hi, indexDeq_bits_readOffset_lo_lo_lo_lo};
  wire [1:0]  indexDeq_bits_readOffset_lo_lo_hi_lo = {indexVec_5_2, indexVec_4_2};
  wire [1:0]  indexDeq_bits_readOffset_lo_lo_hi_hi = {indexVec_7_2, indexVec_6_2};
  wire [3:0]  indexDeq_bits_readOffset_lo_lo_hi = {indexDeq_bits_readOffset_lo_lo_hi_hi, indexDeq_bits_readOffset_lo_lo_hi_lo};
  wire [7:0]  indexDeq_bits_readOffset_lo_lo = {indexDeq_bits_readOffset_lo_lo_hi, indexDeq_bits_readOffset_lo_lo_lo};
  wire [1:0]  indexDeq_bits_readOffset_lo_hi_lo_lo = {indexVec_9_2, indexVec_8_2};
  wire [1:0]  indexDeq_bits_readOffset_lo_hi_lo_hi = {indexVec_11_2, indexVec_10_2};
  wire [3:0]  indexDeq_bits_readOffset_lo_hi_lo = {indexDeq_bits_readOffset_lo_hi_lo_hi, indexDeq_bits_readOffset_lo_hi_lo_lo};
  wire [1:0]  indexDeq_bits_readOffset_lo_hi_hi_lo = {indexVec_13_2, indexVec_12_2};
  wire [1:0]  indexDeq_bits_readOffset_lo_hi_hi_hi = {indexVec_15_2, indexVec_14_2};
  wire [3:0]  indexDeq_bits_readOffset_lo_hi_hi = {indexDeq_bits_readOffset_lo_hi_hi_hi, indexDeq_bits_readOffset_lo_hi_hi_lo};
  wire [7:0]  indexDeq_bits_readOffset_lo_hi = {indexDeq_bits_readOffset_lo_hi_hi, indexDeq_bits_readOffset_lo_hi_lo};
  wire [15:0] indexDeq_bits_readOffset_lo = {indexDeq_bits_readOffset_lo_hi, indexDeq_bits_readOffset_lo_lo};
  wire [1:0]  indexDeq_bits_readOffset_hi_lo_lo_lo = {indexVec_17_2, indexVec_16_2};
  wire [1:0]  indexDeq_bits_readOffset_hi_lo_lo_hi = {indexVec_19_2, indexVec_18_2};
  wire [3:0]  indexDeq_bits_readOffset_hi_lo_lo = {indexDeq_bits_readOffset_hi_lo_lo_hi, indexDeq_bits_readOffset_hi_lo_lo_lo};
  wire [1:0]  indexDeq_bits_readOffset_hi_lo_hi_lo = {indexVec_21_2, indexVec_20_2};
  wire [1:0]  indexDeq_bits_readOffset_hi_lo_hi_hi = {indexVec_23_2, indexVec_22_2};
  wire [3:0]  indexDeq_bits_readOffset_hi_lo_hi = {indexDeq_bits_readOffset_hi_lo_hi_hi, indexDeq_bits_readOffset_hi_lo_hi_lo};
  wire [7:0]  indexDeq_bits_readOffset_hi_lo = {indexDeq_bits_readOffset_hi_lo_hi, indexDeq_bits_readOffset_hi_lo_lo};
  wire [1:0]  indexDeq_bits_readOffset_hi_hi_lo_lo = {indexVec_25_2, indexVec_24_2};
  wire [1:0]  indexDeq_bits_readOffset_hi_hi_lo_hi = {indexVec_27_2, indexVec_26_2};
  wire [3:0]  indexDeq_bits_readOffset_hi_hi_lo = {indexDeq_bits_readOffset_hi_hi_lo_hi, indexDeq_bits_readOffset_hi_hi_lo_lo};
  wire [1:0]  indexDeq_bits_readOffset_hi_hi_hi_lo = {indexVec_29_2, indexVec_28_2};
  wire [1:0]  indexDeq_bits_readOffset_hi_hi_hi_hi = {indexVec_31_2, indexVec_30_2};
  wire [3:0]  indexDeq_bits_readOffset_hi_hi_hi = {indexDeq_bits_readOffset_hi_hi_hi_hi, indexDeq_bits_readOffset_hi_hi_hi_lo};
  wire [7:0]  indexDeq_bits_readOffset_hi_hi = {indexDeq_bits_readOffset_hi_hi_hi, indexDeq_bits_readOffset_hi_hi_lo};
  wire [15:0] indexDeq_bits_readOffset_hi = {indexDeq_bits_readOffset_hi_hi, indexDeq_bits_readOffset_hi_lo};
  wire [31:0] indexDeq_bits_readOffset_0 = {indexDeq_bits_readOffset_hi, indexDeq_bits_readOffset_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_lo_lo_lo = {indexVec_1_0, indexVec_0_0};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_lo_lo_hi = {indexVec_3_0, indexVec_2_0};
  wire [7:0]  indexDeq_bits_readDataOffset_lo_lo_lo = {indexDeq_bits_readDataOffset_lo_lo_lo_hi, indexDeq_bits_readDataOffset_lo_lo_lo_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_lo_hi_lo = {indexVec_5_0, indexVec_4_0};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_lo_hi_hi = {indexVec_7_0, indexVec_6_0};
  wire [7:0]  indexDeq_bits_readDataOffset_lo_lo_hi = {indexDeq_bits_readDataOffset_lo_lo_hi_hi, indexDeq_bits_readDataOffset_lo_lo_hi_lo};
  wire [15:0] indexDeq_bits_readDataOffset_lo_lo = {indexDeq_bits_readDataOffset_lo_lo_hi, indexDeq_bits_readDataOffset_lo_lo_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_hi_lo_lo = {indexVec_9_0, indexVec_8_0};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_hi_lo_hi = {indexVec_11_0, indexVec_10_0};
  wire [7:0]  indexDeq_bits_readDataOffset_lo_hi_lo = {indexDeq_bits_readDataOffset_lo_hi_lo_hi, indexDeq_bits_readDataOffset_lo_hi_lo_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_hi_hi_lo = {indexVec_13_0, indexVec_12_0};
  wire [3:0]  indexDeq_bits_readDataOffset_lo_hi_hi_hi = {indexVec_15_0, indexVec_14_0};
  wire [7:0]  indexDeq_bits_readDataOffset_lo_hi_hi = {indexDeq_bits_readDataOffset_lo_hi_hi_hi, indexDeq_bits_readDataOffset_lo_hi_hi_lo};
  wire [15:0] indexDeq_bits_readDataOffset_lo_hi = {indexDeq_bits_readDataOffset_lo_hi_hi, indexDeq_bits_readDataOffset_lo_hi_lo};
  wire [31:0] indexDeq_bits_readDataOffset_lo = {indexDeq_bits_readDataOffset_lo_hi, indexDeq_bits_readDataOffset_lo_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_lo_lo_lo = {indexVec_17_0, indexVec_16_0};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_lo_lo_hi = {indexVec_19_0, indexVec_18_0};
  wire [7:0]  indexDeq_bits_readDataOffset_hi_lo_lo = {indexDeq_bits_readDataOffset_hi_lo_lo_hi, indexDeq_bits_readDataOffset_hi_lo_lo_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_lo_hi_lo = {indexVec_21_0, indexVec_20_0};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_lo_hi_hi = {indexVec_23_0, indexVec_22_0};
  wire [7:0]  indexDeq_bits_readDataOffset_hi_lo_hi = {indexDeq_bits_readDataOffset_hi_lo_hi_hi, indexDeq_bits_readDataOffset_hi_lo_hi_lo};
  wire [15:0] indexDeq_bits_readDataOffset_hi_lo = {indexDeq_bits_readDataOffset_hi_lo_hi, indexDeq_bits_readDataOffset_hi_lo_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_hi_lo_lo = {indexVec_25_0, indexVec_24_0};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_hi_lo_hi = {indexVec_27_0, indexVec_26_0};
  wire [7:0]  indexDeq_bits_readDataOffset_hi_hi_lo = {indexDeq_bits_readDataOffset_hi_hi_lo_hi, indexDeq_bits_readDataOffset_hi_hi_lo_lo};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_hi_hi_lo = {indexVec_29_0, indexVec_28_0};
  wire [3:0]  indexDeq_bits_readDataOffset_hi_hi_hi_hi = {indexVec_31_0, indexVec_30_0};
  wire [7:0]  indexDeq_bits_readDataOffset_hi_hi_hi = {indexDeq_bits_readDataOffset_hi_hi_hi_hi, indexDeq_bits_readDataOffset_hi_hi_hi_lo};
  wire [15:0] indexDeq_bits_readDataOffset_hi_hi = {indexDeq_bits_readDataOffset_hi_hi_hi, indexDeq_bits_readDataOffset_hi_hi_lo};
  wire [31:0] indexDeq_bits_readDataOffset_hi = {indexDeq_bits_readDataOffset_hi_hi, indexDeq_bits_readDataOffset_hi_lo};
  wire [63:0] indexDeq_bits_readDataOffset_0 = {indexDeq_bits_readDataOffset_hi, indexDeq_bits_readDataOffset_lo};
  always @(posedge clock) begin
    if (reset) begin
      InstructionValid <= 1'h0;
      slideGroup <= 7'h0;
    end
    else begin
      if (newInstruction | lastFire)
        InstructionValid <= newInstruction;
      if (newInstruction | _lastFire_T_1)
        slideGroup <= newInstruction ? 7'h0 : slideGroup + 7'h1;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:0];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        _RANDOM[/*Zero width*/ 1'b0] = `RANDOM;
        InstructionValid = _RANDOM[/*Zero width*/ 1'b0][0];
        slideGroup = _RANDOM[/*Zero width*/ 1'b0][7:1];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  assign indexDeq_valid = indexDeq_valid_0;
  assign indexDeq_bits_needRead = indexDeq_bits_needRead_0;
  assign indexDeq_bits_elementValid = indexDeq_bits_elementValid_0;
  assign indexDeq_bits_replaceVs1 = indexDeq_bits_replaceVs1_0;
  assign indexDeq_bits_readOffset = indexDeq_bits_readOffset_0;
  assign indexDeq_bits_accessLane_0 = indexDeq_bits_accessLane_0_0;
  assign indexDeq_bits_accessLane_1 = indexDeq_bits_accessLane_1_0;
  assign indexDeq_bits_accessLane_2 = indexDeq_bits_accessLane_2_0;
  assign indexDeq_bits_accessLane_3 = indexDeq_bits_accessLane_3_0;
  assign indexDeq_bits_accessLane_4 = indexDeq_bits_accessLane_4_0;
  assign indexDeq_bits_accessLane_5 = indexDeq_bits_accessLane_5_0;
  assign indexDeq_bits_accessLane_6 = indexDeq_bits_accessLane_6_0;
  assign indexDeq_bits_accessLane_7 = indexDeq_bits_accessLane_7_0;
  assign indexDeq_bits_accessLane_8 = indexDeq_bits_accessLane_8_0;
  assign indexDeq_bits_accessLane_9 = indexDeq_bits_accessLane_9_0;
  assign indexDeq_bits_accessLane_10 = indexDeq_bits_accessLane_10_0;
  assign indexDeq_bits_accessLane_11 = indexDeq_bits_accessLane_11_0;
  assign indexDeq_bits_accessLane_12 = indexDeq_bits_accessLane_12_0;
  assign indexDeq_bits_accessLane_13 = indexDeq_bits_accessLane_13_0;
  assign indexDeq_bits_accessLane_14 = indexDeq_bits_accessLane_14_0;
  assign indexDeq_bits_accessLane_15 = indexDeq_bits_accessLane_15_0;
  assign indexDeq_bits_accessLane_16 = indexDeq_bits_accessLane_16_0;
  assign indexDeq_bits_accessLane_17 = indexDeq_bits_accessLane_17_0;
  assign indexDeq_bits_accessLane_18 = indexDeq_bits_accessLane_18_0;
  assign indexDeq_bits_accessLane_19 = indexDeq_bits_accessLane_19_0;
  assign indexDeq_bits_accessLane_20 = indexDeq_bits_accessLane_20_0;
  assign indexDeq_bits_accessLane_21 = indexDeq_bits_accessLane_21_0;
  assign indexDeq_bits_accessLane_22 = indexDeq_bits_accessLane_22_0;
  assign indexDeq_bits_accessLane_23 = indexDeq_bits_accessLane_23_0;
  assign indexDeq_bits_accessLane_24 = indexDeq_bits_accessLane_24_0;
  assign indexDeq_bits_accessLane_25 = indexDeq_bits_accessLane_25_0;
  assign indexDeq_bits_accessLane_26 = indexDeq_bits_accessLane_26_0;
  assign indexDeq_bits_accessLane_27 = indexDeq_bits_accessLane_27_0;
  assign indexDeq_bits_accessLane_28 = indexDeq_bits_accessLane_28_0;
  assign indexDeq_bits_accessLane_29 = indexDeq_bits_accessLane_29_0;
  assign indexDeq_bits_accessLane_30 = indexDeq_bits_accessLane_30_0;
  assign indexDeq_bits_accessLane_31 = indexDeq_bits_accessLane_31_0;
  assign indexDeq_bits_vsGrowth_0 = indexDeq_bits_vsGrowth_0_0;
  assign indexDeq_bits_vsGrowth_1 = indexDeq_bits_vsGrowth_1_0;
  assign indexDeq_bits_vsGrowth_2 = indexDeq_bits_vsGrowth_2_0;
  assign indexDeq_bits_vsGrowth_3 = indexDeq_bits_vsGrowth_3_0;
  assign indexDeq_bits_vsGrowth_4 = indexDeq_bits_vsGrowth_4_0;
  assign indexDeq_bits_vsGrowth_5 = indexDeq_bits_vsGrowth_5_0;
  assign indexDeq_bits_vsGrowth_6 = indexDeq_bits_vsGrowth_6_0;
  assign indexDeq_bits_vsGrowth_7 = indexDeq_bits_vsGrowth_7_0;
  assign indexDeq_bits_vsGrowth_8 = indexDeq_bits_vsGrowth_8_0;
  assign indexDeq_bits_vsGrowth_9 = indexDeq_bits_vsGrowth_9_0;
  assign indexDeq_bits_vsGrowth_10 = indexDeq_bits_vsGrowth_10_0;
  assign indexDeq_bits_vsGrowth_11 = indexDeq_bits_vsGrowth_11_0;
  assign indexDeq_bits_vsGrowth_12 = indexDeq_bits_vsGrowth_12_0;
  assign indexDeq_bits_vsGrowth_13 = indexDeq_bits_vsGrowth_13_0;
  assign indexDeq_bits_vsGrowth_14 = indexDeq_bits_vsGrowth_14_0;
  assign indexDeq_bits_vsGrowth_15 = indexDeq_bits_vsGrowth_15_0;
  assign indexDeq_bits_vsGrowth_16 = indexDeq_bits_vsGrowth_16_0;
  assign indexDeq_bits_vsGrowth_17 = indexDeq_bits_vsGrowth_17_0;
  assign indexDeq_bits_vsGrowth_18 = indexDeq_bits_vsGrowth_18_0;
  assign indexDeq_bits_vsGrowth_19 = indexDeq_bits_vsGrowth_19_0;
  assign indexDeq_bits_vsGrowth_20 = indexDeq_bits_vsGrowth_20_0;
  assign indexDeq_bits_vsGrowth_21 = indexDeq_bits_vsGrowth_21_0;
  assign indexDeq_bits_vsGrowth_22 = indexDeq_bits_vsGrowth_22_0;
  assign indexDeq_bits_vsGrowth_23 = indexDeq_bits_vsGrowth_23_0;
  assign indexDeq_bits_vsGrowth_24 = indexDeq_bits_vsGrowth_24_0;
  assign indexDeq_bits_vsGrowth_25 = indexDeq_bits_vsGrowth_25_0;
  assign indexDeq_bits_vsGrowth_26 = indexDeq_bits_vsGrowth_26_0;
  assign indexDeq_bits_vsGrowth_27 = indexDeq_bits_vsGrowth_27_0;
  assign indexDeq_bits_vsGrowth_28 = indexDeq_bits_vsGrowth_28_0;
  assign indexDeq_bits_vsGrowth_29 = indexDeq_bits_vsGrowth_29_0;
  assign indexDeq_bits_vsGrowth_30 = indexDeq_bits_vsGrowth_30_0;
  assign indexDeq_bits_vsGrowth_31 = indexDeq_bits_vsGrowth_31_0;
  assign indexDeq_bits_executeGroup = indexDeq_bits_executeGroup_0;
  assign indexDeq_bits_readDataOffset = indexDeq_bits_readDataOffset_0;
  assign indexDeq_bits_last = indexDeq_bits_last_0;
  assign slideGroupOut = slideGroup;
endmodule

