
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module MaskUnit(
  input         clock,
                reset,
                instReq_valid,
  input  [2:0]  instReq_bits_instructionIndex,
  input         instReq_bits_decodeResult_specialSlot,
  input  [4:0]  instReq_bits_decodeResult_topUop,
  input         instReq_bits_decodeResult_popCount,
                instReq_bits_decodeResult_ffo,
                instReq_bits_decodeResult_average,
                instReq_bits_decodeResult_reverse,
                instReq_bits_decodeResult_dontNeedExecuteInLane,
                instReq_bits_decodeResult_scheduler,
                instReq_bits_decodeResult_sReadVD,
                instReq_bits_decodeResult_vtype,
                instReq_bits_decodeResult_sWrite,
                instReq_bits_decodeResult_crossRead,
                instReq_bits_decodeResult_crossWrite,
                instReq_bits_decodeResult_maskUnit,
                instReq_bits_decodeResult_special,
                instReq_bits_decodeResult_saturate,
                instReq_bits_decodeResult_vwmacc,
                instReq_bits_decodeResult_readOnly,
                instReq_bits_decodeResult_maskSource,
                instReq_bits_decodeResult_maskDestination,
                instReq_bits_decodeResult_maskLogic,
  input  [3:0]  instReq_bits_decodeResult_uop,
  input         instReq_bits_decodeResult_iota,
                instReq_bits_decodeResult_mv,
                instReq_bits_decodeResult_extend,
                instReq_bits_decodeResult_unOrderWrite,
                instReq_bits_decodeResult_compress,
                instReq_bits_decodeResult_gather16,
                instReq_bits_decodeResult_gather,
                instReq_bits_decodeResult_slid,
                instReq_bits_decodeResult_targetRd,
                instReq_bits_decodeResult_widenReduce,
                instReq_bits_decodeResult_red,
                instReq_bits_decodeResult_nr,
                instReq_bits_decodeResult_itype,
                instReq_bits_decodeResult_unsigned1,
                instReq_bits_decodeResult_unsigned0,
                instReq_bits_decodeResult_other,
                instReq_bits_decodeResult_multiCycle,
                instReq_bits_decodeResult_divider,
                instReq_bits_decodeResult_multiplier,
                instReq_bits_decodeResult_shift,
                instReq_bits_decodeResult_adder,
                instReq_bits_decodeResult_logic,
  input  [31:0] instReq_bits_readFromScala,
  input  [1:0]  instReq_bits_sew,
  input  [2:0]  instReq_bits_vlmul,
  input         instReq_bits_maskType,
  input  [2:0]  instReq_bits_vxrm,
  input  [4:0]  instReq_bits_vs2,
                instReq_bits_vs1,
                instReq_bits_vd,
  input  [11:0] instReq_bits_vl,
  input         exeReq_0_valid,
  input  [31:0] exeReq_0_bits_source1,
                exeReq_0_bits_source2,
  input  [2:0]  exeReq_0_bits_index,
  input         exeReq_0_bits_ffo,
                exeReq_1_valid,
  input  [31:0] exeReq_1_bits_source1,
                exeReq_1_bits_source2,
  input  [2:0]  exeReq_1_bits_index,
  input         exeReq_1_bits_ffo,
                exeReq_2_valid,
  input  [31:0] exeReq_2_bits_source1,
                exeReq_2_bits_source2,
  input  [2:0]  exeReq_2_bits_index,
  input         exeReq_2_bits_ffo,
                exeReq_3_valid,
  input  [31:0] exeReq_3_bits_source1,
                exeReq_3_bits_source2,
  input  [2:0]  exeReq_3_bits_index,
  input         exeReq_3_bits_ffo,
                exeResp_0_ready,
  output        exeResp_0_valid,
  output [4:0]  exeResp_0_bits_vd,
  output [3:0]  exeResp_0_bits_offset,
                exeResp_0_bits_mask,
  output [31:0] exeResp_0_bits_data,
  output [2:0]  exeResp_0_bits_instructionIndex,
  input         exeResp_1_ready,
  output        exeResp_1_valid,
  output [4:0]  exeResp_1_bits_vd,
  output [3:0]  exeResp_1_bits_offset,
                exeResp_1_bits_mask,
  output [31:0] exeResp_1_bits_data,
  output [2:0]  exeResp_1_bits_instructionIndex,
  input         exeResp_2_ready,
  output        exeResp_2_valid,
  output [4:0]  exeResp_2_bits_vd,
  output [3:0]  exeResp_2_bits_offset,
                exeResp_2_bits_mask,
  output [31:0] exeResp_2_bits_data,
  output [2:0]  exeResp_2_bits_instructionIndex,
  input         exeResp_3_ready,
  output        exeResp_3_valid,
  output [4:0]  exeResp_3_bits_vd,
  output [3:0]  exeResp_3_bits_offset,
                exeResp_3_bits_mask,
  output [31:0] exeResp_3_bits_data,
  output [2:0]  exeResp_3_bits_instructionIndex,
  input         writeRelease_0,
                writeRelease_1,
                writeRelease_2,
                writeRelease_3,
  output        tokenIO_0_maskRequestRelease,
                tokenIO_1_maskRequestRelease,
                tokenIO_2_maskRequestRelease,
                tokenIO_3_maskRequestRelease,
  input         readChannel_0_ready,
  output        readChannel_0_valid,
  output [4:0]  readChannel_0_bits_vs,
  output [3:0]  readChannel_0_bits_offset,
  output [2:0]  readChannel_0_bits_instructionIndex,
  input         readChannel_1_ready,
  output        readChannel_1_valid,
  output [4:0]  readChannel_1_bits_vs,
  output [3:0]  readChannel_1_bits_offset,
  output [2:0]  readChannel_1_bits_instructionIndex,
  input         readChannel_2_ready,
  output        readChannel_2_valid,
  output [4:0]  readChannel_2_bits_vs,
  output [3:0]  readChannel_2_bits_offset,
  output [2:0]  readChannel_2_bits_instructionIndex,
  input         readChannel_3_ready,
  output        readChannel_3_valid,
  output [4:0]  readChannel_3_bits_vs,
  output [3:0]  readChannel_3_bits_offset,
  output [2:0]  readChannel_3_bits_instructionIndex,
  input         readResult_0_valid,
  input  [31:0] readResult_0_bits,
  input         readResult_1_valid,
  input  [31:0] readResult_1_bits,
  input         readResult_2_valid,
  input  [31:0] readResult_2_bits,
  input         readResult_3_valid,
  input  [31:0] readResult_3_bits,
  output [7:0]  lastReport,
  output [31:0] laneMaskInput_0,
                laneMaskInput_1,
                laneMaskInput_2,
                laneMaskInput_3,
  input  [5:0]  laneMaskSelect_0,
                laneMaskSelect_1,
                laneMaskSelect_2,
                laneMaskSelect_3,
  input  [1:0]  laneMaskSewSelect_0,
                laneMaskSewSelect_1,
                laneMaskSewSelect_2,
                laneMaskSewSelect_3,
  input         v0UpdateVec_0_valid,
  input  [31:0] v0UpdateVec_0_bits_data,
  input  [3:0]  v0UpdateVec_0_bits_offset,
                v0UpdateVec_0_bits_mask,
  input         v0UpdateVec_1_valid,
  input  [31:0] v0UpdateVec_1_bits_data,
  input  [3:0]  v0UpdateVec_1_bits_offset,
                v0UpdateVec_1_bits_mask,
  input         v0UpdateVec_2_valid,
  input  [31:0] v0UpdateVec_2_bits_data,
  input  [3:0]  v0UpdateVec_2_bits_offset,
                v0UpdateVec_2_bits_mask,
  input         v0UpdateVec_3_valid,
  input  [31:0] v0UpdateVec_3_bits_data,
  input  [3:0]  v0UpdateVec_3_bits_offset,
                v0UpdateVec_3_bits_mask,
  output [31:0] writeRDData,
  input         gatherData_ready,
  output        gatherData_valid,
  output [31:0] gatherData_bits,
  input         gatherRead
);

  wire               readCrossBar_input_3_valid;
  wire               readCrossBar_input_2_valid;
  wire               readCrossBar_input_1_valid;
  wire               readCrossBar_input_0_valid;
  wire               _writeQueue_fifo_3_empty;
  wire               _writeQueue_fifo_3_full;
  wire               _writeQueue_fifo_3_error;
  wire [52:0]        _writeQueue_fifo_3_data_out;
  wire               _writeQueue_fifo_2_empty;
  wire               _writeQueue_fifo_2_full;
  wire               _writeQueue_fifo_2_error;
  wire [52:0]        _writeQueue_fifo_2_data_out;
  wire               _writeQueue_fifo_1_empty;
  wire               _writeQueue_fifo_1_full;
  wire               _writeQueue_fifo_1_error;
  wire [52:0]        _writeQueue_fifo_1_data_out;
  wire               _writeQueue_fifo_empty;
  wire               _writeQueue_fifo_full;
  wire               _writeQueue_fifo_error;
  wire [52:0]        _writeQueue_fifo_data_out;
  wire [127:0]       _extendUnit_out;
  wire               _reduceUnit_in_ready;
  wire               _reduceUnit_out_valid;
  wire [31:0]        _reduceUnit_out_bits_data;
  wire [3:0]         _reduceUnit_out_bits_mask;
  wire               _compressUnit_out_compressValid;
  wire [31:0]        _compressUnit_writeData;
  wire               _compressUnit_stageValid;
  wire               _readData_readDataQueue_fifo_3_empty;
  wire               _readData_readDataQueue_fifo_3_full;
  wire               _readData_readDataQueue_fifo_3_error;
  wire [31:0]        _readData_readDataQueue_fifo_3_data_out;
  wire               _readData_readDataQueue_fifo_2_empty;
  wire               _readData_readDataQueue_fifo_2_full;
  wire               _readData_readDataQueue_fifo_2_error;
  wire [31:0]        _readData_readDataQueue_fifo_2_data_out;
  wire               _readData_readDataQueue_fifo_1_empty;
  wire               _readData_readDataQueue_fifo_1_full;
  wire               _readData_readDataQueue_fifo_1_error;
  wire [31:0]        _readData_readDataQueue_fifo_1_data_out;
  wire               _readData_readDataQueue_fifo_empty;
  wire               _readData_readDataQueue_fifo_full;
  wire               _readData_readDataQueue_fifo_error;
  wire [31:0]        _readData_readDataQueue_fifo_data_out;
  wire               _readMessageQueue_fifo_3_empty;
  wire               _readMessageQueue_fifo_3_full;
  wire               _readMessageQueue_fifo_3_error;
  wire [5:0]         _readMessageQueue_fifo_3_data_out;
  wire               _readMessageQueue_fifo_2_empty;
  wire               _readMessageQueue_fifo_2_full;
  wire               _readMessageQueue_fifo_2_error;
  wire [5:0]         _readMessageQueue_fifo_2_data_out;
  wire               _readMessageQueue_fifo_1_empty;
  wire               _readMessageQueue_fifo_1_full;
  wire               _readMessageQueue_fifo_1_error;
  wire [5:0]         _readMessageQueue_fifo_1_data_out;
  wire               _readMessageQueue_fifo_empty;
  wire               _readMessageQueue_fifo_full;
  wire               _readMessageQueue_fifo_error;
  wire [5:0]         _readMessageQueue_fifo_data_out;
  wire               _reorderQueueVec_fifo_3_empty;
  wire               _reorderQueueVec_fifo_3_full;
  wire               _reorderQueueVec_fifo_3_error;
  wire [35:0]        _reorderQueueVec_fifo_3_data_out;
  wire               _reorderQueueVec_fifo_2_empty;
  wire               _reorderQueueVec_fifo_2_full;
  wire               _reorderQueueVec_fifo_2_error;
  wire [35:0]        _reorderQueueVec_fifo_2_data_out;
  wire               _reorderQueueVec_fifo_1_empty;
  wire               _reorderQueueVec_fifo_1_full;
  wire               _reorderQueueVec_fifo_1_error;
  wire [35:0]        _reorderQueueVec_fifo_1_data_out;
  wire               _reorderQueueVec_fifo_empty;
  wire               _reorderQueueVec_fifo_full;
  wire               _reorderQueueVec_fifo_error;
  wire [35:0]        _reorderQueueVec_fifo_data_out;
  wire               _compressUnitResultQueue_fifo_empty;
  wire               _compressUnitResultQueue_fifo_full;
  wire               _compressUnitResultQueue_fifo_error;
  wire [156:0]       _compressUnitResultQueue_fifo_data_out;
  wire               _readWaitQueue_fifo_empty;
  wire               _readWaitQueue_fifo_full;
  wire               _readWaitQueue_fifo_error;
  wire [22:0]        _readWaitQueue_fifo_data_out;
  wire               _readCrossBar_input_0_ready;
  wire               _readCrossBar_input_1_ready;
  wire               _readCrossBar_input_2_ready;
  wire               _readCrossBar_input_3_ready;
  wire               _readCrossBar_output_0_valid;
  wire [4:0]         _readCrossBar_output_0_bits_vs;
  wire [3:0]         _readCrossBar_output_0_bits_offset;
  wire [1:0]         _readCrossBar_output_0_bits_writeIndex;
  wire               _readCrossBar_output_1_valid;
  wire [4:0]         _readCrossBar_output_1_bits_vs;
  wire [3:0]         _readCrossBar_output_1_bits_offset;
  wire [1:0]         _readCrossBar_output_1_bits_writeIndex;
  wire               _readCrossBar_output_2_valid;
  wire [4:0]         _readCrossBar_output_2_bits_vs;
  wire [3:0]         _readCrossBar_output_2_bits_offset;
  wire [1:0]         _readCrossBar_output_2_bits_writeIndex;
  wire               _readCrossBar_output_3_valid;
  wire [4:0]         _readCrossBar_output_3_bits_vs;
  wire [3:0]         _readCrossBar_output_3_bits_offset;
  wire [1:0]         _readCrossBar_output_3_bits_writeIndex;
  wire               _accessCountQueue_fifo_empty;
  wire               _accessCountQueue_fifo_full;
  wire               _accessCountQueue_fifo_error;
  wire [11:0]        _accessCountQueue_fifo_data_out;
  wire               _slideAddressGen_indexDeq_valid;
  wire [3:0]         _slideAddressGen_indexDeq_bits_needRead;
  wire [3:0]         _slideAddressGen_indexDeq_bits_elementValid;
  wire [3:0]         _slideAddressGen_indexDeq_bits_replaceVs1;
  wire [15:0]        _slideAddressGen_indexDeq_bits_readOffset;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_0;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_1;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_2;
  wire [1:0]         _slideAddressGen_indexDeq_bits_accessLane_3;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_0;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_1;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_2;
  wire [2:0]         _slideAddressGen_indexDeq_bits_vsGrowth_3;
  wire [9:0]         _slideAddressGen_indexDeq_bits_executeGroup;
  wire [7:0]         _slideAddressGen_indexDeq_bits_readDataOffset;
  wire               _slideAddressGen_indexDeq_bits_last;
  wire [9:0]         _slideAddressGen_slideGroupOut;
  wire               _exeRequestQueue_queue_fifo_3_empty;
  wire               _exeRequestQueue_queue_fifo_3_full;
  wire               _exeRequestQueue_queue_fifo_3_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_3_data_out;
  wire               _exeRequestQueue_queue_fifo_2_empty;
  wire               _exeRequestQueue_queue_fifo_2_full;
  wire               _exeRequestQueue_queue_fifo_2_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_2_data_out;
  wire               _exeRequestQueue_queue_fifo_1_empty;
  wire               _exeRequestQueue_queue_fifo_1_full;
  wire               _exeRequestQueue_queue_fifo_1_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_1_data_out;
  wire               _exeRequestQueue_queue_fifo_empty;
  wire               _exeRequestQueue_queue_fifo_full;
  wire               _exeRequestQueue_queue_fifo_error;
  wire [67:0]        _exeRequestQueue_queue_fifo_data_out;
  wire               _maskedWrite_in_0_ready;
  wire               _maskedWrite_in_1_ready;
  wire               _maskedWrite_in_2_ready;
  wire               _maskedWrite_in_3_ready;
  wire               _maskedWrite_out_0_valid;
  wire               _maskedWrite_out_0_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_0_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_0_bits_writeData_mask;
  wire [7:0]         _maskedWrite_out_0_bits_writeData_groupCounter;
  wire               _maskedWrite_out_1_valid;
  wire               _maskedWrite_out_1_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_1_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_1_bits_writeData_mask;
  wire [7:0]         _maskedWrite_out_1_bits_writeData_groupCounter;
  wire               _maskedWrite_out_2_valid;
  wire               _maskedWrite_out_2_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_2_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_2_bits_writeData_mask;
  wire [7:0]         _maskedWrite_out_2_bits_writeData_groupCounter;
  wire               _maskedWrite_out_3_valid;
  wire               _maskedWrite_out_3_bits_ffoByOther;
  wire [31:0]        _maskedWrite_out_3_bits_writeData_data;
  wire [3:0]         _maskedWrite_out_3_bits_writeData_mask;
  wire [7:0]         _maskedWrite_out_3_bits_writeData_groupCounter;
  wire               _maskedWrite_readChannel_0_valid;
  wire [4:0]         _maskedWrite_readChannel_0_bits_vs;
  wire [3:0]         _maskedWrite_readChannel_0_bits_offset;
  wire               _maskedWrite_readChannel_1_valid;
  wire [4:0]         _maskedWrite_readChannel_1_bits_vs;
  wire [3:0]         _maskedWrite_readChannel_1_bits_offset;
  wire               _maskedWrite_readChannel_2_valid;
  wire [4:0]         _maskedWrite_readChannel_2_bits_vs;
  wire [3:0]         _maskedWrite_readChannel_2_bits_offset;
  wire               _maskedWrite_readChannel_3_valid;
  wire [4:0]         _maskedWrite_readChannel_3_bits_vs;
  wire [3:0]         _maskedWrite_readChannel_3_bits_offset;
  wire               _maskedWrite_stageClear;
  wire               writeQueue_3_almostFull;
  wire               writeQueue_3_almostEmpty;
  wire               writeQueue_2_almostFull;
  wire               writeQueue_2_almostEmpty;
  wire               writeQueue_1_almostFull;
  wire               writeQueue_1_almostEmpty;
  wire               writeQueue_0_almostFull;
  wire               writeQueue_0_almostEmpty;
  wire               readData_readDataQueue_3_almostFull;
  wire               readData_readDataQueue_3_almostEmpty;
  wire               readData_readDataQueue_2_almostFull;
  wire               readData_readDataQueue_2_almostEmpty;
  wire               readData_readDataQueue_1_almostFull;
  wire               readData_readDataQueue_1_almostEmpty;
  wire               readData_readDataQueue_almostFull;
  wire               readData_readDataQueue_almostEmpty;
  wire               readMessageQueue_3_almostFull;
  wire               readMessageQueue_3_almostEmpty;
  wire               readMessageQueue_2_almostFull;
  wire               readMessageQueue_2_almostEmpty;
  wire               readMessageQueue_1_almostFull;
  wire               readMessageQueue_1_almostEmpty;
  wire               readMessageQueue_almostFull;
  wire               readMessageQueue_almostEmpty;
  wire               reorderQueueVec_3_almostFull;
  wire               reorderQueueVec_3_almostEmpty;
  wire               reorderQueueVec_2_almostFull;
  wire               reorderQueueVec_2_almostEmpty;
  wire               reorderQueueVec_1_almostFull;
  wire               reorderQueueVec_1_almostEmpty;
  wire               reorderQueueVec_0_almostFull;
  wire               reorderQueueVec_0_almostEmpty;
  wire               compressUnitResultQueue_almostFull;
  wire               compressUnitResultQueue_almostEmpty;
  wire               readWaitQueue_almostFull;
  wire               readWaitQueue_almostEmpty;
  wire               accessCountQueue_almostFull;
  wire               accessCountQueue_almostEmpty;
  wire               exeRequestQueue_3_almostFull;
  wire               exeRequestQueue_3_almostEmpty;
  wire               exeRequestQueue_2_almostFull;
  wire               exeRequestQueue_2_almostEmpty;
  wire               exeRequestQueue_1_almostFull;
  wire               exeRequestQueue_1_almostEmpty;
  wire               exeRequestQueue_0_almostFull;
  wire               exeRequestQueue_0_almostEmpty;
  wire [31:0]        reorderQueueVec_3_deq_bits_data;
  wire [31:0]        reorderQueueVec_2_deq_bits_data;
  wire [31:0]        reorderQueueVec_1_deq_bits_data;
  wire [31:0]        reorderQueueVec_0_deq_bits_data;
  wire [2:0]         accessCountEnq_3;
  wire [2:0]         accessCountEnq_2;
  wire [2:0]         accessCountEnq_1;
  wire [2:0]         accessCountEnq_0;
  wire               exeResp_0_ready_0 = exeResp_0_ready;
  wire               exeResp_1_ready_0 = exeResp_1_ready;
  wire               exeResp_2_ready_0 = exeResp_2_ready;
  wire               exeResp_3_ready_0 = exeResp_3_ready;
  wire               readChannel_0_ready_0 = readChannel_0_ready;
  wire               readChannel_1_ready_0 = readChannel_1_ready;
  wire               readChannel_2_ready_0 = readChannel_2_ready;
  wire               readChannel_3_ready_0 = readChannel_3_ready;
  wire               gatherData_ready_0 = gatherData_ready;
  wire               exeRequestQueue_0_enq_valid = exeReq_0_valid;
  wire [31:0]        exeRequestQueue_0_enq_bits_source1 = exeReq_0_bits_source1;
  wire [31:0]        exeRequestQueue_0_enq_bits_source2 = exeReq_0_bits_source2;
  wire [2:0]         exeRequestQueue_0_enq_bits_index = exeReq_0_bits_index;
  wire               exeRequestQueue_0_enq_bits_ffo = exeReq_0_bits_ffo;
  wire               exeRequestQueue_1_enq_valid = exeReq_1_valid;
  wire [31:0]        exeRequestQueue_1_enq_bits_source1 = exeReq_1_bits_source1;
  wire [31:0]        exeRequestQueue_1_enq_bits_source2 = exeReq_1_bits_source2;
  wire [2:0]         exeRequestQueue_1_enq_bits_index = exeReq_1_bits_index;
  wire               exeRequestQueue_1_enq_bits_ffo = exeReq_1_bits_ffo;
  wire               exeRequestQueue_2_enq_valid = exeReq_2_valid;
  wire [31:0]        exeRequestQueue_2_enq_bits_source1 = exeReq_2_bits_source1;
  wire [31:0]        exeRequestQueue_2_enq_bits_source2 = exeReq_2_bits_source2;
  wire [2:0]         exeRequestQueue_2_enq_bits_index = exeReq_2_bits_index;
  wire               exeRequestQueue_2_enq_bits_ffo = exeReq_2_bits_ffo;
  wire               exeRequestQueue_3_enq_valid = exeReq_3_valid;
  wire [31:0]        exeRequestQueue_3_enq_bits_source1 = exeReq_3_bits_source1;
  wire [31:0]        exeRequestQueue_3_enq_bits_source2 = exeReq_3_bits_source2;
  wire [2:0]         exeRequestQueue_3_enq_bits_index = exeReq_3_bits_index;
  wire               exeRequestQueue_3_enq_bits_ffo = exeReq_3_bits_ffo;
  wire               reorderQueueVec_0_enq_valid = readResult_0_valid;
  wire               reorderQueueVec_1_enq_valid = readResult_1_valid;
  wire               reorderQueueVec_2_enq_valid = readResult_2_valid;
  wire               reorderQueueVec_3_enq_valid = readResult_3_valid;
  wire               readMessageQueue_deq_ready = readResult_0_valid;
  wire               readMessageQueue_1_deq_ready = readResult_1_valid;
  wire               readMessageQueue_2_deq_ready = readResult_2_valid;
  wire               readMessageQueue_3_deq_ready = readResult_3_valid;
  wire [7:0]         checkVec_checkResult_lo_14 = 8'hFF;
  wire [7:0]         checkVec_checkResult_hi_14 = 8'hFF;
  wire [15:0]        checkVec_2_0 = 16'hFFFF;
  wire [7:0]         checkVec_2_1 = 8'h0;
  wire [1:0]         readVS1Req_requestIndex = 2'h0;
  wire [1:0]         checkVec_checkResultVec_0_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_1_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_2_1_2 = 2'h0;
  wire [1:0]         checkVec_checkResultVec_3_1_2 = 2'h0;
  wire [1:0]         selectExecuteReq_0_bits_requestIndex = 2'h0;
  wire [1:0]         selectExecuteReq_1_bits_requestIndex = 2'h1;
  wire [1:0]         selectExecuteReq_3_bits_requestIndex = 2'h3;
  wire [3:0]         checkVec_checkResult_lo_15 = 4'h0;
  wire [3:0]         checkVec_checkResult_hi_15 = 4'h0;
  wire [1:0]         readChannel_0_bits_readSource = 2'h2;
  wire [1:0]         readChannel_1_bits_readSource = 2'h2;
  wire [1:0]         readChannel_2_bits_readSource = 2'h2;
  wire [1:0]         readChannel_3_bits_readSource = 2'h2;
  wire [1:0]         selectExecuteReq_2_bits_requestIndex = 2'h2;
  wire               exeResp_0_bits_last = 1'h0;
  wire               exeResp_1_bits_last = 1'h0;
  wire               exeResp_2_bits_last = 1'h0;
  wire               exeResp_3_bits_last = 1'h0;
  wire               writeRequest_0_ffoByOther = 1'h0;
  wire               writeRequest_1_ffoByOther = 1'h0;
  wire               writeRequest_2_ffoByOther = 1'h0;
  wire               writeRequest_3_ffoByOther = 1'h0;
  wire               writeQueue_0_deq_ready = exeResp_0_ready_0;
  wire               writeQueue_0_deq_valid;
  wire [3:0]         writeQueue_0_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_0_deq_bits_writeData_data;
  wire               writeQueue_1_deq_ready = exeResp_1_ready_0;
  wire               writeQueue_1_deq_valid;
  wire [3:0]         writeQueue_1_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_1_deq_bits_writeData_data;
  wire               writeQueue_2_deq_ready = exeResp_2_ready_0;
  wire               writeQueue_2_deq_valid;
  wire [3:0]         writeQueue_2_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_2_deq_bits_writeData_data;
  wire               writeQueue_3_deq_ready = exeResp_3_ready_0;
  wire               writeQueue_3_deq_valid;
  wire [3:0]         writeQueue_3_deq_bits_writeData_mask;
  wire [31:0]        writeQueue_3_deq_bits_writeData_data;
  wire               gatherResponse;
  reg  [31:0]        v0_0;
  reg  [31:0]        v0_1;
  reg  [31:0]        v0_2;
  reg  [31:0]        v0_3;
  reg  [31:0]        v0_4;
  reg  [31:0]        v0_5;
  reg  [31:0]        v0_6;
  reg  [31:0]        v0_7;
  reg  [31:0]        v0_8;
  reg  [31:0]        v0_9;
  reg  [31:0]        v0_10;
  reg  [31:0]        v0_11;
  reg  [31:0]        v0_12;
  reg  [31:0]        v0_13;
  reg  [31:0]        v0_14;
  reg  [31:0]        v0_15;
  reg  [31:0]        v0_16;
  reg  [31:0]        v0_17;
  reg  [31:0]        v0_18;
  reg  [31:0]        v0_19;
  reg  [31:0]        v0_20;
  reg  [31:0]        v0_21;
  reg  [31:0]        v0_22;
  reg  [31:0]        v0_23;
  reg  [31:0]        v0_24;
  reg  [31:0]        v0_25;
  reg  [31:0]        v0_26;
  reg  [31:0]        v0_27;
  reg  [31:0]        v0_28;
  reg  [31:0]        v0_29;
  reg  [31:0]        v0_30;
  reg  [31:0]        v0_31;
  reg  [31:0]        v0_32;
  reg  [31:0]        v0_33;
  reg  [31:0]        v0_34;
  reg  [31:0]        v0_35;
  reg  [31:0]        v0_36;
  reg  [31:0]        v0_37;
  reg  [31:0]        v0_38;
  reg  [31:0]        v0_39;
  reg  [31:0]        v0_40;
  reg  [31:0]        v0_41;
  reg  [31:0]        v0_42;
  reg  [31:0]        v0_43;
  reg  [31:0]        v0_44;
  reg  [31:0]        v0_45;
  reg  [31:0]        v0_46;
  reg  [31:0]        v0_47;
  reg  [31:0]        v0_48;
  reg  [31:0]        v0_49;
  reg  [31:0]        v0_50;
  reg  [31:0]        v0_51;
  reg  [31:0]        v0_52;
  reg  [31:0]        v0_53;
  reg  [31:0]        v0_54;
  reg  [31:0]        v0_55;
  reg  [31:0]        v0_56;
  reg  [31:0]        v0_57;
  reg  [31:0]        v0_58;
  reg  [31:0]        v0_59;
  reg  [31:0]        v0_60;
  reg  [31:0]        v0_61;
  reg  [31:0]        v0_62;
  reg  [31:0]        v0_63;
  wire [15:0]        maskExt_lo = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt = {maskExt_hi, maskExt_lo};
  wire [15:0]        maskExt_lo_1 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_1 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_1 = {maskExt_hi_1, maskExt_lo_1};
  wire [15:0]        maskExt_lo_2 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_2 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_2 = {maskExt_hi_2, maskExt_lo_2};
  wire [15:0]        maskExt_lo_3 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_3 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_3 = {maskExt_hi_3, maskExt_lo_3};
  wire [15:0]        maskExt_lo_4 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_4 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_4 = {maskExt_hi_4, maskExt_lo_4};
  wire [15:0]        maskExt_lo_5 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_5 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_5 = {maskExt_hi_5, maskExt_lo_5};
  wire [15:0]        maskExt_lo_6 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_6 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_6 = {maskExt_hi_6, maskExt_lo_6};
  wire [15:0]        maskExt_lo_7 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_7 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_7 = {maskExt_hi_7, maskExt_lo_7};
  wire [15:0]        maskExt_lo_8 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_8 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_8 = {maskExt_hi_8, maskExt_lo_8};
  wire [15:0]        maskExt_lo_9 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_9 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_9 = {maskExt_hi_9, maskExt_lo_9};
  wire [15:0]        maskExt_lo_10 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_10 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_10 = {maskExt_hi_10, maskExt_lo_10};
  wire [15:0]        maskExt_lo_11 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_11 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_11 = {maskExt_hi_11, maskExt_lo_11};
  wire [15:0]        maskExt_lo_12 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_12 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_12 = {maskExt_hi_12, maskExt_lo_12};
  wire [15:0]        maskExt_lo_13 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_13 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_13 = {maskExt_hi_13, maskExt_lo_13};
  wire [15:0]        maskExt_lo_14 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_14 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_14 = {maskExt_hi_14, maskExt_lo_14};
  wire [15:0]        maskExt_lo_15 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_15 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_15 = {maskExt_hi_15, maskExt_lo_15};
  wire [15:0]        maskExt_lo_16 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_16 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_16 = {maskExt_hi_16, maskExt_lo_16};
  wire [15:0]        maskExt_lo_17 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_17 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_17 = {maskExt_hi_17, maskExt_lo_17};
  wire [15:0]        maskExt_lo_18 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_18 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_18 = {maskExt_hi_18, maskExt_lo_18};
  wire [15:0]        maskExt_lo_19 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_19 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_19 = {maskExt_hi_19, maskExt_lo_19};
  wire [15:0]        maskExt_lo_20 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_20 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_20 = {maskExt_hi_20, maskExt_lo_20};
  wire [15:0]        maskExt_lo_21 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_21 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_21 = {maskExt_hi_21, maskExt_lo_21};
  wire [15:0]        maskExt_lo_22 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_22 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_22 = {maskExt_hi_22, maskExt_lo_22};
  wire [15:0]        maskExt_lo_23 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_23 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_23 = {maskExt_hi_23, maskExt_lo_23};
  wire [15:0]        maskExt_lo_24 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_24 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_24 = {maskExt_hi_24, maskExt_lo_24};
  wire [15:0]        maskExt_lo_25 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_25 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_25 = {maskExt_hi_25, maskExt_lo_25};
  wire [15:0]        maskExt_lo_26 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_26 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_26 = {maskExt_hi_26, maskExt_lo_26};
  wire [15:0]        maskExt_lo_27 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_27 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_27 = {maskExt_hi_27, maskExt_lo_27};
  wire [15:0]        maskExt_lo_28 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_28 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_28 = {maskExt_hi_28, maskExt_lo_28};
  wire [15:0]        maskExt_lo_29 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_29 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_29 = {maskExt_hi_29, maskExt_lo_29};
  wire [15:0]        maskExt_lo_30 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_30 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_30 = {maskExt_hi_30, maskExt_lo_30};
  wire [15:0]        maskExt_lo_31 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_31 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_31 = {maskExt_hi_31, maskExt_lo_31};
  wire [15:0]        maskExt_lo_32 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_32 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_32 = {maskExt_hi_32, maskExt_lo_32};
  wire [15:0]        maskExt_lo_33 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_33 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_33 = {maskExt_hi_33, maskExt_lo_33};
  wire [15:0]        maskExt_lo_34 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_34 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_34 = {maskExt_hi_34, maskExt_lo_34};
  wire [15:0]        maskExt_lo_35 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_35 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_35 = {maskExt_hi_35, maskExt_lo_35};
  wire [15:0]        maskExt_lo_36 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_36 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_36 = {maskExt_hi_36, maskExt_lo_36};
  wire [15:0]        maskExt_lo_37 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_37 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_37 = {maskExt_hi_37, maskExt_lo_37};
  wire [15:0]        maskExt_lo_38 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_38 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_38 = {maskExt_hi_38, maskExt_lo_38};
  wire [15:0]        maskExt_lo_39 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_39 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_39 = {maskExt_hi_39, maskExt_lo_39};
  wire [15:0]        maskExt_lo_40 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_40 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_40 = {maskExt_hi_40, maskExt_lo_40};
  wire [15:0]        maskExt_lo_41 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_41 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_41 = {maskExt_hi_41, maskExt_lo_41};
  wire [15:0]        maskExt_lo_42 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_42 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_42 = {maskExt_hi_42, maskExt_lo_42};
  wire [15:0]        maskExt_lo_43 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_43 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_43 = {maskExt_hi_43, maskExt_lo_43};
  wire [15:0]        maskExt_lo_44 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_44 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_44 = {maskExt_hi_44, maskExt_lo_44};
  wire [15:0]        maskExt_lo_45 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_45 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_45 = {maskExt_hi_45, maskExt_lo_45};
  wire [15:0]        maskExt_lo_46 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_46 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_46 = {maskExt_hi_46, maskExt_lo_46};
  wire [15:0]        maskExt_lo_47 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_47 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_47 = {maskExt_hi_47, maskExt_lo_47};
  wire [15:0]        maskExt_lo_48 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_48 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_48 = {maskExt_hi_48, maskExt_lo_48};
  wire [15:0]        maskExt_lo_49 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_49 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_49 = {maskExt_hi_49, maskExt_lo_49};
  wire [15:0]        maskExt_lo_50 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_50 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_50 = {maskExt_hi_50, maskExt_lo_50};
  wire [15:0]        maskExt_lo_51 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_51 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_51 = {maskExt_hi_51, maskExt_lo_51};
  wire [15:0]        maskExt_lo_52 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_52 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_52 = {maskExt_hi_52, maskExt_lo_52};
  wire [15:0]        maskExt_lo_53 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_53 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_53 = {maskExt_hi_53, maskExt_lo_53};
  wire [15:0]        maskExt_lo_54 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_54 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_54 = {maskExt_hi_54, maskExt_lo_54};
  wire [15:0]        maskExt_lo_55 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_55 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_55 = {maskExt_hi_55, maskExt_lo_55};
  wire [15:0]        maskExt_lo_56 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_56 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_56 = {maskExt_hi_56, maskExt_lo_56};
  wire [15:0]        maskExt_lo_57 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_57 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_57 = {maskExt_hi_57, maskExt_lo_57};
  wire [15:0]        maskExt_lo_58 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_58 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_58 = {maskExt_hi_58, maskExt_lo_58};
  wire [15:0]        maskExt_lo_59 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_59 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_59 = {maskExt_hi_59, maskExt_lo_59};
  wire [15:0]        maskExt_lo_60 = {{8{v0UpdateVec_0_bits_mask[1]}}, {8{v0UpdateVec_0_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_60 = {{8{v0UpdateVec_0_bits_mask[3]}}, {8{v0UpdateVec_0_bits_mask[2]}}};
  wire [31:0]        maskExt_60 = {maskExt_hi_60, maskExt_lo_60};
  wire [15:0]        maskExt_lo_61 = {{8{v0UpdateVec_1_bits_mask[1]}}, {8{v0UpdateVec_1_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_61 = {{8{v0UpdateVec_1_bits_mask[3]}}, {8{v0UpdateVec_1_bits_mask[2]}}};
  wire [31:0]        maskExt_61 = {maskExt_hi_61, maskExt_lo_61};
  wire [15:0]        maskExt_lo_62 = {{8{v0UpdateVec_2_bits_mask[1]}}, {8{v0UpdateVec_2_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_62 = {{8{v0UpdateVec_2_bits_mask[3]}}, {8{v0UpdateVec_2_bits_mask[2]}}};
  wire [31:0]        maskExt_62 = {maskExt_hi_62, maskExt_lo_62};
  wire [15:0]        maskExt_lo_63 = {{8{v0UpdateVec_3_bits_mask[1]}}, {8{v0UpdateVec_3_bits_mask[0]}}};
  wire [15:0]        maskExt_hi_63 = {{8{v0UpdateVec_3_bits_mask[3]}}, {8{v0UpdateVec_3_bits_mask[2]}}};
  wire [31:0]        maskExt_63 = {maskExt_hi_63, maskExt_lo_63};
  wire [63:0]        _GEN = {v0_1, v0_0};
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo;
  assign regroupV0_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_5;
  assign regroupV0_lo_lo_lo_lo_lo_5 = _GEN;
  wire [63:0]        regroupV0_lo_lo_lo_lo_lo_10;
  assign regroupV0_lo_lo_lo_lo_lo_10 = _GEN;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_lo;
  assign selectReadStageMask_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_1 = _GEN;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_lo_2 = _GEN;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_lo;
  assign maskForDestination_lo_lo_lo_lo_lo = _GEN;
  wire [63:0]        _GEN_0 = {v0_3, v0_2};
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi;
  assign regroupV0_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_5;
  assign regroupV0_lo_lo_lo_lo_hi_5 = _GEN_0;
  wire [63:0]        regroupV0_lo_lo_lo_lo_hi_10;
  assign regroupV0_lo_lo_lo_lo_hi_10 = _GEN_0;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        selectReadStageMask_lo_lo_lo_lo_hi;
  assign selectReadStageMask_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_1 = _GEN_0;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_lo_hi_2 = _GEN_0;
  wire [63:0]        maskForDestination_lo_lo_lo_lo_hi;
  assign maskForDestination_lo_lo_lo_lo_hi = _GEN_0;
  wire [127:0]       regroupV0_lo_lo_lo_lo = {regroupV0_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo};
  wire [63:0]        _GEN_1 = {v0_5, v0_4};
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo;
  assign regroupV0_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_5;
  assign regroupV0_lo_lo_lo_hi_lo_5 = _GEN_1;
  wire [63:0]        regroupV0_lo_lo_lo_hi_lo_10;
  assign regroupV0_lo_lo_lo_hi_lo_10 = _GEN_1;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_lo;
  assign selectReadStageMask_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_1 = _GEN_1;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_lo_2 = _GEN_1;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_lo;
  assign maskForDestination_lo_lo_lo_hi_lo = _GEN_1;
  wire [63:0]        _GEN_2 = {v0_7, v0_6};
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi;
  assign regroupV0_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_5;
  assign regroupV0_lo_lo_lo_hi_hi_5 = _GEN_2;
  wire [63:0]        regroupV0_lo_lo_lo_hi_hi_10;
  assign regroupV0_lo_lo_lo_hi_hi_10 = _GEN_2;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        selectReadStageMask_lo_lo_lo_hi_hi;
  assign selectReadStageMask_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_1 = _GEN_2;
  wire [63:0]        maskSplit_maskSelect_lo_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_lo_hi_hi_2 = _GEN_2;
  wire [63:0]        maskForDestination_lo_lo_lo_hi_hi;
  assign maskForDestination_lo_lo_lo_hi_hi = _GEN_2;
  wire [127:0]       regroupV0_lo_lo_lo_hi = {regroupV0_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo};
  wire [255:0]       regroupV0_lo_lo_lo = {regroupV0_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo};
  wire [63:0]        _GEN_3 = {v0_9, v0_8};
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo;
  assign regroupV0_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_5;
  assign regroupV0_lo_lo_hi_lo_lo_5 = _GEN_3;
  wire [63:0]        regroupV0_lo_lo_hi_lo_lo_10;
  assign regroupV0_lo_lo_hi_lo_lo_10 = _GEN_3;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_lo;
  assign selectReadStageMask_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_1 = _GEN_3;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_lo_2 = _GEN_3;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_lo;
  assign maskForDestination_lo_lo_hi_lo_lo = _GEN_3;
  wire [63:0]        _GEN_4 = {v0_11, v0_10};
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi;
  assign regroupV0_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_5;
  assign regroupV0_lo_lo_hi_lo_hi_5 = _GEN_4;
  wire [63:0]        regroupV0_lo_lo_hi_lo_hi_10;
  assign regroupV0_lo_lo_hi_lo_hi_10 = _GEN_4;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        selectReadStageMask_lo_lo_hi_lo_hi;
  assign selectReadStageMask_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_1 = _GEN_4;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_lo_hi_2 = _GEN_4;
  wire [63:0]        maskForDestination_lo_lo_hi_lo_hi;
  assign maskForDestination_lo_lo_hi_lo_hi = _GEN_4;
  wire [127:0]       regroupV0_lo_lo_hi_lo = {regroupV0_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo};
  wire [63:0]        _GEN_5 = {v0_13, v0_12};
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo;
  assign regroupV0_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_5;
  assign regroupV0_lo_lo_hi_hi_lo_5 = _GEN_5;
  wire [63:0]        regroupV0_lo_lo_hi_hi_lo_10;
  assign regroupV0_lo_lo_hi_hi_lo_10 = _GEN_5;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_lo;
  assign selectReadStageMask_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_1 = _GEN_5;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_lo_2 = _GEN_5;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_lo;
  assign maskForDestination_lo_lo_hi_hi_lo = _GEN_5;
  wire [63:0]        _GEN_6 = {v0_15, v0_14};
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi;
  assign regroupV0_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_5;
  assign regroupV0_lo_lo_hi_hi_hi_5 = _GEN_6;
  wire [63:0]        regroupV0_lo_lo_hi_hi_hi_10;
  assign regroupV0_lo_lo_hi_hi_hi_10 = _GEN_6;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        selectReadStageMask_lo_lo_hi_hi_hi;
  assign selectReadStageMask_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_1 = _GEN_6;
  wire [63:0]        maskSplit_maskSelect_lo_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_lo_hi_hi_hi_2 = _GEN_6;
  wire [63:0]        maskForDestination_lo_lo_hi_hi_hi;
  assign maskForDestination_lo_lo_hi_hi_hi = _GEN_6;
  wire [127:0]       regroupV0_lo_lo_hi_hi = {regroupV0_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo};
  wire [255:0]       regroupV0_lo_lo_hi = {regroupV0_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo};
  wire [511:0]       regroupV0_lo_lo = {regroupV0_lo_lo_hi, regroupV0_lo_lo_lo};
  wire [63:0]        _GEN_7 = {v0_17, v0_16};
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo;
  assign regroupV0_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_5;
  assign regroupV0_lo_hi_lo_lo_lo_5 = _GEN_7;
  wire [63:0]        regroupV0_lo_hi_lo_lo_lo_10;
  assign regroupV0_lo_hi_lo_lo_lo_10 = _GEN_7;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_lo;
  assign selectReadStageMask_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_1 = _GEN_7;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_lo_2 = _GEN_7;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_lo;
  assign maskForDestination_lo_hi_lo_lo_lo = _GEN_7;
  wire [63:0]        _GEN_8 = {v0_19, v0_18};
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi;
  assign regroupV0_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_5;
  assign regroupV0_lo_hi_lo_lo_hi_5 = _GEN_8;
  wire [63:0]        regroupV0_lo_hi_lo_lo_hi_10;
  assign regroupV0_lo_hi_lo_lo_hi_10 = _GEN_8;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        selectReadStageMask_lo_hi_lo_lo_hi;
  assign selectReadStageMask_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_1 = _GEN_8;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_lo_hi_2 = _GEN_8;
  wire [63:0]        maskForDestination_lo_hi_lo_lo_hi;
  assign maskForDestination_lo_hi_lo_lo_hi = _GEN_8;
  wire [127:0]       regroupV0_lo_hi_lo_lo = {regroupV0_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo};
  wire [63:0]        _GEN_9 = {v0_21, v0_20};
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo;
  assign regroupV0_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_5;
  assign regroupV0_lo_hi_lo_hi_lo_5 = _GEN_9;
  wire [63:0]        regroupV0_lo_hi_lo_hi_lo_10;
  assign regroupV0_lo_hi_lo_hi_lo_10 = _GEN_9;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_lo;
  assign selectReadStageMask_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_1 = _GEN_9;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_lo_2 = _GEN_9;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_lo;
  assign maskForDestination_lo_hi_lo_hi_lo = _GEN_9;
  wire [63:0]        _GEN_10 = {v0_23, v0_22};
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi;
  assign regroupV0_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_5;
  assign regroupV0_lo_hi_lo_hi_hi_5 = _GEN_10;
  wire [63:0]        regroupV0_lo_hi_lo_hi_hi_10;
  assign regroupV0_lo_hi_lo_hi_hi_10 = _GEN_10;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        selectReadStageMask_lo_hi_lo_hi_hi;
  assign selectReadStageMask_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_1 = _GEN_10;
  wire [63:0]        maskSplit_maskSelect_lo_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_lo_hi_hi_2 = _GEN_10;
  wire [63:0]        maskForDestination_lo_hi_lo_hi_hi;
  assign maskForDestination_lo_hi_lo_hi_hi = _GEN_10;
  wire [127:0]       regroupV0_lo_hi_lo_hi = {regroupV0_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo};
  wire [255:0]       regroupV0_lo_hi_lo = {regroupV0_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo};
  wire [63:0]        _GEN_11 = {v0_25, v0_24};
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo;
  assign regroupV0_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_5;
  assign regroupV0_lo_hi_hi_lo_lo_5 = _GEN_11;
  wire [63:0]        regroupV0_lo_hi_hi_lo_lo_10;
  assign regroupV0_lo_hi_hi_lo_lo_10 = _GEN_11;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_lo;
  assign selectReadStageMask_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_1 = _GEN_11;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_lo_2 = _GEN_11;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_lo;
  assign maskForDestination_lo_hi_hi_lo_lo = _GEN_11;
  wire [63:0]        _GEN_12 = {v0_27, v0_26};
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi;
  assign regroupV0_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_5;
  assign regroupV0_lo_hi_hi_lo_hi_5 = _GEN_12;
  wire [63:0]        regroupV0_lo_hi_hi_lo_hi_10;
  assign regroupV0_lo_hi_hi_lo_hi_10 = _GEN_12;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        selectReadStageMask_lo_hi_hi_lo_hi;
  assign selectReadStageMask_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_1 = _GEN_12;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_lo_hi_2 = _GEN_12;
  wire [63:0]        maskForDestination_lo_hi_hi_lo_hi;
  assign maskForDestination_lo_hi_hi_lo_hi = _GEN_12;
  wire [127:0]       regroupV0_lo_hi_hi_lo = {regroupV0_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo};
  wire [63:0]        _GEN_13 = {v0_29, v0_28};
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo;
  assign regroupV0_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_5;
  assign regroupV0_lo_hi_hi_hi_lo_5 = _GEN_13;
  wire [63:0]        regroupV0_lo_hi_hi_hi_lo_10;
  assign regroupV0_lo_hi_hi_hi_lo_10 = _GEN_13;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_lo;
  assign selectReadStageMask_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_1 = _GEN_13;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_lo_2 = _GEN_13;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_lo;
  assign maskForDestination_lo_hi_hi_hi_lo = _GEN_13;
  wire [63:0]        _GEN_14 = {v0_31, v0_30};
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi;
  assign regroupV0_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_5;
  assign regroupV0_lo_hi_hi_hi_hi_5 = _GEN_14;
  wire [63:0]        regroupV0_lo_hi_hi_hi_hi_10;
  assign regroupV0_lo_hi_hi_hi_hi_10 = _GEN_14;
  wire [63:0]        slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        selectReadStageMask_lo_hi_hi_hi_hi;
  assign selectReadStageMask_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_1 = _GEN_14;
  wire [63:0]        maskSplit_maskSelect_lo_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_lo_hi_hi_hi_hi_2 = _GEN_14;
  wire [63:0]        maskForDestination_lo_hi_hi_hi_hi;
  assign maskForDestination_lo_hi_hi_hi_hi = _GEN_14;
  wire [127:0]       regroupV0_lo_hi_hi_hi = {regroupV0_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo};
  wire [255:0]       regroupV0_lo_hi_hi = {regroupV0_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo};
  wire [511:0]       regroupV0_lo_hi = {regroupV0_lo_hi_hi, regroupV0_lo_hi_lo};
  wire [1023:0]      regroupV0_lo = {regroupV0_lo_hi, regroupV0_lo_lo};
  wire [63:0]        _GEN_15 = {v0_33, v0_32};
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo;
  assign regroupV0_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_5;
  assign regroupV0_hi_lo_lo_lo_lo_5 = _GEN_15;
  wire [63:0]        regroupV0_hi_lo_lo_lo_lo_10;
  assign regroupV0_hi_lo_lo_lo_lo_10 = _GEN_15;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_lo;
  assign selectReadStageMask_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_1 = _GEN_15;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_lo_2 = _GEN_15;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_lo;
  assign maskForDestination_hi_lo_lo_lo_lo = _GEN_15;
  wire [63:0]        _GEN_16 = {v0_35, v0_34};
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi;
  assign regroupV0_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_5;
  assign regroupV0_hi_lo_lo_lo_hi_5 = _GEN_16;
  wire [63:0]        regroupV0_hi_lo_lo_lo_hi_10;
  assign regroupV0_hi_lo_lo_lo_hi_10 = _GEN_16;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        selectReadStageMask_hi_lo_lo_lo_hi;
  assign selectReadStageMask_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_1 = _GEN_16;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_lo_hi_2 = _GEN_16;
  wire [63:0]        maskForDestination_hi_lo_lo_lo_hi;
  assign maskForDestination_hi_lo_lo_lo_hi = _GEN_16;
  wire [127:0]       regroupV0_hi_lo_lo_lo = {regroupV0_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo};
  wire [63:0]        _GEN_17 = {v0_37, v0_36};
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo;
  assign regroupV0_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_5;
  assign regroupV0_hi_lo_lo_hi_lo_5 = _GEN_17;
  wire [63:0]        regroupV0_hi_lo_lo_hi_lo_10;
  assign regroupV0_hi_lo_lo_hi_lo_10 = _GEN_17;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_lo;
  assign selectReadStageMask_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_1 = _GEN_17;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_lo_2 = _GEN_17;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_lo;
  assign maskForDestination_hi_lo_lo_hi_lo = _GEN_17;
  wire [63:0]        _GEN_18 = {v0_39, v0_38};
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi;
  assign regroupV0_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_5;
  assign regroupV0_hi_lo_lo_hi_hi_5 = _GEN_18;
  wire [63:0]        regroupV0_hi_lo_lo_hi_hi_10;
  assign regroupV0_hi_lo_lo_hi_hi_10 = _GEN_18;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        selectReadStageMask_hi_lo_lo_hi_hi;
  assign selectReadStageMask_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_1 = _GEN_18;
  wire [63:0]        maskSplit_maskSelect_hi_lo_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_lo_hi_hi_2 = _GEN_18;
  wire [63:0]        maskForDestination_hi_lo_lo_hi_hi;
  assign maskForDestination_hi_lo_lo_hi_hi = _GEN_18;
  wire [127:0]       regroupV0_hi_lo_lo_hi = {regroupV0_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo};
  wire [255:0]       regroupV0_hi_lo_lo = {regroupV0_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo};
  wire [63:0]        _GEN_19 = {v0_41, v0_40};
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo;
  assign regroupV0_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_5;
  assign regroupV0_hi_lo_hi_lo_lo_5 = _GEN_19;
  wire [63:0]        regroupV0_hi_lo_hi_lo_lo_10;
  assign regroupV0_hi_lo_hi_lo_lo_10 = _GEN_19;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_lo;
  assign selectReadStageMask_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_1 = _GEN_19;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_lo_2 = _GEN_19;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_lo;
  assign maskForDestination_hi_lo_hi_lo_lo = _GEN_19;
  wire [63:0]        _GEN_20 = {v0_43, v0_42};
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi;
  assign regroupV0_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_5;
  assign regroupV0_hi_lo_hi_lo_hi_5 = _GEN_20;
  wire [63:0]        regroupV0_hi_lo_hi_lo_hi_10;
  assign regroupV0_hi_lo_hi_lo_hi_10 = _GEN_20;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        selectReadStageMask_hi_lo_hi_lo_hi;
  assign selectReadStageMask_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_1 = _GEN_20;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_lo_hi_2 = _GEN_20;
  wire [63:0]        maskForDestination_hi_lo_hi_lo_hi;
  assign maskForDestination_hi_lo_hi_lo_hi = _GEN_20;
  wire [127:0]       regroupV0_hi_lo_hi_lo = {regroupV0_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo};
  wire [63:0]        _GEN_21 = {v0_45, v0_44};
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo;
  assign regroupV0_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_5;
  assign regroupV0_hi_lo_hi_hi_lo_5 = _GEN_21;
  wire [63:0]        regroupV0_hi_lo_hi_hi_lo_10;
  assign regroupV0_hi_lo_hi_hi_lo_10 = _GEN_21;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_lo;
  assign selectReadStageMask_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_1 = _GEN_21;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_lo_2 = _GEN_21;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_lo;
  assign maskForDestination_hi_lo_hi_hi_lo = _GEN_21;
  wire [63:0]        _GEN_22 = {v0_47, v0_46};
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi;
  assign regroupV0_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_5;
  assign regroupV0_hi_lo_hi_hi_hi_5 = _GEN_22;
  wire [63:0]        regroupV0_hi_lo_hi_hi_hi_10;
  assign regroupV0_hi_lo_hi_hi_hi_10 = _GEN_22;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        selectReadStageMask_hi_lo_hi_hi_hi;
  assign selectReadStageMask_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_1 = _GEN_22;
  wire [63:0]        maskSplit_maskSelect_hi_lo_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_lo_hi_hi_hi_2 = _GEN_22;
  wire [63:0]        maskForDestination_hi_lo_hi_hi_hi;
  assign maskForDestination_hi_lo_hi_hi_hi = _GEN_22;
  wire [127:0]       regroupV0_hi_lo_hi_hi = {regroupV0_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo};
  wire [255:0]       regroupV0_hi_lo_hi = {regroupV0_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo};
  wire [511:0]       regroupV0_hi_lo = {regroupV0_hi_lo_hi, regroupV0_hi_lo_lo};
  wire [63:0]        _GEN_23 = {v0_49, v0_48};
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo;
  assign regroupV0_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_5;
  assign regroupV0_hi_hi_lo_lo_lo_5 = _GEN_23;
  wire [63:0]        regroupV0_hi_hi_lo_lo_lo_10;
  assign regroupV0_hi_hi_lo_lo_lo_10 = _GEN_23;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_lo;
  assign selectReadStageMask_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_1 = _GEN_23;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_lo_2 = _GEN_23;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_lo;
  assign maskForDestination_hi_hi_lo_lo_lo = _GEN_23;
  wire [63:0]        _GEN_24 = {v0_51, v0_50};
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi;
  assign regroupV0_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_5;
  assign regroupV0_hi_hi_lo_lo_hi_5 = _GEN_24;
  wire [63:0]        regroupV0_hi_hi_lo_lo_hi_10;
  assign regroupV0_hi_hi_lo_lo_hi_10 = _GEN_24;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        selectReadStageMask_hi_hi_lo_lo_hi;
  assign selectReadStageMask_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_1 = _GEN_24;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_lo_hi_2 = _GEN_24;
  wire [63:0]        maskForDestination_hi_hi_lo_lo_hi;
  assign maskForDestination_hi_hi_lo_lo_hi = _GEN_24;
  wire [127:0]       regroupV0_hi_hi_lo_lo = {regroupV0_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo};
  wire [63:0]        _GEN_25 = {v0_53, v0_52};
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo;
  assign regroupV0_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_5;
  assign regroupV0_hi_hi_lo_hi_lo_5 = _GEN_25;
  wire [63:0]        regroupV0_hi_hi_lo_hi_lo_10;
  assign regroupV0_hi_hi_lo_hi_lo_10 = _GEN_25;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_lo;
  assign selectReadStageMask_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_1 = _GEN_25;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_lo_2 = _GEN_25;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_lo;
  assign maskForDestination_hi_hi_lo_hi_lo = _GEN_25;
  wire [63:0]        _GEN_26 = {v0_55, v0_54};
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi;
  assign regroupV0_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_5;
  assign regroupV0_hi_hi_lo_hi_hi_5 = _GEN_26;
  wire [63:0]        regroupV0_hi_hi_lo_hi_hi_10;
  assign regroupV0_hi_hi_lo_hi_hi_10 = _GEN_26;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        selectReadStageMask_hi_hi_lo_hi_hi;
  assign selectReadStageMask_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_1 = _GEN_26;
  wire [63:0]        maskSplit_maskSelect_hi_hi_lo_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_lo_hi_hi_2 = _GEN_26;
  wire [63:0]        maskForDestination_hi_hi_lo_hi_hi;
  assign maskForDestination_hi_hi_lo_hi_hi = _GEN_26;
  wire [127:0]       regroupV0_hi_hi_lo_hi = {regroupV0_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo};
  wire [255:0]       regroupV0_hi_hi_lo = {regroupV0_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo};
  wire [63:0]        _GEN_27 = {v0_57, v0_56};
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo;
  assign regroupV0_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_5;
  assign regroupV0_hi_hi_hi_lo_lo_5 = _GEN_27;
  wire [63:0]        regroupV0_hi_hi_hi_lo_lo_10;
  assign regroupV0_hi_hi_hi_lo_lo_10 = _GEN_27;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_lo;
  assign selectReadStageMask_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_1 = _GEN_27;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_lo_2 = _GEN_27;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_lo;
  assign maskForDestination_hi_hi_hi_lo_lo = _GEN_27;
  wire [63:0]        _GEN_28 = {v0_59, v0_58};
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi;
  assign regroupV0_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_5;
  assign regroupV0_hi_hi_hi_lo_hi_5 = _GEN_28;
  wire [63:0]        regroupV0_hi_hi_hi_lo_hi_10;
  assign regroupV0_hi_hi_hi_lo_hi_10 = _GEN_28;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        selectReadStageMask_hi_hi_hi_lo_hi;
  assign selectReadStageMask_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_1 = _GEN_28;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_lo_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_lo_hi_2 = _GEN_28;
  wire [63:0]        maskForDestination_hi_hi_hi_lo_hi;
  assign maskForDestination_hi_hi_hi_lo_hi = _GEN_28;
  wire [127:0]       regroupV0_hi_hi_hi_lo = {regroupV0_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo};
  wire [63:0]        _GEN_29 = {v0_61, v0_60};
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo;
  assign regroupV0_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_5;
  assign regroupV0_hi_hi_hi_hi_lo_5 = _GEN_29;
  wire [63:0]        regroupV0_hi_hi_hi_hi_lo_10;
  assign regroupV0_hi_hi_hi_hi_lo_10 = _GEN_29;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_lo;
  assign selectReadStageMask_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_1 = _GEN_29;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_lo_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_lo_2 = _GEN_29;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_lo;
  assign maskForDestination_hi_hi_hi_hi_lo = _GEN_29;
  wire [63:0]        _GEN_30 = {v0_63, v0_62};
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi;
  assign regroupV0_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_5;
  assign regroupV0_hi_hi_hi_hi_hi_5 = _GEN_30;
  wire [63:0]        regroupV0_hi_hi_hi_hi_hi_10;
  assign regroupV0_hi_hi_hi_hi_hi_10 = _GEN_30;
  wire [63:0]        slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi;
  assign slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        selectReadStageMask_hi_hi_hi_hi_hi;
  assign selectReadStageMask_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_1;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_1 = _GEN_30;
  wire [63:0]        maskSplit_maskSelect_hi_hi_hi_hi_hi_2;
  assign maskSplit_maskSelect_hi_hi_hi_hi_hi_2 = _GEN_30;
  wire [63:0]        maskForDestination_hi_hi_hi_hi_hi;
  assign maskForDestination_hi_hi_hi_hi_hi = _GEN_30;
  wire [127:0]       regroupV0_hi_hi_hi_hi = {regroupV0_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo};
  wire [255:0]       regroupV0_hi_hi_hi = {regroupV0_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo};
  wire [511:0]       regroupV0_hi_hi = {regroupV0_hi_hi_hi, regroupV0_hi_hi_lo};
  wire [1023:0]      regroupV0_hi = {regroupV0_hi_hi, regroupV0_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo = {regroupV0_lo[19:16], regroupV0_lo[3:0]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi = {regroupV0_lo[51:48], regroupV0_lo[35:32]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_1 = {regroupV0_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo = {regroupV0_lo[83:80], regroupV0_lo[67:64]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi = {regroupV0_lo[115:112], regroupV0_lo[99:96]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_1 = {regroupV0_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_lo_1 = {regroupV0_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo = {regroupV0_lo[147:144], regroupV0_lo[131:128]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi = {regroupV0_lo[179:176], regroupV0_lo[163:160]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_1 = {regroupV0_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo = {regroupV0_lo[211:208], regroupV0_lo[195:192]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi = {regroupV0_lo[243:240], regroupV0_lo[227:224]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_1 = {regroupV0_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_lo_hi_1 = {regroupV0_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_lo_1 = {regroupV0_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo = {regroupV0_lo[275:272], regroupV0_lo[259:256]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi = {regroupV0_lo[307:304], regroupV0_lo[291:288]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_1 = {regroupV0_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo = {regroupV0_lo[339:336], regroupV0_lo[323:320]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi = {regroupV0_lo[371:368], regroupV0_lo[355:352]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_1 = {regroupV0_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_lo_1 = {regroupV0_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo = {regroupV0_lo[403:400], regroupV0_lo[387:384]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi = {regroupV0_lo[435:432], regroupV0_lo[419:416]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_1 = {regroupV0_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo = {regroupV0_lo[467:464], regroupV0_lo[451:448]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi = {regroupV0_lo[499:496], regroupV0_lo[483:480]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_1 = {regroupV0_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_lo_hi_hi_1 = {regroupV0_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_lo_hi_1 = {regroupV0_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_1};
  wire [127:0]       regroupV0_lo_lo_1 = {regroupV0_lo_lo_hi_1, regroupV0_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo = {regroupV0_lo[531:528], regroupV0_lo[515:512]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi = {regroupV0_lo[563:560], regroupV0_lo[547:544]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_1 = {regroupV0_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo = {regroupV0_lo[595:592], regroupV0_lo[579:576]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi = {regroupV0_lo[627:624], regroupV0_lo[611:608]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_1 = {regroupV0_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_lo_1 = {regroupV0_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo = {regroupV0_lo[659:656], regroupV0_lo[643:640]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi = {regroupV0_lo[691:688], regroupV0_lo[675:672]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_1 = {regroupV0_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo = {regroupV0_lo[723:720], regroupV0_lo[707:704]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi = {regroupV0_lo[755:752], regroupV0_lo[739:736]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_1 = {regroupV0_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_lo_hi_1 = {regroupV0_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_lo_1 = {regroupV0_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo = {regroupV0_lo[787:784], regroupV0_lo[771:768]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi = {regroupV0_lo[819:816], regroupV0_lo[803:800]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_1 = {regroupV0_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo = {regroupV0_lo[851:848], regroupV0_lo[835:832]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi = {regroupV0_lo[883:880], regroupV0_lo[867:864]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_1 = {regroupV0_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_lo_1 = {regroupV0_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo = {regroupV0_lo[915:912], regroupV0_lo[899:896]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi = {regroupV0_lo[947:944], regroupV0_lo[931:928]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_1 = {regroupV0_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo = {regroupV0_lo[979:976], regroupV0_lo[963:960]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi = {regroupV0_lo[1011:1008], regroupV0_lo[995:992]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_1 = {regroupV0_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_lo_hi_hi_hi_1 = {regroupV0_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_lo_hi_hi_1 = {regroupV0_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_1};
  wire [127:0]       regroupV0_lo_hi_1 = {regroupV0_lo_hi_hi_1, regroupV0_lo_hi_lo_1};
  wire [255:0]       regroupV0_lo_1 = {regroupV0_lo_hi_1, regroupV0_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo = {regroupV0_hi[19:16], regroupV0_hi[3:0]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi = {regroupV0_hi[51:48], regroupV0_hi[35:32]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_1 = {regroupV0_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo = {regroupV0_hi[83:80], regroupV0_hi[67:64]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi = {regroupV0_hi[115:112], regroupV0_hi[99:96]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_1 = {regroupV0_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_lo_1 = {regroupV0_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo = {regroupV0_hi[147:144], regroupV0_hi[131:128]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi = {regroupV0_hi[179:176], regroupV0_hi[163:160]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_1 = {regroupV0_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo = {regroupV0_hi[211:208], regroupV0_hi[195:192]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi = {regroupV0_hi[243:240], regroupV0_hi[227:224]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_1 = {regroupV0_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_lo_hi_1 = {regroupV0_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_lo_1 = {regroupV0_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo = {regroupV0_hi[275:272], regroupV0_hi[259:256]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi = {regroupV0_hi[307:304], regroupV0_hi[291:288]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_1 = {regroupV0_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo = {regroupV0_hi[339:336], regroupV0_hi[323:320]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi = {regroupV0_hi[371:368], regroupV0_hi[355:352]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_1 = {regroupV0_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_lo_1 = {regroupV0_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo = {regroupV0_hi[403:400], regroupV0_hi[387:384]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi = {regroupV0_hi[435:432], regroupV0_hi[419:416]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_1 = {regroupV0_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo = {regroupV0_hi[467:464], regroupV0_hi[451:448]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi = {regroupV0_hi[499:496], regroupV0_hi[483:480]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_1 = {regroupV0_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_lo_hi_hi_1 = {regroupV0_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_lo_hi_1 = {regroupV0_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_1};
  wire [127:0]       regroupV0_hi_lo_1 = {regroupV0_hi_lo_hi_1, regroupV0_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo = {regroupV0_hi[531:528], regroupV0_hi[515:512]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi = {regroupV0_hi[563:560], regroupV0_hi[547:544]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_1 = {regroupV0_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo = {regroupV0_hi[595:592], regroupV0_hi[579:576]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi = {regroupV0_hi[627:624], regroupV0_hi[611:608]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_1 = {regroupV0_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_lo_1 = {regroupV0_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo = {regroupV0_hi[659:656], regroupV0_hi[643:640]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi = {regroupV0_hi[691:688], regroupV0_hi[675:672]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_1 = {regroupV0_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo = {regroupV0_hi[723:720], regroupV0_hi[707:704]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi = {regroupV0_hi[755:752], regroupV0_hi[739:736]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_1 = {regroupV0_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_lo_hi_1 = {regroupV0_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_lo_1 = {regroupV0_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo = {regroupV0_hi[787:784], regroupV0_hi[771:768]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi = {regroupV0_hi[819:816], regroupV0_hi[803:800]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_1 = {regroupV0_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo = {regroupV0_hi[851:848], regroupV0_hi[835:832]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi = {regroupV0_hi[883:880], regroupV0_hi[867:864]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_1 = {regroupV0_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_lo_1 = {regroupV0_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo = {regroupV0_hi[915:912], regroupV0_hi[899:896]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi = {regroupV0_hi[947:944], regroupV0_hi[931:928]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_1 = {regroupV0_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo = {regroupV0_hi[979:976], regroupV0_hi[963:960]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi = {regroupV0_hi[1011:1008], regroupV0_hi[995:992]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo};
  wire [31:0]        regroupV0_hi_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_1};
  wire [63:0]        regroupV0_hi_hi_hi_1 = {regroupV0_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_1};
  wire [127:0]       regroupV0_hi_hi_1 = {regroupV0_hi_hi_hi_1, regroupV0_hi_hi_lo_1};
  wire [255:0]       regroupV0_hi_1 = {regroupV0_hi_hi_1, regroupV0_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo[23:20], regroupV0_lo[7:4]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo[55:52], regroupV0_lo[39:36]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_2 = {regroupV0_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo[87:84], regroupV0_lo[71:68]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo[119:116], regroupV0_lo[103:100]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_2 = {regroupV0_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_lo_2 = {regroupV0_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo[151:148], regroupV0_lo[135:132]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo[183:180], regroupV0_lo[167:164]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_2 = {regroupV0_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo[215:212], regroupV0_lo[199:196]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo[247:244], regroupV0_lo[231:228]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_2 = {regroupV0_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_lo_hi_2 = {regroupV0_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_lo_2 = {regroupV0_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo[279:276], regroupV0_lo[263:260]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo[311:308], regroupV0_lo[295:292]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_2 = {regroupV0_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo[343:340], regroupV0_lo[327:324]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo[375:372], regroupV0_lo[359:356]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_2 = {regroupV0_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_lo_2 = {regroupV0_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo[407:404], regroupV0_lo[391:388]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo[439:436], regroupV0_lo[423:420]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_2 = {regroupV0_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo[471:468], regroupV0_lo[455:452]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo[503:500], regroupV0_lo[487:484]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_2 = {regroupV0_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_lo_hi_hi_2 = {regroupV0_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_lo_hi_2 = {regroupV0_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_2};
  wire [127:0]       regroupV0_lo_lo_2 = {regroupV0_lo_lo_hi_2, regroupV0_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo[535:532], regroupV0_lo[519:516]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo[567:564], regroupV0_lo[551:548]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_2 = {regroupV0_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo[599:596], regroupV0_lo[583:580]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo[631:628], regroupV0_lo[615:612]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_2 = {regroupV0_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_lo_2 = {regroupV0_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo[663:660], regroupV0_lo[647:644]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo[695:692], regroupV0_lo[679:676]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_2 = {regroupV0_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo[727:724], regroupV0_lo[711:708]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo[759:756], regroupV0_lo[743:740]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_2 = {regroupV0_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_lo_hi_2 = {regroupV0_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_lo_2 = {regroupV0_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo[791:788], regroupV0_lo[775:772]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo[823:820], regroupV0_lo[807:804]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_2 = {regroupV0_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo[855:852], regroupV0_lo[839:836]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo[887:884], regroupV0_lo[871:868]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_2 = {regroupV0_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_lo_2 = {regroupV0_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo[919:916], regroupV0_lo[903:900]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo[951:948], regroupV0_lo[935:932]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_2 = {regroupV0_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo[983:980], regroupV0_lo[967:964]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo[1015:1012], regroupV0_lo[999:996]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_2 = {regroupV0_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_lo_hi_hi_hi_2 = {regroupV0_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_lo_hi_hi_2 = {regroupV0_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_2};
  wire [127:0]       regroupV0_lo_hi_2 = {regroupV0_lo_hi_hi_2, regroupV0_lo_hi_lo_2};
  wire [255:0]       regroupV0_lo_2 = {regroupV0_lo_hi_2, regroupV0_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi[23:20], regroupV0_hi[7:4]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi[55:52], regroupV0_hi[39:36]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_2 = {regroupV0_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi[87:84], regroupV0_hi[71:68]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi[119:116], regroupV0_hi[103:100]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_2 = {regroupV0_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_lo_2 = {regroupV0_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi[151:148], regroupV0_hi[135:132]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi[183:180], regroupV0_hi[167:164]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_2 = {regroupV0_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi[215:212], regroupV0_hi[199:196]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi[247:244], regroupV0_hi[231:228]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_2 = {regroupV0_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_lo_hi_2 = {regroupV0_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_lo_2 = {regroupV0_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi[279:276], regroupV0_hi[263:260]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi[311:308], regroupV0_hi[295:292]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_2 = {regroupV0_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi[343:340], regroupV0_hi[327:324]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi[375:372], regroupV0_hi[359:356]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_2 = {regroupV0_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_lo_2 = {regroupV0_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi[407:404], regroupV0_hi[391:388]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi[439:436], regroupV0_hi[423:420]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_2 = {regroupV0_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi[471:468], regroupV0_hi[455:452]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi[503:500], regroupV0_hi[487:484]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_2 = {regroupV0_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_lo_hi_hi_2 = {regroupV0_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_lo_hi_2 = {regroupV0_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_2};
  wire [127:0]       regroupV0_hi_lo_2 = {regroupV0_hi_lo_hi_2, regroupV0_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi[535:532], regroupV0_hi[519:516]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi[567:564], regroupV0_hi[551:548]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_2 = {regroupV0_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi[599:596], regroupV0_hi[583:580]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi[631:628], regroupV0_hi[615:612]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_2 = {regroupV0_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_lo_2 = {regroupV0_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi[663:660], regroupV0_hi[647:644]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi[695:692], regroupV0_hi[679:676]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_2 = {regroupV0_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi[727:724], regroupV0_hi[711:708]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi[759:756], regroupV0_hi[743:740]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_2 = {regroupV0_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_lo_hi_2 = {regroupV0_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_lo_2 = {regroupV0_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi[791:788], regroupV0_hi[775:772]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi[823:820], regroupV0_hi[807:804]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_2 = {regroupV0_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi[855:852], regroupV0_hi[839:836]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi[887:884], regroupV0_hi[871:868]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_2 = {regroupV0_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_lo_2 = {regroupV0_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi[919:916], regroupV0_hi[903:900]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi[951:948], regroupV0_hi[935:932]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_2 = {regroupV0_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi[983:980], regroupV0_hi[967:964]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi[1015:1012], regroupV0_hi[999:996]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_1};
  wire [31:0]        regroupV0_hi_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_2};
  wire [63:0]        regroupV0_hi_hi_hi_2 = {regroupV0_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_2};
  wire [127:0]       regroupV0_hi_hi_2 = {regroupV0_hi_hi_hi_2, regroupV0_hi_hi_lo_2};
  wire [255:0]       regroupV0_hi_2 = {regroupV0_hi_hi_2, regroupV0_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo[27:24], regroupV0_lo[11:8]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo[59:56], regroupV0_lo[43:40]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_3 = {regroupV0_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo[91:88], regroupV0_lo[75:72]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo[123:120], regroupV0_lo[107:104]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_3 = {regroupV0_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_lo_3 = {regroupV0_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo[155:152], regroupV0_lo[139:136]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo[187:184], regroupV0_lo[171:168]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_3 = {regroupV0_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo[219:216], regroupV0_lo[203:200]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo[251:248], regroupV0_lo[235:232]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_3 = {regroupV0_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_lo_hi_3 = {regroupV0_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_lo_3 = {regroupV0_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo[283:280], regroupV0_lo[267:264]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo[315:312], regroupV0_lo[299:296]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_3 = {regroupV0_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo[347:344], regroupV0_lo[331:328]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo[379:376], regroupV0_lo[363:360]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_3 = {regroupV0_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_lo_3 = {regroupV0_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo[411:408], regroupV0_lo[395:392]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo[443:440], regroupV0_lo[427:424]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_3 = {regroupV0_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo[475:472], regroupV0_lo[459:456]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo[507:504], regroupV0_lo[491:488]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_3 = {regroupV0_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_lo_hi_hi_3 = {regroupV0_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_lo_hi_3 = {regroupV0_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_3};
  wire [127:0]       regroupV0_lo_lo_3 = {regroupV0_lo_lo_hi_3, regroupV0_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo[539:536], regroupV0_lo[523:520]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo[571:568], regroupV0_lo[555:552]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_3 = {regroupV0_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo[603:600], regroupV0_lo[587:584]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo[635:632], regroupV0_lo[619:616]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_3 = {regroupV0_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_lo_3 = {regroupV0_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo[667:664], regroupV0_lo[651:648]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo[699:696], regroupV0_lo[683:680]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_3 = {regroupV0_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo[731:728], regroupV0_lo[715:712]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo[763:760], regroupV0_lo[747:744]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_3 = {regroupV0_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_lo_hi_3 = {regroupV0_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_lo_3 = {regroupV0_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo[795:792], regroupV0_lo[779:776]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo[827:824], regroupV0_lo[811:808]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_3 = {regroupV0_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo[859:856], regroupV0_lo[843:840]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo[891:888], regroupV0_lo[875:872]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_3 = {regroupV0_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_lo_3 = {regroupV0_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo[923:920], regroupV0_lo[907:904]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo[955:952], regroupV0_lo[939:936]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_3 = {regroupV0_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo[987:984], regroupV0_lo[971:968]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo[1019:1016], regroupV0_lo[1003:1000]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_3 = {regroupV0_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_lo_hi_hi_hi_3 = {regroupV0_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_lo_hi_hi_3 = {regroupV0_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_3};
  wire [127:0]       regroupV0_lo_hi_3 = {regroupV0_lo_hi_hi_3, regroupV0_lo_hi_lo_3};
  wire [255:0]       regroupV0_lo_3 = {regroupV0_lo_hi_3, regroupV0_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi[27:24], regroupV0_hi[11:8]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi[59:56], regroupV0_hi[43:40]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_3 = {regroupV0_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi[91:88], regroupV0_hi[75:72]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi[123:120], regroupV0_hi[107:104]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_3 = {regroupV0_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_lo_3 = {regroupV0_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi[155:152], regroupV0_hi[139:136]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi[187:184], regroupV0_hi[171:168]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_3 = {regroupV0_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi[219:216], regroupV0_hi[203:200]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi[251:248], regroupV0_hi[235:232]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_3 = {regroupV0_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_lo_hi_3 = {regroupV0_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_lo_3 = {regroupV0_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi[283:280], regroupV0_hi[267:264]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi[315:312], regroupV0_hi[299:296]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_3 = {regroupV0_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi[347:344], regroupV0_hi[331:328]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi[379:376], regroupV0_hi[363:360]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_3 = {regroupV0_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_lo_3 = {regroupV0_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi[411:408], regroupV0_hi[395:392]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi[443:440], regroupV0_hi[427:424]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_3 = {regroupV0_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi[475:472], regroupV0_hi[459:456]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi[507:504], regroupV0_hi[491:488]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_3 = {regroupV0_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_lo_hi_hi_3 = {regroupV0_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_lo_hi_3 = {regroupV0_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_3};
  wire [127:0]       regroupV0_hi_lo_3 = {regroupV0_hi_lo_hi_3, regroupV0_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi[539:536], regroupV0_hi[523:520]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi[571:568], regroupV0_hi[555:552]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_3 = {regroupV0_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi[603:600], regroupV0_hi[587:584]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi[635:632], regroupV0_hi[619:616]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_3 = {regroupV0_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_lo_3 = {regroupV0_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi[667:664], regroupV0_hi[651:648]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi[699:696], regroupV0_hi[683:680]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_3 = {regroupV0_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi[731:728], regroupV0_hi[715:712]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi[763:760], regroupV0_hi[747:744]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_3 = {regroupV0_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_lo_hi_3 = {regroupV0_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_lo_3 = {regroupV0_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi[795:792], regroupV0_hi[779:776]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi[827:824], regroupV0_hi[811:808]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_3 = {regroupV0_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi[859:856], regroupV0_hi[843:840]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi[891:888], regroupV0_hi[875:872]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_3 = {regroupV0_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_lo_3 = {regroupV0_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi[923:920], regroupV0_hi[907:904]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi[955:952], regroupV0_hi[939:936]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_3 = {regroupV0_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi[987:984], regroupV0_hi[971:968]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi[1019:1016], regroupV0_hi[1003:1000]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_2};
  wire [31:0]        regroupV0_hi_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_3};
  wire [63:0]        regroupV0_hi_hi_hi_3 = {regroupV0_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_3};
  wire [127:0]       regroupV0_hi_hi_3 = {regroupV0_hi_hi_hi_3, regroupV0_hi_hi_lo_3};
  wire [255:0]       regroupV0_hi_3 = {regroupV0_hi_hi_3, regroupV0_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo[31:28], regroupV0_lo[15:12]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo[63:60], regroupV0_lo[47:44]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo[95:92], regroupV0_lo[79:76]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo[127:124], regroupV0_lo[111:108]};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo[159:156], regroupV0_lo[143:140]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo[191:188], regroupV0_lo[175:172]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo[223:220], regroupV0_lo[207:204]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo[255:252], regroupV0_lo[239:236]};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo[287:284], regroupV0_lo[271:268]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo[319:316], regroupV0_lo[303:300]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo[351:348], regroupV0_lo[335:332]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo[383:380], regroupV0_lo[367:364]};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo[415:412], regroupV0_lo[399:396]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo[447:444], regroupV0_lo[431:428]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo[479:476], regroupV0_lo[463:460]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo[511:508], regroupV0_lo[495:492]};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_4};
  wire [127:0]       regroupV0_lo_lo_4 = {regroupV0_lo_lo_hi_4, regroupV0_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo[543:540], regroupV0_lo[527:524]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo[575:572], regroupV0_lo[559:556]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo[607:604], regroupV0_lo[591:588]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo[639:636], regroupV0_lo[623:620]};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo[671:668], regroupV0_lo[655:652]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo[703:700], regroupV0_lo[687:684]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo[735:732], regroupV0_lo[719:716]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo[767:764], regroupV0_lo[751:748]};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo[799:796], regroupV0_lo[783:780]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo[831:828], regroupV0_lo[815:812]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo[863:860], regroupV0_lo[847:844]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo[895:892], regroupV0_lo[879:876]};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo[927:924], regroupV0_lo[911:908]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo[959:956], regroupV0_lo[943:940]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo[991:988], regroupV0_lo[975:972]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo[1023:1020], regroupV0_lo[1007:1004]};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_4};
  wire [127:0]       regroupV0_lo_hi_4 = {regroupV0_lo_hi_hi_4, regroupV0_lo_hi_lo_4};
  wire [255:0]       regroupV0_lo_4 = {regroupV0_lo_hi_4, regroupV0_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi[31:28], regroupV0_hi[15:12]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi[63:60], regroupV0_hi[47:44]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi[95:92], regroupV0_hi[79:76]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi[127:124], regroupV0_hi[111:108]};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi[159:156], regroupV0_hi[143:140]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi[191:188], regroupV0_hi[175:172]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi[223:220], regroupV0_hi[207:204]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi[255:252], regroupV0_hi[239:236]};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi[287:284], regroupV0_hi[271:268]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi[319:316], regroupV0_hi[303:300]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi[351:348], regroupV0_hi[335:332]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi[383:380], regroupV0_hi[367:364]};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi[415:412], regroupV0_hi[399:396]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi[447:444], regroupV0_hi[431:428]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi[479:476], regroupV0_hi[463:460]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi[511:508], regroupV0_hi[495:492]};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_4};
  wire [127:0]       regroupV0_hi_lo_4 = {regroupV0_hi_lo_hi_4, regroupV0_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi[543:540], regroupV0_hi[527:524]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi[575:572], regroupV0_hi[559:556]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi[607:604], regroupV0_hi[591:588]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi[639:636], regroupV0_hi[623:620]};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi[671:668], regroupV0_hi[655:652]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi[703:700], regroupV0_hi[687:684]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi[735:732], regroupV0_hi[719:716]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi[767:764], regroupV0_hi[751:748]};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi[799:796], regroupV0_hi[783:780]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi[831:828], regroupV0_hi[815:812]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi[863:860], regroupV0_hi[847:844]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi[895:892], regroupV0_hi[879:876]};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_4};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi[927:924], regroupV0_hi[911:908]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi[959:956], regroupV0_hi[943:940]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi[991:988], regroupV0_hi[975:972]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi[1023:1020], regroupV0_hi[1007:1004]};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_3};
  wire [31:0]        regroupV0_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_4};
  wire [63:0]        regroupV0_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_4};
  wire [127:0]       regroupV0_hi_hi_4 = {regroupV0_hi_hi_hi_4, regroupV0_hi_hi_lo_4};
  wire [255:0]       regroupV0_hi_4 = {regroupV0_hi_hi_4, regroupV0_hi_lo_4};
  wire [1023:0]      regroupV0_lo_5 = {regroupV0_hi_2, regroupV0_lo_2, regroupV0_hi_1, regroupV0_lo_1};
  wire [1023:0]      regroupV0_hi_5 = {regroupV0_hi_4, regroupV0_lo_4, regroupV0_hi_3, regroupV0_lo_3};
  wire [2047:0]      regroupV0_0 = {regroupV0_hi_5, regroupV0_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_5};
  wire [511:0]       regroupV0_lo_lo_5 = {regroupV0_lo_lo_hi_5, regroupV0_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_5};
  wire [511:0]       regroupV0_lo_hi_5 = {regroupV0_lo_hi_hi_5, regroupV0_lo_hi_lo_5};
  wire [1023:0]      regroupV0_lo_6 = {regroupV0_lo_hi_5, regroupV0_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_5};
  wire [511:0]       regroupV0_hi_lo_5 = {regroupV0_hi_lo_hi_5, regroupV0_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_5};
  wire [127:0]       regroupV0_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_5};
  wire [255:0]       regroupV0_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_5};
  wire [511:0]       regroupV0_hi_hi_5 = {regroupV0_hi_hi_hi_5, regroupV0_hi_hi_lo_5};
  wire [1023:0]      regroupV0_hi_6 = {regroupV0_hi_hi_5, regroupV0_hi_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_6[9:8], regroupV0_lo_6[1:0]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_6[25:24], regroupV0_lo_6[17:16]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_6[41:40], regroupV0_lo_6[33:32]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_6[57:56], regroupV0_lo_6[49:48]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_6[73:72], regroupV0_lo_6[65:64]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_6[89:88], regroupV0_lo_6[81:80]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_6[105:104], regroupV0_lo_6[97:96]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_6[121:120], regroupV0_lo_6[113:112]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_6[137:136], regroupV0_lo_6[129:128]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_6[153:152], regroupV0_lo_6[145:144]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_6[169:168], regroupV0_lo_6[161:160]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_6[185:184], regroupV0_lo_6[177:176]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_6[201:200], regroupV0_lo_6[193:192]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_6[217:216], regroupV0_lo_6[209:208]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_6[233:232], regroupV0_lo_6[225:224]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_6[249:248], regroupV0_lo_6[241:240]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_6[265:264], regroupV0_lo_6[257:256]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_6[281:280], regroupV0_lo_6[273:272]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_6[297:296], regroupV0_lo_6[289:288]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_6[313:312], regroupV0_lo_6[305:304]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_6[329:328], regroupV0_lo_6[321:320]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_6[345:344], regroupV0_lo_6[337:336]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_6[361:360], regroupV0_lo_6[353:352]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_6[377:376], regroupV0_lo_6[369:368]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_6[393:392], regroupV0_lo_6[385:384]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_6[409:408], regroupV0_lo_6[401:400]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_6[425:424], regroupV0_lo_6[417:416]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_6[441:440], regroupV0_lo_6[433:432]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_6[457:456], regroupV0_lo_6[449:448]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_6[473:472], regroupV0_lo_6[465:464]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_6[489:488], regroupV0_lo_6[481:480]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_6[505:504], regroupV0_lo_6[497:496]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_6};
  wire [127:0]       regroupV0_lo_lo_6 = {regroupV0_lo_lo_hi_6, regroupV0_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_6[521:520], regroupV0_lo_6[513:512]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_6[537:536], regroupV0_lo_6[529:528]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_6[553:552], regroupV0_lo_6[545:544]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_6[569:568], regroupV0_lo_6[561:560]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_6[585:584], regroupV0_lo_6[577:576]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_6[601:600], regroupV0_lo_6[593:592]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_6[617:616], regroupV0_lo_6[609:608]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_6[633:632], regroupV0_lo_6[625:624]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_6[649:648], regroupV0_lo_6[641:640]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_6[665:664], regroupV0_lo_6[657:656]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_6[681:680], regroupV0_lo_6[673:672]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_6[697:696], regroupV0_lo_6[689:688]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_6[713:712], regroupV0_lo_6[705:704]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_6[729:728], regroupV0_lo_6[721:720]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_6[745:744], regroupV0_lo_6[737:736]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_6[761:760], regroupV0_lo_6[753:752]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_6[777:776], regroupV0_lo_6[769:768]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_6[793:792], regroupV0_lo_6[785:784]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_6[809:808], regroupV0_lo_6[801:800]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_6[825:824], regroupV0_lo_6[817:816]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_6[841:840], regroupV0_lo_6[833:832]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_6[857:856], regroupV0_lo_6[849:848]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_6[873:872], regroupV0_lo_6[865:864]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_6[889:888], regroupV0_lo_6[881:880]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_6[905:904], regroupV0_lo_6[897:896]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_6[921:920], regroupV0_lo_6[913:912]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_6[937:936], regroupV0_lo_6[929:928]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_6[953:952], regroupV0_lo_6[945:944]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_6[969:968], regroupV0_lo_6[961:960]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_6[985:984], regroupV0_lo_6[977:976]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_6[1001:1000], regroupV0_lo_6[993:992]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_6[1017:1016], regroupV0_lo_6[1009:1008]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_6};
  wire [127:0]       regroupV0_lo_hi_6 = {regroupV0_lo_hi_hi_6, regroupV0_lo_hi_lo_6};
  wire [255:0]       regroupV0_lo_7 = {regroupV0_lo_hi_6, regroupV0_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_6[9:8], regroupV0_hi_6[1:0]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_6[25:24], regroupV0_hi_6[17:16]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_6[41:40], regroupV0_hi_6[33:32]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_6[57:56], regroupV0_hi_6[49:48]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_6[73:72], regroupV0_hi_6[65:64]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_6[89:88], regroupV0_hi_6[81:80]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_6[105:104], regroupV0_hi_6[97:96]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_6[121:120], regroupV0_hi_6[113:112]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_6[137:136], regroupV0_hi_6[129:128]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_6[153:152], regroupV0_hi_6[145:144]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_6[169:168], regroupV0_hi_6[161:160]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_6[185:184], regroupV0_hi_6[177:176]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_6[201:200], regroupV0_hi_6[193:192]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_6[217:216], regroupV0_hi_6[209:208]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_6[233:232], regroupV0_hi_6[225:224]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_6[249:248], regroupV0_hi_6[241:240]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_6[265:264], regroupV0_hi_6[257:256]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_6[281:280], regroupV0_hi_6[273:272]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_6[297:296], regroupV0_hi_6[289:288]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_6[313:312], regroupV0_hi_6[305:304]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_6[329:328], regroupV0_hi_6[321:320]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_6[345:344], regroupV0_hi_6[337:336]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_6[361:360], regroupV0_hi_6[353:352]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_6[377:376], regroupV0_hi_6[369:368]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_6[393:392], regroupV0_hi_6[385:384]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_6[409:408], regroupV0_hi_6[401:400]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_6[425:424], regroupV0_hi_6[417:416]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_6[441:440], regroupV0_hi_6[433:432]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_6[457:456], regroupV0_hi_6[449:448]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_6[473:472], regroupV0_hi_6[465:464]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_6[489:488], regroupV0_hi_6[481:480]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_6[505:504], regroupV0_hi_6[497:496]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_6};
  wire [127:0]       regroupV0_hi_lo_6 = {regroupV0_hi_lo_hi_6, regroupV0_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_6[521:520], regroupV0_hi_6[513:512]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_6[537:536], regroupV0_hi_6[529:528]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_6[553:552], regroupV0_hi_6[545:544]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_6[569:568], regroupV0_hi_6[561:560]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_6[585:584], regroupV0_hi_6[577:576]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_6[601:600], regroupV0_hi_6[593:592]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_6[617:616], regroupV0_hi_6[609:608]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_6[633:632], regroupV0_hi_6[625:624]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_6[649:648], regroupV0_hi_6[641:640]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_6[665:664], regroupV0_hi_6[657:656]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_6[681:680], regroupV0_hi_6[673:672]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_6[697:696], regroupV0_hi_6[689:688]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_6[713:712], regroupV0_hi_6[705:704]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_6[729:728], regroupV0_hi_6[721:720]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_6[745:744], regroupV0_hi_6[737:736]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_6[761:760], regroupV0_hi_6[753:752]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_6[777:776], regroupV0_hi_6[769:768]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_6[793:792], regroupV0_hi_6[785:784]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_6[809:808], regroupV0_hi_6[801:800]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_6[825:824], regroupV0_hi_6[817:816]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_6[841:840], regroupV0_hi_6[833:832]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_6[857:856], regroupV0_hi_6[849:848]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_6[873:872], regroupV0_hi_6[865:864]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_6[889:888], regroupV0_hi_6[881:880]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_6[905:904], regroupV0_hi_6[897:896]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_6[921:920], regroupV0_hi_6[913:912]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_6[937:936], regroupV0_hi_6[929:928]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_6[953:952], regroupV0_hi_6[945:944]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_4};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_6[969:968], regroupV0_hi_6[961:960]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_6[985:984], regroupV0_hi_6[977:976]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_6[1001:1000], regroupV0_hi_6[993:992]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_6[1017:1016], regroupV0_hi_6[1009:1008]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_4};
  wire [31:0]        regroupV0_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_6};
  wire [63:0]        regroupV0_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_6};
  wire [127:0]       regroupV0_hi_hi_6 = {regroupV0_hi_hi_hi_6, regroupV0_hi_hi_lo_6};
  wire [255:0]       regroupV0_hi_7 = {regroupV0_hi_hi_6, regroupV0_hi_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[11:10], regroupV0_lo_6[3:2]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[27:26], regroupV0_lo_6[19:18]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[43:42], regroupV0_lo_6[35:34]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[59:58], regroupV0_lo_6[51:50]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[75:74], regroupV0_lo_6[67:66]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[91:90], regroupV0_lo_6[83:82]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[107:106], regroupV0_lo_6[99:98]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[123:122], regroupV0_lo_6[115:114]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[139:138], regroupV0_lo_6[131:130]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[155:154], regroupV0_lo_6[147:146]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[171:170], regroupV0_lo_6[163:162]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[187:186], regroupV0_lo_6[179:178]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[203:202], regroupV0_lo_6[195:194]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[219:218], regroupV0_lo_6[211:210]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[235:234], regroupV0_lo_6[227:226]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[251:250], regroupV0_lo_6[243:242]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[267:266], regroupV0_lo_6[259:258]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[283:282], regroupV0_lo_6[275:274]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[299:298], regroupV0_lo_6[291:290]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[315:314], regroupV0_lo_6[307:306]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[331:330], regroupV0_lo_6[323:322]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[347:346], regroupV0_lo_6[339:338]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[363:362], regroupV0_lo_6[355:354]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[379:378], regroupV0_lo_6[371:370]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[395:394], regroupV0_lo_6[387:386]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[411:410], regroupV0_lo_6[403:402]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[427:426], regroupV0_lo_6[419:418]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[443:442], regroupV0_lo_6[435:434]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[459:458], regroupV0_lo_6[451:450]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[475:474], regroupV0_lo_6[467:466]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[491:490], regroupV0_lo_6[483:482]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[507:506], regroupV0_lo_6[499:498]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_7};
  wire [127:0]       regroupV0_lo_lo_7 = {regroupV0_lo_lo_hi_7, regroupV0_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_6[523:522], regroupV0_lo_6[515:514]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_6[539:538], regroupV0_lo_6[531:530]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_6[555:554], regroupV0_lo_6[547:546]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_6[571:570], regroupV0_lo_6[563:562]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_6[587:586], regroupV0_lo_6[579:578]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_6[603:602], regroupV0_lo_6[595:594]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_6[619:618], regroupV0_lo_6[611:610]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_6[635:634], regroupV0_lo_6[627:626]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_6[651:650], regroupV0_lo_6[643:642]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_6[667:666], regroupV0_lo_6[659:658]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_6[683:682], regroupV0_lo_6[675:674]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_6[699:698], regroupV0_lo_6[691:690]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_6[715:714], regroupV0_lo_6[707:706]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_6[731:730], regroupV0_lo_6[723:722]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_6[747:746], regroupV0_lo_6[739:738]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_6[763:762], regroupV0_lo_6[755:754]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_6[779:778], regroupV0_lo_6[771:770]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_6[795:794], regroupV0_lo_6[787:786]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_6[811:810], regroupV0_lo_6[803:802]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_6[827:826], regroupV0_lo_6[819:818]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_6[843:842], regroupV0_lo_6[835:834]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_6[859:858], regroupV0_lo_6[851:850]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_6[875:874], regroupV0_lo_6[867:866]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_6[891:890], regroupV0_lo_6[883:882]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_6[907:906], regroupV0_lo_6[899:898]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_6[923:922], regroupV0_lo_6[915:914]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_6[939:938], regroupV0_lo_6[931:930]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_6[955:954], regroupV0_lo_6[947:946]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_6[971:970], regroupV0_lo_6[963:962]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_6[987:986], regroupV0_lo_6[979:978]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_6[1003:1002], regroupV0_lo_6[995:994]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_6[1019:1018], regroupV0_lo_6[1011:1010]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_7};
  wire [127:0]       regroupV0_lo_hi_7 = {regroupV0_lo_hi_hi_7, regroupV0_lo_hi_lo_7};
  wire [255:0]       regroupV0_lo_8 = {regroupV0_lo_hi_7, regroupV0_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[11:10], regroupV0_hi_6[3:2]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[27:26], regroupV0_hi_6[19:18]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[43:42], regroupV0_hi_6[35:34]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[59:58], regroupV0_hi_6[51:50]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[75:74], regroupV0_hi_6[67:66]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[91:90], regroupV0_hi_6[83:82]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[107:106], regroupV0_hi_6[99:98]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[123:122], regroupV0_hi_6[115:114]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[139:138], regroupV0_hi_6[131:130]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[155:154], regroupV0_hi_6[147:146]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[171:170], regroupV0_hi_6[163:162]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[187:186], regroupV0_hi_6[179:178]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[203:202], regroupV0_hi_6[195:194]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[219:218], regroupV0_hi_6[211:210]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[235:234], regroupV0_hi_6[227:226]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[251:250], regroupV0_hi_6[243:242]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[267:266], regroupV0_hi_6[259:258]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[283:282], regroupV0_hi_6[275:274]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[299:298], regroupV0_hi_6[291:290]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[315:314], regroupV0_hi_6[307:306]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[331:330], regroupV0_hi_6[323:322]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[347:346], regroupV0_hi_6[339:338]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[363:362], regroupV0_hi_6[355:354]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[379:378], regroupV0_hi_6[371:370]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[395:394], regroupV0_hi_6[387:386]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[411:410], regroupV0_hi_6[403:402]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[427:426], regroupV0_hi_6[419:418]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[443:442], regroupV0_hi_6[435:434]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[459:458], regroupV0_hi_6[451:450]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[475:474], regroupV0_hi_6[467:466]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[491:490], regroupV0_hi_6[483:482]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[507:506], regroupV0_hi_6[499:498]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_7};
  wire [127:0]       regroupV0_hi_lo_7 = {regroupV0_hi_lo_hi_7, regroupV0_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_6[523:522], regroupV0_hi_6[515:514]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_6[539:538], regroupV0_hi_6[531:530]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_6[555:554], regroupV0_hi_6[547:546]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_6[571:570], regroupV0_hi_6[563:562]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_6[587:586], regroupV0_hi_6[579:578]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_6[603:602], regroupV0_hi_6[595:594]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_6[619:618], regroupV0_hi_6[611:610]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_6[635:634], regroupV0_hi_6[627:626]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_6[651:650], regroupV0_hi_6[643:642]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_6[667:666], regroupV0_hi_6[659:658]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_6[683:682], regroupV0_hi_6[675:674]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_6[699:698], regroupV0_hi_6[691:690]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_6[715:714], regroupV0_hi_6[707:706]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_6[731:730], regroupV0_hi_6[723:722]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_6[747:746], regroupV0_hi_6[739:738]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_6[763:762], regroupV0_hi_6[755:754]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_6[779:778], regroupV0_hi_6[771:770]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_6[795:794], regroupV0_hi_6[787:786]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_6[811:810], regroupV0_hi_6[803:802]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_6[827:826], regroupV0_hi_6[819:818]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_6[843:842], regroupV0_hi_6[835:834]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_6[859:858], regroupV0_hi_6[851:850]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_6[875:874], regroupV0_hi_6[867:866]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_6[891:890], regroupV0_hi_6[883:882]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_6[907:906], regroupV0_hi_6[899:898]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_6[923:922], regroupV0_hi_6[915:914]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_6[939:938], regroupV0_hi_6[931:930]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_6[955:954], regroupV0_hi_6[947:946]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_5};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_6[971:970], regroupV0_hi_6[963:962]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_6[987:986], regroupV0_hi_6[979:978]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_6[1003:1002], regroupV0_hi_6[995:994]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_6[1019:1018], regroupV0_hi_6[1011:1010]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_5};
  wire [31:0]        regroupV0_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_7};
  wire [63:0]        regroupV0_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_7};
  wire [127:0]       regroupV0_hi_hi_7 = {regroupV0_hi_hi_hi_7, regroupV0_hi_hi_lo_7};
  wire [255:0]       regroupV0_hi_8 = {regroupV0_hi_hi_7, regroupV0_hi_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[13:12], regroupV0_lo_6[5:4]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[29:28], regroupV0_lo_6[21:20]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[45:44], regroupV0_lo_6[37:36]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[61:60], regroupV0_lo_6[53:52]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[77:76], regroupV0_lo_6[69:68]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[93:92], regroupV0_lo_6[85:84]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[109:108], regroupV0_lo_6[101:100]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[125:124], regroupV0_lo_6[117:116]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[141:140], regroupV0_lo_6[133:132]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[157:156], regroupV0_lo_6[149:148]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[173:172], regroupV0_lo_6[165:164]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[189:188], regroupV0_lo_6[181:180]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[205:204], regroupV0_lo_6[197:196]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[221:220], regroupV0_lo_6[213:212]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[237:236], regroupV0_lo_6[229:228]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[253:252], regroupV0_lo_6[245:244]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_lo_8 = {regroupV0_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[269:268], regroupV0_lo_6[261:260]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[285:284], regroupV0_lo_6[277:276]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[301:300], regroupV0_lo_6[293:292]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[317:316], regroupV0_lo_6[309:308]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[333:332], regroupV0_lo_6[325:324]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[349:348], regroupV0_lo_6[341:340]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[365:364], regroupV0_lo_6[357:356]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[381:380], regroupV0_lo_6[373:372]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_lo_8 = {regroupV0_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[397:396], regroupV0_lo_6[389:388]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[413:412], regroupV0_lo_6[405:404]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[429:428], regroupV0_lo_6[421:420]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[445:444], regroupV0_lo_6[437:436]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[461:460], regroupV0_lo_6[453:452]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[477:476], regroupV0_lo_6[469:468]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[493:492], regroupV0_lo_6[485:484]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[509:508], regroupV0_lo_6[501:500]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_lo_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_lo_hi_8 = {regroupV0_lo_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_8};
  wire [127:0]       regroupV0_lo_lo_8 = {regroupV0_lo_lo_hi_8, regroupV0_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_6[525:524], regroupV0_lo_6[517:516]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_6[541:540], regroupV0_lo_6[533:532]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_6[557:556], regroupV0_lo_6[549:548]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_6[573:572], regroupV0_lo_6[565:564]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_6[589:588], regroupV0_lo_6[581:580]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_6[605:604], regroupV0_lo_6[597:596]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_6[621:620], regroupV0_lo_6[613:612]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_6[637:636], regroupV0_lo_6[629:628]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_lo_8 = {regroupV0_lo_hi_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_6[653:652], regroupV0_lo_6[645:644]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_6[669:668], regroupV0_lo_6[661:660]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_6[685:684], regroupV0_lo_6[677:676]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_6[701:700], regroupV0_lo_6[693:692]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_6[717:716], regroupV0_lo_6[709:708]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_6[733:732], regroupV0_lo_6[725:724]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_6[749:748], regroupV0_lo_6[741:740]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_6[765:764], regroupV0_lo_6[757:756]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_lo_hi_8 = {regroupV0_lo_hi_lo_hi_hi_8, regroupV0_lo_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_lo_8 = {regroupV0_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_6[781:780], regroupV0_lo_6[773:772]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_6[797:796], regroupV0_lo_6[789:788]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_6[813:812], regroupV0_lo_6[805:804]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_6[829:828], regroupV0_lo_6[821:820]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_6[845:844], regroupV0_lo_6[837:836]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_6[861:860], regroupV0_lo_6[853:852]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_6[877:876], regroupV0_lo_6[869:868]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_6[893:892], regroupV0_lo_6[885:884]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_lo_8 = {regroupV0_lo_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_6[909:908], regroupV0_lo_6[901:900]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_6[925:924], regroupV0_lo_6[917:916]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_6[941:940], regroupV0_lo_6[933:932]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_6[957:956], regroupV0_lo_6[949:948]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_6[973:972], regroupV0_lo_6[965:964]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_6[989:988], regroupV0_lo_6[981:980]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_6[1005:1004], regroupV0_lo_6[997:996]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_6[1021:1020], regroupV0_lo_6[1013:1012]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_lo_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_lo_hi_hi_8 = {regroupV0_lo_hi_hi_hi_8, regroupV0_lo_hi_hi_lo_8};
  wire [127:0]       regroupV0_lo_hi_8 = {regroupV0_lo_hi_hi_8, regroupV0_lo_hi_lo_8};
  wire [255:0]       regroupV0_lo_9 = {regroupV0_lo_hi_8, regroupV0_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[13:12], regroupV0_hi_6[5:4]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[29:28], regroupV0_hi_6[21:20]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[45:44], regroupV0_hi_6[37:36]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[61:60], regroupV0_hi_6[53:52]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[77:76], regroupV0_hi_6[69:68]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[93:92], regroupV0_hi_6[85:84]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[109:108], regroupV0_hi_6[101:100]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[125:124], regroupV0_hi_6[117:116]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[141:140], regroupV0_hi_6[133:132]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[157:156], regroupV0_hi_6[149:148]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[173:172], regroupV0_hi_6[165:164]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[189:188], regroupV0_hi_6[181:180]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[205:204], regroupV0_hi_6[197:196]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[221:220], regroupV0_hi_6[213:212]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[237:236], regroupV0_hi_6[229:228]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[253:252], regroupV0_hi_6[245:244]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_lo_hi_8 = {regroupV0_hi_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[269:268], regroupV0_hi_6[261:260]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[285:284], regroupV0_hi_6[277:276]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[301:300], regroupV0_hi_6[293:292]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[317:316], regroupV0_hi_6[309:308]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[333:332], regroupV0_hi_6[325:324]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[349:348], regroupV0_hi_6[341:340]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[365:364], regroupV0_hi_6[357:356]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[381:380], regroupV0_hi_6[373:372]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_lo_8 = {regroupV0_hi_lo_hi_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[397:396], regroupV0_hi_6[389:388]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[413:412], regroupV0_hi_6[405:404]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[429:428], regroupV0_hi_6[421:420]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[445:444], regroupV0_hi_6[437:436]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[461:460], regroupV0_hi_6[453:452]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[477:476], regroupV0_hi_6[469:468]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[493:492], regroupV0_hi_6[485:484]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[509:508], regroupV0_hi_6[501:500]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_lo_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_8};
  wire [127:0]       regroupV0_hi_lo_8 = {regroupV0_hi_lo_hi_8, regroupV0_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_6[525:524], regroupV0_hi_6[517:516]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_6[541:540], regroupV0_hi_6[533:532]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_6[557:556], regroupV0_hi_6[549:548]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_6[573:572], regroupV0_hi_6[565:564]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_6[589:588], regroupV0_hi_6[581:580]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_6[605:604], regroupV0_hi_6[597:596]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_6[621:620], regroupV0_hi_6[613:612]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_6[637:636], regroupV0_hi_6[629:628]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_lo_8 = {regroupV0_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_6[653:652], regroupV0_hi_6[645:644]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_6[669:668], regroupV0_hi_6[661:660]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_6[685:684], regroupV0_hi_6[677:676]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_6[701:700], regroupV0_hi_6[693:692]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_6[717:716], regroupV0_hi_6[709:708]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_6[733:732], regroupV0_hi_6[725:724]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_6[749:748], regroupV0_hi_6[741:740]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_6[765:764], regroupV0_hi_6[757:756]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_lo_hi_8 = {regroupV0_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_lo_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_8, regroupV0_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_6[781:780], regroupV0_hi_6[773:772]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_6[797:796], regroupV0_hi_6[789:788]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_6[813:812], regroupV0_hi_6[805:804]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_6[829:828], regroupV0_hi_6[821:820]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_6[845:844], regroupV0_hi_6[837:836]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_6[861:860], regroupV0_hi_6[853:852]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_6[877:876], regroupV0_hi_6[869:868]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_6[893:892], regroupV0_hi_6[885:884]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_8};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_6[909:908], regroupV0_hi_6[901:900]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_6[925:924], regroupV0_hi_6[917:916]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_6[941:940], regroupV0_hi_6[933:932]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_6[957:956], regroupV0_hi_6[949:948]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_6};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_6[973:972], regroupV0_hi_6[965:964]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_6[989:988], regroupV0_hi_6[981:980]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_2};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_6[1005:1004], regroupV0_hi_6[997:996]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_6[1021:1020], regroupV0_hi_6[1013:1012]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_6};
  wire [31:0]        regroupV0_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_lo_8};
  wire [63:0]        regroupV0_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_lo_8};
  wire [127:0]       regroupV0_hi_hi_8 = {regroupV0_hi_hi_hi_8, regroupV0_hi_hi_lo_8};
  wire [255:0]       regroupV0_hi_9 = {regroupV0_hi_hi_8, regroupV0_hi_lo_8};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[15:14], regroupV0_lo_6[7:6]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[31:30], regroupV0_lo_6[23:22]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[47:46], regroupV0_lo_6[39:38]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[63:62], regroupV0_lo_6[55:54]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[79:78], regroupV0_lo_6[71:70]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[95:94], regroupV0_lo_6[87:86]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[111:110], regroupV0_lo_6[103:102]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[127:126], regroupV0_lo_6[119:118]};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[143:142], regroupV0_lo_6[135:134]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[159:158], regroupV0_lo_6[151:150]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[175:174], regroupV0_lo_6[167:166]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[191:190], regroupV0_lo_6[183:182]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[207:206], regroupV0_lo_6[199:198]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[223:222], regroupV0_lo_6[215:214]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[239:238], regroupV0_lo_6[231:230]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[255:254], regroupV0_lo_6[247:246]};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_lo_9 = {regroupV0_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[271:270], regroupV0_lo_6[263:262]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[287:286], regroupV0_lo_6[279:278]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[303:302], regroupV0_lo_6[295:294]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[319:318], regroupV0_lo_6[311:310]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[335:334], regroupV0_lo_6[327:326]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[351:350], regroupV0_lo_6[343:342]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[367:366], regroupV0_lo_6[359:358]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[383:382], regroupV0_lo_6[375:374]};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_lo_9 = {regroupV0_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[399:398], regroupV0_lo_6[391:390]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[415:414], regroupV0_lo_6[407:406]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[431:430], regroupV0_lo_6[423:422]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[447:446], regroupV0_lo_6[439:438]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[463:462], regroupV0_lo_6[455:454]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[479:478], regroupV0_lo_6[471:470]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[495:494], regroupV0_lo_6[487:486]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[511:510], regroupV0_lo_6[503:502]};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_lo_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_lo_hi_9 = {regroupV0_lo_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_9};
  wire [127:0]       regroupV0_lo_lo_9 = {regroupV0_lo_lo_hi_9, regroupV0_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_6[527:526], regroupV0_lo_6[519:518]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_6[543:542], regroupV0_lo_6[535:534]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_6[559:558], regroupV0_lo_6[551:550]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_6[575:574], regroupV0_lo_6[567:566]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_6[591:590], regroupV0_lo_6[583:582]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_6[607:606], regroupV0_lo_6[599:598]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_6[623:622], regroupV0_lo_6[615:614]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_6[639:638], regroupV0_lo_6[631:630]};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_lo_9 = {regroupV0_lo_hi_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_6[655:654], regroupV0_lo_6[647:646]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_6[671:670], regroupV0_lo_6[663:662]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_6[687:686], regroupV0_lo_6[679:678]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_6[703:702], regroupV0_lo_6[695:694]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_6[719:718], regroupV0_lo_6[711:710]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_6[735:734], regroupV0_lo_6[727:726]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_6[751:750], regroupV0_lo_6[743:742]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_6[767:766], regroupV0_lo_6[759:758]};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_lo_hi_9 = {regroupV0_lo_hi_lo_hi_hi_9, regroupV0_lo_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_lo_9 = {regroupV0_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_6[783:782], regroupV0_lo_6[775:774]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_6[799:798], regroupV0_lo_6[791:790]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_6[815:814], regroupV0_lo_6[807:806]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_6[831:830], regroupV0_lo_6[823:822]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_6[847:846], regroupV0_lo_6[839:838]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_6[863:862], regroupV0_lo_6[855:854]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_6[879:878], regroupV0_lo_6[871:870]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_6[895:894], regroupV0_lo_6[887:886]};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_lo_9 = {regroupV0_lo_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_6[911:910], regroupV0_lo_6[903:902]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_6[927:926], regroupV0_lo_6[919:918]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_6[943:942], regroupV0_lo_6[935:934]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_6[959:958], regroupV0_lo_6[951:950]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_6[975:974], regroupV0_lo_6[967:966]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_6[991:990], regroupV0_lo_6[983:982]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_6[1007:1006], regroupV0_lo_6[999:998]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_6[1023:1022], regroupV0_lo_6[1015:1014]};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_lo_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_lo_hi_hi_9 = {regroupV0_lo_hi_hi_hi_9, regroupV0_lo_hi_hi_lo_9};
  wire [127:0]       regroupV0_lo_hi_9 = {regroupV0_lo_hi_hi_9, regroupV0_lo_hi_lo_9};
  wire [255:0]       regroupV0_lo_10 = {regroupV0_lo_hi_9, regroupV0_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[15:14], regroupV0_hi_6[7:6]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[31:30], regroupV0_hi_6[23:22]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[47:46], regroupV0_hi_6[39:38]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[63:62], regroupV0_hi_6[55:54]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[79:78], regroupV0_hi_6[71:70]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[95:94], regroupV0_hi_6[87:86]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[111:110], regroupV0_hi_6[103:102]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[127:126], regroupV0_hi_6[119:118]};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[143:142], regroupV0_hi_6[135:134]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[159:158], regroupV0_hi_6[151:150]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[175:174], regroupV0_hi_6[167:166]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[191:190], regroupV0_hi_6[183:182]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[207:206], regroupV0_hi_6[199:198]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[223:222], regroupV0_hi_6[215:214]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[239:238], regroupV0_hi_6[231:230]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[255:254], regroupV0_hi_6[247:246]};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_lo_hi_9 = {regroupV0_hi_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[271:270], regroupV0_hi_6[263:262]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[287:286], regroupV0_hi_6[279:278]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[303:302], regroupV0_hi_6[295:294]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[319:318], regroupV0_hi_6[311:310]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[335:334], regroupV0_hi_6[327:326]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[351:350], regroupV0_hi_6[343:342]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[367:366], regroupV0_hi_6[359:358]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[383:382], regroupV0_hi_6[375:374]};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_lo_9 = {regroupV0_hi_lo_hi_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[399:398], regroupV0_hi_6[391:390]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[415:414], regroupV0_hi_6[407:406]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[431:430], regroupV0_hi_6[423:422]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[447:446], regroupV0_hi_6[439:438]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[463:462], regroupV0_hi_6[455:454]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[479:478], regroupV0_hi_6[471:470]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[495:494], regroupV0_hi_6[487:486]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[511:510], regroupV0_hi_6[503:502]};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_lo_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_9};
  wire [127:0]       regroupV0_hi_lo_9 = {regroupV0_hi_lo_hi_9, regroupV0_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_6[527:526], regroupV0_hi_6[519:518]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_6[543:542], regroupV0_hi_6[535:534]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_6[559:558], regroupV0_hi_6[551:550]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_6[575:574], regroupV0_hi_6[567:566]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_6[591:590], regroupV0_hi_6[583:582]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_6[607:606], regroupV0_hi_6[599:598]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_6[623:622], regroupV0_hi_6[615:614]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_6[639:638], regroupV0_hi_6[631:630]};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_lo_9 = {regroupV0_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_6[655:654], regroupV0_hi_6[647:646]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_6[671:670], regroupV0_hi_6[663:662]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_6[687:686], regroupV0_hi_6[679:678]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_6[703:702], regroupV0_hi_6[695:694]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_6[719:718], regroupV0_hi_6[711:710]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_6[735:734], regroupV0_hi_6[727:726]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_6[751:750], regroupV0_hi_6[743:742]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_6[767:766], regroupV0_hi_6[759:758]};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_lo_hi_9 = {regroupV0_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_lo_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_9, regroupV0_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_6[783:782], regroupV0_hi_6[775:774]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_6[799:798], regroupV0_hi_6[791:790]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_6[815:814], regroupV0_hi_6[807:806]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_6[831:830], regroupV0_hi_6[823:822]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_6[847:846], regroupV0_hi_6[839:838]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_6[863:862], regroupV0_hi_6[855:854]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_6[879:878], regroupV0_hi_6[871:870]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_6[895:894], regroupV0_hi_6[887:886]};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_9};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_6[911:910], regroupV0_hi_6[903:902]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_6[927:926], regroupV0_hi_6[919:918]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_6[943:942], regroupV0_hi_6[935:934]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_6[959:958], regroupV0_hi_6[951:950]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_7};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_6[975:974], regroupV0_hi_6[967:966]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_6[991:990], regroupV0_hi_6[983:982]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_3};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_6[1007:1006], regroupV0_hi_6[999:998]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_6[1023:1022], regroupV0_hi_6[1015:1014]};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_7};
  wire [31:0]        regroupV0_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_lo_9};
  wire [63:0]        regroupV0_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_lo_9};
  wire [127:0]       regroupV0_hi_hi_9 = {regroupV0_hi_hi_hi_9, regroupV0_hi_hi_lo_9};
  wire [255:0]       regroupV0_hi_10 = {regroupV0_hi_hi_9, regroupV0_hi_lo_9};
  wire [1023:0]      regroupV0_lo_11 = {regroupV0_hi_8, regroupV0_lo_8, regroupV0_hi_7, regroupV0_lo_7};
  wire [1023:0]      regroupV0_hi_11 = {regroupV0_hi_10, regroupV0_lo_10, regroupV0_hi_9, regroupV0_lo_9};
  wire [2047:0]      regroupV0_1 = {regroupV0_hi_11, regroupV0_lo_11};
  wire [127:0]       regroupV0_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_lo_10 = {regroupV0_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_lo_10 = {regroupV0_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_lo_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_lo_hi_10 = {regroupV0_lo_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_10};
  wire [511:0]       regroupV0_lo_lo_10 = {regroupV0_lo_lo_hi_10, regroupV0_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_lo_10 = {regroupV0_lo_hi_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_lo_hi_10 = {regroupV0_lo_hi_lo_hi_hi_10, regroupV0_lo_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_lo_10 = {regroupV0_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_lo_10 = {regroupV0_lo_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_lo_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_lo_hi_hi_10 = {regroupV0_lo_hi_hi_hi_10, regroupV0_lo_hi_hi_lo_10};
  wire [511:0]       regroupV0_lo_hi_10 = {regroupV0_lo_hi_hi_10, regroupV0_lo_hi_lo_10};
  wire [1023:0]      regroupV0_lo_12 = {regroupV0_lo_hi_10, regroupV0_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_lo_hi_10 = {regroupV0_hi_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_lo_10 = {regroupV0_hi_lo_hi_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_lo_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_10};
  wire [511:0]       regroupV0_hi_lo_10 = {regroupV0_hi_lo_hi_10, regroupV0_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_lo_10 = {regroupV0_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_lo_hi_10 = {regroupV0_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_lo_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_10, regroupV0_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_10};
  wire [127:0]       regroupV0_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_lo_10};
  wire [255:0]       regroupV0_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_lo_10};
  wire [511:0]       regroupV0_hi_hi_10 = {regroupV0_hi_hi_hi_10, regroupV0_hi_hi_lo_10};
  wire [1023:0]      regroupV0_hi_12 = {regroupV0_hi_hi_10, regroupV0_hi_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[4], regroupV0_lo_12[0]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[12], regroupV0_lo_12[8]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_4 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[20], regroupV0_lo_12[16]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[28], regroupV0_lo_12[24]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_4 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_8 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_4, regroupV0_lo_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[36], regroupV0_lo_12[32]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[44], regroupV0_lo_12[40]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_4 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[52], regroupV0_lo_12[48]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[60], regroupV0_lo_12[56]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_4 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_8 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_4, regroupV0_lo_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_hi_8, regroupV0_lo_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[68], regroupV0_lo_12[64]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[76], regroupV0_lo_12[72]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_4 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[84], regroupV0_lo_12[80]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[92], regroupV0_lo_12[88]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_4 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_8 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_4, regroupV0_lo_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[100], regroupV0_lo_12[96]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[108], regroupV0_lo_12[104]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_4 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[116], regroupV0_lo_12[112]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[124], regroupV0_lo_12[120]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_4 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_8 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_4, regroupV0_lo_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_8, regroupV0_lo_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[132], regroupV0_lo_12[128]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[140], regroupV0_lo_12[136]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_4 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[148], regroupV0_lo_12[144]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[156], regroupV0_lo_12[152]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_4 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_8 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_4, regroupV0_lo_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[164], regroupV0_lo_12[160]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[172], regroupV0_lo_12[168]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_4 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[180], regroupV0_lo_12[176]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[188], regroupV0_lo_12[184]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_4 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_8 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_4, regroupV0_lo_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_hi_lo_hi_8, regroupV0_lo_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[196], regroupV0_lo_12[192]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[204], regroupV0_lo_12[200]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_4 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[212], regroupV0_lo_12[208]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[220], regroupV0_lo_12[216]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_4 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_8 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_4, regroupV0_lo_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[228], regroupV0_lo_12[224]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[236], regroupV0_lo_12[232]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_4 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[244], regroupV0_lo_12[240]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[252], regroupV0_lo_12[248]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_4 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_8 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_4, regroupV0_lo_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_8, regroupV0_lo_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_lo_11 = {regroupV0_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[260], regroupV0_lo_12[256]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[268], regroupV0_lo_12[264]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_4 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[276], regroupV0_lo_12[272]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[284], regroupV0_lo_12[280]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_4 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_8 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_4, regroupV0_lo_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[292], regroupV0_lo_12[288]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[300], regroupV0_lo_12[296]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_4 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[308], regroupV0_lo_12[304]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[316], regroupV0_lo_12[312]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_4 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_8 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_4, regroupV0_lo_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_hi_8, regroupV0_lo_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[324], regroupV0_lo_12[320]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[332], regroupV0_lo_12[328]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_4 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[340], regroupV0_lo_12[336]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[348], regroupV0_lo_12[344]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_4 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_8 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_4, regroupV0_lo_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[356], regroupV0_lo_12[352]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[364], regroupV0_lo_12[360]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_4 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[372], regroupV0_lo_12[368]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[380], regroupV0_lo_12[376]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_4 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_8 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_4, regroupV0_lo_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_8, regroupV0_lo_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[388], regroupV0_lo_12[384]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[396], regroupV0_lo_12[392]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_4 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[404], regroupV0_lo_12[400]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[412], regroupV0_lo_12[408]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_4 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_8 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_4, regroupV0_lo_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[420], regroupV0_lo_12[416]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[428], regroupV0_lo_12[424]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_4 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[436], regroupV0_lo_12[432]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[444], regroupV0_lo_12[440]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_4 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_8 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_4, regroupV0_lo_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_lo_hi_8, regroupV0_lo_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[452], regroupV0_lo_12[448]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[460], regroupV0_lo_12[456]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_4 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[468], regroupV0_lo_12[464]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[476], regroupV0_lo_12[472]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_4 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_8 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_4, regroupV0_lo_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[484], regroupV0_lo_12[480]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[492], regroupV0_lo_12[488]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_4 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[500], regroupV0_lo_12[496]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[508], regroupV0_lo_12[504]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_4 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_8 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_4, regroupV0_lo_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_8, regroupV0_lo_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_lo_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_lo_hi_11 = {regroupV0_lo_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_11};
  wire [127:0]       regroupV0_lo_lo_11 = {regroupV0_lo_lo_hi_11, regroupV0_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo = {regroupV0_lo_12[516], regroupV0_lo_12[512]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi = {regroupV0_lo_12[524], regroupV0_lo_12[520]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_4 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo = {regroupV0_lo_12[532], regroupV0_lo_12[528]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi = {regroupV0_lo_12[540], regroupV0_lo_12[536]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_4 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_8 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_4, regroupV0_lo_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo = {regroupV0_lo_12[548], regroupV0_lo_12[544]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi = {regroupV0_lo_12[556], regroupV0_lo_12[552]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_4 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo = {regroupV0_lo_12[564], regroupV0_lo_12[560]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi = {regroupV0_lo_12[572], regroupV0_lo_12[568]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_4 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_8 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_4, regroupV0_lo_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_hi_8, regroupV0_lo_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo = {regroupV0_lo_12[580], regroupV0_lo_12[576]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi = {regroupV0_lo_12[588], regroupV0_lo_12[584]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_4 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo = {regroupV0_lo_12[596], regroupV0_lo_12[592]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi = {regroupV0_lo_12[604], regroupV0_lo_12[600]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_4 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_8 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_4, regroupV0_lo_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo = {regroupV0_lo_12[612], regroupV0_lo_12[608]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi = {regroupV0_lo_12[620], regroupV0_lo_12[616]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_4 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo = {regroupV0_lo_12[628], regroupV0_lo_12[624]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi = {regroupV0_lo_12[636], regroupV0_lo_12[632]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_4 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_8 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_4, regroupV0_lo_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_8, regroupV0_lo_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo = {regroupV0_lo_12[644], regroupV0_lo_12[640]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi = {regroupV0_lo_12[652], regroupV0_lo_12[648]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_4 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo = {regroupV0_lo_12[660], regroupV0_lo_12[656]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi = {regroupV0_lo_12[668], regroupV0_lo_12[664]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_4 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_8 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_4, regroupV0_lo_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo = {regroupV0_lo_12[676], regroupV0_lo_12[672]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi = {regroupV0_lo_12[684], regroupV0_lo_12[680]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_4 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo = {regroupV0_lo_12[692], regroupV0_lo_12[688]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi = {regroupV0_lo_12[700], regroupV0_lo_12[696]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_4 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_8 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_4, regroupV0_lo_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_lo_hi_8, regroupV0_lo_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo = {regroupV0_lo_12[708], regroupV0_lo_12[704]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi = {regroupV0_lo_12[716], regroupV0_lo_12[712]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_4 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo = {regroupV0_lo_12[724], regroupV0_lo_12[720]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi = {regroupV0_lo_12[732], regroupV0_lo_12[728]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_4 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_8 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_4, regroupV0_lo_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo = {regroupV0_lo_12[740], regroupV0_lo_12[736]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi = {regroupV0_lo_12[748], regroupV0_lo_12[744]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_4 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo = {regroupV0_lo_12[756], regroupV0_lo_12[752]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi = {regroupV0_lo_12[764], regroupV0_lo_12[760]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_4 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_8 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_4, regroupV0_lo_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_8, regroupV0_lo_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_hi_11, regroupV0_lo_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_lo_11 = {regroupV0_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo = {regroupV0_lo_12[772], regroupV0_lo_12[768]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi = {regroupV0_lo_12[780], regroupV0_lo_12[776]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_4 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo = {regroupV0_lo_12[788], regroupV0_lo_12[784]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi = {regroupV0_lo_12[796], regroupV0_lo_12[792]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_4 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_8 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_4, regroupV0_lo_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo = {regroupV0_lo_12[804], regroupV0_lo_12[800]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi = {regroupV0_lo_12[812], regroupV0_lo_12[808]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_4 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo = {regroupV0_lo_12[820], regroupV0_lo_12[816]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi = {regroupV0_lo_12[828], regroupV0_lo_12[824]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_4 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_8 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_4, regroupV0_lo_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_hi_8, regroupV0_lo_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo = {regroupV0_lo_12[836], regroupV0_lo_12[832]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi = {regroupV0_lo_12[844], regroupV0_lo_12[840]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_4 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo = {regroupV0_lo_12[852], regroupV0_lo_12[848]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi = {regroupV0_lo_12[860], regroupV0_lo_12[856]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_4 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_8 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_4, regroupV0_lo_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo = {regroupV0_lo_12[868], regroupV0_lo_12[864]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi = {regroupV0_lo_12[876], regroupV0_lo_12[872]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_4 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo = {regroupV0_lo_12[884], regroupV0_lo_12[880]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi = {regroupV0_lo_12[892], regroupV0_lo_12[888]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_4 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_8 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_4, regroupV0_lo_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_8, regroupV0_lo_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo = {regroupV0_lo_12[900], regroupV0_lo_12[896]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi = {regroupV0_lo_12[908], regroupV0_lo_12[904]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_4 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo = {regroupV0_lo_12[916], regroupV0_lo_12[912]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi = {regroupV0_lo_12[924], regroupV0_lo_12[920]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_4 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_8 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_4, regroupV0_lo_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo = {regroupV0_lo_12[932], regroupV0_lo_12[928]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi = {regroupV0_lo_12[940], regroupV0_lo_12[936]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_4 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo = {regroupV0_lo_12[948], regroupV0_lo_12[944]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi = {regroupV0_lo_12[956], regroupV0_lo_12[952]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_4 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_8 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_4, regroupV0_lo_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_lo_hi_8, regroupV0_lo_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo = {regroupV0_lo_12[964], regroupV0_lo_12[960]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi = {regroupV0_lo_12[972], regroupV0_lo_12[968]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_4 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo = {regroupV0_lo_12[980], regroupV0_lo_12[976]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi = {regroupV0_lo_12[988], regroupV0_lo_12[984]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_4 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_8 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_4, regroupV0_lo_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo = {regroupV0_lo_12[996], regroupV0_lo_12[992]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi = {regroupV0_lo_12[1004], regroupV0_lo_12[1000]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_4 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo = {regroupV0_lo_12[1012], regroupV0_lo_12[1008]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi = {regroupV0_lo_12[1020], regroupV0_lo_12[1016]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_4 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_8 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_4, regroupV0_lo_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_8, regroupV0_lo_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_lo_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_lo_hi_hi_11 = {regroupV0_lo_hi_hi_hi_11, regroupV0_lo_hi_hi_lo_11};
  wire [127:0]       regroupV0_lo_hi_11 = {regroupV0_lo_hi_hi_11, regroupV0_lo_hi_lo_11};
  wire [255:0]       regroupV0_lo_13 = {regroupV0_lo_hi_11, regroupV0_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[4], regroupV0_hi_12[0]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[12], regroupV0_hi_12[8]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_4 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[20], regroupV0_hi_12[16]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[28], regroupV0_hi_12[24]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_4 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_8 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_4, regroupV0_hi_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[36], regroupV0_hi_12[32]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[44], regroupV0_hi_12[40]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_4 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[52], regroupV0_hi_12[48]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[60], regroupV0_hi_12[56]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_4 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_8 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_4, regroupV0_hi_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_hi_8, regroupV0_hi_lo_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[68], regroupV0_hi_12[64]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[76], regroupV0_hi_12[72]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_4 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[84], regroupV0_hi_12[80]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[92], regroupV0_hi_12[88]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_4 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_8 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_4, regroupV0_hi_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[100], regroupV0_hi_12[96]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[108], regroupV0_hi_12[104]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_4 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[116], regroupV0_hi_12[112]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[124], regroupV0_hi_12[120]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_4 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_8 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_4, regroupV0_hi_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_8, regroupV0_hi_lo_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[132], regroupV0_hi_12[128]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[140], regroupV0_hi_12[136]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_4 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[148], regroupV0_hi_12[144]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[156], regroupV0_hi_12[152]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_4 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_8 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_4, regroupV0_hi_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[164], regroupV0_hi_12[160]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[172], regroupV0_hi_12[168]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_4 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[180], regroupV0_hi_12[176]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[188], regroupV0_hi_12[184]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_4 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_8 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_4, regroupV0_hi_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_hi_lo_hi_8, regroupV0_hi_lo_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[196], regroupV0_hi_12[192]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[204], regroupV0_hi_12[200]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_4 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[212], regroupV0_hi_12[208]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[220], regroupV0_hi_12[216]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_4 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_8 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_4, regroupV0_hi_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[228], regroupV0_hi_12[224]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[236], regroupV0_hi_12[232]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_4 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[244], regroupV0_hi_12[240]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[252], regroupV0_hi_12[248]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_4 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_8 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_4, regroupV0_hi_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_8, regroupV0_hi_lo_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_lo_hi_11 = {regroupV0_hi_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[260], regroupV0_hi_12[256]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[268], regroupV0_hi_12[264]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_4 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[276], regroupV0_hi_12[272]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[284], regroupV0_hi_12[280]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_4 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_8 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_4, regroupV0_hi_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[292], regroupV0_hi_12[288]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[300], regroupV0_hi_12[296]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_4 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[308], regroupV0_hi_12[304]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[316], regroupV0_hi_12[312]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_4 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_8 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_4, regroupV0_hi_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_hi_8, regroupV0_hi_lo_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[324], regroupV0_hi_12[320]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[332], regroupV0_hi_12[328]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_4 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[340], regroupV0_hi_12[336]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[348], regroupV0_hi_12[344]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_4 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_8 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_4, regroupV0_hi_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[356], regroupV0_hi_12[352]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[364], regroupV0_hi_12[360]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_4 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[372], regroupV0_hi_12[368]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[380], regroupV0_hi_12[376]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_4 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_8 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_4, regroupV0_hi_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_8, regroupV0_hi_lo_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[388], regroupV0_hi_12[384]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[396], regroupV0_hi_12[392]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_4 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[404], regroupV0_hi_12[400]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[412], regroupV0_hi_12[408]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_4 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_8 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_4, regroupV0_hi_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[420], regroupV0_hi_12[416]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[428], regroupV0_hi_12[424]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_4 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[436], regroupV0_hi_12[432]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[444], regroupV0_hi_12[440]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_4 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_8 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_4, regroupV0_hi_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_lo_hi_8, regroupV0_hi_lo_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[452], regroupV0_hi_12[448]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[460], regroupV0_hi_12[456]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_4 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[468], regroupV0_hi_12[464]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[476], regroupV0_hi_12[472]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_4 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_8 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_4, regroupV0_hi_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[484], regroupV0_hi_12[480]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[492], regroupV0_hi_12[488]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_4 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[500], regroupV0_hi_12[496]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[508], regroupV0_hi_12[504]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_4 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_8 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_4, regroupV0_hi_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_8, regroupV0_hi_lo_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_11};
  wire [127:0]       regroupV0_hi_lo_11 = {regroupV0_hi_lo_hi_11, regroupV0_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo = {regroupV0_hi_12[516], regroupV0_hi_12[512]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi = {regroupV0_hi_12[524], regroupV0_hi_12[520]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_4 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo = {regroupV0_hi_12[532], regroupV0_hi_12[528]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi = {regroupV0_hi_12[540], regroupV0_hi_12[536]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_4 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_8 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_4, regroupV0_hi_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo = {regroupV0_hi_12[548], regroupV0_hi_12[544]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi = {regroupV0_hi_12[556], regroupV0_hi_12[552]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_4 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo = {regroupV0_hi_12[564], regroupV0_hi_12[560]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi = {regroupV0_hi_12[572], regroupV0_hi_12[568]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_4 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_8 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_4, regroupV0_hi_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_hi_8, regroupV0_hi_hi_lo_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo = {regroupV0_hi_12[580], regroupV0_hi_12[576]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi = {regroupV0_hi_12[588], regroupV0_hi_12[584]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_4 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo = {regroupV0_hi_12[596], regroupV0_hi_12[592]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi = {regroupV0_hi_12[604], regroupV0_hi_12[600]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_4 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_8 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_4, regroupV0_hi_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo = {regroupV0_hi_12[612], regroupV0_hi_12[608]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi = {regroupV0_hi_12[620], regroupV0_hi_12[616]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_4 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo = {regroupV0_hi_12[628], regroupV0_hi_12[624]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi = {regroupV0_hi_12[636], regroupV0_hi_12[632]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_4 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_8 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_4, regroupV0_hi_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_8, regroupV0_hi_hi_lo_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_lo_11 = {regroupV0_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo = {regroupV0_hi_12[644], regroupV0_hi_12[640]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi = {regroupV0_hi_12[652], regroupV0_hi_12[648]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_4 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo = {regroupV0_hi_12[660], regroupV0_hi_12[656]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi = {regroupV0_hi_12[668], regroupV0_hi_12[664]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_4 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_8 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_4, regroupV0_hi_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo = {regroupV0_hi_12[676], regroupV0_hi_12[672]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi = {regroupV0_hi_12[684], regroupV0_hi_12[680]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_4 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo = {regroupV0_hi_12[692], regroupV0_hi_12[688]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi = {regroupV0_hi_12[700], regroupV0_hi_12[696]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_4 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_8 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_4, regroupV0_hi_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_lo_hi_lo_hi_8, regroupV0_hi_hi_lo_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo = {regroupV0_hi_12[708], regroupV0_hi_12[704]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi = {regroupV0_hi_12[716], regroupV0_hi_12[712]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_4 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo = {regroupV0_hi_12[724], regroupV0_hi_12[720]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi = {regroupV0_hi_12[732], regroupV0_hi_12[728]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_4 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_8 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_4, regroupV0_hi_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo = {regroupV0_hi_12[740], regroupV0_hi_12[736]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi = {regroupV0_hi_12[748], regroupV0_hi_12[744]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_4 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo = {regroupV0_hi_12[756], regroupV0_hi_12[752]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi = {regroupV0_hi_12[764], regroupV0_hi_12[760]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_4 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_8 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_4, regroupV0_hi_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_8, regroupV0_hi_hi_lo_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_lo_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_11, regroupV0_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo = {regroupV0_hi_12[772], regroupV0_hi_12[768]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi = {regroupV0_hi_12[780], regroupV0_hi_12[776]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_4 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo = {regroupV0_hi_12[788], regroupV0_hi_12[784]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi = {regroupV0_hi_12[796], regroupV0_hi_12[792]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_4 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_8 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_4, regroupV0_hi_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo = {regroupV0_hi_12[804], regroupV0_hi_12[800]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi = {regroupV0_hi_12[812], regroupV0_hi_12[808]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_4 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo = {regroupV0_hi_12[820], regroupV0_hi_12[816]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi = {regroupV0_hi_12[828], regroupV0_hi_12[824]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_4 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_8 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_4, regroupV0_hi_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_hi_8, regroupV0_hi_hi_hi_lo_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo = {regroupV0_hi_12[836], regroupV0_hi_12[832]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi = {regroupV0_hi_12[844], regroupV0_hi_12[840]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_4 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo = {regroupV0_hi_12[852], regroupV0_hi_12[848]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi = {regroupV0_hi_12[860], regroupV0_hi_12[856]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_4 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_8 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_4, regroupV0_hi_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo = {regroupV0_hi_12[868], regroupV0_hi_12[864]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi = {regroupV0_hi_12[876], regroupV0_hi_12[872]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_4 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo = {regroupV0_hi_12[884], regroupV0_hi_12[880]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi = {regroupV0_hi_12[892], regroupV0_hi_12[888]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_4 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_8 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_4, regroupV0_hi_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_8, regroupV0_hi_hi_hi_lo_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo = {regroupV0_hi_12[900], regroupV0_hi_12[896]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi = {regroupV0_hi_12[908], regroupV0_hi_12[904]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_4 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo = {regroupV0_hi_12[916], regroupV0_hi_12[912]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi = {regroupV0_hi_12[924], regroupV0_hi_12[920]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_4 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_8 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_4, regroupV0_hi_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo = {regroupV0_hi_12[932], regroupV0_hi_12[928]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi = {regroupV0_hi_12[940], regroupV0_hi_12[936]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_4 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo = {regroupV0_hi_12[948], regroupV0_hi_12[944]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi = {regroupV0_hi_12[956], regroupV0_hi_12[952]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_4 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_8 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_4, regroupV0_hi_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_lo_hi_8, regroupV0_hi_hi_hi_hi_lo_lo_8};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo = {regroupV0_hi_12[964], regroupV0_hi_12[960]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi = {regroupV0_hi_12[972], regroupV0_hi_12[968]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_4 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo = {regroupV0_hi_12[980], regroupV0_hi_12[976]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi = {regroupV0_hi_12[988], regroupV0_hi_12[984]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_4 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_8 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_4, regroupV0_hi_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo = {regroupV0_hi_12[996], regroupV0_hi_12[992]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi = {regroupV0_hi_12[1004], regroupV0_hi_12[1000]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_4 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo = {regroupV0_hi_12[1012], regroupV0_hi_12[1008]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi = {regroupV0_hi_12[1020], regroupV0_hi_12[1016]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_4 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_8 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_4, regroupV0_hi_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_8, regroupV0_hi_hi_hi_hi_hi_lo_8};
  wire [31:0]        regroupV0_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_lo_11};
  wire [63:0]        regroupV0_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_lo_11};
  wire [127:0]       regroupV0_hi_hi_11 = {regroupV0_hi_hi_hi_11, regroupV0_hi_hi_lo_11};
  wire [255:0]       regroupV0_hi_13 = {regroupV0_hi_hi_11, regroupV0_hi_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[5], regroupV0_lo_12[1]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[13], regroupV0_lo_12[9]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_5 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[21], regroupV0_lo_12[17]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[29], regroupV0_lo_12[25]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_5 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_9 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_5, regroupV0_lo_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[37], regroupV0_lo_12[33]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[45], regroupV0_lo_12[41]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_5 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[53], regroupV0_lo_12[49]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[61], regroupV0_lo_12[57]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_5 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_9 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_5, regroupV0_lo_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_lo_hi_9, regroupV0_lo_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[69], regroupV0_lo_12[65]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[77], regroupV0_lo_12[73]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_5 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[85], regroupV0_lo_12[81]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[93], regroupV0_lo_12[89]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_5 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_9 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_5, regroupV0_lo_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[101], regroupV0_lo_12[97]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[109], regroupV0_lo_12[105]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_5 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[117], regroupV0_lo_12[113]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[125], regroupV0_lo_12[121]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_5 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_9 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_5, regroupV0_lo_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_lo_hi_hi_9, regroupV0_lo_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_lo_12 = {regroupV0_lo_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[133], regroupV0_lo_12[129]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[141], regroupV0_lo_12[137]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_5 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[149], regroupV0_lo_12[145]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[157], regroupV0_lo_12[153]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_5 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_9 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_5, regroupV0_lo_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[165], regroupV0_lo_12[161]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[173], regroupV0_lo_12[169]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_5 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[181], regroupV0_lo_12[177]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[189], regroupV0_lo_12[185]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_5 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_9 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_5, regroupV0_lo_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_12 = {regroupV0_lo_lo_lo_hi_lo_hi_9, regroupV0_lo_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[197], regroupV0_lo_12[193]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[205], regroupV0_lo_12[201]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_5 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[213], regroupV0_lo_12[209]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[221], regroupV0_lo_12[217]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_5 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_9 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_5, regroupV0_lo_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[229], regroupV0_lo_12[225]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[237], regroupV0_lo_12[233]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_5 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[245], regroupV0_lo_12[241]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[253], regroupV0_lo_12[249]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_5 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_9 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_5, regroupV0_lo_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_12 = {regroupV0_lo_lo_lo_hi_hi_hi_9, regroupV0_lo_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_lo_hi_12 = {regroupV0_lo_lo_lo_hi_hi_12, regroupV0_lo_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_lo_12 = {regroupV0_lo_lo_lo_hi_12, regroupV0_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[261], regroupV0_lo_12[257]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[269], regroupV0_lo_12[265]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_5 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[277], regroupV0_lo_12[273]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[285], regroupV0_lo_12[281]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_5 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_9 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_5, regroupV0_lo_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[293], regroupV0_lo_12[289]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[301], regroupV0_lo_12[297]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_5 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[309], regroupV0_lo_12[305]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[317], regroupV0_lo_12[313]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_5 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_9 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_5, regroupV0_lo_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_12 = {regroupV0_lo_lo_hi_lo_lo_hi_9, regroupV0_lo_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[325], regroupV0_lo_12[321]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[333], regroupV0_lo_12[329]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_5 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[341], regroupV0_lo_12[337]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[349], regroupV0_lo_12[345]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_5 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_9 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_5, regroupV0_lo_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[357], regroupV0_lo_12[353]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[365], regroupV0_lo_12[361]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_5 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[373], regroupV0_lo_12[369]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[381], regroupV0_lo_12[377]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_5 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_9 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_5, regroupV0_lo_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_12 = {regroupV0_lo_lo_hi_lo_hi_hi_9, regroupV0_lo_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_lo_12 = {regroupV0_lo_lo_hi_lo_hi_12, regroupV0_lo_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[389], regroupV0_lo_12[385]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[397], regroupV0_lo_12[393]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_5 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[405], regroupV0_lo_12[401]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[413], regroupV0_lo_12[409]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_5 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_9 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_5, regroupV0_lo_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[421], regroupV0_lo_12[417]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[429], regroupV0_lo_12[425]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_5 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[437], regroupV0_lo_12[433]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[445], regroupV0_lo_12[441]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_5 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_9 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_5, regroupV0_lo_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_12 = {regroupV0_lo_lo_hi_hi_lo_hi_9, regroupV0_lo_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[453], regroupV0_lo_12[449]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[461], regroupV0_lo_12[457]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_5 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[469], regroupV0_lo_12[465]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[477], regroupV0_lo_12[473]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_5 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_9 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_5, regroupV0_lo_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[485], regroupV0_lo_12[481]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[493], regroupV0_lo_12[489]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_5 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[501], regroupV0_lo_12[497]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[509], regroupV0_lo_12[505]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_5 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_9 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_5, regroupV0_lo_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_hi_9, regroupV0_lo_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_lo_hi_hi_12 = {regroupV0_lo_lo_hi_hi_hi_12, regroupV0_lo_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_lo_hi_12 = {regroupV0_lo_lo_hi_hi_12, regroupV0_lo_lo_hi_lo_12};
  wire [127:0]       regroupV0_lo_lo_12 = {regroupV0_lo_lo_hi_12, regroupV0_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[517], regroupV0_lo_12[513]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[525], regroupV0_lo_12[521]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_5 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[533], regroupV0_lo_12[529]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[541], regroupV0_lo_12[537]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_5 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_9 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_5, regroupV0_lo_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[549], regroupV0_lo_12[545]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[557], regroupV0_lo_12[553]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_5 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[565], regroupV0_lo_12[561]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[573], regroupV0_lo_12[569]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_5 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_9 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_5, regroupV0_lo_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_12 = {regroupV0_lo_hi_lo_lo_lo_hi_9, regroupV0_lo_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[581], regroupV0_lo_12[577]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[589], regroupV0_lo_12[585]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_5 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[597], regroupV0_lo_12[593]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[605], regroupV0_lo_12[601]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_5 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_9 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_5, regroupV0_lo_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[613], regroupV0_lo_12[609]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[621], regroupV0_lo_12[617]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_5 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[629], regroupV0_lo_12[625]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[637], regroupV0_lo_12[633]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_5 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_9 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_5, regroupV0_lo_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_12 = {regroupV0_lo_hi_lo_lo_hi_hi_9, regroupV0_lo_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_lo_12 = {regroupV0_lo_hi_lo_lo_hi_12, regroupV0_lo_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[645], regroupV0_lo_12[641]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[653], regroupV0_lo_12[649]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_5 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[661], regroupV0_lo_12[657]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[669], regroupV0_lo_12[665]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_5 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_9 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_5, regroupV0_lo_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[677], regroupV0_lo_12[673]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[685], regroupV0_lo_12[681]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_5 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[693], regroupV0_lo_12[689]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[701], regroupV0_lo_12[697]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_5 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_9 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_5, regroupV0_lo_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_12 = {regroupV0_lo_hi_lo_hi_lo_hi_9, regroupV0_lo_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[709], regroupV0_lo_12[705]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[717], regroupV0_lo_12[713]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_5 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[725], regroupV0_lo_12[721]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[733], regroupV0_lo_12[729]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_5 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_9 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_5, regroupV0_lo_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[741], regroupV0_lo_12[737]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[749], regroupV0_lo_12[745]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_5 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[757], regroupV0_lo_12[753]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[765], regroupV0_lo_12[761]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_5 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_9 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_5, regroupV0_lo_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_12 = {regroupV0_lo_hi_lo_hi_hi_hi_9, regroupV0_lo_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_lo_hi_12 = {regroupV0_lo_hi_lo_hi_hi_12, regroupV0_lo_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_lo_12 = {regroupV0_lo_hi_lo_hi_12, regroupV0_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_lo_12[773], regroupV0_lo_12[769]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_lo_12[781], regroupV0_lo_12[777]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_5 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_lo_12[789], regroupV0_lo_12[785]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_lo_12[797], regroupV0_lo_12[793]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_5 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_9 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_5, regroupV0_lo_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_lo_12[805], regroupV0_lo_12[801]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_lo_12[813], regroupV0_lo_12[809]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_5 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_lo_12[821], regroupV0_lo_12[817]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_lo_12[829], regroupV0_lo_12[825]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_5 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_9 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_5, regroupV0_lo_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_12 = {regroupV0_lo_hi_hi_lo_lo_hi_9, regroupV0_lo_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_lo_12[837], regroupV0_lo_12[833]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_lo_12[845], regroupV0_lo_12[841]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_5 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_lo_12[853], regroupV0_lo_12[849]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_lo_12[861], regroupV0_lo_12[857]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_5 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_9 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_5, regroupV0_lo_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_lo_12[869], regroupV0_lo_12[865]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_lo_12[877], regroupV0_lo_12[873]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_5 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_lo_12[885], regroupV0_lo_12[881]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_lo_12[893], regroupV0_lo_12[889]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_5 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_9 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_5, regroupV0_lo_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_12 = {regroupV0_lo_hi_hi_lo_hi_hi_9, regroupV0_lo_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_lo_12 = {regroupV0_lo_hi_hi_lo_hi_12, regroupV0_lo_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_lo_12[901], regroupV0_lo_12[897]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_lo_12[909], regroupV0_lo_12[905]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_5 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_lo_12[917], regroupV0_lo_12[913]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_lo_12[925], regroupV0_lo_12[921]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_5 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_9 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_5, regroupV0_lo_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_lo_12[933], regroupV0_lo_12[929]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_lo_12[941], regroupV0_lo_12[937]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_5 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_lo_12[949], regroupV0_lo_12[945]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_lo_12[957], regroupV0_lo_12[953]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_5 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_9 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_5, regroupV0_lo_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_12 = {regroupV0_lo_hi_hi_hi_lo_hi_9, regroupV0_lo_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_lo_12[965], regroupV0_lo_12[961]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_lo_12[973], regroupV0_lo_12[969]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_5 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_lo_12[981], regroupV0_lo_12[977]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_lo_12[989], regroupV0_lo_12[985]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_5 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_9 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_5, regroupV0_lo_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_lo_12[997], regroupV0_lo_12[993]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_lo_12[1005], regroupV0_lo_12[1001]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_5 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_lo_12[1013], regroupV0_lo_12[1009]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_lo_12[1021], regroupV0_lo_12[1017]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_5 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_9 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_5, regroupV0_lo_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_hi_9, regroupV0_lo_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_lo_hi_hi_hi_12 = {regroupV0_lo_hi_hi_hi_hi_12, regroupV0_lo_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_lo_hi_hi_12 = {regroupV0_lo_hi_hi_hi_12, regroupV0_lo_hi_hi_lo_12};
  wire [127:0]       regroupV0_lo_hi_12 = {regroupV0_lo_hi_hi_12, regroupV0_lo_hi_lo_12};
  wire [255:0]       regroupV0_lo_14 = {regroupV0_lo_hi_12, regroupV0_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[5], regroupV0_hi_12[1]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[13], regroupV0_hi_12[9]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_5 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[21], regroupV0_hi_12[17]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[29], regroupV0_hi_12[25]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_5 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_9 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_5, regroupV0_hi_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[37], regroupV0_hi_12[33]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[45], regroupV0_hi_12[41]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_5 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[53], regroupV0_hi_12[49]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[61], regroupV0_hi_12[57]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_5 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_9 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_5, regroupV0_hi_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_lo_hi_9, regroupV0_hi_lo_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[69], regroupV0_hi_12[65]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[77], regroupV0_hi_12[73]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_5 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[85], regroupV0_hi_12[81]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[93], regroupV0_hi_12[89]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_5 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_9 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_5, regroupV0_hi_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[101], regroupV0_hi_12[97]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[109], regroupV0_hi_12[105]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_5 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[117], regroupV0_hi_12[113]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[125], regroupV0_hi_12[121]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_5 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_9 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_5, regroupV0_hi_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_12 = {regroupV0_hi_lo_lo_lo_hi_hi_9, regroupV0_hi_lo_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_lo_12 = {regroupV0_hi_lo_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[133], regroupV0_hi_12[129]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[141], regroupV0_hi_12[137]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_5 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[149], regroupV0_hi_12[145]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[157], regroupV0_hi_12[153]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_5 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_9 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_5, regroupV0_hi_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[165], regroupV0_hi_12[161]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[173], regroupV0_hi_12[169]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_5 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[181], regroupV0_hi_12[177]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[189], regroupV0_hi_12[185]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_5 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_9 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_5, regroupV0_hi_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_12 = {regroupV0_hi_lo_lo_hi_lo_hi_9, regroupV0_hi_lo_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[197], regroupV0_hi_12[193]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[205], regroupV0_hi_12[201]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_5 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[213], regroupV0_hi_12[209]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[221], regroupV0_hi_12[217]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_5 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_9 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_5, regroupV0_hi_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[229], regroupV0_hi_12[225]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[237], regroupV0_hi_12[233]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_5 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[245], regroupV0_hi_12[241]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[253], regroupV0_hi_12[249]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_5 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_9 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_5, regroupV0_hi_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_12 = {regroupV0_hi_lo_lo_hi_hi_hi_9, regroupV0_hi_lo_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_lo_hi_12 = {regroupV0_hi_lo_lo_hi_hi_12, regroupV0_hi_lo_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_lo_12 = {regroupV0_hi_lo_lo_hi_12, regroupV0_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[261], regroupV0_hi_12[257]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[269], regroupV0_hi_12[265]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_5 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[277], regroupV0_hi_12[273]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[285], regroupV0_hi_12[281]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_5 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_9 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_5, regroupV0_hi_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[293], regroupV0_hi_12[289]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[301], regroupV0_hi_12[297]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_5 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[309], regroupV0_hi_12[305]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[317], regroupV0_hi_12[313]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_5 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_9 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_5, regroupV0_hi_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_12 = {regroupV0_hi_lo_hi_lo_lo_hi_9, regroupV0_hi_lo_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[325], regroupV0_hi_12[321]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[333], regroupV0_hi_12[329]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_5 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[341], regroupV0_hi_12[337]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[349], regroupV0_hi_12[345]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_5 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_9 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_5, regroupV0_hi_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[357], regroupV0_hi_12[353]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[365], regroupV0_hi_12[361]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_5 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[373], regroupV0_hi_12[369]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[381], regroupV0_hi_12[377]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_5 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_9 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_5, regroupV0_hi_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_12 = {regroupV0_hi_lo_hi_lo_hi_hi_9, regroupV0_hi_lo_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_lo_12 = {regroupV0_hi_lo_hi_lo_hi_12, regroupV0_hi_lo_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[389], regroupV0_hi_12[385]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[397], regroupV0_hi_12[393]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_5 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[405], regroupV0_hi_12[401]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[413], regroupV0_hi_12[409]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_5 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_9 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_5, regroupV0_hi_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[421], regroupV0_hi_12[417]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[429], regroupV0_hi_12[425]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_5 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[437], regroupV0_hi_12[433]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[445], regroupV0_hi_12[441]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_5 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_9 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_5, regroupV0_hi_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_12 = {regroupV0_hi_lo_hi_hi_lo_hi_9, regroupV0_hi_lo_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[453], regroupV0_hi_12[449]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[461], regroupV0_hi_12[457]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_5 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[469], regroupV0_hi_12[465]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[477], regroupV0_hi_12[473]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_5 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_9 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_5, regroupV0_hi_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[485], regroupV0_hi_12[481]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[493], regroupV0_hi_12[489]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_5 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[501], regroupV0_hi_12[497]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[509], regroupV0_hi_12[505]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_5 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_9 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_5, regroupV0_hi_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_hi_9, regroupV0_hi_lo_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_lo_hi_hi_12 = {regroupV0_hi_lo_hi_hi_hi_12, regroupV0_hi_lo_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_lo_hi_12 = {regroupV0_hi_lo_hi_hi_12, regroupV0_hi_lo_hi_lo_12};
  wire [127:0]       regroupV0_hi_lo_12 = {regroupV0_hi_lo_hi_12, regroupV0_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[517], regroupV0_hi_12[513]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[525], regroupV0_hi_12[521]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_5 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[533], regroupV0_hi_12[529]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[541], regroupV0_hi_12[537]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_5 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_9 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_5, regroupV0_hi_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[549], regroupV0_hi_12[545]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[557], regroupV0_hi_12[553]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_5 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[565], regroupV0_hi_12[561]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[573], regroupV0_hi_12[569]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_5 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_9 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_5, regroupV0_hi_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_12 = {regroupV0_hi_hi_lo_lo_lo_hi_9, regroupV0_hi_hi_lo_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[581], regroupV0_hi_12[577]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[589], regroupV0_hi_12[585]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_5 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[597], regroupV0_hi_12[593]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[605], regroupV0_hi_12[601]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_5 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_9 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_5, regroupV0_hi_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[613], regroupV0_hi_12[609]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[621], regroupV0_hi_12[617]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_5 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[629], regroupV0_hi_12[625]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[637], regroupV0_hi_12[633]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_5 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_9 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_5, regroupV0_hi_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_12 = {regroupV0_hi_hi_lo_lo_hi_hi_9, regroupV0_hi_hi_lo_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_lo_12 = {regroupV0_hi_hi_lo_lo_hi_12, regroupV0_hi_hi_lo_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[645], regroupV0_hi_12[641]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[653], regroupV0_hi_12[649]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_5 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[661], regroupV0_hi_12[657]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[669], regroupV0_hi_12[665]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_5 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_9 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_5, regroupV0_hi_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[677], regroupV0_hi_12[673]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[685], regroupV0_hi_12[681]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_5 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[693], regroupV0_hi_12[689]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[701], regroupV0_hi_12[697]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_5 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_9 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_5, regroupV0_hi_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_12 = {regroupV0_hi_hi_lo_hi_lo_hi_9, regroupV0_hi_hi_lo_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[709], regroupV0_hi_12[705]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[717], regroupV0_hi_12[713]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_5 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[725], regroupV0_hi_12[721]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[733], regroupV0_hi_12[729]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_5 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_9 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_5, regroupV0_hi_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[741], regroupV0_hi_12[737]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[749], regroupV0_hi_12[745]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_5 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[757], regroupV0_hi_12[753]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[765], regroupV0_hi_12[761]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_5 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_9 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_5, regroupV0_hi_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_12 = {regroupV0_hi_hi_lo_hi_hi_hi_9, regroupV0_hi_hi_lo_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_lo_hi_12 = {regroupV0_hi_hi_lo_hi_hi_12, regroupV0_hi_hi_lo_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_lo_12 = {regroupV0_hi_hi_lo_hi_12, regroupV0_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_1 = {regroupV0_hi_12[773], regroupV0_hi_12[769]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_1 = {regroupV0_hi_12[781], regroupV0_hi_12[777]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_5 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_1 = {regroupV0_hi_12[789], regroupV0_hi_12[785]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_1 = {regroupV0_hi_12[797], regroupV0_hi_12[793]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_5 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_9 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_5, regroupV0_hi_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_1 = {regroupV0_hi_12[805], regroupV0_hi_12[801]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_1 = {regroupV0_hi_12[813], regroupV0_hi_12[809]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_5 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_1 = {regroupV0_hi_12[821], regroupV0_hi_12[817]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_1 = {regroupV0_hi_12[829], regroupV0_hi_12[825]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_5 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_9 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_5, regroupV0_hi_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_12 = {regroupV0_hi_hi_hi_lo_lo_hi_9, regroupV0_hi_hi_hi_lo_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_1 = {regroupV0_hi_12[837], regroupV0_hi_12[833]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_1 = {regroupV0_hi_12[845], regroupV0_hi_12[841]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_5 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_1 = {regroupV0_hi_12[853], regroupV0_hi_12[849]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_1 = {regroupV0_hi_12[861], regroupV0_hi_12[857]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_5 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_9 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_5, regroupV0_hi_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_1 = {regroupV0_hi_12[869], regroupV0_hi_12[865]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_1 = {regroupV0_hi_12[877], regroupV0_hi_12[873]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_5 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_1 = {regroupV0_hi_12[885], regroupV0_hi_12[881]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_1 = {regroupV0_hi_12[893], regroupV0_hi_12[889]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_5 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_9 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_5, regroupV0_hi_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_12 = {regroupV0_hi_hi_hi_lo_hi_hi_9, regroupV0_hi_hi_hi_lo_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_lo_hi_12, regroupV0_hi_hi_hi_lo_lo_12};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_1 = {regroupV0_hi_12[901], regroupV0_hi_12[897]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_1 = {regroupV0_hi_12[909], regroupV0_hi_12[905]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_5 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_1 = {regroupV0_hi_12[917], regroupV0_hi_12[913]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_1 = {regroupV0_hi_12[925], regroupV0_hi_12[921]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_5 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_9 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_5, regroupV0_hi_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_1 = {regroupV0_hi_12[933], regroupV0_hi_12[929]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_1 = {regroupV0_hi_12[941], regroupV0_hi_12[937]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_5 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_1 = {regroupV0_hi_12[949], regroupV0_hi_12[945]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_1 = {regroupV0_hi_12[957], regroupV0_hi_12[953]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_5 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_9 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_5, regroupV0_hi_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_12 = {regroupV0_hi_hi_hi_hi_lo_hi_9, regroupV0_hi_hi_hi_hi_lo_lo_9};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_1 = {regroupV0_hi_12[965], regroupV0_hi_12[961]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_1 = {regroupV0_hi_12[973], regroupV0_hi_12[969]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_5 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_1 = {regroupV0_hi_12[981], regroupV0_hi_12[977]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_1 = {regroupV0_hi_12[989], regroupV0_hi_12[985]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_5 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_9 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_5, regroupV0_hi_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_1 = {regroupV0_hi_12[997], regroupV0_hi_12[993]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_1 = {regroupV0_hi_12[1005], regroupV0_hi_12[1001]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_5 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_1 = {regroupV0_hi_12[1013], regroupV0_hi_12[1009]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_1 = {regroupV0_hi_12[1021], regroupV0_hi_12[1017]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_5 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_1, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_9 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_5, regroupV0_hi_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_hi_9, regroupV0_hi_hi_hi_hi_hi_lo_9};
  wire [31:0]        regroupV0_hi_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_hi_lo_12};
  wire [63:0]        regroupV0_hi_hi_hi_12 = {regroupV0_hi_hi_hi_hi_12, regroupV0_hi_hi_hi_lo_12};
  wire [127:0]       regroupV0_hi_hi_12 = {regroupV0_hi_hi_hi_12, regroupV0_hi_hi_lo_12};
  wire [255:0]       regroupV0_hi_14 = {regroupV0_hi_hi_12, regroupV0_hi_lo_12};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[6], regroupV0_lo_12[2]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[14], regroupV0_lo_12[10]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_6 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[22], regroupV0_lo_12[18]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[30], regroupV0_lo_12[26]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_6 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_10 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_6, regroupV0_lo_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[38], regroupV0_lo_12[34]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[46], regroupV0_lo_12[42]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_6 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[54], regroupV0_lo_12[50]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[62], regroupV0_lo_12[58]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_6 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_10 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_6, regroupV0_lo_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_lo_hi_10, regroupV0_lo_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[70], regroupV0_lo_12[66]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[78], regroupV0_lo_12[74]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_6 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[86], regroupV0_lo_12[82]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[94], regroupV0_lo_12[90]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_6 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_10 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_6, regroupV0_lo_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[102], regroupV0_lo_12[98]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[110], regroupV0_lo_12[106]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_6 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[118], regroupV0_lo_12[114]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[126], regroupV0_lo_12[122]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_6 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_10 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_6, regroupV0_lo_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_lo_hi_hi_10, regroupV0_lo_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_lo_13 = {regroupV0_lo_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[134], regroupV0_lo_12[130]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[142], regroupV0_lo_12[138]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_6 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[150], regroupV0_lo_12[146]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[158], regroupV0_lo_12[154]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_6 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_10 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_6, regroupV0_lo_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[166], regroupV0_lo_12[162]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[174], regroupV0_lo_12[170]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_6 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[182], regroupV0_lo_12[178]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[190], regroupV0_lo_12[186]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_6 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_10 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_6, regroupV0_lo_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_13 = {regroupV0_lo_lo_lo_hi_lo_hi_10, regroupV0_lo_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[198], regroupV0_lo_12[194]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[206], regroupV0_lo_12[202]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_6 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[214], regroupV0_lo_12[210]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[222], regroupV0_lo_12[218]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_6 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_10 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_6, regroupV0_lo_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[230], regroupV0_lo_12[226]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[238], regroupV0_lo_12[234]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_6 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[246], regroupV0_lo_12[242]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[254], regroupV0_lo_12[250]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_6 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_10 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_6, regroupV0_lo_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_13 = {regroupV0_lo_lo_lo_hi_hi_hi_10, regroupV0_lo_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_lo_hi_13 = {regroupV0_lo_lo_lo_hi_hi_13, regroupV0_lo_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_lo_13 = {regroupV0_lo_lo_lo_hi_13, regroupV0_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[262], regroupV0_lo_12[258]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[270], regroupV0_lo_12[266]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_6 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[278], regroupV0_lo_12[274]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[286], regroupV0_lo_12[282]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_6 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_10 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_6, regroupV0_lo_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[294], regroupV0_lo_12[290]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[302], regroupV0_lo_12[298]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_6 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[310], regroupV0_lo_12[306]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[318], regroupV0_lo_12[314]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_6 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_10 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_6, regroupV0_lo_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_13 = {regroupV0_lo_lo_hi_lo_lo_hi_10, regroupV0_lo_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[326], regroupV0_lo_12[322]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[334], regroupV0_lo_12[330]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_6 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[342], regroupV0_lo_12[338]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[350], regroupV0_lo_12[346]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_6 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_10 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_6, regroupV0_lo_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[358], regroupV0_lo_12[354]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[366], regroupV0_lo_12[362]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_6 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[374], regroupV0_lo_12[370]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[382], regroupV0_lo_12[378]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_6 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_10 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_6, regroupV0_lo_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_13 = {regroupV0_lo_lo_hi_lo_hi_hi_10, regroupV0_lo_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_lo_13 = {regroupV0_lo_lo_hi_lo_hi_13, regroupV0_lo_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[390], regroupV0_lo_12[386]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[398], regroupV0_lo_12[394]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_6 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[406], regroupV0_lo_12[402]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[414], regroupV0_lo_12[410]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_6 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_10 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_6, regroupV0_lo_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[422], regroupV0_lo_12[418]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[430], regroupV0_lo_12[426]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_6 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[438], regroupV0_lo_12[434]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[446], regroupV0_lo_12[442]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_6 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_10 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_6, regroupV0_lo_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_13 = {regroupV0_lo_lo_hi_hi_lo_hi_10, regroupV0_lo_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[454], regroupV0_lo_12[450]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[462], regroupV0_lo_12[458]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_6 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[470], regroupV0_lo_12[466]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[478], regroupV0_lo_12[474]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_6 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_10 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_6, regroupV0_lo_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[486], regroupV0_lo_12[482]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[494], regroupV0_lo_12[490]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_6 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[502], regroupV0_lo_12[498]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[510], regroupV0_lo_12[506]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_6 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_10 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_6, regroupV0_lo_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_hi_10, regroupV0_lo_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_lo_hi_hi_13 = {regroupV0_lo_lo_hi_hi_hi_13, regroupV0_lo_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_lo_hi_13 = {regroupV0_lo_lo_hi_hi_13, regroupV0_lo_lo_hi_lo_13};
  wire [127:0]       regroupV0_lo_lo_13 = {regroupV0_lo_lo_hi_13, regroupV0_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[518], regroupV0_lo_12[514]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[526], regroupV0_lo_12[522]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_6 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[534], regroupV0_lo_12[530]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[542], regroupV0_lo_12[538]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_6 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_10 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_6, regroupV0_lo_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[550], regroupV0_lo_12[546]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[558], regroupV0_lo_12[554]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_6 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[566], regroupV0_lo_12[562]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[574], regroupV0_lo_12[570]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_6 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_10 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_6, regroupV0_lo_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_13 = {regroupV0_lo_hi_lo_lo_lo_hi_10, regroupV0_lo_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[582], regroupV0_lo_12[578]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[590], regroupV0_lo_12[586]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_6 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[598], regroupV0_lo_12[594]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[606], regroupV0_lo_12[602]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_6 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_10 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_6, regroupV0_lo_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[614], regroupV0_lo_12[610]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[622], regroupV0_lo_12[618]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_6 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[630], regroupV0_lo_12[626]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[638], regroupV0_lo_12[634]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_6 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_10 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_6, regroupV0_lo_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_13 = {regroupV0_lo_hi_lo_lo_hi_hi_10, regroupV0_lo_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_lo_13 = {regroupV0_lo_hi_lo_lo_hi_13, regroupV0_lo_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[646], regroupV0_lo_12[642]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[654], regroupV0_lo_12[650]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_6 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[662], regroupV0_lo_12[658]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[670], regroupV0_lo_12[666]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_6 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_10 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_6, regroupV0_lo_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[678], regroupV0_lo_12[674]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[686], regroupV0_lo_12[682]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_6 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[694], regroupV0_lo_12[690]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[702], regroupV0_lo_12[698]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_6 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_10 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_6, regroupV0_lo_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_13 = {regroupV0_lo_hi_lo_hi_lo_hi_10, regroupV0_lo_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[710], regroupV0_lo_12[706]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[718], regroupV0_lo_12[714]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_6 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[726], regroupV0_lo_12[722]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[734], regroupV0_lo_12[730]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_6 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_10 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_6, regroupV0_lo_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[742], regroupV0_lo_12[738]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[750], regroupV0_lo_12[746]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_6 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[758], regroupV0_lo_12[754]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[766], regroupV0_lo_12[762]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_6 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_10 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_6, regroupV0_lo_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_13 = {regroupV0_lo_hi_lo_hi_hi_hi_10, regroupV0_lo_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_lo_hi_13 = {regroupV0_lo_hi_lo_hi_hi_13, regroupV0_lo_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_lo_13 = {regroupV0_lo_hi_lo_hi_13, regroupV0_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_lo_12[774], regroupV0_lo_12[770]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_lo_12[782], regroupV0_lo_12[778]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_6 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_lo_12[790], regroupV0_lo_12[786]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_lo_12[798], regroupV0_lo_12[794]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_6 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_10 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_6, regroupV0_lo_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_lo_12[806], regroupV0_lo_12[802]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_lo_12[814], regroupV0_lo_12[810]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_6 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_lo_12[822], regroupV0_lo_12[818]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_lo_12[830], regroupV0_lo_12[826]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_6 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_10 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_6, regroupV0_lo_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_13 = {regroupV0_lo_hi_hi_lo_lo_hi_10, regroupV0_lo_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_lo_12[838], regroupV0_lo_12[834]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_lo_12[846], regroupV0_lo_12[842]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_6 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_lo_12[854], regroupV0_lo_12[850]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_lo_12[862], regroupV0_lo_12[858]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_6 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_10 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_6, regroupV0_lo_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_lo_12[870], regroupV0_lo_12[866]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_lo_12[878], regroupV0_lo_12[874]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_6 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_lo_12[886], regroupV0_lo_12[882]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_lo_12[894], regroupV0_lo_12[890]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_6 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_10 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_6, regroupV0_lo_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_13 = {regroupV0_lo_hi_hi_lo_hi_hi_10, regroupV0_lo_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_lo_13 = {regroupV0_lo_hi_hi_lo_hi_13, regroupV0_lo_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_lo_12[902], regroupV0_lo_12[898]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_lo_12[910], regroupV0_lo_12[906]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_6 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_lo_12[918], regroupV0_lo_12[914]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_lo_12[926], regroupV0_lo_12[922]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_6 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_10 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_6, regroupV0_lo_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_lo_12[934], regroupV0_lo_12[930]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_lo_12[942], regroupV0_lo_12[938]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_6 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_lo_12[950], regroupV0_lo_12[946]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_lo_12[958], regroupV0_lo_12[954]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_6 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_10 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_6, regroupV0_lo_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_13 = {regroupV0_lo_hi_hi_hi_lo_hi_10, regroupV0_lo_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_lo_12[966], regroupV0_lo_12[962]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_lo_12[974], regroupV0_lo_12[970]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_6 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_lo_12[982], regroupV0_lo_12[978]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_lo_12[990], regroupV0_lo_12[986]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_6 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_10 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_6, regroupV0_lo_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_lo_12[998], regroupV0_lo_12[994]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_lo_12[1006], regroupV0_lo_12[1002]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_6 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_lo_12[1014], regroupV0_lo_12[1010]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_lo_12[1022], regroupV0_lo_12[1018]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_6 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_10 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_6, regroupV0_lo_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_hi_10, regroupV0_lo_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_lo_hi_hi_hi_13 = {regroupV0_lo_hi_hi_hi_hi_13, regroupV0_lo_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_lo_hi_hi_13 = {regroupV0_lo_hi_hi_hi_13, regroupV0_lo_hi_hi_lo_13};
  wire [127:0]       regroupV0_lo_hi_13 = {regroupV0_lo_hi_hi_13, regroupV0_lo_hi_lo_13};
  wire [255:0]       regroupV0_lo_15 = {regroupV0_lo_hi_13, regroupV0_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[6], regroupV0_hi_12[2]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[14], regroupV0_hi_12[10]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_6 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[22], regroupV0_hi_12[18]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[30], regroupV0_hi_12[26]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_6 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_10 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_6, regroupV0_hi_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[38], regroupV0_hi_12[34]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[46], regroupV0_hi_12[42]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_6 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[54], regroupV0_hi_12[50]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[62], regroupV0_hi_12[58]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_6 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_10 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_6, regroupV0_hi_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_lo_hi_10, regroupV0_hi_lo_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[70], regroupV0_hi_12[66]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[78], regroupV0_hi_12[74]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_6 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[86], regroupV0_hi_12[82]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[94], regroupV0_hi_12[90]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_6 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_10 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_6, regroupV0_hi_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[102], regroupV0_hi_12[98]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[110], regroupV0_hi_12[106]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_6 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[118], regroupV0_hi_12[114]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[126], regroupV0_hi_12[122]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_6 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_10 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_6, regroupV0_hi_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_13 = {regroupV0_hi_lo_lo_lo_hi_hi_10, regroupV0_hi_lo_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_lo_13 = {regroupV0_hi_lo_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[134], regroupV0_hi_12[130]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[142], regroupV0_hi_12[138]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_6 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[150], regroupV0_hi_12[146]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[158], regroupV0_hi_12[154]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_6 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_10 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_6, regroupV0_hi_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[166], regroupV0_hi_12[162]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[174], regroupV0_hi_12[170]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_6 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[182], regroupV0_hi_12[178]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[190], regroupV0_hi_12[186]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_6 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_10 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_6, regroupV0_hi_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_13 = {regroupV0_hi_lo_lo_hi_lo_hi_10, regroupV0_hi_lo_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[198], regroupV0_hi_12[194]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[206], regroupV0_hi_12[202]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_6 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[214], regroupV0_hi_12[210]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[222], regroupV0_hi_12[218]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_6 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_10 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_6, regroupV0_hi_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[230], regroupV0_hi_12[226]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[238], regroupV0_hi_12[234]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_6 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[246], regroupV0_hi_12[242]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[254], regroupV0_hi_12[250]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_6 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_10 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_6, regroupV0_hi_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_13 = {regroupV0_hi_lo_lo_hi_hi_hi_10, regroupV0_hi_lo_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_lo_hi_13 = {regroupV0_hi_lo_lo_hi_hi_13, regroupV0_hi_lo_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_lo_13 = {regroupV0_hi_lo_lo_hi_13, regroupV0_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[262], regroupV0_hi_12[258]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[270], regroupV0_hi_12[266]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_6 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[278], regroupV0_hi_12[274]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[286], regroupV0_hi_12[282]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_6 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_10 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_6, regroupV0_hi_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[294], regroupV0_hi_12[290]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[302], regroupV0_hi_12[298]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_6 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[310], regroupV0_hi_12[306]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[318], regroupV0_hi_12[314]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_6 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_10 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_6, regroupV0_hi_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_13 = {regroupV0_hi_lo_hi_lo_lo_hi_10, regroupV0_hi_lo_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[326], regroupV0_hi_12[322]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[334], regroupV0_hi_12[330]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_6 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[342], regroupV0_hi_12[338]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[350], regroupV0_hi_12[346]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_6 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_10 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_6, regroupV0_hi_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[358], regroupV0_hi_12[354]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[366], regroupV0_hi_12[362]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_6 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[374], regroupV0_hi_12[370]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[382], regroupV0_hi_12[378]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_6 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_10 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_6, regroupV0_hi_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_13 = {regroupV0_hi_lo_hi_lo_hi_hi_10, regroupV0_hi_lo_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_lo_13 = {regroupV0_hi_lo_hi_lo_hi_13, regroupV0_hi_lo_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[390], regroupV0_hi_12[386]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[398], regroupV0_hi_12[394]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_6 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[406], regroupV0_hi_12[402]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[414], regroupV0_hi_12[410]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_6 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_10 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_6, regroupV0_hi_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[422], regroupV0_hi_12[418]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[430], regroupV0_hi_12[426]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_6 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[438], regroupV0_hi_12[434]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[446], regroupV0_hi_12[442]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_6 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_10 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_6, regroupV0_hi_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_13 = {regroupV0_hi_lo_hi_hi_lo_hi_10, regroupV0_hi_lo_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[454], regroupV0_hi_12[450]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[462], regroupV0_hi_12[458]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_6 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[470], regroupV0_hi_12[466]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[478], regroupV0_hi_12[474]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_6 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_10 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_6, regroupV0_hi_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[486], regroupV0_hi_12[482]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[494], regroupV0_hi_12[490]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_6 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[502], regroupV0_hi_12[498]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[510], regroupV0_hi_12[506]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_6 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_10 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_6, regroupV0_hi_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_hi_10, regroupV0_hi_lo_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_lo_hi_hi_13 = {regroupV0_hi_lo_hi_hi_hi_13, regroupV0_hi_lo_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_lo_hi_13 = {regroupV0_hi_lo_hi_hi_13, regroupV0_hi_lo_hi_lo_13};
  wire [127:0]       regroupV0_hi_lo_13 = {regroupV0_hi_lo_hi_13, regroupV0_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[518], regroupV0_hi_12[514]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[526], regroupV0_hi_12[522]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_6 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[534], regroupV0_hi_12[530]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[542], regroupV0_hi_12[538]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_6 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_10 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_6, regroupV0_hi_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[550], regroupV0_hi_12[546]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[558], regroupV0_hi_12[554]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_6 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[566], regroupV0_hi_12[562]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[574], regroupV0_hi_12[570]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_6 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_10 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_6, regroupV0_hi_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_13 = {regroupV0_hi_hi_lo_lo_lo_hi_10, regroupV0_hi_hi_lo_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[582], regroupV0_hi_12[578]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[590], regroupV0_hi_12[586]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_6 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[598], regroupV0_hi_12[594]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[606], regroupV0_hi_12[602]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_6 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_10 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_6, regroupV0_hi_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[614], regroupV0_hi_12[610]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[622], regroupV0_hi_12[618]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_6 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[630], regroupV0_hi_12[626]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[638], regroupV0_hi_12[634]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_6 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_10 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_6, regroupV0_hi_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_13 = {regroupV0_hi_hi_lo_lo_hi_hi_10, regroupV0_hi_hi_lo_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_lo_13 = {regroupV0_hi_hi_lo_lo_hi_13, regroupV0_hi_hi_lo_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[646], regroupV0_hi_12[642]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[654], regroupV0_hi_12[650]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_6 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[662], regroupV0_hi_12[658]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[670], regroupV0_hi_12[666]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_6 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_10 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_6, regroupV0_hi_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[678], regroupV0_hi_12[674]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[686], regroupV0_hi_12[682]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_6 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[694], regroupV0_hi_12[690]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[702], regroupV0_hi_12[698]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_6 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_10 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_6, regroupV0_hi_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_13 = {regroupV0_hi_hi_lo_hi_lo_hi_10, regroupV0_hi_hi_lo_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[710], regroupV0_hi_12[706]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[718], regroupV0_hi_12[714]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_6 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[726], regroupV0_hi_12[722]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[734], regroupV0_hi_12[730]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_6 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_10 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_6, regroupV0_hi_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[742], regroupV0_hi_12[738]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[750], regroupV0_hi_12[746]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_6 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[758], regroupV0_hi_12[754]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[766], regroupV0_hi_12[762]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_6 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_10 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_6, regroupV0_hi_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_13 = {regroupV0_hi_hi_lo_hi_hi_hi_10, regroupV0_hi_hi_lo_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_lo_hi_13 = {regroupV0_hi_hi_lo_hi_hi_13, regroupV0_hi_hi_lo_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_lo_13 = {regroupV0_hi_hi_lo_hi_13, regroupV0_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_2 = {regroupV0_hi_12[774], regroupV0_hi_12[770]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_2 = {regroupV0_hi_12[782], regroupV0_hi_12[778]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_6 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_2 = {regroupV0_hi_12[790], regroupV0_hi_12[786]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_2 = {regroupV0_hi_12[798], regroupV0_hi_12[794]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_6 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_10 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_6, regroupV0_hi_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_2 = {regroupV0_hi_12[806], regroupV0_hi_12[802]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_2 = {regroupV0_hi_12[814], regroupV0_hi_12[810]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_6 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_2 = {regroupV0_hi_12[822], regroupV0_hi_12[818]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_2 = {regroupV0_hi_12[830], regroupV0_hi_12[826]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_6 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_10 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_6, regroupV0_hi_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_13 = {regroupV0_hi_hi_hi_lo_lo_hi_10, regroupV0_hi_hi_hi_lo_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_2 = {regroupV0_hi_12[838], regroupV0_hi_12[834]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_2 = {regroupV0_hi_12[846], regroupV0_hi_12[842]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_6 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_2 = {regroupV0_hi_12[854], regroupV0_hi_12[850]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_2 = {regroupV0_hi_12[862], regroupV0_hi_12[858]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_6 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_10 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_6, regroupV0_hi_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_2 = {regroupV0_hi_12[870], regroupV0_hi_12[866]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_2 = {regroupV0_hi_12[878], regroupV0_hi_12[874]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_6 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_2 = {regroupV0_hi_12[886], regroupV0_hi_12[882]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_2 = {regroupV0_hi_12[894], regroupV0_hi_12[890]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_6 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_10 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_6, regroupV0_hi_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_13 = {regroupV0_hi_hi_hi_lo_hi_hi_10, regroupV0_hi_hi_hi_lo_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_lo_hi_13, regroupV0_hi_hi_hi_lo_lo_13};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_2 = {regroupV0_hi_12[902], regroupV0_hi_12[898]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_2 = {regroupV0_hi_12[910], regroupV0_hi_12[906]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_6 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_2 = {regroupV0_hi_12[918], regroupV0_hi_12[914]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_2 = {regroupV0_hi_12[926], regroupV0_hi_12[922]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_6 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_10 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_6, regroupV0_hi_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_2 = {regroupV0_hi_12[934], regroupV0_hi_12[930]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_2 = {regroupV0_hi_12[942], regroupV0_hi_12[938]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_6 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_2 = {regroupV0_hi_12[950], regroupV0_hi_12[946]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_2 = {regroupV0_hi_12[958], regroupV0_hi_12[954]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_6 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_10 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_6, regroupV0_hi_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_13 = {regroupV0_hi_hi_hi_hi_lo_hi_10, regroupV0_hi_hi_hi_hi_lo_lo_10};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_2 = {regroupV0_hi_12[966], regroupV0_hi_12[962]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_2 = {regroupV0_hi_12[974], regroupV0_hi_12[970]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_6 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_2 = {regroupV0_hi_12[982], regroupV0_hi_12[978]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_2 = {regroupV0_hi_12[990], regroupV0_hi_12[986]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_6 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_10 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_6, regroupV0_hi_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_2 = {regroupV0_hi_12[998], regroupV0_hi_12[994]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_2 = {regroupV0_hi_12[1006], regroupV0_hi_12[1002]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_6 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_2 = {regroupV0_hi_12[1014], regroupV0_hi_12[1010]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_2 = {regroupV0_hi_12[1022], regroupV0_hi_12[1018]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_6 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_2, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_10 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_6, regroupV0_hi_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_hi_10, regroupV0_hi_hi_hi_hi_hi_lo_10};
  wire [31:0]        regroupV0_hi_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_hi_lo_13};
  wire [63:0]        regroupV0_hi_hi_hi_13 = {regroupV0_hi_hi_hi_hi_13, regroupV0_hi_hi_hi_lo_13};
  wire [127:0]       regroupV0_hi_hi_13 = {regroupV0_hi_hi_hi_13, regroupV0_hi_hi_lo_13};
  wire [255:0]       regroupV0_hi_15 = {regroupV0_hi_hi_13, regroupV0_hi_lo_13};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[7], regroupV0_lo_12[3]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[15], regroupV0_lo_12[11]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_lo_7 = {regroupV0_lo_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[23], regroupV0_lo_12[19]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[31], regroupV0_lo_12[27]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_lo_hi_7 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_lo_11 = {regroupV0_lo_lo_lo_lo_lo_lo_hi_7, regroupV0_lo_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[39], regroupV0_lo_12[35]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[47], regroupV0_lo_12[43]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_lo_7 = {regroupV0_lo_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[55], regroupV0_lo_12[51]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[63], regroupV0_lo_12[59]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_lo_hi_hi_7 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_lo_hi_11 = {regroupV0_lo_lo_lo_lo_lo_hi_hi_7, regroupV0_lo_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_lo_hi_11, regroupV0_lo_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[71], regroupV0_lo_12[67]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[79], regroupV0_lo_12[75]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_lo_7 = {regroupV0_lo_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[87], regroupV0_lo_12[83]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[95], regroupV0_lo_12[91]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_lo_hi_7 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_lo_11 = {regroupV0_lo_lo_lo_lo_hi_lo_hi_7, regroupV0_lo_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[103], regroupV0_lo_12[99]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[111], regroupV0_lo_12[107]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_lo_7 = {regroupV0_lo_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[119], regroupV0_lo_12[115]};
  wire [1:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[127], regroupV0_lo_12[123]};
  wire [3:0]         regroupV0_lo_lo_lo_lo_hi_hi_hi_7 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_lo_hi_hi_11 = {regroupV0_lo_lo_lo_lo_hi_hi_hi_7, regroupV0_lo_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_lo_hi_hi_11, regroupV0_lo_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_lo_14 = {regroupV0_lo_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[135], regroupV0_lo_12[131]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[143], regroupV0_lo_12[139]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_lo_7 = {regroupV0_lo_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[151], regroupV0_lo_12[147]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[159], regroupV0_lo_12[155]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_lo_hi_7 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_lo_11 = {regroupV0_lo_lo_lo_hi_lo_lo_hi_7, regroupV0_lo_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[167], regroupV0_lo_12[163]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[175], regroupV0_lo_12[171]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_lo_7 = {regroupV0_lo_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[183], regroupV0_lo_12[179]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[191], regroupV0_lo_12[187]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_lo_hi_hi_7 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_lo_hi_11 = {regroupV0_lo_lo_lo_hi_lo_hi_hi_7, regroupV0_lo_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_lo_14 = {regroupV0_lo_lo_lo_hi_lo_hi_11, regroupV0_lo_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[199], regroupV0_lo_12[195]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[207], regroupV0_lo_12[203]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_lo_7 = {regroupV0_lo_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[215], regroupV0_lo_12[211]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[223], regroupV0_lo_12[219]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_lo_hi_7 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_lo_11 = {regroupV0_lo_lo_lo_hi_hi_lo_hi_7, regroupV0_lo_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[231], regroupV0_lo_12[227]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[239], regroupV0_lo_12[235]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_lo_7 = {regroupV0_lo_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[247], regroupV0_lo_12[243]};
  wire [1:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[255], regroupV0_lo_12[251]};
  wire [3:0]         regroupV0_lo_lo_lo_hi_hi_hi_hi_7 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_lo_hi_hi_hi_11 = {regroupV0_lo_lo_lo_hi_hi_hi_hi_7, regroupV0_lo_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_lo_hi_hi_14 = {regroupV0_lo_lo_lo_hi_hi_hi_11, regroupV0_lo_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_lo_hi_14 = {regroupV0_lo_lo_lo_hi_hi_14, regroupV0_lo_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_lo_14 = {regroupV0_lo_lo_lo_hi_14, regroupV0_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[263], regroupV0_lo_12[259]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[271], regroupV0_lo_12[267]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_lo_7 = {regroupV0_lo_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[279], regroupV0_lo_12[275]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[287], regroupV0_lo_12[283]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_lo_hi_7 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_lo_11 = {regroupV0_lo_lo_hi_lo_lo_lo_hi_7, regroupV0_lo_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[295], regroupV0_lo_12[291]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[303], regroupV0_lo_12[299]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_lo_7 = {regroupV0_lo_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[311], regroupV0_lo_12[307]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[319], regroupV0_lo_12[315]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_lo_hi_hi_7 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_lo_hi_11 = {regroupV0_lo_lo_hi_lo_lo_hi_hi_7, regroupV0_lo_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_lo_14 = {regroupV0_lo_lo_hi_lo_lo_hi_11, regroupV0_lo_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[327], regroupV0_lo_12[323]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[335], regroupV0_lo_12[331]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_lo_7 = {regroupV0_lo_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[343], regroupV0_lo_12[339]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[351], regroupV0_lo_12[347]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_lo_hi_7 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_lo_11 = {regroupV0_lo_lo_hi_lo_hi_lo_hi_7, regroupV0_lo_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[359], regroupV0_lo_12[355]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[367], regroupV0_lo_12[363]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_lo_7 = {regroupV0_lo_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[375], regroupV0_lo_12[371]};
  wire [1:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[383], regroupV0_lo_12[379]};
  wire [3:0]         regroupV0_lo_lo_hi_lo_hi_hi_hi_7 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_lo_hi_hi_11 = {regroupV0_lo_lo_hi_lo_hi_hi_hi_7, regroupV0_lo_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_lo_hi_14 = {regroupV0_lo_lo_hi_lo_hi_hi_11, regroupV0_lo_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_lo_14 = {regroupV0_lo_lo_hi_lo_hi_14, regroupV0_lo_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[391], regroupV0_lo_12[387]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[399], regroupV0_lo_12[395]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_lo_7 = {regroupV0_lo_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[407], regroupV0_lo_12[403]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[415], regroupV0_lo_12[411]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_lo_hi_7 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_lo_11 = {regroupV0_lo_lo_hi_hi_lo_lo_hi_7, regroupV0_lo_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[423], regroupV0_lo_12[419]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[431], regroupV0_lo_12[427]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_lo_7 = {regroupV0_lo_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[439], regroupV0_lo_12[435]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[447], regroupV0_lo_12[443]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_lo_hi_hi_7 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_lo_hi_11 = {regroupV0_lo_lo_hi_hi_lo_hi_hi_7, regroupV0_lo_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_lo_14 = {regroupV0_lo_lo_hi_hi_lo_hi_11, regroupV0_lo_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[455], regroupV0_lo_12[451]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[463], regroupV0_lo_12[459]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_lo_7 = {regroupV0_lo_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[471], regroupV0_lo_12[467]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[479], regroupV0_lo_12[475]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_lo_hi_7 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_lo_11 = {regroupV0_lo_lo_hi_hi_hi_lo_hi_7, regroupV0_lo_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[487], regroupV0_lo_12[483]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[495], regroupV0_lo_12[491]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_lo_7 = {regroupV0_lo_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[503], regroupV0_lo_12[499]};
  wire [1:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[511], regroupV0_lo_12[507]};
  wire [3:0]         regroupV0_lo_lo_hi_hi_hi_hi_hi_7 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_lo_hi_hi_hi_hi_11 = {regroupV0_lo_lo_hi_hi_hi_hi_hi_7, regroupV0_lo_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_lo_hi_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_hi_11, regroupV0_lo_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_lo_hi_hi_14 = {regroupV0_lo_lo_hi_hi_hi_14, regroupV0_lo_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_lo_hi_14 = {regroupV0_lo_lo_hi_hi_14, regroupV0_lo_lo_hi_lo_14};
  wire [127:0]       regroupV0_lo_lo_14 = {regroupV0_lo_lo_hi_14, regroupV0_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[519], regroupV0_lo_12[515]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[527], regroupV0_lo_12[523]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_lo_7 = {regroupV0_lo_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[535], regroupV0_lo_12[531]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[543], regroupV0_lo_12[539]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_lo_hi_7 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_lo_11 = {regroupV0_lo_hi_lo_lo_lo_lo_hi_7, regroupV0_lo_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[551], regroupV0_lo_12[547]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[559], regroupV0_lo_12[555]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_lo_7 = {regroupV0_lo_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[567], regroupV0_lo_12[563]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[575], regroupV0_lo_12[571]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_lo_hi_hi_7 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_lo_hi_11 = {regroupV0_lo_hi_lo_lo_lo_hi_hi_7, regroupV0_lo_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_lo_14 = {regroupV0_lo_hi_lo_lo_lo_hi_11, regroupV0_lo_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[583], regroupV0_lo_12[579]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[591], regroupV0_lo_12[587]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_lo_7 = {regroupV0_lo_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[599], regroupV0_lo_12[595]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[607], regroupV0_lo_12[603]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_lo_hi_7 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_lo_11 = {regroupV0_lo_hi_lo_lo_hi_lo_hi_7, regroupV0_lo_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[615], regroupV0_lo_12[611]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[623], regroupV0_lo_12[619]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_lo_7 = {regroupV0_lo_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[631], regroupV0_lo_12[627]};
  wire [1:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[639], regroupV0_lo_12[635]};
  wire [3:0]         regroupV0_lo_hi_lo_lo_hi_hi_hi_7 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_lo_hi_hi_11 = {regroupV0_lo_hi_lo_lo_hi_hi_hi_7, regroupV0_lo_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_lo_hi_14 = {regroupV0_lo_hi_lo_lo_hi_hi_11, regroupV0_lo_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_lo_14 = {regroupV0_lo_hi_lo_lo_hi_14, regroupV0_lo_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[647], regroupV0_lo_12[643]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[655], regroupV0_lo_12[651]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_lo_7 = {regroupV0_lo_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[663], regroupV0_lo_12[659]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[671], regroupV0_lo_12[667]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_lo_hi_7 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_lo_11 = {regroupV0_lo_hi_lo_hi_lo_lo_hi_7, regroupV0_lo_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[679], regroupV0_lo_12[675]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[687], regroupV0_lo_12[683]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_lo_7 = {regroupV0_lo_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[695], regroupV0_lo_12[691]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[703], regroupV0_lo_12[699]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_lo_hi_hi_7 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_lo_hi_11 = {regroupV0_lo_hi_lo_hi_lo_hi_hi_7, regroupV0_lo_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_lo_14 = {regroupV0_lo_hi_lo_hi_lo_hi_11, regroupV0_lo_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[711], regroupV0_lo_12[707]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[719], regroupV0_lo_12[715]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_lo_7 = {regroupV0_lo_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[727], regroupV0_lo_12[723]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[735], regroupV0_lo_12[731]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_lo_hi_7 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_lo_11 = {regroupV0_lo_hi_lo_hi_hi_lo_hi_7, regroupV0_lo_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[743], regroupV0_lo_12[739]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[751], regroupV0_lo_12[747]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_lo_7 = {regroupV0_lo_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[759], regroupV0_lo_12[755]};
  wire [1:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[767], regroupV0_lo_12[763]};
  wire [3:0]         regroupV0_lo_hi_lo_hi_hi_hi_hi_7 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_lo_hi_hi_hi_11 = {regroupV0_lo_hi_lo_hi_hi_hi_hi_7, regroupV0_lo_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_lo_hi_hi_14 = {regroupV0_lo_hi_lo_hi_hi_hi_11, regroupV0_lo_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_lo_hi_14 = {regroupV0_lo_hi_lo_hi_hi_14, regroupV0_lo_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_lo_14 = {regroupV0_lo_hi_lo_hi_14, regroupV0_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_lo_12[775], regroupV0_lo_12[771]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_lo_12[783], regroupV0_lo_12[779]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_lo_7 = {regroupV0_lo_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_lo_12[791], regroupV0_lo_12[787]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_lo_12[799], regroupV0_lo_12[795]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_lo_hi_7 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_lo_11 = {regroupV0_lo_hi_hi_lo_lo_lo_hi_7, regroupV0_lo_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_lo_12[807], regroupV0_lo_12[803]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_lo_12[815], regroupV0_lo_12[811]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_lo_7 = {regroupV0_lo_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_lo_12[823], regroupV0_lo_12[819]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_lo_12[831], regroupV0_lo_12[827]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_lo_hi_hi_7 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_lo_hi_11 = {regroupV0_lo_hi_hi_lo_lo_hi_hi_7, regroupV0_lo_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_lo_14 = {regroupV0_lo_hi_hi_lo_lo_hi_11, regroupV0_lo_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_lo_12[839], regroupV0_lo_12[835]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_lo_12[847], regroupV0_lo_12[843]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_lo_7 = {regroupV0_lo_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_lo_12[855], regroupV0_lo_12[851]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_lo_12[863], regroupV0_lo_12[859]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_lo_hi_7 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_lo_11 = {regroupV0_lo_hi_hi_lo_hi_lo_hi_7, regroupV0_lo_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_lo_12[871], regroupV0_lo_12[867]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_lo_12[879], regroupV0_lo_12[875]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_lo_7 = {regroupV0_lo_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_lo_12[887], regroupV0_lo_12[883]};
  wire [1:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_lo_12[895], regroupV0_lo_12[891]};
  wire [3:0]         regroupV0_lo_hi_hi_lo_hi_hi_hi_7 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_lo_hi_hi_11 = {regroupV0_lo_hi_hi_lo_hi_hi_hi_7, regroupV0_lo_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_lo_hi_14 = {regroupV0_lo_hi_hi_lo_hi_hi_11, regroupV0_lo_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_lo_14 = {regroupV0_lo_hi_hi_lo_hi_14, regroupV0_lo_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_lo_12[903], regroupV0_lo_12[899]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_lo_12[911], regroupV0_lo_12[907]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_lo_7 = {regroupV0_lo_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_lo_12[919], regroupV0_lo_12[915]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_lo_12[927], regroupV0_lo_12[923]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_lo_hi_7 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_lo_11 = {regroupV0_lo_hi_hi_hi_lo_lo_hi_7, regroupV0_lo_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_lo_12[935], regroupV0_lo_12[931]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_lo_12[943], regroupV0_lo_12[939]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_lo_7 = {regroupV0_lo_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_lo_12[951], regroupV0_lo_12[947]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_lo_12[959], regroupV0_lo_12[955]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_lo_hi_hi_7 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_lo_hi_11 = {regroupV0_lo_hi_hi_hi_lo_hi_hi_7, regroupV0_lo_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_lo_14 = {regroupV0_lo_hi_hi_hi_lo_hi_11, regroupV0_lo_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_lo_12[967], regroupV0_lo_12[963]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_lo_12[975], regroupV0_lo_12[971]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_lo_7 = {regroupV0_lo_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_lo_12[983], regroupV0_lo_12[979]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_lo_12[991], regroupV0_lo_12[987]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_lo_hi_7 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_lo_11 = {regroupV0_lo_hi_hi_hi_hi_lo_hi_7, regroupV0_lo_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_lo_12[999], regroupV0_lo_12[995]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_lo_12[1007], regroupV0_lo_12[1003]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_lo_7 = {regroupV0_lo_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_lo_12[1015], regroupV0_lo_12[1011]};
  wire [1:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_lo_12[1023], regroupV0_lo_12[1019]};
  wire [3:0]         regroupV0_lo_hi_hi_hi_hi_hi_hi_7 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_lo_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_lo_hi_hi_hi_hi_hi_11 = {regroupV0_lo_hi_hi_hi_hi_hi_hi_7, regroupV0_lo_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_lo_hi_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_hi_11, regroupV0_lo_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_lo_hi_hi_hi_14 = {regroupV0_lo_hi_hi_hi_hi_14, regroupV0_lo_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_lo_hi_hi_14 = {regroupV0_lo_hi_hi_hi_14, regroupV0_lo_hi_hi_lo_14};
  wire [127:0]       regroupV0_lo_hi_14 = {regroupV0_lo_hi_hi_14, regroupV0_lo_hi_lo_14};
  wire [255:0]       regroupV0_lo_16 = {regroupV0_lo_hi_14, regroupV0_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[7], regroupV0_hi_12[3]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[15], regroupV0_hi_12[11]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_lo_7 = {regroupV0_hi_lo_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[23], regroupV0_hi_12[19]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[31], regroupV0_hi_12[27]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_lo_hi_7 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_lo_11 = {regroupV0_hi_lo_lo_lo_lo_lo_hi_7, regroupV0_hi_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[39], regroupV0_hi_12[35]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[47], regroupV0_hi_12[43]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_lo_7 = {regroupV0_hi_lo_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[55], regroupV0_hi_12[51]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[63], regroupV0_hi_12[59]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_lo_hi_hi_7 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_lo_hi_11 = {regroupV0_hi_lo_lo_lo_lo_hi_hi_7, regroupV0_hi_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_lo_hi_11, regroupV0_hi_lo_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[71], regroupV0_hi_12[67]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[79], regroupV0_hi_12[75]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_lo_7 = {regroupV0_hi_lo_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[87], regroupV0_hi_12[83]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[95], regroupV0_hi_12[91]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_lo_hi_7 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_lo_11 = {regroupV0_hi_lo_lo_lo_hi_lo_hi_7, regroupV0_hi_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[103], regroupV0_hi_12[99]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[111], regroupV0_hi_12[107]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_lo_7 = {regroupV0_hi_lo_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[119], regroupV0_hi_12[115]};
  wire [1:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[127], regroupV0_hi_12[123]};
  wire [3:0]         regroupV0_hi_lo_lo_lo_hi_hi_hi_7 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_lo_hi_hi_11 = {regroupV0_hi_lo_lo_lo_hi_hi_hi_7, regroupV0_hi_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_lo_hi_14 = {regroupV0_hi_lo_lo_lo_hi_hi_11, regroupV0_hi_lo_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_lo_14 = {regroupV0_hi_lo_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[135], regroupV0_hi_12[131]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[143], regroupV0_hi_12[139]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_lo_7 = {regroupV0_hi_lo_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[151], regroupV0_hi_12[147]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[159], regroupV0_hi_12[155]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_lo_hi_7 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_lo_11 = {regroupV0_hi_lo_lo_hi_lo_lo_hi_7, regroupV0_hi_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[167], regroupV0_hi_12[163]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[175], regroupV0_hi_12[171]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_lo_7 = {regroupV0_hi_lo_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[183], regroupV0_hi_12[179]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[191], regroupV0_hi_12[187]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_lo_hi_hi_7 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_lo_hi_11 = {regroupV0_hi_lo_lo_hi_lo_hi_hi_7, regroupV0_hi_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_lo_14 = {regroupV0_hi_lo_lo_hi_lo_hi_11, regroupV0_hi_lo_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[199], regroupV0_hi_12[195]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[207], regroupV0_hi_12[203]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_lo_7 = {regroupV0_hi_lo_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[215], regroupV0_hi_12[211]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[223], regroupV0_hi_12[219]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_lo_hi_7 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_lo_11 = {regroupV0_hi_lo_lo_hi_hi_lo_hi_7, regroupV0_hi_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[231], regroupV0_hi_12[227]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[239], regroupV0_hi_12[235]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_lo_7 = {regroupV0_hi_lo_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[247], regroupV0_hi_12[243]};
  wire [1:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[255], regroupV0_hi_12[251]};
  wire [3:0]         regroupV0_hi_lo_lo_hi_hi_hi_hi_7 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_lo_hi_hi_hi_11 = {regroupV0_hi_lo_lo_hi_hi_hi_hi_7, regroupV0_hi_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_lo_hi_hi_14 = {regroupV0_hi_lo_lo_hi_hi_hi_11, regroupV0_hi_lo_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_lo_hi_14 = {regroupV0_hi_lo_lo_hi_hi_14, regroupV0_hi_lo_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_lo_14 = {regroupV0_hi_lo_lo_hi_14, regroupV0_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[263], regroupV0_hi_12[259]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[271], regroupV0_hi_12[267]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_lo_7 = {regroupV0_hi_lo_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[279], regroupV0_hi_12[275]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[287], regroupV0_hi_12[283]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_lo_hi_7 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_lo_11 = {regroupV0_hi_lo_hi_lo_lo_lo_hi_7, regroupV0_hi_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[295], regroupV0_hi_12[291]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[303], regroupV0_hi_12[299]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_lo_7 = {regroupV0_hi_lo_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[311], regroupV0_hi_12[307]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[319], regroupV0_hi_12[315]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_lo_hi_hi_7 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_lo_hi_11 = {regroupV0_hi_lo_hi_lo_lo_hi_hi_7, regroupV0_hi_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_lo_14 = {regroupV0_hi_lo_hi_lo_lo_hi_11, regroupV0_hi_lo_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[327], regroupV0_hi_12[323]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[335], regroupV0_hi_12[331]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_lo_7 = {regroupV0_hi_lo_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[343], regroupV0_hi_12[339]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[351], regroupV0_hi_12[347]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_lo_hi_7 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_lo_11 = {regroupV0_hi_lo_hi_lo_hi_lo_hi_7, regroupV0_hi_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[359], regroupV0_hi_12[355]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[367], regroupV0_hi_12[363]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_lo_7 = {regroupV0_hi_lo_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[375], regroupV0_hi_12[371]};
  wire [1:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[383], regroupV0_hi_12[379]};
  wire [3:0]         regroupV0_hi_lo_hi_lo_hi_hi_hi_7 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_lo_hi_hi_11 = {regroupV0_hi_lo_hi_lo_hi_hi_hi_7, regroupV0_hi_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_lo_hi_14 = {regroupV0_hi_lo_hi_lo_hi_hi_11, regroupV0_hi_lo_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_lo_14 = {regroupV0_hi_lo_hi_lo_hi_14, regroupV0_hi_lo_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[391], regroupV0_hi_12[387]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[399], regroupV0_hi_12[395]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_lo_7 = {regroupV0_hi_lo_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[407], regroupV0_hi_12[403]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[415], regroupV0_hi_12[411]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_lo_hi_7 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_lo_11 = {regroupV0_hi_lo_hi_hi_lo_lo_hi_7, regroupV0_hi_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[423], regroupV0_hi_12[419]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[431], regroupV0_hi_12[427]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_lo_7 = {regroupV0_hi_lo_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[439], regroupV0_hi_12[435]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[447], regroupV0_hi_12[443]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_lo_hi_hi_7 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_lo_hi_11 = {regroupV0_hi_lo_hi_hi_lo_hi_hi_7, regroupV0_hi_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_lo_14 = {regroupV0_hi_lo_hi_hi_lo_hi_11, regroupV0_hi_lo_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[455], regroupV0_hi_12[451]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[463], regroupV0_hi_12[459]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_lo_7 = {regroupV0_hi_lo_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[471], regroupV0_hi_12[467]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[479], regroupV0_hi_12[475]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_lo_hi_7 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_lo_11 = {regroupV0_hi_lo_hi_hi_hi_lo_hi_7, regroupV0_hi_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[487], regroupV0_hi_12[483]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[495], regroupV0_hi_12[491]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_lo_7 = {regroupV0_hi_lo_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[503], regroupV0_hi_12[499]};
  wire [1:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[511], regroupV0_hi_12[507]};
  wire [3:0]         regroupV0_hi_lo_hi_hi_hi_hi_hi_7 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_lo_hi_hi_hi_hi_11 = {regroupV0_hi_lo_hi_hi_hi_hi_hi_7, regroupV0_hi_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_lo_hi_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_hi_11, regroupV0_hi_lo_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_lo_hi_hi_14 = {regroupV0_hi_lo_hi_hi_hi_14, regroupV0_hi_lo_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_lo_hi_14 = {regroupV0_hi_lo_hi_hi_14, regroupV0_hi_lo_hi_lo_14};
  wire [127:0]       regroupV0_hi_lo_14 = {regroupV0_hi_lo_hi_14, regroupV0_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[519], regroupV0_hi_12[515]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[527], regroupV0_hi_12[523]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_lo_7 = {regroupV0_hi_hi_lo_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[535], regroupV0_hi_12[531]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[543], regroupV0_hi_12[539]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_lo_hi_7 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_lo_11 = {regroupV0_hi_hi_lo_lo_lo_lo_hi_7, regroupV0_hi_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[551], regroupV0_hi_12[547]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[559], regroupV0_hi_12[555]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_lo_7 = {regroupV0_hi_hi_lo_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[567], regroupV0_hi_12[563]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[575], regroupV0_hi_12[571]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_lo_hi_hi_7 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_lo_hi_11 = {regroupV0_hi_hi_lo_lo_lo_hi_hi_7, regroupV0_hi_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_lo_14 = {regroupV0_hi_hi_lo_lo_lo_hi_11, regroupV0_hi_hi_lo_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[583], regroupV0_hi_12[579]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[591], regroupV0_hi_12[587]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_lo_7 = {regroupV0_hi_hi_lo_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[599], regroupV0_hi_12[595]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[607], regroupV0_hi_12[603]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_lo_hi_7 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_lo_11 = {regroupV0_hi_hi_lo_lo_hi_lo_hi_7, regroupV0_hi_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[615], regroupV0_hi_12[611]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[623], regroupV0_hi_12[619]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_lo_7 = {regroupV0_hi_hi_lo_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[631], regroupV0_hi_12[627]};
  wire [1:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[639], regroupV0_hi_12[635]};
  wire [3:0]         regroupV0_hi_hi_lo_lo_hi_hi_hi_7 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_lo_hi_hi_11 = {regroupV0_hi_hi_lo_lo_hi_hi_hi_7, regroupV0_hi_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_lo_hi_14 = {regroupV0_hi_hi_lo_lo_hi_hi_11, regroupV0_hi_hi_lo_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_lo_14 = {regroupV0_hi_hi_lo_lo_hi_14, regroupV0_hi_hi_lo_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[647], regroupV0_hi_12[643]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[655], regroupV0_hi_12[651]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_lo_7 = {regroupV0_hi_hi_lo_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[663], regroupV0_hi_12[659]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[671], regroupV0_hi_12[667]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_lo_hi_7 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_lo_11 = {regroupV0_hi_hi_lo_hi_lo_lo_hi_7, regroupV0_hi_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[679], regroupV0_hi_12[675]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[687], regroupV0_hi_12[683]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_lo_7 = {regroupV0_hi_hi_lo_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[695], regroupV0_hi_12[691]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[703], regroupV0_hi_12[699]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_lo_hi_hi_7 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_lo_hi_11 = {regroupV0_hi_hi_lo_hi_lo_hi_hi_7, regroupV0_hi_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_lo_14 = {regroupV0_hi_hi_lo_hi_lo_hi_11, regroupV0_hi_hi_lo_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[711], regroupV0_hi_12[707]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[719], regroupV0_hi_12[715]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_lo_7 = {regroupV0_hi_hi_lo_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[727], regroupV0_hi_12[723]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[735], regroupV0_hi_12[731]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_lo_hi_7 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_lo_11 = {regroupV0_hi_hi_lo_hi_hi_lo_hi_7, regroupV0_hi_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[743], regroupV0_hi_12[739]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[751], regroupV0_hi_12[747]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_lo_7 = {regroupV0_hi_hi_lo_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[759], regroupV0_hi_12[755]};
  wire [1:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[767], regroupV0_hi_12[763]};
  wire [3:0]         regroupV0_hi_hi_lo_hi_hi_hi_hi_7 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_lo_hi_hi_hi_11 = {regroupV0_hi_hi_lo_hi_hi_hi_hi_7, regroupV0_hi_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_lo_hi_hi_14 = {regroupV0_hi_hi_lo_hi_hi_hi_11, regroupV0_hi_hi_lo_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_lo_hi_14 = {regroupV0_hi_hi_lo_hi_hi_14, regroupV0_hi_hi_lo_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_lo_14 = {regroupV0_hi_hi_lo_hi_14, regroupV0_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_3 = {regroupV0_hi_12[775], regroupV0_hi_12[771]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_3 = {regroupV0_hi_12[783], regroupV0_hi_12[779]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_lo_7 = {regroupV0_hi_hi_hi_lo_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_3 = {regroupV0_hi_12[791], regroupV0_hi_12[787]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_3 = {regroupV0_hi_12[799], regroupV0_hi_12[795]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_lo_hi_7 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_lo_11 = {regroupV0_hi_hi_hi_lo_lo_lo_hi_7, regroupV0_hi_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_3 = {regroupV0_hi_12[807], regroupV0_hi_12[803]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_3 = {regroupV0_hi_12[815], regroupV0_hi_12[811]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_lo_7 = {regroupV0_hi_hi_hi_lo_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_3 = {regroupV0_hi_12[823], regroupV0_hi_12[819]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_3 = {regroupV0_hi_12[831], regroupV0_hi_12[827]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_lo_hi_hi_7 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_lo_hi_11 = {regroupV0_hi_hi_hi_lo_lo_hi_hi_7, regroupV0_hi_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_lo_14 = {regroupV0_hi_hi_hi_lo_lo_hi_11, regroupV0_hi_hi_hi_lo_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_3 = {regroupV0_hi_12[839], regroupV0_hi_12[835]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_3 = {regroupV0_hi_12[847], regroupV0_hi_12[843]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_lo_7 = {regroupV0_hi_hi_hi_lo_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_3 = {regroupV0_hi_12[855], regroupV0_hi_12[851]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_3 = {regroupV0_hi_12[863], regroupV0_hi_12[859]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_lo_hi_7 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_lo_11 = {regroupV0_hi_hi_hi_lo_hi_lo_hi_7, regroupV0_hi_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_3 = {regroupV0_hi_12[871], regroupV0_hi_12[867]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_3 = {regroupV0_hi_12[879], regroupV0_hi_12[875]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_lo_7 = {regroupV0_hi_hi_hi_lo_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_3 = {regroupV0_hi_12[887], regroupV0_hi_12[883]};
  wire [1:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_3 = {regroupV0_hi_12[895], regroupV0_hi_12[891]};
  wire [3:0]         regroupV0_hi_hi_hi_lo_hi_hi_hi_7 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_lo_hi_hi_11 = {regroupV0_hi_hi_hi_lo_hi_hi_hi_7, regroupV0_hi_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_lo_hi_14 = {regroupV0_hi_hi_hi_lo_hi_hi_11, regroupV0_hi_hi_hi_lo_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_lo_hi_14, regroupV0_hi_hi_hi_lo_lo_14};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_3 = {regroupV0_hi_12[903], regroupV0_hi_12[899]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_3 = {regroupV0_hi_12[911], regroupV0_hi_12[907]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_lo_7 = {regroupV0_hi_hi_hi_hi_lo_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_3 = {regroupV0_hi_12[919], regroupV0_hi_12[915]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_3 = {regroupV0_hi_12[927], regroupV0_hi_12[923]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_lo_hi_7 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_lo_11 = {regroupV0_hi_hi_hi_hi_lo_lo_hi_7, regroupV0_hi_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_3 = {regroupV0_hi_12[935], regroupV0_hi_12[931]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_3 = {regroupV0_hi_12[943], regroupV0_hi_12[939]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_lo_7 = {regroupV0_hi_hi_hi_hi_lo_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_3 = {regroupV0_hi_12[951], regroupV0_hi_12[947]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_3 = {regroupV0_hi_12[959], regroupV0_hi_12[955]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_lo_hi_hi_7 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_lo_hi_11 = {regroupV0_hi_hi_hi_hi_lo_hi_hi_7, regroupV0_hi_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_lo_14 = {regroupV0_hi_hi_hi_hi_lo_hi_11, regroupV0_hi_hi_hi_hi_lo_lo_11};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_3 = {regroupV0_hi_12[967], regroupV0_hi_12[963]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_3 = {regroupV0_hi_12[975], regroupV0_hi_12[971]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_lo_7 = {regroupV0_hi_hi_hi_hi_hi_lo_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_3 = {regroupV0_hi_12[983], regroupV0_hi_12[979]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_3 = {regroupV0_hi_12[991], regroupV0_hi_12[987]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_lo_hi_7 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_lo_11 = {regroupV0_hi_hi_hi_hi_hi_lo_hi_7, regroupV0_hi_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_3 = {regroupV0_hi_12[999], regroupV0_hi_12[995]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_3 = {regroupV0_hi_12[1007], regroupV0_hi_12[1003]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_lo_7 = {regroupV0_hi_hi_hi_hi_hi_hi_lo_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_3 = {regroupV0_hi_12[1015], regroupV0_hi_12[1011]};
  wire [1:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_3 = {regroupV0_hi_12[1023], regroupV0_hi_12[1019]};
  wire [3:0]         regroupV0_hi_hi_hi_hi_hi_hi_hi_7 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_hi_3, regroupV0_hi_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]         regroupV0_hi_hi_hi_hi_hi_hi_11 = {regroupV0_hi_hi_hi_hi_hi_hi_hi_7, regroupV0_hi_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]        regroupV0_hi_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_hi_11, regroupV0_hi_hi_hi_hi_hi_lo_11};
  wire [31:0]        regroupV0_hi_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_hi_lo_14};
  wire [63:0]        regroupV0_hi_hi_hi_14 = {regroupV0_hi_hi_hi_hi_14, regroupV0_hi_hi_hi_lo_14};
  wire [127:0]       regroupV0_hi_hi_14 = {regroupV0_hi_hi_hi_14, regroupV0_hi_hi_lo_14};
  wire [255:0]       regroupV0_hi_16 = {regroupV0_hi_hi_14, regroupV0_hi_lo_14};
  wire [1023:0]      regroupV0_lo_17 = {regroupV0_hi_14, regroupV0_lo_14, regroupV0_hi_13, regroupV0_lo_13};
  wire [1023:0]      regroupV0_hi_17 = {regroupV0_hi_16, regroupV0_lo_16, regroupV0_hi_15, regroupV0_lo_15};
  wire [2047:0]      regroupV0_2 = {regroupV0_hi_17, regroupV0_lo_17};
  wire [3:0]         _v0SelectBySew_T = 4'h1 << laneMaskSewSelect_0;
  wire [511:0]       v0SelectBySew = (_v0SelectBySew_T[0] ? regroupV0_0[511:0] : 512'h0) | (_v0SelectBySew_T[1] ? regroupV0_1[511:0] : 512'h0) | (_v0SelectBySew_T[2] ? regroupV0_2[511:0] : 512'h0);
  wire [15:0][31:0]  _GEN_31 =
    {{v0SelectBySew[511:480]},
     {v0SelectBySew[479:448]},
     {v0SelectBySew[447:416]},
     {v0SelectBySew[415:384]},
     {v0SelectBySew[383:352]},
     {v0SelectBySew[351:320]},
     {v0SelectBySew[319:288]},
     {v0SelectBySew[287:256]},
     {v0SelectBySew[255:224]},
     {v0SelectBySew[223:192]},
     {v0SelectBySew[191:160]},
     {v0SelectBySew[159:128]},
     {v0SelectBySew[127:96]},
     {v0SelectBySew[95:64]},
     {v0SelectBySew[63:32]},
     {v0SelectBySew[31:0]}};
  wire [3:0]         _v0SelectBySew_T_9 = 4'h1 << laneMaskSewSelect_1;
  wire [511:0]       v0SelectBySew_1 = (_v0SelectBySew_T_9[0] ? regroupV0_0[1023:512] : 512'h0) | (_v0SelectBySew_T_9[1] ? regroupV0_1[1023:512] : 512'h0) | (_v0SelectBySew_T_9[2] ? regroupV0_2[1023:512] : 512'h0);
  wire [15:0][31:0]  _GEN_32 =
    {{v0SelectBySew_1[511:480]},
     {v0SelectBySew_1[479:448]},
     {v0SelectBySew_1[447:416]},
     {v0SelectBySew_1[415:384]},
     {v0SelectBySew_1[383:352]},
     {v0SelectBySew_1[351:320]},
     {v0SelectBySew_1[319:288]},
     {v0SelectBySew_1[287:256]},
     {v0SelectBySew_1[255:224]},
     {v0SelectBySew_1[223:192]},
     {v0SelectBySew_1[191:160]},
     {v0SelectBySew_1[159:128]},
     {v0SelectBySew_1[127:96]},
     {v0SelectBySew_1[95:64]},
     {v0SelectBySew_1[63:32]},
     {v0SelectBySew_1[31:0]}};
  wire [3:0]         _v0SelectBySew_T_18 = 4'h1 << laneMaskSewSelect_2;
  wire [511:0]       v0SelectBySew_2 = (_v0SelectBySew_T_18[0] ? regroupV0_0[1535:1024] : 512'h0) | (_v0SelectBySew_T_18[1] ? regroupV0_1[1535:1024] : 512'h0) | (_v0SelectBySew_T_18[2] ? regroupV0_2[1535:1024] : 512'h0);
  wire [15:0][31:0]  _GEN_33 =
    {{v0SelectBySew_2[511:480]},
     {v0SelectBySew_2[479:448]},
     {v0SelectBySew_2[447:416]},
     {v0SelectBySew_2[415:384]},
     {v0SelectBySew_2[383:352]},
     {v0SelectBySew_2[351:320]},
     {v0SelectBySew_2[319:288]},
     {v0SelectBySew_2[287:256]},
     {v0SelectBySew_2[255:224]},
     {v0SelectBySew_2[223:192]},
     {v0SelectBySew_2[191:160]},
     {v0SelectBySew_2[159:128]},
     {v0SelectBySew_2[127:96]},
     {v0SelectBySew_2[95:64]},
     {v0SelectBySew_2[63:32]},
     {v0SelectBySew_2[31:0]}};
  wire [3:0]         _v0SelectBySew_T_27 = 4'h1 << laneMaskSewSelect_3;
  wire [511:0]       v0SelectBySew_3 = (_v0SelectBySew_T_27[0] ? regroupV0_0[2047:1536] : 512'h0) | (_v0SelectBySew_T_27[1] ? regroupV0_1[2047:1536] : 512'h0) | (_v0SelectBySew_T_27[2] ? regroupV0_2[2047:1536] : 512'h0);
  wire [15:0][31:0]  _GEN_34 =
    {{v0SelectBySew_3[511:480]},
     {v0SelectBySew_3[479:448]},
     {v0SelectBySew_3[447:416]},
     {v0SelectBySew_3[415:384]},
     {v0SelectBySew_3[383:352]},
     {v0SelectBySew_3[351:320]},
     {v0SelectBySew_3[319:288]},
     {v0SelectBySew_3[287:256]},
     {v0SelectBySew_3[255:224]},
     {v0SelectBySew_3[223:192]},
     {v0SelectBySew_3[191:160]},
     {v0SelectBySew_3[159:128]},
     {v0SelectBySew_3[127:96]},
     {v0SelectBySew_3[95:64]},
     {v0SelectBySew_3[63:32]},
     {v0SelectBySew_3[31:0]}};
  wire [3:0]         intLMULInput = 4'h1 << instReq_bits_vlmul[1:0];
  wire [13:0]        _dataPosition_T_1 = {3'h0, instReq_bits_readFromScala[10:0]} << instReq_bits_sew;
  wire [10:0]        dataPosition = _dataPosition_T_1[10:0];
  wire [3:0]         _sewOHInput_T = 4'h1 << instReq_bits_sew;
  wire [2:0]         sewOHInput = _sewOHInput_T[2:0];
  wire [1:0]         dataOffset = {dataPosition[1] & (|(sewOHInput[1:0])), dataPosition[0] & sewOHInput[0]};
  wire [1:0]         accessLane = dataPosition[3:2];
  wire [6:0]         dataGroup = dataPosition[10:4];
  wire [3:0]         offset = dataGroup[3:0];
  wire [2:0]         accessRegGrowth = dataGroup[6:4];
  wire [2:0]         reallyGrowth = accessRegGrowth;
  wire [5:0]         decimalProportion = {offset, accessLane};
  wire [2:0]         decimal = decimalProportion[5:3];
  wire               notNeedRead = |{instReq_bits_vlmul[2] & decimal >= intLMULInput[3:1] | ~(instReq_bits_vlmul[2]) & {1'h0, accessRegGrowth} >= intLMULInput, instReq_bits_readFromScala[31:11]};
  reg  [1:0]         gatherReadState;
  wire               gatherSRead = gatherReadState == 2'h1;
  wire               gatherWaiteRead = gatherReadState == 2'h2;
  assign gatherResponse = &gatherReadState;
  wire               gatherData_valid_0 = gatherResponse;
  reg  [1:0]         gatherDatOffset;
  reg  [1:0]         gatherLane;
  reg  [3:0]         gatherOffset;
  reg  [2:0]         gatherGrowth;
  reg  [2:0]         instReg_instructionIndex;
  wire [2:0]         exeResp_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         exeResp_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_0_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_1_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_2_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         readChannel_3_bits_instructionIndex_0 = instReg_instructionIndex;
  wire [2:0]         writeRequest_0_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_1_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_2_index = instReg_instructionIndex;
  wire [2:0]         writeRequest_3_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_0_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_1_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_2_enq_bits_index = instReg_instructionIndex;
  wire [2:0]         writeQueue_3_enq_bits_index = instReg_instructionIndex;
  reg                instReg_decodeResult_specialSlot;
  reg  [4:0]         instReg_decodeResult_topUop;
  reg                instReg_decodeResult_popCount;
  reg                instReg_decodeResult_ffo;
  reg                instReg_decodeResult_average;
  reg                instReg_decodeResult_reverse;
  reg                instReg_decodeResult_dontNeedExecuteInLane;
  reg                instReg_decodeResult_scheduler;
  reg                instReg_decodeResult_sReadVD;
  reg                instReg_decodeResult_vtype;
  reg                instReg_decodeResult_sWrite;
  reg                instReg_decodeResult_crossRead;
  reg                instReg_decodeResult_crossWrite;
  reg                instReg_decodeResult_maskUnit;
  reg                instReg_decodeResult_special;
  reg                instReg_decodeResult_saturate;
  reg                instReg_decodeResult_vwmacc;
  reg                instReg_decodeResult_readOnly;
  reg                instReg_decodeResult_maskSource;
  reg                instReg_decodeResult_maskDestination;
  reg                instReg_decodeResult_maskLogic;
  reg  [3:0]         instReg_decodeResult_uop;
  reg                instReg_decodeResult_iota;
  reg                instReg_decodeResult_mv;
  reg                instReg_decodeResult_extend;
  reg                instReg_decodeResult_unOrderWrite;
  reg                instReg_decodeResult_compress;
  reg                instReg_decodeResult_gather16;
  reg                instReg_decodeResult_gather;
  reg                instReg_decodeResult_slid;
  reg                instReg_decodeResult_targetRd;
  reg                instReg_decodeResult_widenReduce;
  reg                instReg_decodeResult_red;
  reg                instReg_decodeResult_nr;
  reg                instReg_decodeResult_itype;
  reg                instReg_decodeResult_unsigned1;
  reg                instReg_decodeResult_unsigned0;
  reg                instReg_decodeResult_other;
  reg                instReg_decodeResult_multiCycle;
  reg                instReg_decodeResult_divider;
  reg                instReg_decodeResult_multiplier;
  reg                instReg_decodeResult_shift;
  reg                instReg_decodeResult_adder;
  reg                instReg_decodeResult_logic;
  reg  [31:0]        instReg_readFromScala;
  reg  [1:0]         instReg_sew;
  reg  [2:0]         instReg_vlmul;
  reg                instReg_maskType;
  reg  [2:0]         instReg_vxrm;
  reg  [4:0]         instReg_vs2;
  reg  [4:0]         instReg_vs1;
  reg  [4:0]         instReg_vd;
  wire [4:0]         writeRequest_0_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_1_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_2_writeData_vd = instReg_vd;
  wire [4:0]         writeRequest_3_writeData_vd = instReg_vd;
  reg  [11:0]        instReg_vl;
  wire [11:0]        reduceLastDataNeed_byteForVl = instReg_vl;
  wire               enqMvRD = instReq_bits_decodeResult_topUop == 5'hB;
  reg                instVlValid;
  wire               gatherRequestFire = gatherReadState == 2'h0 & gatherRead & ~instVlValid;
  wire               viotaReq = instReq_bits_decodeResult_topUop == 5'h8;
  reg                readVS1Reg_dataValid;
  reg                readVS1Reg_requestSend;
  reg                readVS1Reg_sendToExecution;
  reg  [31:0]        readVS1Reg_data;
  reg  [6:0]         readVS1Reg_readIndex;
  wire [3:0]         _sew1H_T = 4'h1 << instReg_sew;
  wire [2:0]         sew1H = _sew1H_T[2:0];
  wire [3:0]         unitType = 4'h1 << instReg_decodeResult_topUop[4:3];
  wire [3:0]         subType = 4'h1 << instReg_decodeResult_topUop[2:1];
  wire               readType = unitType[0];
  wire               gather16 = instReg_decodeResult_topUop == 5'h5;
  wire               maskDestinationType = instReg_decodeResult_topUop == 5'h18;
  wire               compress = instReg_decodeResult_topUop[4:1] == 4'h4;
  wire               viota = instReg_decodeResult_topUop == 5'h8;
  wire               mv = instReg_decodeResult_topUop[4:1] == 4'h5;
  wire               mvRd = instReg_decodeResult_topUop == 5'hB;
  wire               mvVd = instReg_decodeResult_topUop == 5'hA;
  wire               orderReduce = {instReg_decodeResult_topUop[4:2], instReg_decodeResult_topUop[0]} == 4'hB;
  wire               ffo = instReg_decodeResult_topUop[4:1] == 4'h7;
  wire               extendType = unitType[3] & (subType[2] | subType[1]);
  wire               readValid = readType & instVlValid;
  wire               noSource = mv | viota;
  wire               allGroupExecute = maskDestinationType | unitType[2] | compress | ffo;
  wire               useDefaultSew = readType & ~gather16;
  wire [1:0]         _dataSplitSew_T_11 = useDefaultSew ? instReg_sew : 2'h0;
  wire [1:0]         dataSplitSew = {_dataSplitSew_T_11[1], _dataSplitSew_T_11[0] | unitType[3] & subType[1] | gather16} | {allGroupExecute, 1'h0};
  wire               sourceDataUseDefaultSew = ~(unitType[3] | gather16);
  wire [1:0]         _sourceDataEEW_T_6 = (sourceDataUseDefaultSew ? instReg_sew : 2'h0) | (unitType[3] ? instReg_sew >> subType[2:1] : 2'h0);
  wire [1:0]         sourceDataEEW = {_sourceDataEEW_T_6[1], _sourceDataEEW_T_6[0] | gather16};
  wire [3:0]         executeIndexGrowth = 4'h1 << dataSplitSew;
  wire [1:0]         lastExecuteIndex = {2{executeIndexGrowth[0]}} | {executeIndexGrowth[1], 1'h0};
  wire [3:0]         _sourceDataEEW1H_T = 4'h1 << sourceDataEEW;
  wire [2:0]         sourceDataEEW1H = _sourceDataEEW1H_T[2:0];
  wire [10:0]        lastElementIndex = instReg_vl[10:0] - {10'h0, |instReg_vl};
  wire [10:0]        processingVl_lastByteIndex = lastElementIndex;
  wire               maskFormatSource = ffo | maskDestinationType;
  wire [3:0]         processingVl_lastGroupRemaining = processingVl_lastByteIndex[3:0];
  wire [6:0]         processingVl_0_1 = processingVl_lastByteIndex[10:4];
  wire [1:0]         processingVl_lastLaneIndex = processingVl_lastGroupRemaining[3:2];
  wire [3:0]         _processingVl_lastGroupDataNeed_T = 4'h1 << processingVl_lastLaneIndex;
  wire [2:0]         _GEN_35 = _processingVl_lastGroupDataNeed_T[2:0] | _processingVl_lastGroupDataNeed_T[3:1];
  wire [3:0]         processingVl_0_2 = {_processingVl_lastGroupDataNeed_T[3], _GEN_35[2], _GEN_35[1:0] | {_processingVl_lastGroupDataNeed_T[3], _GEN_35[2]}};
  wire [11:0]        processingVl_lastByteIndex_1 = {lastElementIndex, 1'h0};
  wire [3:0]         processingVl_lastGroupRemaining_1 = processingVl_lastByteIndex_1[3:0];
  wire [7:0]         processingVl_1_1 = processingVl_lastByteIndex_1[11:4];
  wire [1:0]         processingVl_lastLaneIndex_1 = processingVl_lastGroupRemaining_1[3:2];
  wire [3:0]         _processingVl_lastGroupDataNeed_T_5 = 4'h1 << processingVl_lastLaneIndex_1;
  wire [2:0]         _GEN_36 = _processingVl_lastGroupDataNeed_T_5[2:0] | _processingVl_lastGroupDataNeed_T_5[3:1];
  wire [3:0]         processingVl_1_2 = {_processingVl_lastGroupDataNeed_T_5[3], _GEN_36[2], _GEN_36[1:0] | {_processingVl_lastGroupDataNeed_T_5[3], _GEN_36[2]}};
  wire [12:0]        processingVl_lastByteIndex_2 = {lastElementIndex, 2'h0};
  wire [3:0]         processingVl_lastGroupRemaining_2 = processingVl_lastByteIndex_2[3:0];
  wire [8:0]         processingVl_2_1 = processingVl_lastByteIndex_2[12:4];
  wire [1:0]         processingVl_lastLaneIndex_2 = processingVl_lastGroupRemaining_2[3:2];
  wire [3:0]         _processingVl_lastGroupDataNeed_T_10 = 4'h1 << processingVl_lastLaneIndex_2;
  wire [2:0]         _GEN_37 = _processingVl_lastGroupDataNeed_T_10[2:0] | _processingVl_lastGroupDataNeed_T_10[3:1];
  wire [3:0]         processingVl_2_2 = {_processingVl_lastGroupDataNeed_T_10[3], _GEN_37[2], _GEN_37[1:0] | {_processingVl_lastGroupDataNeed_T_10[3], _GEN_37[2]}};
  wire [6:0]         processingMaskVl_lastGroupRemaining = lastElementIndex[6:0];
  wire [6:0]         elementTailForMaskDestination = lastElementIndex[6:0];
  wire               processingMaskVl_lastGroupMisAlign = |processingMaskVl_lastGroupRemaining;
  wire [3:0]         processingMaskVl_0_1 = lastElementIndex[10:7];
  wire [1:0]         processingMaskVl_lastLaneIndex = processingMaskVl_lastGroupRemaining[6:5] - {1'h0, processingMaskVl_lastGroupRemaining[4:0] == 5'h0};
  wire [3:0]         _processingMaskVl_dataNeedForPL_T = 4'h1 << processingMaskVl_lastLaneIndex;
  wire [2:0]         _GEN_38 = _processingMaskVl_dataNeedForPL_T[2:0] | _processingMaskVl_dataNeedForPL_T[3:1];
  wire [3:0]         processingMaskVl_dataNeedForPL = {_processingMaskVl_dataNeedForPL_T[3], _GEN_38[2], _GEN_38[1:0] | {_processingMaskVl_dataNeedForPL_T[3], _GEN_38[2]}};
  wire               processingMaskVl_dataNeedForNPL_misAlign = |(processingMaskVl_lastGroupRemaining[1:0]);
  wire [5:0]         processingMaskVl_dataNeedForNPL_datapathSize = {1'h0, processingMaskVl_lastGroupRemaining[6:2]} + {5'h0, processingMaskVl_dataNeedForNPL_misAlign};
  wire               processingMaskVl_dataNeedForNPL_allNeed = |(processingMaskVl_dataNeedForNPL_datapathSize[5:2]);
  wire [1:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex = processingMaskVl_dataNeedForNPL_datapathSize[1:0];
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex;
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_3 = _processingMaskVl_dataNeedForNPL_dataNeed_T | {_processingMaskVl_dataNeedForNPL_dataNeed_T[2:0], 1'h0};
  wire [3:0]         processingMaskVl_dataNeedForNPL_dataNeed = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_3 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_3[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed}};
  wire               processingMaskVl_dataNeedForNPL_misAlign_1 = processingMaskVl_lastGroupRemaining[0];
  wire [6:0]         processingMaskVl_dataNeedForNPL_datapathSize_1 = {1'h0, processingMaskVl_lastGroupRemaining[6:1]} + {6'h0, processingMaskVl_dataNeedForNPL_misAlign_1};
  wire               processingMaskVl_dataNeedForNPL_allNeed_1 = |(processingMaskVl_dataNeedForNPL_datapathSize_1[6:2]);
  wire [1:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex_1 = processingMaskVl_dataNeedForNPL_datapathSize_1[1:0];
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_10 = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_1;
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_13 = _processingMaskVl_dataNeedForNPL_dataNeed_T_10 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_10[2:0], 1'h0};
  wire [3:0]         processingMaskVl_dataNeedForNPL_dataNeed_1 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_13 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_13[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed_1}};
  wire [7:0]         processingMaskVl_dataNeedForNPL_datapathSize_2 = {1'h0, processingMaskVl_lastGroupRemaining};
  wire               processingMaskVl_dataNeedForNPL_allNeed_2 = |(processingMaskVl_dataNeedForNPL_datapathSize_2[7:2]);
  wire [1:0]         processingMaskVl_dataNeedForNPL_lastLaneIndex_2 = processingMaskVl_dataNeedForNPL_datapathSize_2[1:0];
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_20 = 4'h1 << processingMaskVl_dataNeedForNPL_lastLaneIndex_2;
  wire [3:0]         _processingMaskVl_dataNeedForNPL_dataNeed_T_23 = _processingMaskVl_dataNeedForNPL_dataNeed_T_20 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_20[2:0], 1'h0};
  wire [3:0]         processingMaskVl_dataNeedForNPL_dataNeed_2 = ~(_processingMaskVl_dataNeedForNPL_dataNeed_T_23 | {_processingMaskVl_dataNeedForNPL_dataNeed_T_23[1:0], 2'h0}) | {4{processingMaskVl_dataNeedForNPL_allNeed_2}};
  wire [3:0]         processingMaskVl_dataNeedForNPL =
    (sew1H[0] ? processingMaskVl_dataNeedForNPL_dataNeed : 4'h0) | (sew1H[1] ? processingMaskVl_dataNeedForNPL_dataNeed_1 : 4'h0) | (sew1H[2] ? processingMaskVl_dataNeedForNPL_dataNeed_2 : 4'h0);
  wire [3:0]         processingMaskVl_0_2 = ffo ? processingMaskVl_dataNeedForPL : processingMaskVl_dataNeedForNPL;
  wire               reduceLastDataNeed_vlMSB = |(reduceLastDataNeed_byteForVl[11:4]);
  wire [3:0]         reduceLastDataNeed_vlLSB = instReg_vl[3:0];
  wire [3:0]         reduceLastDataNeed_vlLSB_1 = instReg_vl[3:0];
  wire [3:0]         reduceLastDataNeed_vlLSB_2 = instReg_vl[3:0];
  wire [1:0]         reduceLastDataNeed_lsbDSize = reduceLastDataNeed_vlLSB[3:2] - {1'h0, reduceLastDataNeed_vlLSB[1:0] == 2'h0};
  wire [3:0]         _reduceLastDataNeed_T = 4'h1 << reduceLastDataNeed_lsbDSize;
  wire [2:0]         _GEN_39 = _reduceLastDataNeed_T[2:0] | _reduceLastDataNeed_T[3:1];
  wire [12:0]        reduceLastDataNeed_byteForVl_1 = {instReg_vl, 1'h0};
  wire               reduceLastDataNeed_vlMSB_1 = |(reduceLastDataNeed_byteForVl_1[12:4]);
  wire [1:0]         reduceLastDataNeed_lsbDSize_1 = reduceLastDataNeed_vlLSB_1[3:2] - {1'h0, reduceLastDataNeed_vlLSB_1[1:0] == 2'h0};
  wire [3:0]         _reduceLastDataNeed_T_8 = 4'h1 << reduceLastDataNeed_lsbDSize_1;
  wire [2:0]         _GEN_40 = _reduceLastDataNeed_T_8[2:0] | _reduceLastDataNeed_T_8[3:1];
  wire [13:0]        reduceLastDataNeed_byteForVl_2 = {instReg_vl, 2'h0};
  wire               reduceLastDataNeed_vlMSB_2 = |(reduceLastDataNeed_byteForVl_2[13:4]);
  wire [1:0]         reduceLastDataNeed_lsbDSize_2 = reduceLastDataNeed_vlLSB_2[3:2] - {1'h0, reduceLastDataNeed_vlLSB_2[1:0] == 2'h0};
  wire [3:0]         _reduceLastDataNeed_T_16 = 4'h1 << reduceLastDataNeed_lsbDSize_2;
  wire [2:0]         _GEN_41 = _reduceLastDataNeed_T_16[2:0] | _reduceLastDataNeed_T_16[3:1];
  wire [3:0]         reduceLastDataNeed =
    (sew1H[0] ? {_reduceLastDataNeed_T[3], _GEN_39[2], _GEN_39[1:0] | {_reduceLastDataNeed_T[3], _GEN_39[2]}} | {4{reduceLastDataNeed_vlMSB}} : 4'h0)
    | (sew1H[1] ? {_reduceLastDataNeed_T_8[3], _GEN_40[2], _GEN_40[1:0] | {_reduceLastDataNeed_T_8[3], _GEN_40[2]}} | {4{reduceLastDataNeed_vlMSB_1}} : 4'h0)
    | (sew1H[2] ? {_reduceLastDataNeed_T_16[3], _GEN_41[2], _GEN_41[1:0] | {_reduceLastDataNeed_T_16[3], _GEN_41[2]}} | {4{reduceLastDataNeed_vlMSB_2}} : 4'h0);
  wire [1:0]         dataSourceSew = unitType[3] ? instReg_sew - instReg_decodeResult_topUop[2:1] : gather16 ? 2'h1 : instReg_sew;
  wire [3:0]         _dataSourceSew1H_T = 4'h1 << dataSourceSew;
  wire [2:0]         dataSourceSew1H = _dataSourceSew1H_T[2:0];
  wire               unorderReduce = ~orderReduce & unitType[2];
  wire               normalFormat = ~maskFormatSource & ~unorderReduce & ~mv;
  wire [8:0]         lastGroupForInstruction =
    {1'h0, {1'h0, {3'h0, maskFormatSource ? processingMaskVl_0_1 : 4'h0} | (normalFormat & dataSourceSew1H[0] ? processingVl_0_1 : 7'h0)} | (normalFormat & dataSourceSew1H[1] ? processingVl_1_1 : 8'h0)}
    | (normalFormat & dataSourceSew1H[2] ? processingVl_2_1 : 9'h0);
  wire [5:0]         popDataNeed_dataPathGroups = lastElementIndex[10:5];
  wire [1:0]         popDataNeed_lastLaneIndex = popDataNeed_dataPathGroups[1:0];
  wire               popDataNeed_lagerThanDLen = |(popDataNeed_dataPathGroups[5:2]);
  wire [3:0]         _popDataNeed_T = 4'h1 << popDataNeed_lastLaneIndex;
  wire [2:0]         _GEN_42 = _popDataNeed_T[2:0] | _popDataNeed_T[3:1];
  wire [3:0]         popDataNeed = {_popDataNeed_T[3], _GEN_42[2], _GEN_42[1:0] | {_popDataNeed_T[3], _GEN_42[2]}} | {4{popDataNeed_lagerThanDLen}};
  wire [3:0]         lastGroupDataNeed =
    (unorderReduce & instReg_decodeResult_popCount ? popDataNeed : 4'h0) | (unorderReduce & ~instReg_decodeResult_popCount ? reduceLastDataNeed : 4'h0) | (maskFormatSource ? processingMaskVl_0_2 : 4'h0)
    | (normalFormat & dataSourceSew1H[0] ? processingVl_0_2 : 4'h0) | (normalFormat & dataSourceSew1H[1] ? processingVl_1_2 : 4'h0) | (normalFormat & dataSourceSew1H[2] ? processingVl_2_2 : 4'h0);
  wire [3:0]         exeRequestQueue_queue_dataIn_lo = {exeRequestQueue_0_enq_bits_index, exeRequestQueue_0_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi = {exeRequestQueue_0_enq_bits_source1, exeRequestQueue_0_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn = {exeRequestQueue_queue_dataIn_hi, exeRequestQueue_queue_dataIn_lo};
  wire               exeRequestQueue_queue_dataOut_ffo = _exeRequestQueue_queue_fifo_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_index = _exeRequestQueue_queue_fifo_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_source2 = _exeRequestQueue_queue_fifo_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_source1 = _exeRequestQueue_queue_fifo_data_out[67:36];
  wire               exeRequestQueue_0_enq_ready = ~_exeRequestQueue_queue_fifo_full;
  wire               exeRequestQueue_0_deq_ready;
  wire               exeRequestQueue_0_deq_valid = ~_exeRequestQueue_queue_fifo_empty | exeRequestQueue_0_enq_valid;
  wire [31:0]        exeRequestQueue_0_deq_bits_source1 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source1 : exeRequestQueue_queue_dataOut_source1;
  wire [31:0]        exeRequestQueue_0_deq_bits_source2 = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_source2 : exeRequestQueue_queue_dataOut_source2;
  wire [2:0]         exeRequestQueue_0_deq_bits_index = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_index : exeRequestQueue_queue_dataOut_index;
  wire               exeRequestQueue_0_deq_bits_ffo = _exeRequestQueue_queue_fifo_empty ? exeRequestQueue_0_enq_bits_ffo : exeRequestQueue_queue_dataOut_ffo;
  wire               tokenIO_0_maskRequestRelease_0 = exeRequestQueue_0_deq_ready & exeRequestQueue_0_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_1 = {exeRequestQueue_1_enq_bits_index, exeRequestQueue_1_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_1 = {exeRequestQueue_1_enq_bits_source1, exeRequestQueue_1_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_1 = {exeRequestQueue_queue_dataIn_hi_1, exeRequestQueue_queue_dataIn_lo_1};
  wire               exeRequestQueue_queue_dataOut_1_ffo = _exeRequestQueue_queue_fifo_1_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_1_index = _exeRequestQueue_queue_fifo_1_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_1_source2 = _exeRequestQueue_queue_fifo_1_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_1_source1 = _exeRequestQueue_queue_fifo_1_data_out[67:36];
  wire               exeRequestQueue_1_enq_ready = ~_exeRequestQueue_queue_fifo_1_full;
  wire               exeRequestQueue_1_deq_ready;
  wire               exeRequestQueue_1_deq_valid = ~_exeRequestQueue_queue_fifo_1_empty | exeRequestQueue_1_enq_valid;
  wire [31:0]        exeRequestQueue_1_deq_bits_source1 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source1 : exeRequestQueue_queue_dataOut_1_source1;
  wire [31:0]        exeRequestQueue_1_deq_bits_source2 = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_source2 : exeRequestQueue_queue_dataOut_1_source2;
  wire [2:0]         exeRequestQueue_1_deq_bits_index = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_index : exeRequestQueue_queue_dataOut_1_index;
  wire               exeRequestQueue_1_deq_bits_ffo = _exeRequestQueue_queue_fifo_1_empty ? exeRequestQueue_1_enq_bits_ffo : exeRequestQueue_queue_dataOut_1_ffo;
  wire               tokenIO_1_maskRequestRelease_0 = exeRequestQueue_1_deq_ready & exeRequestQueue_1_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_2 = {exeRequestQueue_2_enq_bits_index, exeRequestQueue_2_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_2 = {exeRequestQueue_2_enq_bits_source1, exeRequestQueue_2_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_2 = {exeRequestQueue_queue_dataIn_hi_2, exeRequestQueue_queue_dataIn_lo_2};
  wire               exeRequestQueue_queue_dataOut_2_ffo = _exeRequestQueue_queue_fifo_2_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_2_index = _exeRequestQueue_queue_fifo_2_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_2_source2 = _exeRequestQueue_queue_fifo_2_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_2_source1 = _exeRequestQueue_queue_fifo_2_data_out[67:36];
  wire               exeRequestQueue_2_enq_ready = ~_exeRequestQueue_queue_fifo_2_full;
  wire               exeRequestQueue_2_deq_ready;
  wire               exeRequestQueue_2_deq_valid = ~_exeRequestQueue_queue_fifo_2_empty | exeRequestQueue_2_enq_valid;
  wire [31:0]        exeRequestQueue_2_deq_bits_source1 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source1 : exeRequestQueue_queue_dataOut_2_source1;
  wire [31:0]        exeRequestQueue_2_deq_bits_source2 = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_source2 : exeRequestQueue_queue_dataOut_2_source2;
  wire [2:0]         exeRequestQueue_2_deq_bits_index = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_index : exeRequestQueue_queue_dataOut_2_index;
  wire               exeRequestQueue_2_deq_bits_ffo = _exeRequestQueue_queue_fifo_2_empty ? exeRequestQueue_2_enq_bits_ffo : exeRequestQueue_queue_dataOut_2_ffo;
  wire               tokenIO_2_maskRequestRelease_0 = exeRequestQueue_2_deq_ready & exeRequestQueue_2_deq_valid;
  wire [3:0]         exeRequestQueue_queue_dataIn_lo_3 = {exeRequestQueue_3_enq_bits_index, exeRequestQueue_3_enq_bits_ffo};
  wire [63:0]        exeRequestQueue_queue_dataIn_hi_3 = {exeRequestQueue_3_enq_bits_source1, exeRequestQueue_3_enq_bits_source2};
  wire [67:0]        exeRequestQueue_queue_dataIn_3 = {exeRequestQueue_queue_dataIn_hi_3, exeRequestQueue_queue_dataIn_lo_3};
  wire               exeRequestQueue_queue_dataOut_3_ffo = _exeRequestQueue_queue_fifo_3_data_out[0];
  wire [2:0]         exeRequestQueue_queue_dataOut_3_index = _exeRequestQueue_queue_fifo_3_data_out[3:1];
  wire [31:0]        exeRequestQueue_queue_dataOut_3_source2 = _exeRequestQueue_queue_fifo_3_data_out[35:4];
  wire [31:0]        exeRequestQueue_queue_dataOut_3_source1 = _exeRequestQueue_queue_fifo_3_data_out[67:36];
  wire               exeRequestQueue_3_enq_ready = ~_exeRequestQueue_queue_fifo_3_full;
  wire               exeRequestQueue_3_deq_ready;
  wire               exeRequestQueue_3_deq_valid = ~_exeRequestQueue_queue_fifo_3_empty | exeRequestQueue_3_enq_valid;
  wire [31:0]        exeRequestQueue_3_deq_bits_source1 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source1 : exeRequestQueue_queue_dataOut_3_source1;
  wire [31:0]        exeRequestQueue_3_deq_bits_source2 = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_source2 : exeRequestQueue_queue_dataOut_3_source2;
  wire [2:0]         exeRequestQueue_3_deq_bits_index = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_index : exeRequestQueue_queue_dataOut_3_index;
  wire               exeRequestQueue_3_deq_bits_ffo = _exeRequestQueue_queue_fifo_3_empty ? exeRequestQueue_3_enq_bits_ffo : exeRequestQueue_queue_dataOut_3_ffo;
  wire               tokenIO_3_maskRequestRelease_0 = exeRequestQueue_3_deq_ready & exeRequestQueue_3_deq_valid;
  reg                exeReqReg_0_valid;
  reg  [31:0]        exeReqReg_0_bits_source1;
  reg  [31:0]        exeReqReg_0_bits_source2;
  reg  [2:0]         exeReqReg_0_bits_index;
  reg                exeReqReg_0_bits_ffo;
  reg                exeReqReg_1_valid;
  reg  [31:0]        exeReqReg_1_bits_source1;
  reg  [31:0]        exeReqReg_1_bits_source2;
  reg  [2:0]         exeReqReg_1_bits_index;
  reg                exeReqReg_1_bits_ffo;
  reg                exeReqReg_2_valid;
  reg  [31:0]        exeReqReg_2_bits_source1;
  reg  [31:0]        exeReqReg_2_bits_source2;
  reg  [2:0]         exeReqReg_2_bits_index;
  reg                exeReqReg_2_bits_ffo;
  reg                exeReqReg_3_valid;
  reg  [31:0]        exeReqReg_3_bits_source1;
  reg  [31:0]        exeReqReg_3_bits_source2;
  reg  [2:0]         exeReqReg_3_bits_index;
  reg                exeReqReg_3_bits_ffo;
  reg  [7:0]         requestCounter;
  wire [8:0]         _GEN_43 = {1'h0, requestCounter};
  wire               counterValid = _GEN_43 <= lastGroupForInstruction;
  wire               lastGroup = _GEN_43 == lastGroupForInstruction | ~orderReduce & unitType[2] | mv;
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_lo_hi = {slideAddressGen_slideMaskInput_lo_lo_hi_hi, slideAddressGen_slideMaskInput_lo_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_lo = {slideAddressGen_slideMaskInput_lo_lo_hi, slideAddressGen_slideMaskInput_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_lo = {slideAddressGen_slideMaskInput_lo_hi_hi_lo_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_lo_hi_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_lo_hi_hi = {slideAddressGen_slideMaskInput_lo_hi_hi_hi, slideAddressGen_slideMaskInput_lo_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_lo_hi = {slideAddressGen_slideMaskInput_lo_hi_hi, slideAddressGen_slideMaskInput_lo_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_lo = {slideAddressGen_slideMaskInput_lo_hi, slideAddressGen_slideMaskInput_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_lo_hi_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_lo_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_lo = {slideAddressGen_slideMaskInput_hi_lo_hi, slideAddressGen_slideMaskInput_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_lo_hi = {slideAddressGen_slideMaskInput_hi_hi_lo_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_lo = {slideAddressGen_slideMaskInput_hi_hi_hi_lo_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo_lo};
  wire [127:0]       slideAddressGen_slideMaskInput_hi_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_hi_lo};
  wire [255:0]       slideAddressGen_slideMaskInput_hi_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_hi_lo};
  wire [511:0]       slideAddressGen_slideMaskInput_hi_hi = {slideAddressGen_slideMaskInput_hi_hi_hi, slideAddressGen_slideMaskInput_hi_hi_lo};
  wire [1023:0]      slideAddressGen_slideMaskInput_hi = {slideAddressGen_slideMaskInput_hi_hi, slideAddressGen_slideMaskInput_hi_lo};
  wire [511:0][3:0]  _GEN_44 =
    {{slideAddressGen_slideMaskInput_hi[1023:1020]},
     {slideAddressGen_slideMaskInput_hi[1019:1016]},
     {slideAddressGen_slideMaskInput_hi[1015:1012]},
     {slideAddressGen_slideMaskInput_hi[1011:1008]},
     {slideAddressGen_slideMaskInput_hi[1007:1004]},
     {slideAddressGen_slideMaskInput_hi[1003:1000]},
     {slideAddressGen_slideMaskInput_hi[999:996]},
     {slideAddressGen_slideMaskInput_hi[995:992]},
     {slideAddressGen_slideMaskInput_hi[991:988]},
     {slideAddressGen_slideMaskInput_hi[987:984]},
     {slideAddressGen_slideMaskInput_hi[983:980]},
     {slideAddressGen_slideMaskInput_hi[979:976]},
     {slideAddressGen_slideMaskInput_hi[975:972]},
     {slideAddressGen_slideMaskInput_hi[971:968]},
     {slideAddressGen_slideMaskInput_hi[967:964]},
     {slideAddressGen_slideMaskInput_hi[963:960]},
     {slideAddressGen_slideMaskInput_hi[959:956]},
     {slideAddressGen_slideMaskInput_hi[955:952]},
     {slideAddressGen_slideMaskInput_hi[951:948]},
     {slideAddressGen_slideMaskInput_hi[947:944]},
     {slideAddressGen_slideMaskInput_hi[943:940]},
     {slideAddressGen_slideMaskInput_hi[939:936]},
     {slideAddressGen_slideMaskInput_hi[935:932]},
     {slideAddressGen_slideMaskInput_hi[931:928]},
     {slideAddressGen_slideMaskInput_hi[927:924]},
     {slideAddressGen_slideMaskInput_hi[923:920]},
     {slideAddressGen_slideMaskInput_hi[919:916]},
     {slideAddressGen_slideMaskInput_hi[915:912]},
     {slideAddressGen_slideMaskInput_hi[911:908]},
     {slideAddressGen_slideMaskInput_hi[907:904]},
     {slideAddressGen_slideMaskInput_hi[903:900]},
     {slideAddressGen_slideMaskInput_hi[899:896]},
     {slideAddressGen_slideMaskInput_hi[895:892]},
     {slideAddressGen_slideMaskInput_hi[891:888]},
     {slideAddressGen_slideMaskInput_hi[887:884]},
     {slideAddressGen_slideMaskInput_hi[883:880]},
     {slideAddressGen_slideMaskInput_hi[879:876]},
     {slideAddressGen_slideMaskInput_hi[875:872]},
     {slideAddressGen_slideMaskInput_hi[871:868]},
     {slideAddressGen_slideMaskInput_hi[867:864]},
     {slideAddressGen_slideMaskInput_hi[863:860]},
     {slideAddressGen_slideMaskInput_hi[859:856]},
     {slideAddressGen_slideMaskInput_hi[855:852]},
     {slideAddressGen_slideMaskInput_hi[851:848]},
     {slideAddressGen_slideMaskInput_hi[847:844]},
     {slideAddressGen_slideMaskInput_hi[843:840]},
     {slideAddressGen_slideMaskInput_hi[839:836]},
     {slideAddressGen_slideMaskInput_hi[835:832]},
     {slideAddressGen_slideMaskInput_hi[831:828]},
     {slideAddressGen_slideMaskInput_hi[827:824]},
     {slideAddressGen_slideMaskInput_hi[823:820]},
     {slideAddressGen_slideMaskInput_hi[819:816]},
     {slideAddressGen_slideMaskInput_hi[815:812]},
     {slideAddressGen_slideMaskInput_hi[811:808]},
     {slideAddressGen_slideMaskInput_hi[807:804]},
     {slideAddressGen_slideMaskInput_hi[803:800]},
     {slideAddressGen_slideMaskInput_hi[799:796]},
     {slideAddressGen_slideMaskInput_hi[795:792]},
     {slideAddressGen_slideMaskInput_hi[791:788]},
     {slideAddressGen_slideMaskInput_hi[787:784]},
     {slideAddressGen_slideMaskInput_hi[783:780]},
     {slideAddressGen_slideMaskInput_hi[779:776]},
     {slideAddressGen_slideMaskInput_hi[775:772]},
     {slideAddressGen_slideMaskInput_hi[771:768]},
     {slideAddressGen_slideMaskInput_hi[767:764]},
     {slideAddressGen_slideMaskInput_hi[763:760]},
     {slideAddressGen_slideMaskInput_hi[759:756]},
     {slideAddressGen_slideMaskInput_hi[755:752]},
     {slideAddressGen_slideMaskInput_hi[751:748]},
     {slideAddressGen_slideMaskInput_hi[747:744]},
     {slideAddressGen_slideMaskInput_hi[743:740]},
     {slideAddressGen_slideMaskInput_hi[739:736]},
     {slideAddressGen_slideMaskInput_hi[735:732]},
     {slideAddressGen_slideMaskInput_hi[731:728]},
     {slideAddressGen_slideMaskInput_hi[727:724]},
     {slideAddressGen_slideMaskInput_hi[723:720]},
     {slideAddressGen_slideMaskInput_hi[719:716]},
     {slideAddressGen_slideMaskInput_hi[715:712]},
     {slideAddressGen_slideMaskInput_hi[711:708]},
     {slideAddressGen_slideMaskInput_hi[707:704]},
     {slideAddressGen_slideMaskInput_hi[703:700]},
     {slideAddressGen_slideMaskInput_hi[699:696]},
     {slideAddressGen_slideMaskInput_hi[695:692]},
     {slideAddressGen_slideMaskInput_hi[691:688]},
     {slideAddressGen_slideMaskInput_hi[687:684]},
     {slideAddressGen_slideMaskInput_hi[683:680]},
     {slideAddressGen_slideMaskInput_hi[679:676]},
     {slideAddressGen_slideMaskInput_hi[675:672]},
     {slideAddressGen_slideMaskInput_hi[671:668]},
     {slideAddressGen_slideMaskInput_hi[667:664]},
     {slideAddressGen_slideMaskInput_hi[663:660]},
     {slideAddressGen_slideMaskInput_hi[659:656]},
     {slideAddressGen_slideMaskInput_hi[655:652]},
     {slideAddressGen_slideMaskInput_hi[651:648]},
     {slideAddressGen_slideMaskInput_hi[647:644]},
     {slideAddressGen_slideMaskInput_hi[643:640]},
     {slideAddressGen_slideMaskInput_hi[639:636]},
     {slideAddressGen_slideMaskInput_hi[635:632]},
     {slideAddressGen_slideMaskInput_hi[631:628]},
     {slideAddressGen_slideMaskInput_hi[627:624]},
     {slideAddressGen_slideMaskInput_hi[623:620]},
     {slideAddressGen_slideMaskInput_hi[619:616]},
     {slideAddressGen_slideMaskInput_hi[615:612]},
     {slideAddressGen_slideMaskInput_hi[611:608]},
     {slideAddressGen_slideMaskInput_hi[607:604]},
     {slideAddressGen_slideMaskInput_hi[603:600]},
     {slideAddressGen_slideMaskInput_hi[599:596]},
     {slideAddressGen_slideMaskInput_hi[595:592]},
     {slideAddressGen_slideMaskInput_hi[591:588]},
     {slideAddressGen_slideMaskInput_hi[587:584]},
     {slideAddressGen_slideMaskInput_hi[583:580]},
     {slideAddressGen_slideMaskInput_hi[579:576]},
     {slideAddressGen_slideMaskInput_hi[575:572]},
     {slideAddressGen_slideMaskInput_hi[571:568]},
     {slideAddressGen_slideMaskInput_hi[567:564]},
     {slideAddressGen_slideMaskInput_hi[563:560]},
     {slideAddressGen_slideMaskInput_hi[559:556]},
     {slideAddressGen_slideMaskInput_hi[555:552]},
     {slideAddressGen_slideMaskInput_hi[551:548]},
     {slideAddressGen_slideMaskInput_hi[547:544]},
     {slideAddressGen_slideMaskInput_hi[543:540]},
     {slideAddressGen_slideMaskInput_hi[539:536]},
     {slideAddressGen_slideMaskInput_hi[535:532]},
     {slideAddressGen_slideMaskInput_hi[531:528]},
     {slideAddressGen_slideMaskInput_hi[527:524]},
     {slideAddressGen_slideMaskInput_hi[523:520]},
     {slideAddressGen_slideMaskInput_hi[519:516]},
     {slideAddressGen_slideMaskInput_hi[515:512]},
     {slideAddressGen_slideMaskInput_hi[511:508]},
     {slideAddressGen_slideMaskInput_hi[507:504]},
     {slideAddressGen_slideMaskInput_hi[503:500]},
     {slideAddressGen_slideMaskInput_hi[499:496]},
     {slideAddressGen_slideMaskInput_hi[495:492]},
     {slideAddressGen_slideMaskInput_hi[491:488]},
     {slideAddressGen_slideMaskInput_hi[487:484]},
     {slideAddressGen_slideMaskInput_hi[483:480]},
     {slideAddressGen_slideMaskInput_hi[479:476]},
     {slideAddressGen_slideMaskInput_hi[475:472]},
     {slideAddressGen_slideMaskInput_hi[471:468]},
     {slideAddressGen_slideMaskInput_hi[467:464]},
     {slideAddressGen_slideMaskInput_hi[463:460]},
     {slideAddressGen_slideMaskInput_hi[459:456]},
     {slideAddressGen_slideMaskInput_hi[455:452]},
     {slideAddressGen_slideMaskInput_hi[451:448]},
     {slideAddressGen_slideMaskInput_hi[447:444]},
     {slideAddressGen_slideMaskInput_hi[443:440]},
     {slideAddressGen_slideMaskInput_hi[439:436]},
     {slideAddressGen_slideMaskInput_hi[435:432]},
     {slideAddressGen_slideMaskInput_hi[431:428]},
     {slideAddressGen_slideMaskInput_hi[427:424]},
     {slideAddressGen_slideMaskInput_hi[423:420]},
     {slideAddressGen_slideMaskInput_hi[419:416]},
     {slideAddressGen_slideMaskInput_hi[415:412]},
     {slideAddressGen_slideMaskInput_hi[411:408]},
     {slideAddressGen_slideMaskInput_hi[407:404]},
     {slideAddressGen_slideMaskInput_hi[403:400]},
     {slideAddressGen_slideMaskInput_hi[399:396]},
     {slideAddressGen_slideMaskInput_hi[395:392]},
     {slideAddressGen_slideMaskInput_hi[391:388]},
     {slideAddressGen_slideMaskInput_hi[387:384]},
     {slideAddressGen_slideMaskInput_hi[383:380]},
     {slideAddressGen_slideMaskInput_hi[379:376]},
     {slideAddressGen_slideMaskInput_hi[375:372]},
     {slideAddressGen_slideMaskInput_hi[371:368]},
     {slideAddressGen_slideMaskInput_hi[367:364]},
     {slideAddressGen_slideMaskInput_hi[363:360]},
     {slideAddressGen_slideMaskInput_hi[359:356]},
     {slideAddressGen_slideMaskInput_hi[355:352]},
     {slideAddressGen_slideMaskInput_hi[351:348]},
     {slideAddressGen_slideMaskInput_hi[347:344]},
     {slideAddressGen_slideMaskInput_hi[343:340]},
     {slideAddressGen_slideMaskInput_hi[339:336]},
     {slideAddressGen_slideMaskInput_hi[335:332]},
     {slideAddressGen_slideMaskInput_hi[331:328]},
     {slideAddressGen_slideMaskInput_hi[327:324]},
     {slideAddressGen_slideMaskInput_hi[323:320]},
     {slideAddressGen_slideMaskInput_hi[319:316]},
     {slideAddressGen_slideMaskInput_hi[315:312]},
     {slideAddressGen_slideMaskInput_hi[311:308]},
     {slideAddressGen_slideMaskInput_hi[307:304]},
     {slideAddressGen_slideMaskInput_hi[303:300]},
     {slideAddressGen_slideMaskInput_hi[299:296]},
     {slideAddressGen_slideMaskInput_hi[295:292]},
     {slideAddressGen_slideMaskInput_hi[291:288]},
     {slideAddressGen_slideMaskInput_hi[287:284]},
     {slideAddressGen_slideMaskInput_hi[283:280]},
     {slideAddressGen_slideMaskInput_hi[279:276]},
     {slideAddressGen_slideMaskInput_hi[275:272]},
     {slideAddressGen_slideMaskInput_hi[271:268]},
     {slideAddressGen_slideMaskInput_hi[267:264]},
     {slideAddressGen_slideMaskInput_hi[263:260]},
     {slideAddressGen_slideMaskInput_hi[259:256]},
     {slideAddressGen_slideMaskInput_hi[255:252]},
     {slideAddressGen_slideMaskInput_hi[251:248]},
     {slideAddressGen_slideMaskInput_hi[247:244]},
     {slideAddressGen_slideMaskInput_hi[243:240]},
     {slideAddressGen_slideMaskInput_hi[239:236]},
     {slideAddressGen_slideMaskInput_hi[235:232]},
     {slideAddressGen_slideMaskInput_hi[231:228]},
     {slideAddressGen_slideMaskInput_hi[227:224]},
     {slideAddressGen_slideMaskInput_hi[223:220]},
     {slideAddressGen_slideMaskInput_hi[219:216]},
     {slideAddressGen_slideMaskInput_hi[215:212]},
     {slideAddressGen_slideMaskInput_hi[211:208]},
     {slideAddressGen_slideMaskInput_hi[207:204]},
     {slideAddressGen_slideMaskInput_hi[203:200]},
     {slideAddressGen_slideMaskInput_hi[199:196]},
     {slideAddressGen_slideMaskInput_hi[195:192]},
     {slideAddressGen_slideMaskInput_hi[191:188]},
     {slideAddressGen_slideMaskInput_hi[187:184]},
     {slideAddressGen_slideMaskInput_hi[183:180]},
     {slideAddressGen_slideMaskInput_hi[179:176]},
     {slideAddressGen_slideMaskInput_hi[175:172]},
     {slideAddressGen_slideMaskInput_hi[171:168]},
     {slideAddressGen_slideMaskInput_hi[167:164]},
     {slideAddressGen_slideMaskInput_hi[163:160]},
     {slideAddressGen_slideMaskInput_hi[159:156]},
     {slideAddressGen_slideMaskInput_hi[155:152]},
     {slideAddressGen_slideMaskInput_hi[151:148]},
     {slideAddressGen_slideMaskInput_hi[147:144]},
     {slideAddressGen_slideMaskInput_hi[143:140]},
     {slideAddressGen_slideMaskInput_hi[139:136]},
     {slideAddressGen_slideMaskInput_hi[135:132]},
     {slideAddressGen_slideMaskInput_hi[131:128]},
     {slideAddressGen_slideMaskInput_hi[127:124]},
     {slideAddressGen_slideMaskInput_hi[123:120]},
     {slideAddressGen_slideMaskInput_hi[119:116]},
     {slideAddressGen_slideMaskInput_hi[115:112]},
     {slideAddressGen_slideMaskInput_hi[111:108]},
     {slideAddressGen_slideMaskInput_hi[107:104]},
     {slideAddressGen_slideMaskInput_hi[103:100]},
     {slideAddressGen_slideMaskInput_hi[99:96]},
     {slideAddressGen_slideMaskInput_hi[95:92]},
     {slideAddressGen_slideMaskInput_hi[91:88]},
     {slideAddressGen_slideMaskInput_hi[87:84]},
     {slideAddressGen_slideMaskInput_hi[83:80]},
     {slideAddressGen_slideMaskInput_hi[79:76]},
     {slideAddressGen_slideMaskInput_hi[75:72]},
     {slideAddressGen_slideMaskInput_hi[71:68]},
     {slideAddressGen_slideMaskInput_hi[67:64]},
     {slideAddressGen_slideMaskInput_hi[63:60]},
     {slideAddressGen_slideMaskInput_hi[59:56]},
     {slideAddressGen_slideMaskInput_hi[55:52]},
     {slideAddressGen_slideMaskInput_hi[51:48]},
     {slideAddressGen_slideMaskInput_hi[47:44]},
     {slideAddressGen_slideMaskInput_hi[43:40]},
     {slideAddressGen_slideMaskInput_hi[39:36]},
     {slideAddressGen_slideMaskInput_hi[35:32]},
     {slideAddressGen_slideMaskInput_hi[31:28]},
     {slideAddressGen_slideMaskInput_hi[27:24]},
     {slideAddressGen_slideMaskInput_hi[23:20]},
     {slideAddressGen_slideMaskInput_hi[19:16]},
     {slideAddressGen_slideMaskInput_hi[15:12]},
     {slideAddressGen_slideMaskInput_hi[11:8]},
     {slideAddressGen_slideMaskInput_hi[7:4]},
     {slideAddressGen_slideMaskInput_hi[3:0]},
     {slideAddressGen_slideMaskInput_lo[1023:1020]},
     {slideAddressGen_slideMaskInput_lo[1019:1016]},
     {slideAddressGen_slideMaskInput_lo[1015:1012]},
     {slideAddressGen_slideMaskInput_lo[1011:1008]},
     {slideAddressGen_slideMaskInput_lo[1007:1004]},
     {slideAddressGen_slideMaskInput_lo[1003:1000]},
     {slideAddressGen_slideMaskInput_lo[999:996]},
     {slideAddressGen_slideMaskInput_lo[995:992]},
     {slideAddressGen_slideMaskInput_lo[991:988]},
     {slideAddressGen_slideMaskInput_lo[987:984]},
     {slideAddressGen_slideMaskInput_lo[983:980]},
     {slideAddressGen_slideMaskInput_lo[979:976]},
     {slideAddressGen_slideMaskInput_lo[975:972]},
     {slideAddressGen_slideMaskInput_lo[971:968]},
     {slideAddressGen_slideMaskInput_lo[967:964]},
     {slideAddressGen_slideMaskInput_lo[963:960]},
     {slideAddressGen_slideMaskInput_lo[959:956]},
     {slideAddressGen_slideMaskInput_lo[955:952]},
     {slideAddressGen_slideMaskInput_lo[951:948]},
     {slideAddressGen_slideMaskInput_lo[947:944]},
     {slideAddressGen_slideMaskInput_lo[943:940]},
     {slideAddressGen_slideMaskInput_lo[939:936]},
     {slideAddressGen_slideMaskInput_lo[935:932]},
     {slideAddressGen_slideMaskInput_lo[931:928]},
     {slideAddressGen_slideMaskInput_lo[927:924]},
     {slideAddressGen_slideMaskInput_lo[923:920]},
     {slideAddressGen_slideMaskInput_lo[919:916]},
     {slideAddressGen_slideMaskInput_lo[915:912]},
     {slideAddressGen_slideMaskInput_lo[911:908]},
     {slideAddressGen_slideMaskInput_lo[907:904]},
     {slideAddressGen_slideMaskInput_lo[903:900]},
     {slideAddressGen_slideMaskInput_lo[899:896]},
     {slideAddressGen_slideMaskInput_lo[895:892]},
     {slideAddressGen_slideMaskInput_lo[891:888]},
     {slideAddressGen_slideMaskInput_lo[887:884]},
     {slideAddressGen_slideMaskInput_lo[883:880]},
     {slideAddressGen_slideMaskInput_lo[879:876]},
     {slideAddressGen_slideMaskInput_lo[875:872]},
     {slideAddressGen_slideMaskInput_lo[871:868]},
     {slideAddressGen_slideMaskInput_lo[867:864]},
     {slideAddressGen_slideMaskInput_lo[863:860]},
     {slideAddressGen_slideMaskInput_lo[859:856]},
     {slideAddressGen_slideMaskInput_lo[855:852]},
     {slideAddressGen_slideMaskInput_lo[851:848]},
     {slideAddressGen_slideMaskInput_lo[847:844]},
     {slideAddressGen_slideMaskInput_lo[843:840]},
     {slideAddressGen_slideMaskInput_lo[839:836]},
     {slideAddressGen_slideMaskInput_lo[835:832]},
     {slideAddressGen_slideMaskInput_lo[831:828]},
     {slideAddressGen_slideMaskInput_lo[827:824]},
     {slideAddressGen_slideMaskInput_lo[823:820]},
     {slideAddressGen_slideMaskInput_lo[819:816]},
     {slideAddressGen_slideMaskInput_lo[815:812]},
     {slideAddressGen_slideMaskInput_lo[811:808]},
     {slideAddressGen_slideMaskInput_lo[807:804]},
     {slideAddressGen_slideMaskInput_lo[803:800]},
     {slideAddressGen_slideMaskInput_lo[799:796]},
     {slideAddressGen_slideMaskInput_lo[795:792]},
     {slideAddressGen_slideMaskInput_lo[791:788]},
     {slideAddressGen_slideMaskInput_lo[787:784]},
     {slideAddressGen_slideMaskInput_lo[783:780]},
     {slideAddressGen_slideMaskInput_lo[779:776]},
     {slideAddressGen_slideMaskInput_lo[775:772]},
     {slideAddressGen_slideMaskInput_lo[771:768]},
     {slideAddressGen_slideMaskInput_lo[767:764]},
     {slideAddressGen_slideMaskInput_lo[763:760]},
     {slideAddressGen_slideMaskInput_lo[759:756]},
     {slideAddressGen_slideMaskInput_lo[755:752]},
     {slideAddressGen_slideMaskInput_lo[751:748]},
     {slideAddressGen_slideMaskInput_lo[747:744]},
     {slideAddressGen_slideMaskInput_lo[743:740]},
     {slideAddressGen_slideMaskInput_lo[739:736]},
     {slideAddressGen_slideMaskInput_lo[735:732]},
     {slideAddressGen_slideMaskInput_lo[731:728]},
     {slideAddressGen_slideMaskInput_lo[727:724]},
     {slideAddressGen_slideMaskInput_lo[723:720]},
     {slideAddressGen_slideMaskInput_lo[719:716]},
     {slideAddressGen_slideMaskInput_lo[715:712]},
     {slideAddressGen_slideMaskInput_lo[711:708]},
     {slideAddressGen_slideMaskInput_lo[707:704]},
     {slideAddressGen_slideMaskInput_lo[703:700]},
     {slideAddressGen_slideMaskInput_lo[699:696]},
     {slideAddressGen_slideMaskInput_lo[695:692]},
     {slideAddressGen_slideMaskInput_lo[691:688]},
     {slideAddressGen_slideMaskInput_lo[687:684]},
     {slideAddressGen_slideMaskInput_lo[683:680]},
     {slideAddressGen_slideMaskInput_lo[679:676]},
     {slideAddressGen_slideMaskInput_lo[675:672]},
     {slideAddressGen_slideMaskInput_lo[671:668]},
     {slideAddressGen_slideMaskInput_lo[667:664]},
     {slideAddressGen_slideMaskInput_lo[663:660]},
     {slideAddressGen_slideMaskInput_lo[659:656]},
     {slideAddressGen_slideMaskInput_lo[655:652]},
     {slideAddressGen_slideMaskInput_lo[651:648]},
     {slideAddressGen_slideMaskInput_lo[647:644]},
     {slideAddressGen_slideMaskInput_lo[643:640]},
     {slideAddressGen_slideMaskInput_lo[639:636]},
     {slideAddressGen_slideMaskInput_lo[635:632]},
     {slideAddressGen_slideMaskInput_lo[631:628]},
     {slideAddressGen_slideMaskInput_lo[627:624]},
     {slideAddressGen_slideMaskInput_lo[623:620]},
     {slideAddressGen_slideMaskInput_lo[619:616]},
     {slideAddressGen_slideMaskInput_lo[615:612]},
     {slideAddressGen_slideMaskInput_lo[611:608]},
     {slideAddressGen_slideMaskInput_lo[607:604]},
     {slideAddressGen_slideMaskInput_lo[603:600]},
     {slideAddressGen_slideMaskInput_lo[599:596]},
     {slideAddressGen_slideMaskInput_lo[595:592]},
     {slideAddressGen_slideMaskInput_lo[591:588]},
     {slideAddressGen_slideMaskInput_lo[587:584]},
     {slideAddressGen_slideMaskInput_lo[583:580]},
     {slideAddressGen_slideMaskInput_lo[579:576]},
     {slideAddressGen_slideMaskInput_lo[575:572]},
     {slideAddressGen_slideMaskInput_lo[571:568]},
     {slideAddressGen_slideMaskInput_lo[567:564]},
     {slideAddressGen_slideMaskInput_lo[563:560]},
     {slideAddressGen_slideMaskInput_lo[559:556]},
     {slideAddressGen_slideMaskInput_lo[555:552]},
     {slideAddressGen_slideMaskInput_lo[551:548]},
     {slideAddressGen_slideMaskInput_lo[547:544]},
     {slideAddressGen_slideMaskInput_lo[543:540]},
     {slideAddressGen_slideMaskInput_lo[539:536]},
     {slideAddressGen_slideMaskInput_lo[535:532]},
     {slideAddressGen_slideMaskInput_lo[531:528]},
     {slideAddressGen_slideMaskInput_lo[527:524]},
     {slideAddressGen_slideMaskInput_lo[523:520]},
     {slideAddressGen_slideMaskInput_lo[519:516]},
     {slideAddressGen_slideMaskInput_lo[515:512]},
     {slideAddressGen_slideMaskInput_lo[511:508]},
     {slideAddressGen_slideMaskInput_lo[507:504]},
     {slideAddressGen_slideMaskInput_lo[503:500]},
     {slideAddressGen_slideMaskInput_lo[499:496]},
     {slideAddressGen_slideMaskInput_lo[495:492]},
     {slideAddressGen_slideMaskInput_lo[491:488]},
     {slideAddressGen_slideMaskInput_lo[487:484]},
     {slideAddressGen_slideMaskInput_lo[483:480]},
     {slideAddressGen_slideMaskInput_lo[479:476]},
     {slideAddressGen_slideMaskInput_lo[475:472]},
     {slideAddressGen_slideMaskInput_lo[471:468]},
     {slideAddressGen_slideMaskInput_lo[467:464]},
     {slideAddressGen_slideMaskInput_lo[463:460]},
     {slideAddressGen_slideMaskInput_lo[459:456]},
     {slideAddressGen_slideMaskInput_lo[455:452]},
     {slideAddressGen_slideMaskInput_lo[451:448]},
     {slideAddressGen_slideMaskInput_lo[447:444]},
     {slideAddressGen_slideMaskInput_lo[443:440]},
     {slideAddressGen_slideMaskInput_lo[439:436]},
     {slideAddressGen_slideMaskInput_lo[435:432]},
     {slideAddressGen_slideMaskInput_lo[431:428]},
     {slideAddressGen_slideMaskInput_lo[427:424]},
     {slideAddressGen_slideMaskInput_lo[423:420]},
     {slideAddressGen_slideMaskInput_lo[419:416]},
     {slideAddressGen_slideMaskInput_lo[415:412]},
     {slideAddressGen_slideMaskInput_lo[411:408]},
     {slideAddressGen_slideMaskInput_lo[407:404]},
     {slideAddressGen_slideMaskInput_lo[403:400]},
     {slideAddressGen_slideMaskInput_lo[399:396]},
     {slideAddressGen_slideMaskInput_lo[395:392]},
     {slideAddressGen_slideMaskInput_lo[391:388]},
     {slideAddressGen_slideMaskInput_lo[387:384]},
     {slideAddressGen_slideMaskInput_lo[383:380]},
     {slideAddressGen_slideMaskInput_lo[379:376]},
     {slideAddressGen_slideMaskInput_lo[375:372]},
     {slideAddressGen_slideMaskInput_lo[371:368]},
     {slideAddressGen_slideMaskInput_lo[367:364]},
     {slideAddressGen_slideMaskInput_lo[363:360]},
     {slideAddressGen_slideMaskInput_lo[359:356]},
     {slideAddressGen_slideMaskInput_lo[355:352]},
     {slideAddressGen_slideMaskInput_lo[351:348]},
     {slideAddressGen_slideMaskInput_lo[347:344]},
     {slideAddressGen_slideMaskInput_lo[343:340]},
     {slideAddressGen_slideMaskInput_lo[339:336]},
     {slideAddressGen_slideMaskInput_lo[335:332]},
     {slideAddressGen_slideMaskInput_lo[331:328]},
     {slideAddressGen_slideMaskInput_lo[327:324]},
     {slideAddressGen_slideMaskInput_lo[323:320]},
     {slideAddressGen_slideMaskInput_lo[319:316]},
     {slideAddressGen_slideMaskInput_lo[315:312]},
     {slideAddressGen_slideMaskInput_lo[311:308]},
     {slideAddressGen_slideMaskInput_lo[307:304]},
     {slideAddressGen_slideMaskInput_lo[303:300]},
     {slideAddressGen_slideMaskInput_lo[299:296]},
     {slideAddressGen_slideMaskInput_lo[295:292]},
     {slideAddressGen_slideMaskInput_lo[291:288]},
     {slideAddressGen_slideMaskInput_lo[287:284]},
     {slideAddressGen_slideMaskInput_lo[283:280]},
     {slideAddressGen_slideMaskInput_lo[279:276]},
     {slideAddressGen_slideMaskInput_lo[275:272]},
     {slideAddressGen_slideMaskInput_lo[271:268]},
     {slideAddressGen_slideMaskInput_lo[267:264]},
     {slideAddressGen_slideMaskInput_lo[263:260]},
     {slideAddressGen_slideMaskInput_lo[259:256]},
     {slideAddressGen_slideMaskInput_lo[255:252]},
     {slideAddressGen_slideMaskInput_lo[251:248]},
     {slideAddressGen_slideMaskInput_lo[247:244]},
     {slideAddressGen_slideMaskInput_lo[243:240]},
     {slideAddressGen_slideMaskInput_lo[239:236]},
     {slideAddressGen_slideMaskInput_lo[235:232]},
     {slideAddressGen_slideMaskInput_lo[231:228]},
     {slideAddressGen_slideMaskInput_lo[227:224]},
     {slideAddressGen_slideMaskInput_lo[223:220]},
     {slideAddressGen_slideMaskInput_lo[219:216]},
     {slideAddressGen_slideMaskInput_lo[215:212]},
     {slideAddressGen_slideMaskInput_lo[211:208]},
     {slideAddressGen_slideMaskInput_lo[207:204]},
     {slideAddressGen_slideMaskInput_lo[203:200]},
     {slideAddressGen_slideMaskInput_lo[199:196]},
     {slideAddressGen_slideMaskInput_lo[195:192]},
     {slideAddressGen_slideMaskInput_lo[191:188]},
     {slideAddressGen_slideMaskInput_lo[187:184]},
     {slideAddressGen_slideMaskInput_lo[183:180]},
     {slideAddressGen_slideMaskInput_lo[179:176]},
     {slideAddressGen_slideMaskInput_lo[175:172]},
     {slideAddressGen_slideMaskInput_lo[171:168]},
     {slideAddressGen_slideMaskInput_lo[167:164]},
     {slideAddressGen_slideMaskInput_lo[163:160]},
     {slideAddressGen_slideMaskInput_lo[159:156]},
     {slideAddressGen_slideMaskInput_lo[155:152]},
     {slideAddressGen_slideMaskInput_lo[151:148]},
     {slideAddressGen_slideMaskInput_lo[147:144]},
     {slideAddressGen_slideMaskInput_lo[143:140]},
     {slideAddressGen_slideMaskInput_lo[139:136]},
     {slideAddressGen_slideMaskInput_lo[135:132]},
     {slideAddressGen_slideMaskInput_lo[131:128]},
     {slideAddressGen_slideMaskInput_lo[127:124]},
     {slideAddressGen_slideMaskInput_lo[123:120]},
     {slideAddressGen_slideMaskInput_lo[119:116]},
     {slideAddressGen_slideMaskInput_lo[115:112]},
     {slideAddressGen_slideMaskInput_lo[111:108]},
     {slideAddressGen_slideMaskInput_lo[107:104]},
     {slideAddressGen_slideMaskInput_lo[103:100]},
     {slideAddressGen_slideMaskInput_lo[99:96]},
     {slideAddressGen_slideMaskInput_lo[95:92]},
     {slideAddressGen_slideMaskInput_lo[91:88]},
     {slideAddressGen_slideMaskInput_lo[87:84]},
     {slideAddressGen_slideMaskInput_lo[83:80]},
     {slideAddressGen_slideMaskInput_lo[79:76]},
     {slideAddressGen_slideMaskInput_lo[75:72]},
     {slideAddressGen_slideMaskInput_lo[71:68]},
     {slideAddressGen_slideMaskInput_lo[67:64]},
     {slideAddressGen_slideMaskInput_lo[63:60]},
     {slideAddressGen_slideMaskInput_lo[59:56]},
     {slideAddressGen_slideMaskInput_lo[55:52]},
     {slideAddressGen_slideMaskInput_lo[51:48]},
     {slideAddressGen_slideMaskInput_lo[47:44]},
     {slideAddressGen_slideMaskInput_lo[43:40]},
     {slideAddressGen_slideMaskInput_lo[39:36]},
     {slideAddressGen_slideMaskInput_lo[35:32]},
     {slideAddressGen_slideMaskInput_lo[31:28]},
     {slideAddressGen_slideMaskInput_lo[27:24]},
     {slideAddressGen_slideMaskInput_lo[23:20]},
     {slideAddressGen_slideMaskInput_lo[19:16]},
     {slideAddressGen_slideMaskInput_lo[15:12]},
     {slideAddressGen_slideMaskInput_lo[11:8]},
     {slideAddressGen_slideMaskInput_lo[7:4]},
     {slideAddressGen_slideMaskInput_lo[3:0]}};
  wire               lastExecuteGroupDeq;
  wire               viotaCounterAdd;
  wire               groupCounterAdd = noSource ? viotaCounterAdd : lastExecuteGroupDeq;
  wire [3:0]         groupDataNeed = lastGroup ? lastGroupDataNeed : 4'hF;
  reg  [1:0]         executeIndex;
  reg  [3:0]         readIssueStageState_groupReadState;
  reg  [3:0]         readIssueStageState_needRead;
  wire [3:0]         readWaitQueue_enq_bits_needRead = readIssueStageState_needRead;
  reg  [3:0]         readIssueStageState_elementValid;
  wire [3:0]         readWaitQueue_enq_bits_sourceValid = readIssueStageState_elementValid;
  reg  [3:0]         readIssueStageState_replaceVs1;
  wire [3:0]         readWaitQueue_enq_bits_replaceVs1 = readIssueStageState_replaceVs1;
  reg  [15:0]        readIssueStageState_readOffset;
  reg  [1:0]         readIssueStageState_accessLane_0;
  reg  [1:0]         readIssueStageState_accessLane_1;
  wire [1:0]         selectExecuteReq_1_bits_readLane = readIssueStageState_accessLane_1;
  reg  [1:0]         readIssueStageState_accessLane_2;
  wire [1:0]         selectExecuteReq_2_bits_readLane = readIssueStageState_accessLane_2;
  reg  [1:0]         readIssueStageState_accessLane_3;
  wire [1:0]         selectExecuteReq_3_bits_readLane = readIssueStageState_accessLane_3;
  reg  [2:0]         readIssueStageState_vsGrowth_0;
  reg  [2:0]         readIssueStageState_vsGrowth_1;
  reg  [2:0]         readIssueStageState_vsGrowth_2;
  reg  [2:0]         readIssueStageState_vsGrowth_3;
  reg  [9:0]         readIssueStageState_executeGroup;
  wire [9:0]         readWaitQueue_enq_bits_executeGroup = readIssueStageState_executeGroup;
  reg  [7:0]         readIssueStageState_readDataOffset;
  reg                readIssueStageState_last;
  wire               readWaitQueue_enq_bits_last = readIssueStageState_last;
  reg                readIssueStageValid;
  wire [2:0]         accessCountQueue_enq_bits_0 = accessCountEnq_0;
  wire [2:0]         accessCountQueue_enq_bits_1 = accessCountEnq_1;
  wire [2:0]         accessCountQueue_enq_bits_2 = accessCountEnq_2;
  wire [2:0]         accessCountQueue_enq_bits_3 = accessCountEnq_3;
  wire               readIssueStageEnq;
  wire               accessCountQueue_deq_valid;
  assign accessCountQueue_deq_valid = ~_accessCountQueue_fifo_empty;
  wire [2:0]         accessCountQueue_dataOut_0;
  wire [2:0]         accessCountQueue_dataOut_1;
  wire [2:0]         accessCountQueue_dataOut_2;
  wire [2:0]         accessCountQueue_dataOut_3;
  wire [5:0]         accessCountQueue_dataIn_lo = {accessCountQueue_enq_bits_1, accessCountQueue_enq_bits_0};
  wire [5:0]         accessCountQueue_dataIn_hi = {accessCountQueue_enq_bits_3, accessCountQueue_enq_bits_2};
  wire [11:0]        accessCountQueue_dataIn = {accessCountQueue_dataIn_hi, accessCountQueue_dataIn_lo};
  assign accessCountQueue_dataOut_0 = _accessCountQueue_fifo_data_out[2:0];
  assign accessCountQueue_dataOut_1 = _accessCountQueue_fifo_data_out[5:3];
  assign accessCountQueue_dataOut_2 = _accessCountQueue_fifo_data_out[8:6];
  assign accessCountQueue_dataOut_3 = _accessCountQueue_fifo_data_out[11:9];
  wire [2:0]         accessCountQueue_deq_bits_0 = accessCountQueue_dataOut_0;
  wire [2:0]         accessCountQueue_deq_bits_1 = accessCountQueue_dataOut_1;
  wire [2:0]         accessCountQueue_deq_bits_2 = accessCountQueue_dataOut_2;
  wire [2:0]         accessCountQueue_deq_bits_3 = accessCountQueue_dataOut_3;
  wire               accessCountQueue_enq_ready = ~_accessCountQueue_fifo_full;
  wire               accessCountQueue_enq_valid;
  wire               accessCountQueue_deq_ready;
  wire [9:0]         _extendGroupCount_T_1 = {requestCounter, executeIndex};
  wire [9:0]         _executeGroup_T_8 = executeIndexGrowth[0] ? _extendGroupCount_T_1 : 10'h0;
  wire [8:0]         _GEN_45 = _executeGroup_T_8[8:0] | (executeIndexGrowth[1] ? {requestCounter, executeIndex[1]} : 9'h0);
  wire [9:0]         executeGroup = {_executeGroup_T_8[9], _GEN_45[8], _GEN_45[7:0] | (executeIndexGrowth[2] ? requestCounter : 8'h0)};
  wire               vlMisAlign;
  assign vlMisAlign = |(instReg_vl[1:0]);
  wire [9:0]         lastexecuteGroup = instReg_vl[11:2] - {9'h0, ~vlMisAlign};
  wire               isVlBoundary = executeGroup == lastexecuteGroup;
  wire               validExecuteGroup = executeGroup <= lastexecuteGroup;
  wire [3:0]         _maskSplit_vlBoundaryCorrection_T_37 = 4'h1 << instReg_vl[1:0];
  wire [3:0]         _vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_37 | {_maskSplit_vlBoundaryCorrection_T_37[2:0], 1'h0};
  wire [3:0]         vlBoundaryCorrection = ~({4{vlMisAlign & isVlBoundary}} & (_vlBoundaryCorrection_T_5 | {_vlBoundaryCorrection_T_5[1:0], 2'h0})) & {4{validExecuteGroup}};
  wire [127:0]       selectReadStageMask_lo_lo_lo_lo = {selectReadStageMask_lo_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_lo_hi = {selectReadStageMask_lo_lo_lo_hi_hi, selectReadStageMask_lo_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_lo = {selectReadStageMask_lo_lo_lo_hi, selectReadStageMask_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_lo = {selectReadStageMask_lo_lo_hi_lo_hi, selectReadStageMask_lo_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_lo_hi_hi = {selectReadStageMask_lo_lo_hi_hi_hi, selectReadStageMask_lo_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_lo_hi = {selectReadStageMask_lo_lo_hi_hi, selectReadStageMask_lo_lo_hi_lo};
  wire [511:0]       selectReadStageMask_lo_lo = {selectReadStageMask_lo_lo_hi, selectReadStageMask_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_lo = {selectReadStageMask_lo_hi_lo_lo_hi, selectReadStageMask_lo_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_lo_hi = {selectReadStageMask_lo_hi_lo_hi_hi, selectReadStageMask_lo_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_lo = {selectReadStageMask_lo_hi_lo_hi, selectReadStageMask_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_lo = {selectReadStageMask_lo_hi_hi_lo_hi, selectReadStageMask_lo_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_lo_hi_hi_hi = {selectReadStageMask_lo_hi_hi_hi_hi, selectReadStageMask_lo_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_lo_hi_hi = {selectReadStageMask_lo_hi_hi_hi, selectReadStageMask_lo_hi_hi_lo};
  wire [511:0]       selectReadStageMask_lo_hi = {selectReadStageMask_lo_hi_hi, selectReadStageMask_lo_hi_lo};
  wire [1023:0]      selectReadStageMask_lo = {selectReadStageMask_lo_hi, selectReadStageMask_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_lo = {selectReadStageMask_hi_lo_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_lo_hi = {selectReadStageMask_hi_lo_lo_hi_hi, selectReadStageMask_hi_lo_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_lo = {selectReadStageMask_hi_lo_lo_hi, selectReadStageMask_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_lo = {selectReadStageMask_hi_lo_hi_lo_hi, selectReadStageMask_hi_lo_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_lo_hi_hi = {selectReadStageMask_hi_lo_hi_hi_hi, selectReadStageMask_hi_lo_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_lo_hi = {selectReadStageMask_hi_lo_hi_hi, selectReadStageMask_hi_lo_hi_lo};
  wire [511:0]       selectReadStageMask_hi_lo = {selectReadStageMask_hi_lo_hi, selectReadStageMask_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_lo = {selectReadStageMask_hi_hi_lo_lo_hi, selectReadStageMask_hi_hi_lo_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_lo_hi = {selectReadStageMask_hi_hi_lo_hi_hi, selectReadStageMask_hi_hi_lo_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_lo = {selectReadStageMask_hi_hi_lo_hi, selectReadStageMask_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_lo = {selectReadStageMask_hi_hi_hi_lo_hi, selectReadStageMask_hi_hi_hi_lo_lo};
  wire [127:0]       selectReadStageMask_hi_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_hi_lo};
  wire [255:0]       selectReadStageMask_hi_hi_hi = {selectReadStageMask_hi_hi_hi_hi, selectReadStageMask_hi_hi_hi_lo};
  wire [511:0]       selectReadStageMask_hi_hi = {selectReadStageMask_hi_hi_hi, selectReadStageMask_hi_hi_lo};
  wire [1023:0]      selectReadStageMask_hi = {selectReadStageMask_hi_hi, selectReadStageMask_hi_lo};
  wire [511:0][3:0]  _GEN_46 =
    {{selectReadStageMask_hi[1023:1020]},
     {selectReadStageMask_hi[1019:1016]},
     {selectReadStageMask_hi[1015:1012]},
     {selectReadStageMask_hi[1011:1008]},
     {selectReadStageMask_hi[1007:1004]},
     {selectReadStageMask_hi[1003:1000]},
     {selectReadStageMask_hi[999:996]},
     {selectReadStageMask_hi[995:992]},
     {selectReadStageMask_hi[991:988]},
     {selectReadStageMask_hi[987:984]},
     {selectReadStageMask_hi[983:980]},
     {selectReadStageMask_hi[979:976]},
     {selectReadStageMask_hi[975:972]},
     {selectReadStageMask_hi[971:968]},
     {selectReadStageMask_hi[967:964]},
     {selectReadStageMask_hi[963:960]},
     {selectReadStageMask_hi[959:956]},
     {selectReadStageMask_hi[955:952]},
     {selectReadStageMask_hi[951:948]},
     {selectReadStageMask_hi[947:944]},
     {selectReadStageMask_hi[943:940]},
     {selectReadStageMask_hi[939:936]},
     {selectReadStageMask_hi[935:932]},
     {selectReadStageMask_hi[931:928]},
     {selectReadStageMask_hi[927:924]},
     {selectReadStageMask_hi[923:920]},
     {selectReadStageMask_hi[919:916]},
     {selectReadStageMask_hi[915:912]},
     {selectReadStageMask_hi[911:908]},
     {selectReadStageMask_hi[907:904]},
     {selectReadStageMask_hi[903:900]},
     {selectReadStageMask_hi[899:896]},
     {selectReadStageMask_hi[895:892]},
     {selectReadStageMask_hi[891:888]},
     {selectReadStageMask_hi[887:884]},
     {selectReadStageMask_hi[883:880]},
     {selectReadStageMask_hi[879:876]},
     {selectReadStageMask_hi[875:872]},
     {selectReadStageMask_hi[871:868]},
     {selectReadStageMask_hi[867:864]},
     {selectReadStageMask_hi[863:860]},
     {selectReadStageMask_hi[859:856]},
     {selectReadStageMask_hi[855:852]},
     {selectReadStageMask_hi[851:848]},
     {selectReadStageMask_hi[847:844]},
     {selectReadStageMask_hi[843:840]},
     {selectReadStageMask_hi[839:836]},
     {selectReadStageMask_hi[835:832]},
     {selectReadStageMask_hi[831:828]},
     {selectReadStageMask_hi[827:824]},
     {selectReadStageMask_hi[823:820]},
     {selectReadStageMask_hi[819:816]},
     {selectReadStageMask_hi[815:812]},
     {selectReadStageMask_hi[811:808]},
     {selectReadStageMask_hi[807:804]},
     {selectReadStageMask_hi[803:800]},
     {selectReadStageMask_hi[799:796]},
     {selectReadStageMask_hi[795:792]},
     {selectReadStageMask_hi[791:788]},
     {selectReadStageMask_hi[787:784]},
     {selectReadStageMask_hi[783:780]},
     {selectReadStageMask_hi[779:776]},
     {selectReadStageMask_hi[775:772]},
     {selectReadStageMask_hi[771:768]},
     {selectReadStageMask_hi[767:764]},
     {selectReadStageMask_hi[763:760]},
     {selectReadStageMask_hi[759:756]},
     {selectReadStageMask_hi[755:752]},
     {selectReadStageMask_hi[751:748]},
     {selectReadStageMask_hi[747:744]},
     {selectReadStageMask_hi[743:740]},
     {selectReadStageMask_hi[739:736]},
     {selectReadStageMask_hi[735:732]},
     {selectReadStageMask_hi[731:728]},
     {selectReadStageMask_hi[727:724]},
     {selectReadStageMask_hi[723:720]},
     {selectReadStageMask_hi[719:716]},
     {selectReadStageMask_hi[715:712]},
     {selectReadStageMask_hi[711:708]},
     {selectReadStageMask_hi[707:704]},
     {selectReadStageMask_hi[703:700]},
     {selectReadStageMask_hi[699:696]},
     {selectReadStageMask_hi[695:692]},
     {selectReadStageMask_hi[691:688]},
     {selectReadStageMask_hi[687:684]},
     {selectReadStageMask_hi[683:680]},
     {selectReadStageMask_hi[679:676]},
     {selectReadStageMask_hi[675:672]},
     {selectReadStageMask_hi[671:668]},
     {selectReadStageMask_hi[667:664]},
     {selectReadStageMask_hi[663:660]},
     {selectReadStageMask_hi[659:656]},
     {selectReadStageMask_hi[655:652]},
     {selectReadStageMask_hi[651:648]},
     {selectReadStageMask_hi[647:644]},
     {selectReadStageMask_hi[643:640]},
     {selectReadStageMask_hi[639:636]},
     {selectReadStageMask_hi[635:632]},
     {selectReadStageMask_hi[631:628]},
     {selectReadStageMask_hi[627:624]},
     {selectReadStageMask_hi[623:620]},
     {selectReadStageMask_hi[619:616]},
     {selectReadStageMask_hi[615:612]},
     {selectReadStageMask_hi[611:608]},
     {selectReadStageMask_hi[607:604]},
     {selectReadStageMask_hi[603:600]},
     {selectReadStageMask_hi[599:596]},
     {selectReadStageMask_hi[595:592]},
     {selectReadStageMask_hi[591:588]},
     {selectReadStageMask_hi[587:584]},
     {selectReadStageMask_hi[583:580]},
     {selectReadStageMask_hi[579:576]},
     {selectReadStageMask_hi[575:572]},
     {selectReadStageMask_hi[571:568]},
     {selectReadStageMask_hi[567:564]},
     {selectReadStageMask_hi[563:560]},
     {selectReadStageMask_hi[559:556]},
     {selectReadStageMask_hi[555:552]},
     {selectReadStageMask_hi[551:548]},
     {selectReadStageMask_hi[547:544]},
     {selectReadStageMask_hi[543:540]},
     {selectReadStageMask_hi[539:536]},
     {selectReadStageMask_hi[535:532]},
     {selectReadStageMask_hi[531:528]},
     {selectReadStageMask_hi[527:524]},
     {selectReadStageMask_hi[523:520]},
     {selectReadStageMask_hi[519:516]},
     {selectReadStageMask_hi[515:512]},
     {selectReadStageMask_hi[511:508]},
     {selectReadStageMask_hi[507:504]},
     {selectReadStageMask_hi[503:500]},
     {selectReadStageMask_hi[499:496]},
     {selectReadStageMask_hi[495:492]},
     {selectReadStageMask_hi[491:488]},
     {selectReadStageMask_hi[487:484]},
     {selectReadStageMask_hi[483:480]},
     {selectReadStageMask_hi[479:476]},
     {selectReadStageMask_hi[475:472]},
     {selectReadStageMask_hi[471:468]},
     {selectReadStageMask_hi[467:464]},
     {selectReadStageMask_hi[463:460]},
     {selectReadStageMask_hi[459:456]},
     {selectReadStageMask_hi[455:452]},
     {selectReadStageMask_hi[451:448]},
     {selectReadStageMask_hi[447:444]},
     {selectReadStageMask_hi[443:440]},
     {selectReadStageMask_hi[439:436]},
     {selectReadStageMask_hi[435:432]},
     {selectReadStageMask_hi[431:428]},
     {selectReadStageMask_hi[427:424]},
     {selectReadStageMask_hi[423:420]},
     {selectReadStageMask_hi[419:416]},
     {selectReadStageMask_hi[415:412]},
     {selectReadStageMask_hi[411:408]},
     {selectReadStageMask_hi[407:404]},
     {selectReadStageMask_hi[403:400]},
     {selectReadStageMask_hi[399:396]},
     {selectReadStageMask_hi[395:392]},
     {selectReadStageMask_hi[391:388]},
     {selectReadStageMask_hi[387:384]},
     {selectReadStageMask_hi[383:380]},
     {selectReadStageMask_hi[379:376]},
     {selectReadStageMask_hi[375:372]},
     {selectReadStageMask_hi[371:368]},
     {selectReadStageMask_hi[367:364]},
     {selectReadStageMask_hi[363:360]},
     {selectReadStageMask_hi[359:356]},
     {selectReadStageMask_hi[355:352]},
     {selectReadStageMask_hi[351:348]},
     {selectReadStageMask_hi[347:344]},
     {selectReadStageMask_hi[343:340]},
     {selectReadStageMask_hi[339:336]},
     {selectReadStageMask_hi[335:332]},
     {selectReadStageMask_hi[331:328]},
     {selectReadStageMask_hi[327:324]},
     {selectReadStageMask_hi[323:320]},
     {selectReadStageMask_hi[319:316]},
     {selectReadStageMask_hi[315:312]},
     {selectReadStageMask_hi[311:308]},
     {selectReadStageMask_hi[307:304]},
     {selectReadStageMask_hi[303:300]},
     {selectReadStageMask_hi[299:296]},
     {selectReadStageMask_hi[295:292]},
     {selectReadStageMask_hi[291:288]},
     {selectReadStageMask_hi[287:284]},
     {selectReadStageMask_hi[283:280]},
     {selectReadStageMask_hi[279:276]},
     {selectReadStageMask_hi[275:272]},
     {selectReadStageMask_hi[271:268]},
     {selectReadStageMask_hi[267:264]},
     {selectReadStageMask_hi[263:260]},
     {selectReadStageMask_hi[259:256]},
     {selectReadStageMask_hi[255:252]},
     {selectReadStageMask_hi[251:248]},
     {selectReadStageMask_hi[247:244]},
     {selectReadStageMask_hi[243:240]},
     {selectReadStageMask_hi[239:236]},
     {selectReadStageMask_hi[235:232]},
     {selectReadStageMask_hi[231:228]},
     {selectReadStageMask_hi[227:224]},
     {selectReadStageMask_hi[223:220]},
     {selectReadStageMask_hi[219:216]},
     {selectReadStageMask_hi[215:212]},
     {selectReadStageMask_hi[211:208]},
     {selectReadStageMask_hi[207:204]},
     {selectReadStageMask_hi[203:200]},
     {selectReadStageMask_hi[199:196]},
     {selectReadStageMask_hi[195:192]},
     {selectReadStageMask_hi[191:188]},
     {selectReadStageMask_hi[187:184]},
     {selectReadStageMask_hi[183:180]},
     {selectReadStageMask_hi[179:176]},
     {selectReadStageMask_hi[175:172]},
     {selectReadStageMask_hi[171:168]},
     {selectReadStageMask_hi[167:164]},
     {selectReadStageMask_hi[163:160]},
     {selectReadStageMask_hi[159:156]},
     {selectReadStageMask_hi[155:152]},
     {selectReadStageMask_hi[151:148]},
     {selectReadStageMask_hi[147:144]},
     {selectReadStageMask_hi[143:140]},
     {selectReadStageMask_hi[139:136]},
     {selectReadStageMask_hi[135:132]},
     {selectReadStageMask_hi[131:128]},
     {selectReadStageMask_hi[127:124]},
     {selectReadStageMask_hi[123:120]},
     {selectReadStageMask_hi[119:116]},
     {selectReadStageMask_hi[115:112]},
     {selectReadStageMask_hi[111:108]},
     {selectReadStageMask_hi[107:104]},
     {selectReadStageMask_hi[103:100]},
     {selectReadStageMask_hi[99:96]},
     {selectReadStageMask_hi[95:92]},
     {selectReadStageMask_hi[91:88]},
     {selectReadStageMask_hi[87:84]},
     {selectReadStageMask_hi[83:80]},
     {selectReadStageMask_hi[79:76]},
     {selectReadStageMask_hi[75:72]},
     {selectReadStageMask_hi[71:68]},
     {selectReadStageMask_hi[67:64]},
     {selectReadStageMask_hi[63:60]},
     {selectReadStageMask_hi[59:56]},
     {selectReadStageMask_hi[55:52]},
     {selectReadStageMask_hi[51:48]},
     {selectReadStageMask_hi[47:44]},
     {selectReadStageMask_hi[43:40]},
     {selectReadStageMask_hi[39:36]},
     {selectReadStageMask_hi[35:32]},
     {selectReadStageMask_hi[31:28]},
     {selectReadStageMask_hi[27:24]},
     {selectReadStageMask_hi[23:20]},
     {selectReadStageMask_hi[19:16]},
     {selectReadStageMask_hi[15:12]},
     {selectReadStageMask_hi[11:8]},
     {selectReadStageMask_hi[7:4]},
     {selectReadStageMask_hi[3:0]},
     {selectReadStageMask_lo[1023:1020]},
     {selectReadStageMask_lo[1019:1016]},
     {selectReadStageMask_lo[1015:1012]},
     {selectReadStageMask_lo[1011:1008]},
     {selectReadStageMask_lo[1007:1004]},
     {selectReadStageMask_lo[1003:1000]},
     {selectReadStageMask_lo[999:996]},
     {selectReadStageMask_lo[995:992]},
     {selectReadStageMask_lo[991:988]},
     {selectReadStageMask_lo[987:984]},
     {selectReadStageMask_lo[983:980]},
     {selectReadStageMask_lo[979:976]},
     {selectReadStageMask_lo[975:972]},
     {selectReadStageMask_lo[971:968]},
     {selectReadStageMask_lo[967:964]},
     {selectReadStageMask_lo[963:960]},
     {selectReadStageMask_lo[959:956]},
     {selectReadStageMask_lo[955:952]},
     {selectReadStageMask_lo[951:948]},
     {selectReadStageMask_lo[947:944]},
     {selectReadStageMask_lo[943:940]},
     {selectReadStageMask_lo[939:936]},
     {selectReadStageMask_lo[935:932]},
     {selectReadStageMask_lo[931:928]},
     {selectReadStageMask_lo[927:924]},
     {selectReadStageMask_lo[923:920]},
     {selectReadStageMask_lo[919:916]},
     {selectReadStageMask_lo[915:912]},
     {selectReadStageMask_lo[911:908]},
     {selectReadStageMask_lo[907:904]},
     {selectReadStageMask_lo[903:900]},
     {selectReadStageMask_lo[899:896]},
     {selectReadStageMask_lo[895:892]},
     {selectReadStageMask_lo[891:888]},
     {selectReadStageMask_lo[887:884]},
     {selectReadStageMask_lo[883:880]},
     {selectReadStageMask_lo[879:876]},
     {selectReadStageMask_lo[875:872]},
     {selectReadStageMask_lo[871:868]},
     {selectReadStageMask_lo[867:864]},
     {selectReadStageMask_lo[863:860]},
     {selectReadStageMask_lo[859:856]},
     {selectReadStageMask_lo[855:852]},
     {selectReadStageMask_lo[851:848]},
     {selectReadStageMask_lo[847:844]},
     {selectReadStageMask_lo[843:840]},
     {selectReadStageMask_lo[839:836]},
     {selectReadStageMask_lo[835:832]},
     {selectReadStageMask_lo[831:828]},
     {selectReadStageMask_lo[827:824]},
     {selectReadStageMask_lo[823:820]},
     {selectReadStageMask_lo[819:816]},
     {selectReadStageMask_lo[815:812]},
     {selectReadStageMask_lo[811:808]},
     {selectReadStageMask_lo[807:804]},
     {selectReadStageMask_lo[803:800]},
     {selectReadStageMask_lo[799:796]},
     {selectReadStageMask_lo[795:792]},
     {selectReadStageMask_lo[791:788]},
     {selectReadStageMask_lo[787:784]},
     {selectReadStageMask_lo[783:780]},
     {selectReadStageMask_lo[779:776]},
     {selectReadStageMask_lo[775:772]},
     {selectReadStageMask_lo[771:768]},
     {selectReadStageMask_lo[767:764]},
     {selectReadStageMask_lo[763:760]},
     {selectReadStageMask_lo[759:756]},
     {selectReadStageMask_lo[755:752]},
     {selectReadStageMask_lo[751:748]},
     {selectReadStageMask_lo[747:744]},
     {selectReadStageMask_lo[743:740]},
     {selectReadStageMask_lo[739:736]},
     {selectReadStageMask_lo[735:732]},
     {selectReadStageMask_lo[731:728]},
     {selectReadStageMask_lo[727:724]},
     {selectReadStageMask_lo[723:720]},
     {selectReadStageMask_lo[719:716]},
     {selectReadStageMask_lo[715:712]},
     {selectReadStageMask_lo[711:708]},
     {selectReadStageMask_lo[707:704]},
     {selectReadStageMask_lo[703:700]},
     {selectReadStageMask_lo[699:696]},
     {selectReadStageMask_lo[695:692]},
     {selectReadStageMask_lo[691:688]},
     {selectReadStageMask_lo[687:684]},
     {selectReadStageMask_lo[683:680]},
     {selectReadStageMask_lo[679:676]},
     {selectReadStageMask_lo[675:672]},
     {selectReadStageMask_lo[671:668]},
     {selectReadStageMask_lo[667:664]},
     {selectReadStageMask_lo[663:660]},
     {selectReadStageMask_lo[659:656]},
     {selectReadStageMask_lo[655:652]},
     {selectReadStageMask_lo[651:648]},
     {selectReadStageMask_lo[647:644]},
     {selectReadStageMask_lo[643:640]},
     {selectReadStageMask_lo[639:636]},
     {selectReadStageMask_lo[635:632]},
     {selectReadStageMask_lo[631:628]},
     {selectReadStageMask_lo[627:624]},
     {selectReadStageMask_lo[623:620]},
     {selectReadStageMask_lo[619:616]},
     {selectReadStageMask_lo[615:612]},
     {selectReadStageMask_lo[611:608]},
     {selectReadStageMask_lo[607:604]},
     {selectReadStageMask_lo[603:600]},
     {selectReadStageMask_lo[599:596]},
     {selectReadStageMask_lo[595:592]},
     {selectReadStageMask_lo[591:588]},
     {selectReadStageMask_lo[587:584]},
     {selectReadStageMask_lo[583:580]},
     {selectReadStageMask_lo[579:576]},
     {selectReadStageMask_lo[575:572]},
     {selectReadStageMask_lo[571:568]},
     {selectReadStageMask_lo[567:564]},
     {selectReadStageMask_lo[563:560]},
     {selectReadStageMask_lo[559:556]},
     {selectReadStageMask_lo[555:552]},
     {selectReadStageMask_lo[551:548]},
     {selectReadStageMask_lo[547:544]},
     {selectReadStageMask_lo[543:540]},
     {selectReadStageMask_lo[539:536]},
     {selectReadStageMask_lo[535:532]},
     {selectReadStageMask_lo[531:528]},
     {selectReadStageMask_lo[527:524]},
     {selectReadStageMask_lo[523:520]},
     {selectReadStageMask_lo[519:516]},
     {selectReadStageMask_lo[515:512]},
     {selectReadStageMask_lo[511:508]},
     {selectReadStageMask_lo[507:504]},
     {selectReadStageMask_lo[503:500]},
     {selectReadStageMask_lo[499:496]},
     {selectReadStageMask_lo[495:492]},
     {selectReadStageMask_lo[491:488]},
     {selectReadStageMask_lo[487:484]},
     {selectReadStageMask_lo[483:480]},
     {selectReadStageMask_lo[479:476]},
     {selectReadStageMask_lo[475:472]},
     {selectReadStageMask_lo[471:468]},
     {selectReadStageMask_lo[467:464]},
     {selectReadStageMask_lo[463:460]},
     {selectReadStageMask_lo[459:456]},
     {selectReadStageMask_lo[455:452]},
     {selectReadStageMask_lo[451:448]},
     {selectReadStageMask_lo[447:444]},
     {selectReadStageMask_lo[443:440]},
     {selectReadStageMask_lo[439:436]},
     {selectReadStageMask_lo[435:432]},
     {selectReadStageMask_lo[431:428]},
     {selectReadStageMask_lo[427:424]},
     {selectReadStageMask_lo[423:420]},
     {selectReadStageMask_lo[419:416]},
     {selectReadStageMask_lo[415:412]},
     {selectReadStageMask_lo[411:408]},
     {selectReadStageMask_lo[407:404]},
     {selectReadStageMask_lo[403:400]},
     {selectReadStageMask_lo[399:396]},
     {selectReadStageMask_lo[395:392]},
     {selectReadStageMask_lo[391:388]},
     {selectReadStageMask_lo[387:384]},
     {selectReadStageMask_lo[383:380]},
     {selectReadStageMask_lo[379:376]},
     {selectReadStageMask_lo[375:372]},
     {selectReadStageMask_lo[371:368]},
     {selectReadStageMask_lo[367:364]},
     {selectReadStageMask_lo[363:360]},
     {selectReadStageMask_lo[359:356]},
     {selectReadStageMask_lo[355:352]},
     {selectReadStageMask_lo[351:348]},
     {selectReadStageMask_lo[347:344]},
     {selectReadStageMask_lo[343:340]},
     {selectReadStageMask_lo[339:336]},
     {selectReadStageMask_lo[335:332]},
     {selectReadStageMask_lo[331:328]},
     {selectReadStageMask_lo[327:324]},
     {selectReadStageMask_lo[323:320]},
     {selectReadStageMask_lo[319:316]},
     {selectReadStageMask_lo[315:312]},
     {selectReadStageMask_lo[311:308]},
     {selectReadStageMask_lo[307:304]},
     {selectReadStageMask_lo[303:300]},
     {selectReadStageMask_lo[299:296]},
     {selectReadStageMask_lo[295:292]},
     {selectReadStageMask_lo[291:288]},
     {selectReadStageMask_lo[287:284]},
     {selectReadStageMask_lo[283:280]},
     {selectReadStageMask_lo[279:276]},
     {selectReadStageMask_lo[275:272]},
     {selectReadStageMask_lo[271:268]},
     {selectReadStageMask_lo[267:264]},
     {selectReadStageMask_lo[263:260]},
     {selectReadStageMask_lo[259:256]},
     {selectReadStageMask_lo[255:252]},
     {selectReadStageMask_lo[251:248]},
     {selectReadStageMask_lo[247:244]},
     {selectReadStageMask_lo[243:240]},
     {selectReadStageMask_lo[239:236]},
     {selectReadStageMask_lo[235:232]},
     {selectReadStageMask_lo[231:228]},
     {selectReadStageMask_lo[227:224]},
     {selectReadStageMask_lo[223:220]},
     {selectReadStageMask_lo[219:216]},
     {selectReadStageMask_lo[215:212]},
     {selectReadStageMask_lo[211:208]},
     {selectReadStageMask_lo[207:204]},
     {selectReadStageMask_lo[203:200]},
     {selectReadStageMask_lo[199:196]},
     {selectReadStageMask_lo[195:192]},
     {selectReadStageMask_lo[191:188]},
     {selectReadStageMask_lo[187:184]},
     {selectReadStageMask_lo[183:180]},
     {selectReadStageMask_lo[179:176]},
     {selectReadStageMask_lo[175:172]},
     {selectReadStageMask_lo[171:168]},
     {selectReadStageMask_lo[167:164]},
     {selectReadStageMask_lo[163:160]},
     {selectReadStageMask_lo[159:156]},
     {selectReadStageMask_lo[155:152]},
     {selectReadStageMask_lo[151:148]},
     {selectReadStageMask_lo[147:144]},
     {selectReadStageMask_lo[143:140]},
     {selectReadStageMask_lo[139:136]},
     {selectReadStageMask_lo[135:132]},
     {selectReadStageMask_lo[131:128]},
     {selectReadStageMask_lo[127:124]},
     {selectReadStageMask_lo[123:120]},
     {selectReadStageMask_lo[119:116]},
     {selectReadStageMask_lo[115:112]},
     {selectReadStageMask_lo[111:108]},
     {selectReadStageMask_lo[107:104]},
     {selectReadStageMask_lo[103:100]},
     {selectReadStageMask_lo[99:96]},
     {selectReadStageMask_lo[95:92]},
     {selectReadStageMask_lo[91:88]},
     {selectReadStageMask_lo[87:84]},
     {selectReadStageMask_lo[83:80]},
     {selectReadStageMask_lo[79:76]},
     {selectReadStageMask_lo[75:72]},
     {selectReadStageMask_lo[71:68]},
     {selectReadStageMask_lo[67:64]},
     {selectReadStageMask_lo[63:60]},
     {selectReadStageMask_lo[59:56]},
     {selectReadStageMask_lo[55:52]},
     {selectReadStageMask_lo[51:48]},
     {selectReadStageMask_lo[47:44]},
     {selectReadStageMask_lo[43:40]},
     {selectReadStageMask_lo[39:36]},
     {selectReadStageMask_lo[35:32]},
     {selectReadStageMask_lo[31:28]},
     {selectReadStageMask_lo[27:24]},
     {selectReadStageMask_lo[23:20]},
     {selectReadStageMask_lo[19:16]},
     {selectReadStageMask_lo[15:12]},
     {selectReadStageMask_lo[11:8]},
     {selectReadStageMask_lo[7:4]},
     {selectReadStageMask_lo[3:0]}};
  wire [3:0]         readMaskCorrection = (instReg_maskType ? _GEN_46[executeGroup[8:0]] : 4'hF) & vlBoundaryCorrection;
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi = {maskSplit_maskSelect_lo_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo = {maskSplit_maskSelect_lo_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo = {maskSplit_maskSelect_lo_lo_hi_lo_hi, maskSplit_maskSelect_lo_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi = {maskSplit_maskSelect_lo_lo_hi_hi_hi, maskSplit_maskSelect_lo_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi = {maskSplit_maskSelect_lo_lo_hi_hi, maskSplit_maskSelect_lo_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_lo = {maskSplit_maskSelect_lo_lo_hi, maskSplit_maskSelect_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo = {maskSplit_maskSelect_lo_hi_lo_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi = {maskSplit_maskSelect_lo_hi_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo = {maskSplit_maskSelect_lo_hi_lo_hi, maskSplit_maskSelect_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo = {maskSplit_maskSelect_lo_hi_hi_lo_hi, maskSplit_maskSelect_lo_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi = {maskSplit_maskSelect_lo_hi_hi_hi, maskSplit_maskSelect_lo_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_lo_hi = {maskSplit_maskSelect_lo_hi_hi, maskSplit_maskSelect_lo_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_lo = {maskSplit_maskSelect_lo_hi, maskSplit_maskSelect_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo = {maskSplit_maskSelect_hi_lo_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi = {maskSplit_maskSelect_hi_lo_lo_hi_hi, maskSplit_maskSelect_hi_lo_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo = {maskSplit_maskSelect_hi_lo_lo_hi, maskSplit_maskSelect_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo = {maskSplit_maskSelect_hi_lo_hi_lo_hi, maskSplit_maskSelect_hi_lo_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi = {maskSplit_maskSelect_hi_lo_hi_hi_hi, maskSplit_maskSelect_hi_lo_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi = {maskSplit_maskSelect_hi_lo_hi_hi, maskSplit_maskSelect_hi_lo_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_lo = {maskSplit_maskSelect_hi_lo_hi, maskSplit_maskSelect_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo = {maskSplit_maskSelect_hi_hi_lo_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi = {maskSplit_maskSelect_hi_hi_lo_hi_hi, maskSplit_maskSelect_hi_hi_lo_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo = {maskSplit_maskSelect_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo = {maskSplit_maskSelect_hi_hi_hi_lo_hi, maskSplit_maskSelect_hi_hi_hi_lo_lo};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_hi_lo};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi = {maskSplit_maskSelect_hi_hi_hi_hi, maskSplit_maskSelect_hi_hi_hi_lo};
  wire [511:0]       maskSplit_maskSelect_hi_hi = {maskSplit_maskSelect_hi_hi_hi, maskSplit_maskSelect_hi_hi_lo};
  wire [1023:0]      maskSplit_maskSelect_hi = {maskSplit_maskSelect_hi_hi, maskSplit_maskSelect_hi_lo};
  wire [7:0]         executeGroupCounter;
  wire               maskSplit_vlMisAlign = |(instReg_vl[3:0]);
  wire [7:0]         maskSplit_lastexecuteGroup = instReg_vl[11:4] - {7'h0, ~maskSplit_vlMisAlign};
  wire               maskSplit_isVlBoundary = executeGroupCounter == maskSplit_lastexecuteGroup;
  wire               maskSplit_validExecuteGroup = executeGroupCounter <= maskSplit_lastexecuteGroup;
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_2 = 16'h1 << instReg_vl[3:0];
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_5 = _maskSplit_vlBoundaryCorrection_T_2 | {_maskSplit_vlBoundaryCorrection_T_2[14:0], 1'h0};
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_8 = _maskSplit_vlBoundaryCorrection_T_5 | {_maskSplit_vlBoundaryCorrection_T_5[13:0], 2'h0};
  wire [15:0]        _maskSplit_vlBoundaryCorrection_T_11 = _maskSplit_vlBoundaryCorrection_T_8 | {_maskSplit_vlBoundaryCorrection_T_8[11:0], 4'h0};
  wire [15:0]        maskSplit_vlBoundaryCorrection = ~({16{maskSplit_vlMisAlign & maskSplit_isVlBoundary}} & (_maskSplit_vlBoundaryCorrection_T_11 | {_maskSplit_vlBoundaryCorrection_T_11[7:0], 8'h0})) & {16{maskSplit_validExecuteGroup}};
  wire [127:0][15:0] _GEN_47 =
    {{maskSplit_maskSelect_hi[1023:1008]},
     {maskSplit_maskSelect_hi[1007:992]},
     {maskSplit_maskSelect_hi[991:976]},
     {maskSplit_maskSelect_hi[975:960]},
     {maskSplit_maskSelect_hi[959:944]},
     {maskSplit_maskSelect_hi[943:928]},
     {maskSplit_maskSelect_hi[927:912]},
     {maskSplit_maskSelect_hi[911:896]},
     {maskSplit_maskSelect_hi[895:880]},
     {maskSplit_maskSelect_hi[879:864]},
     {maskSplit_maskSelect_hi[863:848]},
     {maskSplit_maskSelect_hi[847:832]},
     {maskSplit_maskSelect_hi[831:816]},
     {maskSplit_maskSelect_hi[815:800]},
     {maskSplit_maskSelect_hi[799:784]},
     {maskSplit_maskSelect_hi[783:768]},
     {maskSplit_maskSelect_hi[767:752]},
     {maskSplit_maskSelect_hi[751:736]},
     {maskSplit_maskSelect_hi[735:720]},
     {maskSplit_maskSelect_hi[719:704]},
     {maskSplit_maskSelect_hi[703:688]},
     {maskSplit_maskSelect_hi[687:672]},
     {maskSplit_maskSelect_hi[671:656]},
     {maskSplit_maskSelect_hi[655:640]},
     {maskSplit_maskSelect_hi[639:624]},
     {maskSplit_maskSelect_hi[623:608]},
     {maskSplit_maskSelect_hi[607:592]},
     {maskSplit_maskSelect_hi[591:576]},
     {maskSplit_maskSelect_hi[575:560]},
     {maskSplit_maskSelect_hi[559:544]},
     {maskSplit_maskSelect_hi[543:528]},
     {maskSplit_maskSelect_hi[527:512]},
     {maskSplit_maskSelect_hi[511:496]},
     {maskSplit_maskSelect_hi[495:480]},
     {maskSplit_maskSelect_hi[479:464]},
     {maskSplit_maskSelect_hi[463:448]},
     {maskSplit_maskSelect_hi[447:432]},
     {maskSplit_maskSelect_hi[431:416]},
     {maskSplit_maskSelect_hi[415:400]},
     {maskSplit_maskSelect_hi[399:384]},
     {maskSplit_maskSelect_hi[383:368]},
     {maskSplit_maskSelect_hi[367:352]},
     {maskSplit_maskSelect_hi[351:336]},
     {maskSplit_maskSelect_hi[335:320]},
     {maskSplit_maskSelect_hi[319:304]},
     {maskSplit_maskSelect_hi[303:288]},
     {maskSplit_maskSelect_hi[287:272]},
     {maskSplit_maskSelect_hi[271:256]},
     {maskSplit_maskSelect_hi[255:240]},
     {maskSplit_maskSelect_hi[239:224]},
     {maskSplit_maskSelect_hi[223:208]},
     {maskSplit_maskSelect_hi[207:192]},
     {maskSplit_maskSelect_hi[191:176]},
     {maskSplit_maskSelect_hi[175:160]},
     {maskSplit_maskSelect_hi[159:144]},
     {maskSplit_maskSelect_hi[143:128]},
     {maskSplit_maskSelect_hi[127:112]},
     {maskSplit_maskSelect_hi[111:96]},
     {maskSplit_maskSelect_hi[95:80]},
     {maskSplit_maskSelect_hi[79:64]},
     {maskSplit_maskSelect_hi[63:48]},
     {maskSplit_maskSelect_hi[47:32]},
     {maskSplit_maskSelect_hi[31:16]},
     {maskSplit_maskSelect_hi[15:0]},
     {maskSplit_maskSelect_lo[1023:1008]},
     {maskSplit_maskSelect_lo[1007:992]},
     {maskSplit_maskSelect_lo[991:976]},
     {maskSplit_maskSelect_lo[975:960]},
     {maskSplit_maskSelect_lo[959:944]},
     {maskSplit_maskSelect_lo[943:928]},
     {maskSplit_maskSelect_lo[927:912]},
     {maskSplit_maskSelect_lo[911:896]},
     {maskSplit_maskSelect_lo[895:880]},
     {maskSplit_maskSelect_lo[879:864]},
     {maskSplit_maskSelect_lo[863:848]},
     {maskSplit_maskSelect_lo[847:832]},
     {maskSplit_maskSelect_lo[831:816]},
     {maskSplit_maskSelect_lo[815:800]},
     {maskSplit_maskSelect_lo[799:784]},
     {maskSplit_maskSelect_lo[783:768]},
     {maskSplit_maskSelect_lo[767:752]},
     {maskSplit_maskSelect_lo[751:736]},
     {maskSplit_maskSelect_lo[735:720]},
     {maskSplit_maskSelect_lo[719:704]},
     {maskSplit_maskSelect_lo[703:688]},
     {maskSplit_maskSelect_lo[687:672]},
     {maskSplit_maskSelect_lo[671:656]},
     {maskSplit_maskSelect_lo[655:640]},
     {maskSplit_maskSelect_lo[639:624]},
     {maskSplit_maskSelect_lo[623:608]},
     {maskSplit_maskSelect_lo[607:592]},
     {maskSplit_maskSelect_lo[591:576]},
     {maskSplit_maskSelect_lo[575:560]},
     {maskSplit_maskSelect_lo[559:544]},
     {maskSplit_maskSelect_lo[543:528]},
     {maskSplit_maskSelect_lo[527:512]},
     {maskSplit_maskSelect_lo[511:496]},
     {maskSplit_maskSelect_lo[495:480]},
     {maskSplit_maskSelect_lo[479:464]},
     {maskSplit_maskSelect_lo[463:448]},
     {maskSplit_maskSelect_lo[447:432]},
     {maskSplit_maskSelect_lo[431:416]},
     {maskSplit_maskSelect_lo[415:400]},
     {maskSplit_maskSelect_lo[399:384]},
     {maskSplit_maskSelect_lo[383:368]},
     {maskSplit_maskSelect_lo[367:352]},
     {maskSplit_maskSelect_lo[351:336]},
     {maskSplit_maskSelect_lo[335:320]},
     {maskSplit_maskSelect_lo[319:304]},
     {maskSplit_maskSelect_lo[303:288]},
     {maskSplit_maskSelect_lo[287:272]},
     {maskSplit_maskSelect_lo[271:256]},
     {maskSplit_maskSelect_lo[255:240]},
     {maskSplit_maskSelect_lo[239:224]},
     {maskSplit_maskSelect_lo[223:208]},
     {maskSplit_maskSelect_lo[207:192]},
     {maskSplit_maskSelect_lo[191:176]},
     {maskSplit_maskSelect_lo[175:160]},
     {maskSplit_maskSelect_lo[159:144]},
     {maskSplit_maskSelect_lo[143:128]},
     {maskSplit_maskSelect_lo[127:112]},
     {maskSplit_maskSelect_lo[111:96]},
     {maskSplit_maskSelect_lo[95:80]},
     {maskSplit_maskSelect_lo[79:64]},
     {maskSplit_maskSelect_lo[63:48]},
     {maskSplit_maskSelect_lo[47:32]},
     {maskSplit_maskSelect_lo[31:16]},
     {maskSplit_maskSelect_lo[15:0]}};
  wire [15:0]        maskSplit_0_2 = (instReg_maskType ? _GEN_47[executeGroupCounter[6:0]] : 16'hFFFF) & maskSplit_vlBoundaryCorrection;
  wire [1:0]         maskSplit_byteMask_lo_lo_lo = maskSplit_0_2[1:0];
  wire [1:0]         maskSplit_byteMask_lo_lo_hi = maskSplit_0_2[3:2];
  wire [3:0]         maskSplit_byteMask_lo_lo = {maskSplit_byteMask_lo_lo_hi, maskSplit_byteMask_lo_lo_lo};
  wire [1:0]         maskSplit_byteMask_lo_hi_lo = maskSplit_0_2[5:4];
  wire [1:0]         maskSplit_byteMask_lo_hi_hi = maskSplit_0_2[7:6];
  wire [3:0]         maskSplit_byteMask_lo_hi = {maskSplit_byteMask_lo_hi_hi, maskSplit_byteMask_lo_hi_lo};
  wire [7:0]         maskSplit_byteMask_lo = {maskSplit_byteMask_lo_hi, maskSplit_byteMask_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_lo_lo = maskSplit_0_2[9:8];
  wire [1:0]         maskSplit_byteMask_hi_lo_hi = maskSplit_0_2[11:10];
  wire [3:0]         maskSplit_byteMask_hi_lo = {maskSplit_byteMask_hi_lo_hi, maskSplit_byteMask_hi_lo_lo};
  wire [1:0]         maskSplit_byteMask_hi_hi_lo = maskSplit_0_2[13:12];
  wire [1:0]         maskSplit_byteMask_hi_hi_hi = maskSplit_0_2[15:14];
  wire [3:0]         maskSplit_byteMask_hi_hi = {maskSplit_byteMask_hi_hi_hi, maskSplit_byteMask_hi_hi_lo};
  wire [7:0]         maskSplit_byteMask_hi = {maskSplit_byteMask_hi_hi, maskSplit_byteMask_hi_lo};
  wire [15:0]        maskSplit_0_1 = {maskSplit_byteMask_hi, maskSplit_byteMask_lo};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_1 = {maskSplit_maskSelect_lo_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_1 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_1 = {maskSplit_maskSelect_lo_lo_hi_hi_1, maskSplit_maskSelect_lo_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_lo_1 = {maskSplit_maskSelect_lo_lo_hi_1, maskSplit_maskSelect_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_1 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_1 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_1 = {maskSplit_maskSelect_lo_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_1 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_1 = {maskSplit_maskSelect_lo_hi_hi_hi_1, maskSplit_maskSelect_lo_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_lo_hi_1 = {maskSplit_maskSelect_lo_hi_hi_1, maskSplit_maskSelect_lo_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_lo_1 = {maskSplit_maskSelect_lo_hi_1, maskSplit_maskSelect_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_1 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_1 = {maskSplit_maskSelect_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_1 = {maskSplit_maskSelect_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_lo_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_lo_1 = {maskSplit_maskSelect_hi_lo_hi_1, maskSplit_maskSelect_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_1 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_1 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_1 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_lo_1};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_hi_lo_1};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_hi_lo_1};
  wire [511:0]       maskSplit_maskSelect_hi_hi_1 = {maskSplit_maskSelect_hi_hi_hi_1, maskSplit_maskSelect_hi_hi_lo_1};
  wire [1023:0]      maskSplit_maskSelect_hi_1 = {maskSplit_maskSelect_hi_hi_1, maskSplit_maskSelect_hi_lo_1};
  wire               maskSplit_vlMisAlign_1 = |(instReg_vl[2:0]);
  wire [8:0]         maskSplit_lastexecuteGroup_1 = instReg_vl[11:3] - {8'h0, ~maskSplit_vlMisAlign_1};
  wire [8:0]         _GEN_48 = {1'h0, executeGroupCounter};
  wire               maskSplit_isVlBoundary_1 = _GEN_48 == maskSplit_lastexecuteGroup_1;
  wire               maskSplit_validExecuteGroup_1 = _GEN_48 <= maskSplit_lastexecuteGroup_1;
  wire [7:0]         _maskSplit_vlBoundaryCorrection_T_21 = 8'h1 << instReg_vl[2:0];
  wire [7:0]         _maskSplit_vlBoundaryCorrection_T_24 = _maskSplit_vlBoundaryCorrection_T_21 | {_maskSplit_vlBoundaryCorrection_T_21[6:0], 1'h0};
  wire [7:0]         _maskSplit_vlBoundaryCorrection_T_27 = _maskSplit_vlBoundaryCorrection_T_24 | {_maskSplit_vlBoundaryCorrection_T_24[5:0], 2'h0};
  wire [7:0]         maskSplit_vlBoundaryCorrection_1 =
    ~({8{maskSplit_vlMisAlign_1 & maskSplit_isVlBoundary_1}} & (_maskSplit_vlBoundaryCorrection_T_27 | {_maskSplit_vlBoundaryCorrection_T_27[3:0], 4'h0})) & {8{maskSplit_validExecuteGroup_1}};
  wire [255:0][7:0]  _GEN_49 =
    {{maskSplit_maskSelect_hi_1[1023:1016]},
     {maskSplit_maskSelect_hi_1[1015:1008]},
     {maskSplit_maskSelect_hi_1[1007:1000]},
     {maskSplit_maskSelect_hi_1[999:992]},
     {maskSplit_maskSelect_hi_1[991:984]},
     {maskSplit_maskSelect_hi_1[983:976]},
     {maskSplit_maskSelect_hi_1[975:968]},
     {maskSplit_maskSelect_hi_1[967:960]},
     {maskSplit_maskSelect_hi_1[959:952]},
     {maskSplit_maskSelect_hi_1[951:944]},
     {maskSplit_maskSelect_hi_1[943:936]},
     {maskSplit_maskSelect_hi_1[935:928]},
     {maskSplit_maskSelect_hi_1[927:920]},
     {maskSplit_maskSelect_hi_1[919:912]},
     {maskSplit_maskSelect_hi_1[911:904]},
     {maskSplit_maskSelect_hi_1[903:896]},
     {maskSplit_maskSelect_hi_1[895:888]},
     {maskSplit_maskSelect_hi_1[887:880]},
     {maskSplit_maskSelect_hi_1[879:872]},
     {maskSplit_maskSelect_hi_1[871:864]},
     {maskSplit_maskSelect_hi_1[863:856]},
     {maskSplit_maskSelect_hi_1[855:848]},
     {maskSplit_maskSelect_hi_1[847:840]},
     {maskSplit_maskSelect_hi_1[839:832]},
     {maskSplit_maskSelect_hi_1[831:824]},
     {maskSplit_maskSelect_hi_1[823:816]},
     {maskSplit_maskSelect_hi_1[815:808]},
     {maskSplit_maskSelect_hi_1[807:800]},
     {maskSplit_maskSelect_hi_1[799:792]},
     {maskSplit_maskSelect_hi_1[791:784]},
     {maskSplit_maskSelect_hi_1[783:776]},
     {maskSplit_maskSelect_hi_1[775:768]},
     {maskSplit_maskSelect_hi_1[767:760]},
     {maskSplit_maskSelect_hi_1[759:752]},
     {maskSplit_maskSelect_hi_1[751:744]},
     {maskSplit_maskSelect_hi_1[743:736]},
     {maskSplit_maskSelect_hi_1[735:728]},
     {maskSplit_maskSelect_hi_1[727:720]},
     {maskSplit_maskSelect_hi_1[719:712]},
     {maskSplit_maskSelect_hi_1[711:704]},
     {maskSplit_maskSelect_hi_1[703:696]},
     {maskSplit_maskSelect_hi_1[695:688]},
     {maskSplit_maskSelect_hi_1[687:680]},
     {maskSplit_maskSelect_hi_1[679:672]},
     {maskSplit_maskSelect_hi_1[671:664]},
     {maskSplit_maskSelect_hi_1[663:656]},
     {maskSplit_maskSelect_hi_1[655:648]},
     {maskSplit_maskSelect_hi_1[647:640]},
     {maskSplit_maskSelect_hi_1[639:632]},
     {maskSplit_maskSelect_hi_1[631:624]},
     {maskSplit_maskSelect_hi_1[623:616]},
     {maskSplit_maskSelect_hi_1[615:608]},
     {maskSplit_maskSelect_hi_1[607:600]},
     {maskSplit_maskSelect_hi_1[599:592]},
     {maskSplit_maskSelect_hi_1[591:584]},
     {maskSplit_maskSelect_hi_1[583:576]},
     {maskSplit_maskSelect_hi_1[575:568]},
     {maskSplit_maskSelect_hi_1[567:560]},
     {maskSplit_maskSelect_hi_1[559:552]},
     {maskSplit_maskSelect_hi_1[551:544]},
     {maskSplit_maskSelect_hi_1[543:536]},
     {maskSplit_maskSelect_hi_1[535:528]},
     {maskSplit_maskSelect_hi_1[527:520]},
     {maskSplit_maskSelect_hi_1[519:512]},
     {maskSplit_maskSelect_hi_1[511:504]},
     {maskSplit_maskSelect_hi_1[503:496]},
     {maskSplit_maskSelect_hi_1[495:488]},
     {maskSplit_maskSelect_hi_1[487:480]},
     {maskSplit_maskSelect_hi_1[479:472]},
     {maskSplit_maskSelect_hi_1[471:464]},
     {maskSplit_maskSelect_hi_1[463:456]},
     {maskSplit_maskSelect_hi_1[455:448]},
     {maskSplit_maskSelect_hi_1[447:440]},
     {maskSplit_maskSelect_hi_1[439:432]},
     {maskSplit_maskSelect_hi_1[431:424]},
     {maskSplit_maskSelect_hi_1[423:416]},
     {maskSplit_maskSelect_hi_1[415:408]},
     {maskSplit_maskSelect_hi_1[407:400]},
     {maskSplit_maskSelect_hi_1[399:392]},
     {maskSplit_maskSelect_hi_1[391:384]},
     {maskSplit_maskSelect_hi_1[383:376]},
     {maskSplit_maskSelect_hi_1[375:368]},
     {maskSplit_maskSelect_hi_1[367:360]},
     {maskSplit_maskSelect_hi_1[359:352]},
     {maskSplit_maskSelect_hi_1[351:344]},
     {maskSplit_maskSelect_hi_1[343:336]},
     {maskSplit_maskSelect_hi_1[335:328]},
     {maskSplit_maskSelect_hi_1[327:320]},
     {maskSplit_maskSelect_hi_1[319:312]},
     {maskSplit_maskSelect_hi_1[311:304]},
     {maskSplit_maskSelect_hi_1[303:296]},
     {maskSplit_maskSelect_hi_1[295:288]},
     {maskSplit_maskSelect_hi_1[287:280]},
     {maskSplit_maskSelect_hi_1[279:272]},
     {maskSplit_maskSelect_hi_1[271:264]},
     {maskSplit_maskSelect_hi_1[263:256]},
     {maskSplit_maskSelect_hi_1[255:248]},
     {maskSplit_maskSelect_hi_1[247:240]},
     {maskSplit_maskSelect_hi_1[239:232]},
     {maskSplit_maskSelect_hi_1[231:224]},
     {maskSplit_maskSelect_hi_1[223:216]},
     {maskSplit_maskSelect_hi_1[215:208]},
     {maskSplit_maskSelect_hi_1[207:200]},
     {maskSplit_maskSelect_hi_1[199:192]},
     {maskSplit_maskSelect_hi_1[191:184]},
     {maskSplit_maskSelect_hi_1[183:176]},
     {maskSplit_maskSelect_hi_1[175:168]},
     {maskSplit_maskSelect_hi_1[167:160]},
     {maskSplit_maskSelect_hi_1[159:152]},
     {maskSplit_maskSelect_hi_1[151:144]},
     {maskSplit_maskSelect_hi_1[143:136]},
     {maskSplit_maskSelect_hi_1[135:128]},
     {maskSplit_maskSelect_hi_1[127:120]},
     {maskSplit_maskSelect_hi_1[119:112]},
     {maskSplit_maskSelect_hi_1[111:104]},
     {maskSplit_maskSelect_hi_1[103:96]},
     {maskSplit_maskSelect_hi_1[95:88]},
     {maskSplit_maskSelect_hi_1[87:80]},
     {maskSplit_maskSelect_hi_1[79:72]},
     {maskSplit_maskSelect_hi_1[71:64]},
     {maskSplit_maskSelect_hi_1[63:56]},
     {maskSplit_maskSelect_hi_1[55:48]},
     {maskSplit_maskSelect_hi_1[47:40]},
     {maskSplit_maskSelect_hi_1[39:32]},
     {maskSplit_maskSelect_hi_1[31:24]},
     {maskSplit_maskSelect_hi_1[23:16]},
     {maskSplit_maskSelect_hi_1[15:8]},
     {maskSplit_maskSelect_hi_1[7:0]},
     {maskSplit_maskSelect_lo_1[1023:1016]},
     {maskSplit_maskSelect_lo_1[1015:1008]},
     {maskSplit_maskSelect_lo_1[1007:1000]},
     {maskSplit_maskSelect_lo_1[999:992]},
     {maskSplit_maskSelect_lo_1[991:984]},
     {maskSplit_maskSelect_lo_1[983:976]},
     {maskSplit_maskSelect_lo_1[975:968]},
     {maskSplit_maskSelect_lo_1[967:960]},
     {maskSplit_maskSelect_lo_1[959:952]},
     {maskSplit_maskSelect_lo_1[951:944]},
     {maskSplit_maskSelect_lo_1[943:936]},
     {maskSplit_maskSelect_lo_1[935:928]},
     {maskSplit_maskSelect_lo_1[927:920]},
     {maskSplit_maskSelect_lo_1[919:912]},
     {maskSplit_maskSelect_lo_1[911:904]},
     {maskSplit_maskSelect_lo_1[903:896]},
     {maskSplit_maskSelect_lo_1[895:888]},
     {maskSplit_maskSelect_lo_1[887:880]},
     {maskSplit_maskSelect_lo_1[879:872]},
     {maskSplit_maskSelect_lo_1[871:864]},
     {maskSplit_maskSelect_lo_1[863:856]},
     {maskSplit_maskSelect_lo_1[855:848]},
     {maskSplit_maskSelect_lo_1[847:840]},
     {maskSplit_maskSelect_lo_1[839:832]},
     {maskSplit_maskSelect_lo_1[831:824]},
     {maskSplit_maskSelect_lo_1[823:816]},
     {maskSplit_maskSelect_lo_1[815:808]},
     {maskSplit_maskSelect_lo_1[807:800]},
     {maskSplit_maskSelect_lo_1[799:792]},
     {maskSplit_maskSelect_lo_1[791:784]},
     {maskSplit_maskSelect_lo_1[783:776]},
     {maskSplit_maskSelect_lo_1[775:768]},
     {maskSplit_maskSelect_lo_1[767:760]},
     {maskSplit_maskSelect_lo_1[759:752]},
     {maskSplit_maskSelect_lo_1[751:744]},
     {maskSplit_maskSelect_lo_1[743:736]},
     {maskSplit_maskSelect_lo_1[735:728]},
     {maskSplit_maskSelect_lo_1[727:720]},
     {maskSplit_maskSelect_lo_1[719:712]},
     {maskSplit_maskSelect_lo_1[711:704]},
     {maskSplit_maskSelect_lo_1[703:696]},
     {maskSplit_maskSelect_lo_1[695:688]},
     {maskSplit_maskSelect_lo_1[687:680]},
     {maskSplit_maskSelect_lo_1[679:672]},
     {maskSplit_maskSelect_lo_1[671:664]},
     {maskSplit_maskSelect_lo_1[663:656]},
     {maskSplit_maskSelect_lo_1[655:648]},
     {maskSplit_maskSelect_lo_1[647:640]},
     {maskSplit_maskSelect_lo_1[639:632]},
     {maskSplit_maskSelect_lo_1[631:624]},
     {maskSplit_maskSelect_lo_1[623:616]},
     {maskSplit_maskSelect_lo_1[615:608]},
     {maskSplit_maskSelect_lo_1[607:600]},
     {maskSplit_maskSelect_lo_1[599:592]},
     {maskSplit_maskSelect_lo_1[591:584]},
     {maskSplit_maskSelect_lo_1[583:576]},
     {maskSplit_maskSelect_lo_1[575:568]},
     {maskSplit_maskSelect_lo_1[567:560]},
     {maskSplit_maskSelect_lo_1[559:552]},
     {maskSplit_maskSelect_lo_1[551:544]},
     {maskSplit_maskSelect_lo_1[543:536]},
     {maskSplit_maskSelect_lo_1[535:528]},
     {maskSplit_maskSelect_lo_1[527:520]},
     {maskSplit_maskSelect_lo_1[519:512]},
     {maskSplit_maskSelect_lo_1[511:504]},
     {maskSplit_maskSelect_lo_1[503:496]},
     {maskSplit_maskSelect_lo_1[495:488]},
     {maskSplit_maskSelect_lo_1[487:480]},
     {maskSplit_maskSelect_lo_1[479:472]},
     {maskSplit_maskSelect_lo_1[471:464]},
     {maskSplit_maskSelect_lo_1[463:456]},
     {maskSplit_maskSelect_lo_1[455:448]},
     {maskSplit_maskSelect_lo_1[447:440]},
     {maskSplit_maskSelect_lo_1[439:432]},
     {maskSplit_maskSelect_lo_1[431:424]},
     {maskSplit_maskSelect_lo_1[423:416]},
     {maskSplit_maskSelect_lo_1[415:408]},
     {maskSplit_maskSelect_lo_1[407:400]},
     {maskSplit_maskSelect_lo_1[399:392]},
     {maskSplit_maskSelect_lo_1[391:384]},
     {maskSplit_maskSelect_lo_1[383:376]},
     {maskSplit_maskSelect_lo_1[375:368]},
     {maskSplit_maskSelect_lo_1[367:360]},
     {maskSplit_maskSelect_lo_1[359:352]},
     {maskSplit_maskSelect_lo_1[351:344]},
     {maskSplit_maskSelect_lo_1[343:336]},
     {maskSplit_maskSelect_lo_1[335:328]},
     {maskSplit_maskSelect_lo_1[327:320]},
     {maskSplit_maskSelect_lo_1[319:312]},
     {maskSplit_maskSelect_lo_1[311:304]},
     {maskSplit_maskSelect_lo_1[303:296]},
     {maskSplit_maskSelect_lo_1[295:288]},
     {maskSplit_maskSelect_lo_1[287:280]},
     {maskSplit_maskSelect_lo_1[279:272]},
     {maskSplit_maskSelect_lo_1[271:264]},
     {maskSplit_maskSelect_lo_1[263:256]},
     {maskSplit_maskSelect_lo_1[255:248]},
     {maskSplit_maskSelect_lo_1[247:240]},
     {maskSplit_maskSelect_lo_1[239:232]},
     {maskSplit_maskSelect_lo_1[231:224]},
     {maskSplit_maskSelect_lo_1[223:216]},
     {maskSplit_maskSelect_lo_1[215:208]},
     {maskSplit_maskSelect_lo_1[207:200]},
     {maskSplit_maskSelect_lo_1[199:192]},
     {maskSplit_maskSelect_lo_1[191:184]},
     {maskSplit_maskSelect_lo_1[183:176]},
     {maskSplit_maskSelect_lo_1[175:168]},
     {maskSplit_maskSelect_lo_1[167:160]},
     {maskSplit_maskSelect_lo_1[159:152]},
     {maskSplit_maskSelect_lo_1[151:144]},
     {maskSplit_maskSelect_lo_1[143:136]},
     {maskSplit_maskSelect_lo_1[135:128]},
     {maskSplit_maskSelect_lo_1[127:120]},
     {maskSplit_maskSelect_lo_1[119:112]},
     {maskSplit_maskSelect_lo_1[111:104]},
     {maskSplit_maskSelect_lo_1[103:96]},
     {maskSplit_maskSelect_lo_1[95:88]},
     {maskSplit_maskSelect_lo_1[87:80]},
     {maskSplit_maskSelect_lo_1[79:72]},
     {maskSplit_maskSelect_lo_1[71:64]},
     {maskSplit_maskSelect_lo_1[63:56]},
     {maskSplit_maskSelect_lo_1[55:48]},
     {maskSplit_maskSelect_lo_1[47:40]},
     {maskSplit_maskSelect_lo_1[39:32]},
     {maskSplit_maskSelect_lo_1[31:24]},
     {maskSplit_maskSelect_lo_1[23:16]},
     {maskSplit_maskSelect_lo_1[15:8]},
     {maskSplit_maskSelect_lo_1[7:0]}};
  wire [7:0]         maskSplit_1_2 = (instReg_maskType ? _GEN_49[executeGroupCounter] : 8'hFF) & maskSplit_vlBoundaryCorrection_1;
  wire [3:0]         maskSplit_byteMask_lo_lo_1 = {{2{maskSplit_1_2[1]}}, {2{maskSplit_1_2[0]}}};
  wire [3:0]         maskSplit_byteMask_lo_hi_1 = {{2{maskSplit_1_2[3]}}, {2{maskSplit_1_2[2]}}};
  wire [7:0]         maskSplit_byteMask_lo_1 = {maskSplit_byteMask_lo_hi_1, maskSplit_byteMask_lo_lo_1};
  wire [3:0]         maskSplit_byteMask_hi_lo_1 = {{2{maskSplit_1_2[5]}}, {2{maskSplit_1_2[4]}}};
  wire [3:0]         maskSplit_byteMask_hi_hi_1 = {{2{maskSplit_1_2[7]}}, {2{maskSplit_1_2[6]}}};
  wire [7:0]         maskSplit_byteMask_hi_1 = {maskSplit_byteMask_hi_hi_1, maskSplit_byteMask_hi_lo_1};
  wire [15:0]        maskSplit_1_1 = {maskSplit_byteMask_hi_1, maskSplit_byteMask_lo_1};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_lo_2 = {maskSplit_maskSelect_lo_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_lo_2 = {maskSplit_maskSelect_lo_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_lo_hi_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_lo_hi_2 = {maskSplit_maskSelect_lo_lo_hi_hi_2, maskSplit_maskSelect_lo_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_lo_2 = {maskSplit_maskSelect_lo_lo_hi_2, maskSplit_maskSelect_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_lo_2 = {maskSplit_maskSelect_lo_hi_lo_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_lo_hi_2 = {maskSplit_maskSelect_lo_hi_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_lo_2 = {maskSplit_maskSelect_lo_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_lo_2 = {maskSplit_maskSelect_lo_hi_hi_lo_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_lo_hi_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_lo_hi_hi_2 = {maskSplit_maskSelect_lo_hi_hi_hi_2, maskSplit_maskSelect_lo_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_lo_hi_2 = {maskSplit_maskSelect_lo_hi_hi_2, maskSplit_maskSelect_lo_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_lo_2 = {maskSplit_maskSelect_lo_hi_2, maskSplit_maskSelect_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_lo_hi_2 = {maskSplit_maskSelect_hi_lo_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_lo_2 = {maskSplit_maskSelect_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_lo_hi_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_lo_hi_2 = {maskSplit_maskSelect_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_lo_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_lo_2 = {maskSplit_maskSelect_hi_lo_hi_2, maskSplit_maskSelect_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_lo_2 = {maskSplit_maskSelect_hi_hi_lo_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_lo_hi_2 = {maskSplit_maskSelect_hi_hi_lo_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_lo_2 = {maskSplit_maskSelect_hi_hi_hi_lo_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_lo_2};
  wire [127:0]       maskSplit_maskSelect_hi_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_hi_lo_2};
  wire [255:0]       maskSplit_maskSelect_hi_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_hi_lo_2};
  wire [511:0]       maskSplit_maskSelect_hi_hi_2 = {maskSplit_maskSelect_hi_hi_hi_2, maskSplit_maskSelect_hi_hi_lo_2};
  wire [1023:0]      maskSplit_maskSelect_hi_2 = {maskSplit_maskSelect_hi_hi_2, maskSplit_maskSelect_hi_lo_2};
  wire               maskSplit_vlMisAlign_2;
  assign maskSplit_vlMisAlign_2 = |(instReg_vl[1:0]);
  wire [9:0]         maskSplit_lastexecuteGroup_2 = instReg_vl[11:2] - {9'h0, ~maskSplit_vlMisAlign_2};
  wire [9:0]         _GEN_50 = {2'h0, executeGroupCounter};
  wire               maskSplit_isVlBoundary_2 = _GEN_50 == maskSplit_lastexecuteGroup_2;
  wire               maskSplit_validExecuteGroup_2 = _GEN_50 <= maskSplit_lastexecuteGroup_2;
  wire [3:0]         _maskSplit_vlBoundaryCorrection_T_40 = _maskSplit_vlBoundaryCorrection_T_37 | {_maskSplit_vlBoundaryCorrection_T_37[2:0], 1'h0};
  wire [3:0]         maskSplit_vlBoundaryCorrection_2 =
    ~({4{maskSplit_vlMisAlign_2 & maskSplit_isVlBoundary_2}} & (_maskSplit_vlBoundaryCorrection_T_40 | {_maskSplit_vlBoundaryCorrection_T_40[1:0], 2'h0})) & {4{maskSplit_validExecuteGroup_2}};
  wire [255:0][3:0]  _GEN_51 =
    {{maskSplit_maskSelect_lo_2[1023:1020]},
     {maskSplit_maskSelect_lo_2[1019:1016]},
     {maskSplit_maskSelect_lo_2[1015:1012]},
     {maskSplit_maskSelect_lo_2[1011:1008]},
     {maskSplit_maskSelect_lo_2[1007:1004]},
     {maskSplit_maskSelect_lo_2[1003:1000]},
     {maskSplit_maskSelect_lo_2[999:996]},
     {maskSplit_maskSelect_lo_2[995:992]},
     {maskSplit_maskSelect_lo_2[991:988]},
     {maskSplit_maskSelect_lo_2[987:984]},
     {maskSplit_maskSelect_lo_2[983:980]},
     {maskSplit_maskSelect_lo_2[979:976]},
     {maskSplit_maskSelect_lo_2[975:972]},
     {maskSplit_maskSelect_lo_2[971:968]},
     {maskSplit_maskSelect_lo_2[967:964]},
     {maskSplit_maskSelect_lo_2[963:960]},
     {maskSplit_maskSelect_lo_2[959:956]},
     {maskSplit_maskSelect_lo_2[955:952]},
     {maskSplit_maskSelect_lo_2[951:948]},
     {maskSplit_maskSelect_lo_2[947:944]},
     {maskSplit_maskSelect_lo_2[943:940]},
     {maskSplit_maskSelect_lo_2[939:936]},
     {maskSplit_maskSelect_lo_2[935:932]},
     {maskSplit_maskSelect_lo_2[931:928]},
     {maskSplit_maskSelect_lo_2[927:924]},
     {maskSplit_maskSelect_lo_2[923:920]},
     {maskSplit_maskSelect_lo_2[919:916]},
     {maskSplit_maskSelect_lo_2[915:912]},
     {maskSplit_maskSelect_lo_2[911:908]},
     {maskSplit_maskSelect_lo_2[907:904]},
     {maskSplit_maskSelect_lo_2[903:900]},
     {maskSplit_maskSelect_lo_2[899:896]},
     {maskSplit_maskSelect_lo_2[895:892]},
     {maskSplit_maskSelect_lo_2[891:888]},
     {maskSplit_maskSelect_lo_2[887:884]},
     {maskSplit_maskSelect_lo_2[883:880]},
     {maskSplit_maskSelect_lo_2[879:876]},
     {maskSplit_maskSelect_lo_2[875:872]},
     {maskSplit_maskSelect_lo_2[871:868]},
     {maskSplit_maskSelect_lo_2[867:864]},
     {maskSplit_maskSelect_lo_2[863:860]},
     {maskSplit_maskSelect_lo_2[859:856]},
     {maskSplit_maskSelect_lo_2[855:852]},
     {maskSplit_maskSelect_lo_2[851:848]},
     {maskSplit_maskSelect_lo_2[847:844]},
     {maskSplit_maskSelect_lo_2[843:840]},
     {maskSplit_maskSelect_lo_2[839:836]},
     {maskSplit_maskSelect_lo_2[835:832]},
     {maskSplit_maskSelect_lo_2[831:828]},
     {maskSplit_maskSelect_lo_2[827:824]},
     {maskSplit_maskSelect_lo_2[823:820]},
     {maskSplit_maskSelect_lo_2[819:816]},
     {maskSplit_maskSelect_lo_2[815:812]},
     {maskSplit_maskSelect_lo_2[811:808]},
     {maskSplit_maskSelect_lo_2[807:804]},
     {maskSplit_maskSelect_lo_2[803:800]},
     {maskSplit_maskSelect_lo_2[799:796]},
     {maskSplit_maskSelect_lo_2[795:792]},
     {maskSplit_maskSelect_lo_2[791:788]},
     {maskSplit_maskSelect_lo_2[787:784]},
     {maskSplit_maskSelect_lo_2[783:780]},
     {maskSplit_maskSelect_lo_2[779:776]},
     {maskSplit_maskSelect_lo_2[775:772]},
     {maskSplit_maskSelect_lo_2[771:768]},
     {maskSplit_maskSelect_lo_2[767:764]},
     {maskSplit_maskSelect_lo_2[763:760]},
     {maskSplit_maskSelect_lo_2[759:756]},
     {maskSplit_maskSelect_lo_2[755:752]},
     {maskSplit_maskSelect_lo_2[751:748]},
     {maskSplit_maskSelect_lo_2[747:744]},
     {maskSplit_maskSelect_lo_2[743:740]},
     {maskSplit_maskSelect_lo_2[739:736]},
     {maskSplit_maskSelect_lo_2[735:732]},
     {maskSplit_maskSelect_lo_2[731:728]},
     {maskSplit_maskSelect_lo_2[727:724]},
     {maskSplit_maskSelect_lo_2[723:720]},
     {maskSplit_maskSelect_lo_2[719:716]},
     {maskSplit_maskSelect_lo_2[715:712]},
     {maskSplit_maskSelect_lo_2[711:708]},
     {maskSplit_maskSelect_lo_2[707:704]},
     {maskSplit_maskSelect_lo_2[703:700]},
     {maskSplit_maskSelect_lo_2[699:696]},
     {maskSplit_maskSelect_lo_2[695:692]},
     {maskSplit_maskSelect_lo_2[691:688]},
     {maskSplit_maskSelect_lo_2[687:684]},
     {maskSplit_maskSelect_lo_2[683:680]},
     {maskSplit_maskSelect_lo_2[679:676]},
     {maskSplit_maskSelect_lo_2[675:672]},
     {maskSplit_maskSelect_lo_2[671:668]},
     {maskSplit_maskSelect_lo_2[667:664]},
     {maskSplit_maskSelect_lo_2[663:660]},
     {maskSplit_maskSelect_lo_2[659:656]},
     {maskSplit_maskSelect_lo_2[655:652]},
     {maskSplit_maskSelect_lo_2[651:648]},
     {maskSplit_maskSelect_lo_2[647:644]},
     {maskSplit_maskSelect_lo_2[643:640]},
     {maskSplit_maskSelect_lo_2[639:636]},
     {maskSplit_maskSelect_lo_2[635:632]},
     {maskSplit_maskSelect_lo_2[631:628]},
     {maskSplit_maskSelect_lo_2[627:624]},
     {maskSplit_maskSelect_lo_2[623:620]},
     {maskSplit_maskSelect_lo_2[619:616]},
     {maskSplit_maskSelect_lo_2[615:612]},
     {maskSplit_maskSelect_lo_2[611:608]},
     {maskSplit_maskSelect_lo_2[607:604]},
     {maskSplit_maskSelect_lo_2[603:600]},
     {maskSplit_maskSelect_lo_2[599:596]},
     {maskSplit_maskSelect_lo_2[595:592]},
     {maskSplit_maskSelect_lo_2[591:588]},
     {maskSplit_maskSelect_lo_2[587:584]},
     {maskSplit_maskSelect_lo_2[583:580]},
     {maskSplit_maskSelect_lo_2[579:576]},
     {maskSplit_maskSelect_lo_2[575:572]},
     {maskSplit_maskSelect_lo_2[571:568]},
     {maskSplit_maskSelect_lo_2[567:564]},
     {maskSplit_maskSelect_lo_2[563:560]},
     {maskSplit_maskSelect_lo_2[559:556]},
     {maskSplit_maskSelect_lo_2[555:552]},
     {maskSplit_maskSelect_lo_2[551:548]},
     {maskSplit_maskSelect_lo_2[547:544]},
     {maskSplit_maskSelect_lo_2[543:540]},
     {maskSplit_maskSelect_lo_2[539:536]},
     {maskSplit_maskSelect_lo_2[535:532]},
     {maskSplit_maskSelect_lo_2[531:528]},
     {maskSplit_maskSelect_lo_2[527:524]},
     {maskSplit_maskSelect_lo_2[523:520]},
     {maskSplit_maskSelect_lo_2[519:516]},
     {maskSplit_maskSelect_lo_2[515:512]},
     {maskSplit_maskSelect_lo_2[511:508]},
     {maskSplit_maskSelect_lo_2[507:504]},
     {maskSplit_maskSelect_lo_2[503:500]},
     {maskSplit_maskSelect_lo_2[499:496]},
     {maskSplit_maskSelect_lo_2[495:492]},
     {maskSplit_maskSelect_lo_2[491:488]},
     {maskSplit_maskSelect_lo_2[487:484]},
     {maskSplit_maskSelect_lo_2[483:480]},
     {maskSplit_maskSelect_lo_2[479:476]},
     {maskSplit_maskSelect_lo_2[475:472]},
     {maskSplit_maskSelect_lo_2[471:468]},
     {maskSplit_maskSelect_lo_2[467:464]},
     {maskSplit_maskSelect_lo_2[463:460]},
     {maskSplit_maskSelect_lo_2[459:456]},
     {maskSplit_maskSelect_lo_2[455:452]},
     {maskSplit_maskSelect_lo_2[451:448]},
     {maskSplit_maskSelect_lo_2[447:444]},
     {maskSplit_maskSelect_lo_2[443:440]},
     {maskSplit_maskSelect_lo_2[439:436]},
     {maskSplit_maskSelect_lo_2[435:432]},
     {maskSplit_maskSelect_lo_2[431:428]},
     {maskSplit_maskSelect_lo_2[427:424]},
     {maskSplit_maskSelect_lo_2[423:420]},
     {maskSplit_maskSelect_lo_2[419:416]},
     {maskSplit_maskSelect_lo_2[415:412]},
     {maskSplit_maskSelect_lo_2[411:408]},
     {maskSplit_maskSelect_lo_2[407:404]},
     {maskSplit_maskSelect_lo_2[403:400]},
     {maskSplit_maskSelect_lo_2[399:396]},
     {maskSplit_maskSelect_lo_2[395:392]},
     {maskSplit_maskSelect_lo_2[391:388]},
     {maskSplit_maskSelect_lo_2[387:384]},
     {maskSplit_maskSelect_lo_2[383:380]},
     {maskSplit_maskSelect_lo_2[379:376]},
     {maskSplit_maskSelect_lo_2[375:372]},
     {maskSplit_maskSelect_lo_2[371:368]},
     {maskSplit_maskSelect_lo_2[367:364]},
     {maskSplit_maskSelect_lo_2[363:360]},
     {maskSplit_maskSelect_lo_2[359:356]},
     {maskSplit_maskSelect_lo_2[355:352]},
     {maskSplit_maskSelect_lo_2[351:348]},
     {maskSplit_maskSelect_lo_2[347:344]},
     {maskSplit_maskSelect_lo_2[343:340]},
     {maskSplit_maskSelect_lo_2[339:336]},
     {maskSplit_maskSelect_lo_2[335:332]},
     {maskSplit_maskSelect_lo_2[331:328]},
     {maskSplit_maskSelect_lo_2[327:324]},
     {maskSplit_maskSelect_lo_2[323:320]},
     {maskSplit_maskSelect_lo_2[319:316]},
     {maskSplit_maskSelect_lo_2[315:312]},
     {maskSplit_maskSelect_lo_2[311:308]},
     {maskSplit_maskSelect_lo_2[307:304]},
     {maskSplit_maskSelect_lo_2[303:300]},
     {maskSplit_maskSelect_lo_2[299:296]},
     {maskSplit_maskSelect_lo_2[295:292]},
     {maskSplit_maskSelect_lo_2[291:288]},
     {maskSplit_maskSelect_lo_2[287:284]},
     {maskSplit_maskSelect_lo_2[283:280]},
     {maskSplit_maskSelect_lo_2[279:276]},
     {maskSplit_maskSelect_lo_2[275:272]},
     {maskSplit_maskSelect_lo_2[271:268]},
     {maskSplit_maskSelect_lo_2[267:264]},
     {maskSplit_maskSelect_lo_2[263:260]},
     {maskSplit_maskSelect_lo_2[259:256]},
     {maskSplit_maskSelect_lo_2[255:252]},
     {maskSplit_maskSelect_lo_2[251:248]},
     {maskSplit_maskSelect_lo_2[247:244]},
     {maskSplit_maskSelect_lo_2[243:240]},
     {maskSplit_maskSelect_lo_2[239:236]},
     {maskSplit_maskSelect_lo_2[235:232]},
     {maskSplit_maskSelect_lo_2[231:228]},
     {maskSplit_maskSelect_lo_2[227:224]},
     {maskSplit_maskSelect_lo_2[223:220]},
     {maskSplit_maskSelect_lo_2[219:216]},
     {maskSplit_maskSelect_lo_2[215:212]},
     {maskSplit_maskSelect_lo_2[211:208]},
     {maskSplit_maskSelect_lo_2[207:204]},
     {maskSplit_maskSelect_lo_2[203:200]},
     {maskSplit_maskSelect_lo_2[199:196]},
     {maskSplit_maskSelect_lo_2[195:192]},
     {maskSplit_maskSelect_lo_2[191:188]},
     {maskSplit_maskSelect_lo_2[187:184]},
     {maskSplit_maskSelect_lo_2[183:180]},
     {maskSplit_maskSelect_lo_2[179:176]},
     {maskSplit_maskSelect_lo_2[175:172]},
     {maskSplit_maskSelect_lo_2[171:168]},
     {maskSplit_maskSelect_lo_2[167:164]},
     {maskSplit_maskSelect_lo_2[163:160]},
     {maskSplit_maskSelect_lo_2[159:156]},
     {maskSplit_maskSelect_lo_2[155:152]},
     {maskSplit_maskSelect_lo_2[151:148]},
     {maskSplit_maskSelect_lo_2[147:144]},
     {maskSplit_maskSelect_lo_2[143:140]},
     {maskSplit_maskSelect_lo_2[139:136]},
     {maskSplit_maskSelect_lo_2[135:132]},
     {maskSplit_maskSelect_lo_2[131:128]},
     {maskSplit_maskSelect_lo_2[127:124]},
     {maskSplit_maskSelect_lo_2[123:120]},
     {maskSplit_maskSelect_lo_2[119:116]},
     {maskSplit_maskSelect_lo_2[115:112]},
     {maskSplit_maskSelect_lo_2[111:108]},
     {maskSplit_maskSelect_lo_2[107:104]},
     {maskSplit_maskSelect_lo_2[103:100]},
     {maskSplit_maskSelect_lo_2[99:96]},
     {maskSplit_maskSelect_lo_2[95:92]},
     {maskSplit_maskSelect_lo_2[91:88]},
     {maskSplit_maskSelect_lo_2[87:84]},
     {maskSplit_maskSelect_lo_2[83:80]},
     {maskSplit_maskSelect_lo_2[79:76]},
     {maskSplit_maskSelect_lo_2[75:72]},
     {maskSplit_maskSelect_lo_2[71:68]},
     {maskSplit_maskSelect_lo_2[67:64]},
     {maskSplit_maskSelect_lo_2[63:60]},
     {maskSplit_maskSelect_lo_2[59:56]},
     {maskSplit_maskSelect_lo_2[55:52]},
     {maskSplit_maskSelect_lo_2[51:48]},
     {maskSplit_maskSelect_lo_2[47:44]},
     {maskSplit_maskSelect_lo_2[43:40]},
     {maskSplit_maskSelect_lo_2[39:36]},
     {maskSplit_maskSelect_lo_2[35:32]},
     {maskSplit_maskSelect_lo_2[31:28]},
     {maskSplit_maskSelect_lo_2[27:24]},
     {maskSplit_maskSelect_lo_2[23:20]},
     {maskSplit_maskSelect_lo_2[19:16]},
     {maskSplit_maskSelect_lo_2[15:12]},
     {maskSplit_maskSelect_lo_2[11:8]},
     {maskSplit_maskSelect_lo_2[7:4]},
     {maskSplit_maskSelect_lo_2[3:0]}};
  wire [3:0]         maskSplit_2_2 = (instReg_maskType ? _GEN_51[executeGroupCounter] : 4'hF) & maskSplit_vlBoundaryCorrection_2;
  wire [7:0]         maskSplit_byteMask_lo_2 = {{4{maskSplit_2_2[1]}}, {4{maskSplit_2_2[0]}}};
  wire [7:0]         maskSplit_byteMask_hi_2 = {{4{maskSplit_2_2[3]}}, {4{maskSplit_2_2[2]}}};
  wire [15:0]        maskSplit_2_1 = {maskSplit_byteMask_hi_2, maskSplit_byteMask_lo_2};
  wire [15:0]        executeByteMask = (sew1H[0] ? maskSplit_0_1 : 16'h0) | (sew1H[1] ? maskSplit_1_1 : 16'h0) | (sew1H[2] ? maskSplit_2_1 : 16'h0);
  wire [15:0]        _executeElementMask_T_3 = sew1H[0] ? maskSplit_0_2 : 16'h0;
  wire [7:0]         _GEN_52 = _executeElementMask_T_3[7:0] | (sew1H[1] ? maskSplit_1_2 : 8'h0);
  wire [15:0]        executeElementMask = {_executeElementMask_T_3[15:8], _GEN_52[7:4], _GEN_52[3:0] | (sew1H[2] ? maskSplit_2_2 : 4'h0)};
  wire [127:0]       maskForDestination_lo_lo_lo_lo = {maskForDestination_lo_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_lo_hi = {maskForDestination_lo_lo_lo_hi_hi, maskForDestination_lo_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_lo = {maskForDestination_lo_lo_lo_hi, maskForDestination_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_lo = {maskForDestination_lo_lo_hi_lo_hi, maskForDestination_lo_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_lo_hi_hi = {maskForDestination_lo_lo_hi_hi_hi, maskForDestination_lo_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_lo_hi = {maskForDestination_lo_lo_hi_hi, maskForDestination_lo_lo_hi_lo};
  wire [511:0]       maskForDestination_lo_lo = {maskForDestination_lo_lo_hi, maskForDestination_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_lo = {maskForDestination_lo_hi_lo_lo_hi, maskForDestination_lo_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_lo_hi = {maskForDestination_lo_hi_lo_hi_hi, maskForDestination_lo_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_lo = {maskForDestination_lo_hi_lo_hi, maskForDestination_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_lo = {maskForDestination_lo_hi_hi_lo_hi, maskForDestination_lo_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_lo_hi_hi_hi = {maskForDestination_lo_hi_hi_hi_hi, maskForDestination_lo_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_lo_hi_hi = {maskForDestination_lo_hi_hi_hi, maskForDestination_lo_hi_hi_lo};
  wire [511:0]       maskForDestination_lo_hi = {maskForDestination_lo_hi_hi, maskForDestination_lo_hi_lo};
  wire [1023:0]      maskForDestination_lo = {maskForDestination_lo_hi, maskForDestination_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_lo = {maskForDestination_hi_lo_lo_lo_hi, maskForDestination_hi_lo_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_lo_hi = {maskForDestination_hi_lo_lo_hi_hi, maskForDestination_hi_lo_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_lo = {maskForDestination_hi_lo_lo_hi, maskForDestination_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_lo = {maskForDestination_hi_lo_hi_lo_hi, maskForDestination_hi_lo_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_lo_hi_hi = {maskForDestination_hi_lo_hi_hi_hi, maskForDestination_hi_lo_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_lo_hi = {maskForDestination_hi_lo_hi_hi, maskForDestination_hi_lo_hi_lo};
  wire [511:0]       maskForDestination_hi_lo = {maskForDestination_hi_lo_hi, maskForDestination_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_lo = {maskForDestination_hi_hi_lo_lo_hi, maskForDestination_hi_hi_lo_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_lo_hi = {maskForDestination_hi_hi_lo_hi_hi, maskForDestination_hi_hi_lo_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_lo = {maskForDestination_hi_hi_lo_hi, maskForDestination_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_lo = {maskForDestination_hi_hi_hi_lo_hi, maskForDestination_hi_hi_hi_lo_lo};
  wire [127:0]       maskForDestination_hi_hi_hi_hi = {maskForDestination_hi_hi_hi_hi_hi, maskForDestination_hi_hi_hi_hi_lo};
  wire [255:0]       maskForDestination_hi_hi_hi = {maskForDestination_hi_hi_hi_hi, maskForDestination_hi_hi_hi_lo};
  wire [511:0]       maskForDestination_hi_hi = {maskForDestination_hi_hi_hi, maskForDestination_hi_hi_lo};
  wire [1023:0]      maskForDestination_hi = {maskForDestination_hi_hi, maskForDestination_hi_lo};
  wire [127:0]       _lastGroupMask_T = 128'h1 << elementTailForMaskDestination;
  wire [126:0]       _GEN_53 = _lastGroupMask_T[126:0] | _lastGroupMask_T[127:1];
  wire [125:0]       _GEN_54 = _GEN_53[125:0] | {_lastGroupMask_T[127], _GEN_53[126:2]};
  wire [123:0]       _GEN_55 = _GEN_54[123:0] | {_lastGroupMask_T[127], _GEN_53[126], _GEN_54[125:4]};
  wire [119:0]       _GEN_56 = _GEN_55[119:0] | {_lastGroupMask_T[127], _GEN_53[126], _GEN_54[125:124], _GEN_55[123:8]};
  wire [111:0]       _GEN_57 = _GEN_56[111:0] | {_lastGroupMask_T[127], _GEN_53[126], _GEN_54[125:124], _GEN_55[123:120], _GEN_56[119:16]};
  wire [95:0]        _GEN_58 = _GEN_57[95:0] | {_lastGroupMask_T[127], _GEN_53[126], _GEN_54[125:124], _GEN_55[123:120], _GEN_56[119:112], _GEN_57[111:32]};
  wire [127:0]       lastGroupMask =
    {_lastGroupMask_T[127],
     _GEN_53[126],
     _GEN_54[125:124],
     _GEN_55[123:120],
     _GEN_56[119:112],
     _GEN_57[111:96],
     _GEN_58[95:64],
     _GEN_58[63:0] | {_lastGroupMask_T[127], _GEN_53[126], _GEN_54[125:124], _GEN_55[123:120], _GEN_56[119:112], _GEN_57[111:96], _GEN_58[95:64]}};
  wire [15:0][127:0] _GEN_59 =
    {{maskForDestination_hi[1023:896]},
     {maskForDestination_hi[895:768]},
     {maskForDestination_hi[767:640]},
     {maskForDestination_hi[639:512]},
     {maskForDestination_hi[511:384]},
     {maskForDestination_hi[383:256]},
     {maskForDestination_hi[255:128]},
     {maskForDestination_hi[127:0]},
     {maskForDestination_lo[1023:896]},
     {maskForDestination_lo[895:768]},
     {maskForDestination_lo[767:640]},
     {maskForDestination_lo[639:512]},
     {maskForDestination_lo[511:384]},
     {maskForDestination_lo[383:256]},
     {maskForDestination_lo[255:128]},
     {maskForDestination_lo[127:0]}};
  wire [127:0]       currentMaskGroupForDestination =
    (lastGroup ? lastGroupMask : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF) & (instReg_maskType & ~instReg_decodeResult_maskSource ? _GEN_59[requestCounter[3:0]] : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF);
  wire [63:0]        _GEN_60 = {exeReqReg_1_bits_source1, exeReqReg_0_bits_source1};
  wire [63:0]        groupSourceData_lo;
  assign groupSourceData_lo = _GEN_60;
  wire [63:0]        source1_lo;
  assign source1_lo = _GEN_60;
  wire [63:0]        _GEN_61 = {exeReqReg_3_bits_source1, exeReqReg_2_bits_source1};
  wire [63:0]        groupSourceData_hi;
  assign groupSourceData_hi = _GEN_61;
  wire [63:0]        source1_hi;
  assign source1_hi = _GEN_61;
  wire [127:0]       groupSourceData = {groupSourceData_hi, groupSourceData_lo};
  wire [1:0]         _GEN_62 = {exeReqReg_1_valid, exeReqReg_0_valid};
  wire [1:0]         groupSourceValid_lo;
  assign groupSourceValid_lo = _GEN_62;
  wire [1:0]         view__in_bits_validInput_lo;
  assign view__in_bits_validInput_lo = _GEN_62;
  wire [1:0]         view__in_bits_sourceValid_lo;
  assign view__in_bits_sourceValid_lo = _GEN_62;
  wire [1:0]         _GEN_63 = {exeReqReg_3_valid, exeReqReg_2_valid};
  wire [1:0]         groupSourceValid_hi;
  assign groupSourceValid_hi = _GEN_63;
  wire [1:0]         view__in_bits_validInput_hi;
  assign view__in_bits_validInput_hi = _GEN_63;
  wire [1:0]         view__in_bits_sourceValid_hi;
  assign view__in_bits_sourceValid_hi = _GEN_63;
  wire [3:0]         groupSourceValid = {groupSourceValid_hi, groupSourceValid_lo};
  wire [1:0]         shifterSize = (sourceDataEEW1H[0] ? executeIndex : 2'h0) | (sourceDataEEW1H[1] ? {executeIndex[1], 1'h0} : 2'h0);
  wire [3:0]         _shifterSource_T = 4'h1 << shifterSize;
  wire [127:0]       _shifterSource_T_8 = _shifterSource_T[0] ? groupSourceData : 128'h0;
  wire [95:0]        _GEN_64 = _shifterSource_T_8[95:0] | (_shifterSource_T[1] ? groupSourceData[127:32] : 96'h0);
  wire [63:0]        _GEN_65 = _GEN_64[63:0] | (_shifterSource_T[2] ? groupSourceData[127:64] : 64'h0);
  wire [127:0]       shifterSource = {_shifterSource_T_8[127:96], _GEN_64[95:64], _GEN_65[63:32], _GEN_65[31:0] | (_shifterSource_T[3] ? groupSourceData[127:96] : 32'h0)};
  wire [7:0]         selectValid_lo = {{4{groupSourceValid[1]}}, {4{groupSourceValid[0]}}};
  wire [7:0]         selectValid_hi = {{4{groupSourceValid[3]}}, {4{groupSourceValid[2]}}};
  wire [3:0]         selectValid_lo_1 = {{2{groupSourceValid[1]}}, {2{groupSourceValid[0]}}};
  wire [3:0]         selectValid_hi_1 = {{2{groupSourceValid[3]}}, {2{groupSourceValid[2]}}};
  wire [3:0][3:0]    _GEN_66 = {{selectValid_hi[7:4]}, {selectValid_hi[3:0]}, {selectValid_lo[7:4]}, {selectValid_lo[3:0]}};
  wire [3:0]         selectValid = (sourceDataEEW1H[0] ? _GEN_66[executeIndex] : 4'h0) | (sourceDataEEW1H[1] ? (executeIndex[1] ? selectValid_hi_1 : selectValid_lo_1) : 4'h0) | (sourceDataEEW1H[2] ? groupSourceValid : 4'h0);
  wire [31:0]        source_0 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[7:0] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[15:0] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[31:0] : 32'h0);
  wire [31:0]        source_1 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[15:8] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[31:16] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[63:32] : 32'h0);
  wire [31:0]        source_2 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[23:16] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[47:32] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[95:64] : 32'h0);
  wire [31:0]        source_3 = {16'h0, {8'h0, sourceDataEEW1H[0] ? shifterSource[31:24] : 8'h0} | (sourceDataEEW1H[1] ? shifterSource[63:48] : 16'h0)} | (sourceDataEEW1H[2] ? shifterSource[127:96] : 32'h0);
  wire [3:0]         _GEN_67 = selectValid & readMaskCorrection;
  wire [3:0]         checkVec_validVec;
  assign checkVec_validVec = _GEN_67;
  wire [3:0]         checkVec_validVec_1;
  assign checkVec_validVec_1 = _GEN_67;
  wire [3:0]         checkVec_validVec_2;
  assign checkVec_validVec_2 = _GEN_67;
  wire               checkVec_checkResultVec_0_6 = checkVec_validVec[0];
  wire [3:0]         _GEN_68 = 4'h1 << instReg_vlmul[1:0];
  wire [3:0]         checkVec_checkResultVec_intLMULInput;
  assign checkVec_checkResultVec_intLMULInput = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_1;
  assign checkVec_checkResultVec_intLMULInput_1 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_2;
  assign checkVec_checkResultVec_intLMULInput_2 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_3;
  assign checkVec_checkResultVec_intLMULInput_3 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_4;
  assign checkVec_checkResultVec_intLMULInput_4 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_5;
  assign checkVec_checkResultVec_intLMULInput_5 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_6;
  assign checkVec_checkResultVec_intLMULInput_6 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_7;
  assign checkVec_checkResultVec_intLMULInput_7 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_8;
  assign checkVec_checkResultVec_intLMULInput_8 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_9;
  assign checkVec_checkResultVec_intLMULInput_9 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_10;
  assign checkVec_checkResultVec_intLMULInput_10 = _GEN_68;
  wire [3:0]         checkVec_checkResultVec_intLMULInput_11;
  assign checkVec_checkResultVec_intLMULInput_11 = _GEN_68;
  wire [10:0]        checkVec_checkResultVec_dataPosition = source_0[10:0];
  wire [3:0]         checkVec_checkResultVec_0_0 = 4'h1 << checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]         checkVec_checkResultVec_0_1 = checkVec_checkResultVec_dataPosition[1:0];
  wire [1:0]         checkVec_checkResultVec_0_2 = checkVec_checkResultVec_dataPosition[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup = checkVec_checkResultVec_dataPosition[10:4];
  wire [3:0]         checkVec_checkResultVec_0_3 = checkVec_checkResultVec_dataGroup[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth = checkVec_checkResultVec_dataGroup[6:4];
  wire [2:0]         checkVec_checkResultVec_0_4 = checkVec_checkResultVec_accessRegGrowth;
  wire [5:0]         checkVec_checkResultVec_decimalProportion = {checkVec_checkResultVec_0_3, checkVec_checkResultVec_0_2};
  wire [2:0]         checkVec_checkResultVec_decimal = checkVec_checkResultVec_decimalProportion[5:3];
  wire               checkVec_checkResultVec_overlap =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal >= checkVec_checkResultVec_intLMULInput[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth} >= checkVec_checkResultVec_intLMULInput, source_0[31:11]};
  wire               checkVec_checkResultVec_0_5 = checkVec_checkResultVec_overlap | ~checkVec_checkResultVec_0_6;
  wire               checkVec_checkResultVec_1_6 = checkVec_validVec[1];
  wire [10:0]        checkVec_checkResultVec_dataPosition_1 = source_1[10:0];
  wire [3:0]         checkVec_checkResultVec_1_0 = 4'h1 << checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]         checkVec_checkResultVec_1_1 = checkVec_checkResultVec_dataPosition_1[1:0];
  wire [1:0]         checkVec_checkResultVec_1_2 = checkVec_checkResultVec_dataPosition_1[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_1 = checkVec_checkResultVec_dataPosition_1[10:4];
  wire [3:0]         checkVec_checkResultVec_1_3 = checkVec_checkResultVec_dataGroup_1[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_1 = checkVec_checkResultVec_dataGroup_1[6:4];
  wire [2:0]         checkVec_checkResultVec_1_4 = checkVec_checkResultVec_accessRegGrowth_1;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_1 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_1_2};
  wire [2:0]         checkVec_checkResultVec_decimal_1 = checkVec_checkResultVec_decimalProportion_1[5:3];
  wire               checkVec_checkResultVec_overlap_1 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_1 >= checkVec_checkResultVec_intLMULInput_1[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_1} >= checkVec_checkResultVec_intLMULInput_1, source_1[31:11]};
  wire               checkVec_checkResultVec_1_5 = checkVec_checkResultVec_overlap_1 | ~checkVec_checkResultVec_1_6;
  wire               checkVec_checkResultVec_2_6 = checkVec_validVec[2];
  wire [10:0]        checkVec_checkResultVec_dataPosition_2 = source_2[10:0];
  wire [3:0]         checkVec_checkResultVec_2_0 = 4'h1 << checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]         checkVec_checkResultVec_2_1 = checkVec_checkResultVec_dataPosition_2[1:0];
  wire [1:0]         checkVec_checkResultVec_2_2 = checkVec_checkResultVec_dataPosition_2[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_2 = checkVec_checkResultVec_dataPosition_2[10:4];
  wire [3:0]         checkVec_checkResultVec_2_3 = checkVec_checkResultVec_dataGroup_2[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_2 = checkVec_checkResultVec_dataGroup_2[6:4];
  wire [2:0]         checkVec_checkResultVec_2_4 = checkVec_checkResultVec_accessRegGrowth_2;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_2 = {checkVec_checkResultVec_2_3, checkVec_checkResultVec_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_2 = checkVec_checkResultVec_decimalProportion_2[5:3];
  wire               checkVec_checkResultVec_overlap_2 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_2 >= checkVec_checkResultVec_intLMULInput_2[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_2} >= checkVec_checkResultVec_intLMULInput_2, source_2[31:11]};
  wire               checkVec_checkResultVec_2_5 = checkVec_checkResultVec_overlap_2 | ~checkVec_checkResultVec_2_6;
  wire               checkVec_checkResultVec_3_6 = checkVec_validVec[3];
  wire [10:0]        checkVec_checkResultVec_dataPosition_3 = source_3[10:0];
  wire [3:0]         checkVec_checkResultVec_3_0 = 4'h1 << checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]         checkVec_checkResultVec_3_1 = checkVec_checkResultVec_dataPosition_3[1:0];
  wire [1:0]         checkVec_checkResultVec_3_2 = checkVec_checkResultVec_dataPosition_3[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_3 = checkVec_checkResultVec_dataPosition_3[10:4];
  wire [3:0]         checkVec_checkResultVec_3_3 = checkVec_checkResultVec_dataGroup_3[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_3 = checkVec_checkResultVec_dataGroup_3[6:4];
  wire [2:0]         checkVec_checkResultVec_3_4 = checkVec_checkResultVec_accessRegGrowth_3;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_3_2};
  wire [2:0]         checkVec_checkResultVec_decimal_3 = checkVec_checkResultVec_decimalProportion_3[5:3];
  wire               checkVec_checkResultVec_overlap_3 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_3 >= checkVec_checkResultVec_intLMULInput_3[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_3} >= checkVec_checkResultVec_intLMULInput_3, source_3[31:11]};
  wire               checkVec_checkResultVec_3_5 = checkVec_checkResultVec_overlap_3 | ~checkVec_checkResultVec_3_6;
  wire [7:0]         checkVec_checkResult_lo = {checkVec_checkResultVec_1_0, checkVec_checkResultVec_0_0};
  wire [7:0]         checkVec_checkResult_hi = {checkVec_checkResultVec_3_0, checkVec_checkResultVec_2_0};
  wire [15:0]        checkVec_0_0 = {checkVec_checkResult_hi, checkVec_checkResult_lo};
  wire [3:0]         checkVec_checkResult_lo_1 = {checkVec_checkResultVec_1_1, checkVec_checkResultVec_0_1};
  wire [3:0]         checkVec_checkResult_hi_1 = {checkVec_checkResultVec_3_1, checkVec_checkResultVec_2_1};
  wire [7:0]         checkVec_0_1 = {checkVec_checkResult_hi_1, checkVec_checkResult_lo_1};
  wire [3:0]         checkVec_checkResult_lo_2 = {checkVec_checkResultVec_1_2, checkVec_checkResultVec_0_2};
  wire [3:0]         checkVec_checkResult_hi_2 = {checkVec_checkResultVec_3_2, checkVec_checkResultVec_2_2};
  wire [7:0]         checkVec_0_2 = {checkVec_checkResult_hi_2, checkVec_checkResult_lo_2};
  wire [7:0]         checkVec_checkResult_lo_3 = {checkVec_checkResultVec_1_3, checkVec_checkResultVec_0_3};
  wire [7:0]         checkVec_checkResult_hi_3 = {checkVec_checkResultVec_3_3, checkVec_checkResultVec_2_3};
  wire [15:0]        checkVec_0_3 = {checkVec_checkResult_hi_3, checkVec_checkResult_lo_3};
  wire [5:0]         checkVec_checkResult_lo_4 = {checkVec_checkResultVec_1_4, checkVec_checkResultVec_0_4};
  wire [5:0]         checkVec_checkResult_hi_4 = {checkVec_checkResultVec_3_4, checkVec_checkResultVec_2_4};
  wire [11:0]        checkVec_0_4 = {checkVec_checkResult_hi_4, checkVec_checkResult_lo_4};
  wire [1:0]         checkVec_checkResult_lo_5 = {checkVec_checkResultVec_1_5, checkVec_checkResultVec_0_5};
  wire [1:0]         checkVec_checkResult_hi_5 = {checkVec_checkResultVec_3_5, checkVec_checkResultVec_2_5};
  wire [3:0]         checkVec_0_5 = {checkVec_checkResult_hi_5, checkVec_checkResult_lo_5};
  wire [1:0]         checkVec_checkResult_lo_6 = {checkVec_checkResultVec_1_6, checkVec_checkResultVec_0_6};
  wire [1:0]         checkVec_checkResult_hi_6 = {checkVec_checkResultVec_3_6, checkVec_checkResultVec_2_6};
  wire [3:0]         checkVec_0_6 = {checkVec_checkResult_hi_6, checkVec_checkResult_lo_6};
  wire               checkVec_checkResultVec_0_6_1 = checkVec_validVec_1[0];
  wire [10:0]        checkVec_checkResultVec_dataPosition_4 = {source_0[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_35 = 2'h1 << checkVec_checkResultVec_dataPosition_4[1];
  wire [3:0]         checkVec_checkResultVec_0_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_35[1]}}, {2{_checkVec_checkResultVec_accessMask_T_35[0]}}};
  wire [1:0]         checkVec_checkResultVec_0_1_1 = {checkVec_checkResultVec_dataPosition_4[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_0_2_1 = checkVec_checkResultVec_dataPosition_4[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_4 = checkVec_checkResultVec_dataPosition_4[10:4];
  wire [3:0]         checkVec_checkResultVec_0_3_1 = checkVec_checkResultVec_dataGroup_4[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_4 = checkVec_checkResultVec_dataGroup_4[6:4];
  wire [2:0]         checkVec_checkResultVec_0_4_1 = checkVec_checkResultVec_accessRegGrowth_4;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_4 = {checkVec_checkResultVec_0_3_1, checkVec_checkResultVec_0_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_4 = checkVec_checkResultVec_decimalProportion_4[5:3];
  wire               checkVec_checkResultVec_overlap_4 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_4 >= checkVec_checkResultVec_intLMULInput_4[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_4} >= checkVec_checkResultVec_intLMULInput_4, source_0[31:11]};
  wire               checkVec_checkResultVec_0_5_1 = checkVec_checkResultVec_overlap_4 | ~checkVec_checkResultVec_0_6_1;
  wire               checkVec_checkResultVec_1_6_1 = checkVec_validVec_1[1];
  wire [10:0]        checkVec_checkResultVec_dataPosition_5 = {source_1[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_43 = 2'h1 << checkVec_checkResultVec_dataPosition_5[1];
  wire [3:0]         checkVec_checkResultVec_1_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_43[1]}}, {2{_checkVec_checkResultVec_accessMask_T_43[0]}}};
  wire [1:0]         checkVec_checkResultVec_1_1_1 = {checkVec_checkResultVec_dataPosition_5[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_1_2_1 = checkVec_checkResultVec_dataPosition_5[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_5 = checkVec_checkResultVec_dataPosition_5[10:4];
  wire [3:0]         checkVec_checkResultVec_1_3_1 = checkVec_checkResultVec_dataGroup_5[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_5 = checkVec_checkResultVec_dataGroup_5[6:4];
  wire [2:0]         checkVec_checkResultVec_1_4_1 = checkVec_checkResultVec_accessRegGrowth_5;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_5 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_1_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_5 = checkVec_checkResultVec_decimalProportion_5[5:3];
  wire               checkVec_checkResultVec_overlap_5 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_5 >= checkVec_checkResultVec_intLMULInput_5[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_5} >= checkVec_checkResultVec_intLMULInput_5, source_1[31:11]};
  wire               checkVec_checkResultVec_1_5_1 = checkVec_checkResultVec_overlap_5 | ~checkVec_checkResultVec_1_6_1;
  wire               checkVec_checkResultVec_2_6_1 = checkVec_validVec_1[2];
  wire [10:0]        checkVec_checkResultVec_dataPosition_6 = {source_2[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_51 = 2'h1 << checkVec_checkResultVec_dataPosition_6[1];
  wire [3:0]         checkVec_checkResultVec_2_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_51[1]}}, {2{_checkVec_checkResultVec_accessMask_T_51[0]}}};
  wire [1:0]         checkVec_checkResultVec_2_1_1 = {checkVec_checkResultVec_dataPosition_6[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_2_2_1 = checkVec_checkResultVec_dataPosition_6[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_6 = checkVec_checkResultVec_dataPosition_6[10:4];
  wire [3:0]         checkVec_checkResultVec_2_3_1 = checkVec_checkResultVec_dataGroup_6[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_6 = checkVec_checkResultVec_dataGroup_6[6:4];
  wire [2:0]         checkVec_checkResultVec_2_4_1 = checkVec_checkResultVec_accessRegGrowth_6;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_6 = {checkVec_checkResultVec_2_3_1, checkVec_checkResultVec_2_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_6 = checkVec_checkResultVec_decimalProportion_6[5:3];
  wire               checkVec_checkResultVec_overlap_6 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_6 >= checkVec_checkResultVec_intLMULInput_6[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_6} >= checkVec_checkResultVec_intLMULInput_6, source_2[31:11]};
  wire               checkVec_checkResultVec_2_5_1 = checkVec_checkResultVec_overlap_6 | ~checkVec_checkResultVec_2_6_1;
  wire               checkVec_checkResultVec_3_6_1 = checkVec_validVec_1[3];
  wire [10:0]        checkVec_checkResultVec_dataPosition_7 = {source_3[9:0], 1'h0};
  wire [1:0]         _checkVec_checkResultVec_accessMask_T_59 = 2'h1 << checkVec_checkResultVec_dataPosition_7[1];
  wire [3:0]         checkVec_checkResultVec_3_0_1 = {{2{_checkVec_checkResultVec_accessMask_T_59[1]}}, {2{_checkVec_checkResultVec_accessMask_T_59[0]}}};
  wire [1:0]         checkVec_checkResultVec_3_1_1 = {checkVec_checkResultVec_dataPosition_7[1], 1'h0};
  wire [1:0]         checkVec_checkResultVec_3_2_1 = checkVec_checkResultVec_dataPosition_7[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_7 = checkVec_checkResultVec_dataPosition_7[10:4];
  wire [3:0]         checkVec_checkResultVec_3_3_1 = checkVec_checkResultVec_dataGroup_7[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_7 = checkVec_checkResultVec_dataGroup_7[6:4];
  wire [2:0]         checkVec_checkResultVec_3_4_1 = checkVec_checkResultVec_accessRegGrowth_7;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_7 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_3_2_1};
  wire [2:0]         checkVec_checkResultVec_decimal_7 = checkVec_checkResultVec_decimalProportion_7[5:3];
  wire               checkVec_checkResultVec_overlap_7 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_7 >= checkVec_checkResultVec_intLMULInput_7[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_7} >= checkVec_checkResultVec_intLMULInput_7, source_3[31:11]};
  wire               checkVec_checkResultVec_3_5_1 = checkVec_checkResultVec_overlap_7 | ~checkVec_checkResultVec_3_6_1;
  wire [7:0]         checkVec_checkResult_lo_7 = {checkVec_checkResultVec_1_0_1, checkVec_checkResultVec_0_0_1};
  wire [7:0]         checkVec_checkResult_hi_7 = {checkVec_checkResultVec_3_0_1, checkVec_checkResultVec_2_0_1};
  wire [15:0]        checkVec_1_0 = {checkVec_checkResult_hi_7, checkVec_checkResult_lo_7};
  wire [3:0]         checkVec_checkResult_lo_8 = {checkVec_checkResultVec_1_1_1, checkVec_checkResultVec_0_1_1};
  wire [3:0]         checkVec_checkResult_hi_8 = {checkVec_checkResultVec_3_1_1, checkVec_checkResultVec_2_1_1};
  wire [7:0]         checkVec_1_1 = {checkVec_checkResult_hi_8, checkVec_checkResult_lo_8};
  wire [3:0]         checkVec_checkResult_lo_9 = {checkVec_checkResultVec_1_2_1, checkVec_checkResultVec_0_2_1};
  wire [3:0]         checkVec_checkResult_hi_9 = {checkVec_checkResultVec_3_2_1, checkVec_checkResultVec_2_2_1};
  wire [7:0]         checkVec_1_2 = {checkVec_checkResult_hi_9, checkVec_checkResult_lo_9};
  wire [7:0]         checkVec_checkResult_lo_10 = {checkVec_checkResultVec_1_3_1, checkVec_checkResultVec_0_3_1};
  wire [7:0]         checkVec_checkResult_hi_10 = {checkVec_checkResultVec_3_3_1, checkVec_checkResultVec_2_3_1};
  wire [15:0]        checkVec_1_3 = {checkVec_checkResult_hi_10, checkVec_checkResult_lo_10};
  wire [5:0]         checkVec_checkResult_lo_11 = {checkVec_checkResultVec_1_4_1, checkVec_checkResultVec_0_4_1};
  wire [5:0]         checkVec_checkResult_hi_11 = {checkVec_checkResultVec_3_4_1, checkVec_checkResultVec_2_4_1};
  wire [11:0]        checkVec_1_4 = {checkVec_checkResult_hi_11, checkVec_checkResult_lo_11};
  wire [1:0]         checkVec_checkResult_lo_12 = {checkVec_checkResultVec_1_5_1, checkVec_checkResultVec_0_5_1};
  wire [1:0]         checkVec_checkResult_hi_12 = {checkVec_checkResultVec_3_5_1, checkVec_checkResultVec_2_5_1};
  wire [3:0]         checkVec_1_5 = {checkVec_checkResult_hi_12, checkVec_checkResult_lo_12};
  wire [1:0]         checkVec_checkResult_lo_13 = {checkVec_checkResultVec_1_6_1, checkVec_checkResultVec_0_6_1};
  wire [1:0]         checkVec_checkResult_hi_13 = {checkVec_checkResultVec_3_6_1, checkVec_checkResultVec_2_6_1};
  wire [3:0]         checkVec_1_6 = {checkVec_checkResult_hi_13, checkVec_checkResult_lo_13};
  wire               checkVec_checkResultVec_0_6_2 = checkVec_validVec_2[0];
  wire [10:0]        checkVec_checkResultVec_dataPosition_8 = {source_0[8:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_0_2_2 = checkVec_checkResultVec_dataPosition_8[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_8 = checkVec_checkResultVec_dataPosition_8[10:4];
  wire [3:0]         checkVec_checkResultVec_0_3_2 = checkVec_checkResultVec_dataGroup_8[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_8 = checkVec_checkResultVec_dataGroup_8[6:4];
  wire [2:0]         checkVec_checkResultVec_0_4_2 = checkVec_checkResultVec_accessRegGrowth_8;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_8 = {checkVec_checkResultVec_0_3_2, checkVec_checkResultVec_0_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_8 = checkVec_checkResultVec_decimalProportion_8[5:3];
  wire               checkVec_checkResultVec_overlap_8 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_8 >= checkVec_checkResultVec_intLMULInput_8[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_8} >= checkVec_checkResultVec_intLMULInput_8, source_0[31:11]};
  wire               checkVec_checkResultVec_0_5_2 = checkVec_checkResultVec_overlap_8 | ~checkVec_checkResultVec_0_6_2;
  wire               checkVec_checkResultVec_1_6_2 = checkVec_validVec_2[1];
  wire [10:0]        checkVec_checkResultVec_dataPosition_9 = {source_1[8:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_1_2_2 = checkVec_checkResultVec_dataPosition_9[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_9 = checkVec_checkResultVec_dataPosition_9[10:4];
  wire [3:0]         checkVec_checkResultVec_1_3_2 = checkVec_checkResultVec_dataGroup_9[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_9 = checkVec_checkResultVec_dataGroup_9[6:4];
  wire [2:0]         checkVec_checkResultVec_1_4_2 = checkVec_checkResultVec_accessRegGrowth_9;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_9 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_1_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_9 = checkVec_checkResultVec_decimalProportion_9[5:3];
  wire               checkVec_checkResultVec_overlap_9 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_9 >= checkVec_checkResultVec_intLMULInput_9[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_9} >= checkVec_checkResultVec_intLMULInput_9, source_1[31:11]};
  wire               checkVec_checkResultVec_1_5_2 = checkVec_checkResultVec_overlap_9 | ~checkVec_checkResultVec_1_6_2;
  wire               checkVec_checkResultVec_2_6_2 = checkVec_validVec_2[2];
  wire [10:0]        checkVec_checkResultVec_dataPosition_10 = {source_2[8:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_2_2_2 = checkVec_checkResultVec_dataPosition_10[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_10 = checkVec_checkResultVec_dataPosition_10[10:4];
  wire [3:0]         checkVec_checkResultVec_2_3_2 = checkVec_checkResultVec_dataGroup_10[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_10 = checkVec_checkResultVec_dataGroup_10[6:4];
  wire [2:0]         checkVec_checkResultVec_2_4_2 = checkVec_checkResultVec_accessRegGrowth_10;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_10 = {checkVec_checkResultVec_2_3_2, checkVec_checkResultVec_2_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_10 = checkVec_checkResultVec_decimalProportion_10[5:3];
  wire               checkVec_checkResultVec_overlap_10 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_10 >= checkVec_checkResultVec_intLMULInput_10[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_10} >= checkVec_checkResultVec_intLMULInput_10,
      source_2[31:11]};
  wire               checkVec_checkResultVec_2_5_2 = checkVec_checkResultVec_overlap_10 | ~checkVec_checkResultVec_2_6_2;
  wire               checkVec_checkResultVec_3_6_2 = checkVec_validVec_2[3];
  wire [10:0]        checkVec_checkResultVec_dataPosition_11 = {source_3[8:0], 2'h0};
  wire [1:0]         checkVec_checkResultVec_3_2_2 = checkVec_checkResultVec_dataPosition_11[3:2];
  wire [6:0]         checkVec_checkResultVec_dataGroup_11 = checkVec_checkResultVec_dataPosition_11[10:4];
  wire [3:0]         checkVec_checkResultVec_3_3_2 = checkVec_checkResultVec_dataGroup_11[3:0];
  wire [2:0]         checkVec_checkResultVec_accessRegGrowth_11 = checkVec_checkResultVec_dataGroup_11[6:4];
  wire [2:0]         checkVec_checkResultVec_3_4_2 = checkVec_checkResultVec_accessRegGrowth_11;
  wire [5:0]         checkVec_checkResultVec_decimalProportion_11 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_3_2_2};
  wire [2:0]         checkVec_checkResultVec_decimal_11 = checkVec_checkResultVec_decimalProportion_11[5:3];
  wire               checkVec_checkResultVec_overlap_11 =
    |{instReg_vlmul[2] & checkVec_checkResultVec_decimal_11 >= checkVec_checkResultVec_intLMULInput_11[3:1] | ~(instReg_vlmul[2]) & {1'h0, checkVec_checkResultVec_accessRegGrowth_11} >= checkVec_checkResultVec_intLMULInput_11,
      source_3[31:11]};
  wire               checkVec_checkResultVec_3_5_2 = checkVec_checkResultVec_overlap_11 | ~checkVec_checkResultVec_3_6_2;
  wire [3:0]         checkVec_checkResult_lo_16 = {checkVec_checkResultVec_1_2_2, checkVec_checkResultVec_0_2_2};
  wire [3:0]         checkVec_checkResult_hi_16 = {checkVec_checkResultVec_3_2_2, checkVec_checkResultVec_2_2_2};
  wire [7:0]         checkVec_2_2 = {checkVec_checkResult_hi_16, checkVec_checkResult_lo_16};
  wire [7:0]         checkVec_checkResult_lo_17 = {checkVec_checkResultVec_1_3_2, checkVec_checkResultVec_0_3_2};
  wire [7:0]         checkVec_checkResult_hi_17 = {checkVec_checkResultVec_3_3_2, checkVec_checkResultVec_2_3_2};
  wire [15:0]        checkVec_2_3 = {checkVec_checkResult_hi_17, checkVec_checkResult_lo_17};
  wire [5:0]         checkVec_checkResult_lo_18 = {checkVec_checkResultVec_1_4_2, checkVec_checkResultVec_0_4_2};
  wire [5:0]         checkVec_checkResult_hi_18 = {checkVec_checkResultVec_3_4_2, checkVec_checkResultVec_2_4_2};
  wire [11:0]        checkVec_2_4 = {checkVec_checkResult_hi_18, checkVec_checkResult_lo_18};
  wire [1:0]         checkVec_checkResult_lo_19 = {checkVec_checkResultVec_1_5_2, checkVec_checkResultVec_0_5_2};
  wire [1:0]         checkVec_checkResult_hi_19 = {checkVec_checkResultVec_3_5_2, checkVec_checkResultVec_2_5_2};
  wire [3:0]         checkVec_2_5 = {checkVec_checkResult_hi_19, checkVec_checkResult_lo_19};
  wire [1:0]         checkVec_checkResult_lo_20 = {checkVec_checkResultVec_1_6_2, checkVec_checkResultVec_0_6_2};
  wire [1:0]         checkVec_checkResult_hi_20 = {checkVec_checkResultVec_3_6_2, checkVec_checkResultVec_2_6_2};
  wire [3:0]         checkVec_2_6 = {checkVec_checkResult_hi_20, checkVec_checkResult_lo_20};
  wire [7:0]         dataOffsetSelect = (sew1H[0] ? checkVec_0_1 : 8'h0) | (sew1H[1] ? checkVec_1_1 : 8'h0);
  wire [7:0]         accessLaneSelect = (sew1H[0] ? checkVec_0_2 : 8'h0) | (sew1H[1] ? checkVec_1_2 : 8'h0) | (sew1H[2] ? checkVec_2_2 : 8'h0);
  wire [15:0]        offsetSelect = (sew1H[0] ? checkVec_0_3 : 16'h0) | (sew1H[1] ? checkVec_1_3 : 16'h0) | (sew1H[2] ? checkVec_2_3 : 16'h0);
  wire [11:0]        growthSelect = (sew1H[0] ? checkVec_0_4 : 12'h0) | (sew1H[1] ? checkVec_1_4 : 12'h0) | (sew1H[2] ? checkVec_2_4 : 12'h0);
  wire [3:0]         notReadSelect = (sew1H[0] ? checkVec_0_5 : 4'h0) | (sew1H[1] ? checkVec_1_5 : 4'h0) | (sew1H[2] ? checkVec_2_5 : 4'h0);
  wire [3:0]         elementValidSelect = (sew1H[0] ? checkVec_0_6 : 4'h0) | (sew1H[1] ? checkVec_1_6 : 4'h0) | (sew1H[2] ? checkVec_2_6 : 4'h0);
  wire               readTypeRequestDeq;
  wire               waiteStageEnqReady;
  wire               readWaitQueue_deq_valid;
  assign readWaitQueue_deq_valid = ~_readWaitQueue_fifo_empty;
  wire [9:0]         readWaitQueue_dataOut_executeGroup;
  wire [3:0]         readWaitQueue_dataOut_sourceValid;
  wire [3:0]         readWaitQueue_dataOut_replaceVs1;
  wire [3:0]         readWaitQueue_dataOut_needRead;
  wire               readWaitQueue_dataOut_last;
  wire [4:0]         readWaitQueue_dataIn_lo = {readWaitQueue_enq_bits_needRead, readWaitQueue_enq_bits_last};
  wire [13:0]        readWaitQueue_dataIn_hi_hi = {readWaitQueue_enq_bits_executeGroup, readWaitQueue_enq_bits_sourceValid};
  wire [17:0]        readWaitQueue_dataIn_hi = {readWaitQueue_dataIn_hi_hi, readWaitQueue_enq_bits_replaceVs1};
  wire [22:0]        readWaitQueue_dataIn = {readWaitQueue_dataIn_hi, readWaitQueue_dataIn_lo};
  assign readWaitQueue_dataOut_last = _readWaitQueue_fifo_data_out[0];
  assign readWaitQueue_dataOut_needRead = _readWaitQueue_fifo_data_out[4:1];
  assign readWaitQueue_dataOut_replaceVs1 = _readWaitQueue_fifo_data_out[8:5];
  assign readWaitQueue_dataOut_sourceValid = _readWaitQueue_fifo_data_out[12:9];
  assign readWaitQueue_dataOut_executeGroup = _readWaitQueue_fifo_data_out[22:13];
  wire [9:0]         readWaitQueue_deq_bits_executeGroup = readWaitQueue_dataOut_executeGroup;
  wire [3:0]         readWaitQueue_deq_bits_sourceValid = readWaitQueue_dataOut_sourceValid;
  wire [3:0]         readWaitQueue_deq_bits_replaceVs1 = readWaitQueue_dataOut_replaceVs1;
  wire [3:0]         readWaitQueue_deq_bits_needRead = readWaitQueue_dataOut_needRead;
  wire               readWaitQueue_deq_bits_last = readWaitQueue_dataOut_last;
  wire               readWaitQueue_enq_ready = ~_readWaitQueue_fifo_full;
  wire               readWaitQueue_enq_valid;
  wire               readWaitQueue_deq_ready;
  wire               _GEN_69 = lastExecuteGroupDeq | viota;
  assign exeRequestQueue_0_deq_ready = ~exeReqReg_0_valid | _GEN_69;
  assign exeRequestQueue_1_deq_ready = ~exeReqReg_1_valid | _GEN_69;
  assign exeRequestQueue_2_deq_ready = ~exeReqReg_2_valid | _GEN_69;
  assign exeRequestQueue_3_deq_ready = ~exeReqReg_3_valid | _GEN_69;
  wire               isLastExecuteGroup = executeIndex == lastExecuteIndex;
  wire               allDataValid = (exeReqReg_0_valid | ~(groupDataNeed[0])) & (exeReqReg_1_valid | ~(groupDataNeed[1])) & (exeReqReg_2_valid | ~(groupDataNeed[2])) & (exeReqReg_3_valid | ~(groupDataNeed[3]));
  wire               anyDataValid = exeReqReg_0_valid | exeReqReg_1_valid | exeReqReg_2_valid | exeReqReg_3_valid;
  wire               _GEN_70 = compress | mvRd;
  wire               readVs1Valid = (unitType[2] | _GEN_70) & ~readVS1Reg_requestSend | gatherSRead;
  wire [4:0]         readVS1Req_vs = compress ? instReg_vs1 + {4'h0, readVS1Reg_readIndex[6]} : gatherSRead ? instReg_vs1 + {2'h0, gatherGrowth} : instReg_vs1;
  wire [3:0]         readVS1Req_offset = compress ? readVS1Reg_readIndex[5:2] : gatherSRead ? gatherOffset : 4'h0;
  wire [1:0]         readVS1Req_readLane = compress ? readVS1Reg_readIndex[1:0] : gatherSRead ? gatherLane : 2'h0;
  wire [1:0]         readVS1Req_dataOffset = compress | ~gatherSRead ? 2'h0 : gatherDatOffset;
  wire [3:0]         selectExecuteReq_1_bits_offset = readIssueStageState_readOffset[7:4];
  wire [3:0]         selectExecuteReq_2_bits_offset = readIssueStageState_readOffset[11:8];
  wire [3:0]         selectExecuteReq_3_bits_offset = readIssueStageState_readOffset[15:12];
  wire [1:0]         selectExecuteReq_1_bits_dataOffset = readIssueStageState_readDataOffset[3:2];
  wire [1:0]         selectExecuteReq_2_bits_dataOffset = readIssueStageState_readDataOffset[5:4];
  wire [1:0]         selectExecuteReq_3_bits_dataOffset = readIssueStageState_readDataOffset[7:6];
  wire               selectExecuteReq_0_valid = readVs1Valid | readIssueStageValid & ~(readIssueStageState_groupReadState[0]) & readIssueStageState_needRead[0] & readType;
  wire [4:0]         selectExecuteReq_0_bits_vs = readVs1Valid ? readVS1Req_vs : instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_0};
  wire [3:0]         selectExecuteReq_0_bits_offset = readVs1Valid ? readVS1Req_offset : readIssueStageState_readOffset[3:0];
  wire [1:0]         selectExecuteReq_0_bits_readLane = readVs1Valid ? readVS1Req_readLane : readIssueStageState_accessLane_0;
  wire [1:0]         selectExecuteReq_0_bits_dataOffset = readVs1Valid ? readVS1Req_dataOffset : readIssueStageState_readDataOffset[1:0];
  wire               _tokenCheck_T = _readCrossBar_input_0_ready & readCrossBar_input_0_valid;
  wire               pipeReadFire_0 = ~readVs1Valid & _tokenCheck_T;
  wire [4:0]         selectExecuteReq_1_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_1};
  wire               selectExecuteReq_1_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[1]) & readIssueStageState_needRead[1] & readType;
  wire               pipeReadFire_1 = _readCrossBar_input_1_ready & readCrossBar_input_1_valid;
  wire [4:0]         selectExecuteReq_2_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_2};
  wire               selectExecuteReq_2_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[2]) & readIssueStageState_needRead[2] & readType;
  wire               pipeReadFire_2 = _readCrossBar_input_2_ready & readCrossBar_input_2_valid;
  wire [4:0]         selectExecuteReq_3_bits_vs = instReg_vs2 + {2'h0, readIssueStageState_vsGrowth_3};
  wire               selectExecuteReq_3_valid = readIssueStageValid & ~(readIssueStageState_groupReadState[3]) & readIssueStageState_needRead[3] & readType;
  wire               pipeReadFire_3 = _readCrossBar_input_3_ready & readCrossBar_input_3_valid;
  reg  [3:0]         tokenCheck_counter;
  wire [3:0]         tokenCheck_counterChange = _tokenCheck_T ? 4'h1 : 4'hF;
  wire               tokenCheck = ~(tokenCheck_counter[3]);
  assign readCrossBar_input_0_valid = selectExecuteReq_0_valid & tokenCheck;
  reg  [3:0]         tokenCheck_counter_1;
  wire [3:0]         tokenCheck_counterChange_1 = pipeReadFire_1 ? 4'h1 : 4'hF;
  wire               tokenCheck_1 = ~(tokenCheck_counter_1[3]);
  assign readCrossBar_input_1_valid = selectExecuteReq_1_valid & tokenCheck_1;
  reg  [3:0]         tokenCheck_counter_2;
  wire [3:0]         tokenCheck_counterChange_2 = pipeReadFire_2 ? 4'h1 : 4'hF;
  wire               tokenCheck_2 = ~(tokenCheck_counter_2[3]);
  assign readCrossBar_input_2_valid = selectExecuteReq_2_valid & tokenCheck_2;
  reg  [3:0]         tokenCheck_counter_3;
  wire [3:0]         tokenCheck_counterChange_3 = pipeReadFire_3 ? 4'h1 : 4'hF;
  wire               tokenCheck_3 = ~(tokenCheck_counter_3[3]);
  assign readCrossBar_input_3_valid = selectExecuteReq_3_valid & tokenCheck_3;
  wire [1:0]         readFire_lo = {pipeReadFire_1, pipeReadFire_0};
  wire [1:0]         readFire_hi = {pipeReadFire_3, pipeReadFire_2};
  wire [3:0]         readFire = {readFire_hi, readFire_lo};
  wire               anyReadFire = |readFire;
  wire [3:0]         readStateUpdate = readFire | readIssueStageState_groupReadState;
  wire               groupReadFinish = readStateUpdate == readIssueStageState_needRead;
  assign readTypeRequestDeq = anyReadFire & groupReadFinish | readIssueStageValid & readIssueStageState_needRead == 4'h0;
  assign readWaitQueue_enq_valid = readTypeRequestDeq;
  wire [3:0]         compressUnitResultQueue_enq_bits_ffoOutput;
  wire               compressUnitResultQueue_enq_bits_compressValid;
  wire [4:0]         compressUnitResultQueue_dataIn_lo = {compressUnitResultQueue_enq_bits_ffoOutput, compressUnitResultQueue_enq_bits_compressValid};
  wire [127:0]       compressUnitResultQueue_enq_bits_data;
  wire [15:0]        compressUnitResultQueue_enq_bits_mask;
  wire [143:0]       compressUnitResultQueue_dataIn_hi_hi = {compressUnitResultQueue_enq_bits_data, compressUnitResultQueue_enq_bits_mask};
  wire [7:0]         compressUnitResultQueue_enq_bits_groupCounter;
  wire [151:0]       compressUnitResultQueue_dataIn_hi = {compressUnitResultQueue_dataIn_hi_hi, compressUnitResultQueue_enq_bits_groupCounter};
  wire [156:0]       compressUnitResultQueue_dataIn = {compressUnitResultQueue_dataIn_hi, compressUnitResultQueue_dataIn_lo};
  wire               compressUnitResultQueue_dataOut_compressValid = _compressUnitResultQueue_fifo_data_out[0];
  wire [3:0]         compressUnitResultQueue_dataOut_ffoOutput = _compressUnitResultQueue_fifo_data_out[4:1];
  wire [7:0]         compressUnitResultQueue_dataOut_groupCounter = _compressUnitResultQueue_fifo_data_out[12:5];
  wire [15:0]        compressUnitResultQueue_dataOut_mask = _compressUnitResultQueue_fifo_data_out[28:13];
  wire [127:0]       compressUnitResultQueue_dataOut_data = _compressUnitResultQueue_fifo_data_out[156:29];
  wire               compressUnitResultQueue_enq_ready = ~_compressUnitResultQueue_fifo_full;
  wire               compressUnitResultQueue_deq_ready;
  wire               compressUnitResultQueue_enq_valid;
  wire               compressUnitResultQueue_deq_valid = ~_compressUnitResultQueue_fifo_empty | compressUnitResultQueue_enq_valid;
  wire [127:0]       compressUnitResultQueue_deq_bits_data = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_data : compressUnitResultQueue_dataOut_data;
  wire [15:0]        compressUnitResultQueue_deq_bits_mask = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_mask : compressUnitResultQueue_dataOut_mask;
  wire [7:0]         compressUnitResultQueue_deq_bits_groupCounter = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_groupCounter : compressUnitResultQueue_dataOut_groupCounter;
  wire [3:0]         compressUnitResultQueue_deq_bits_ffoOutput = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_ffoOutput : compressUnitResultQueue_dataOut_ffoOutput;
  wire               compressUnitResultQueue_deq_bits_compressValid = _compressUnitResultQueue_fifo_empty ? compressUnitResultQueue_enq_bits_compressValid : compressUnitResultQueue_dataOut_compressValid;
  wire               noSourceValid = noSource & counterValid & ((|instReg_vl) | mvRd & ~readVS1Reg_sendToExecution);
  wire               vs1DataValid = readVS1Reg_dataValid | ~(unitType[2] | _GEN_70);
  wire [1:0]         _GEN_71 = {_maskedWrite_in_1_ready, _maskedWrite_in_0_ready};
  wire [1:0]         executeDeqReady_lo;
  assign executeDeqReady_lo = _GEN_71;
  wire [1:0]         compressUnitResultQueue_deq_ready_lo;
  assign compressUnitResultQueue_deq_ready_lo = _GEN_71;
  wire [1:0]         _GEN_72 = {_maskedWrite_in_3_ready, _maskedWrite_in_2_ready};
  wire [1:0]         executeDeqReady_hi;
  assign executeDeqReady_hi = _GEN_72;
  wire [1:0]         compressUnitResultQueue_deq_ready_hi;
  assign compressUnitResultQueue_deq_ready_hi = _GEN_72;
  wire               compressUnitResultQueue_empty;
  wire               executeDeqReady = (&{executeDeqReady_hi, executeDeqReady_lo}) & compressUnitResultQueue_empty;
  wire               otherTypeRequestDeq = (noSource ? noSourceValid : allDataValid) & vs1DataValid & instVlValid & executeDeqReady;
  wire               reorderQueueAllocate;
  wire               _GEN_73 = accessCountQueue_enq_ready & reorderQueueAllocate;
  assign readIssueStageEnq = (allDataValid | _slideAddressGen_indexDeq_valid) & (readTypeRequestDeq | ~readIssueStageValid) & instVlValid & readType & _GEN_73;
  assign accessCountQueue_enq_valid = readIssueStageEnq;
  wire               executeReady;
  wire               requestStageDeq = readType ? readIssueStageEnq : otherTypeRequestDeq & executeReady;
  wire               slideAddressGen_indexDeq_ready = (readTypeRequestDeq | ~readIssueStageValid) & _GEN_73;
  wire               _GEN_74 = slideAddressGen_indexDeq_ready & _slideAddressGen_indexDeq_valid;
  wire               _GEN_75 = readIssueStageEnq & _GEN_74;
  assign accessCountEnq_0 =
    _GEN_75
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h0 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h0 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h0 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h0 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h0 & ~(notReadSelect[3])}};
  assign accessCountEnq_1 =
    _GEN_75
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h1 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h1 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h1 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h1 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h1 & ~(notReadSelect[3])}};
  assign accessCountEnq_2 =
    _GEN_75
      ? {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_0 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_1 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, _slideAddressGen_indexDeq_bits_accessLane_2 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, _slideAddressGen_indexDeq_bits_accessLane_3 == 2'h2 & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, accessLaneSelect[1:0] == 2'h2 & ~(notReadSelect[0])} + {1'h0, accessLaneSelect[3:2] == 2'h2 & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, accessLaneSelect[5:4] == 2'h2 & ~(notReadSelect[2])} + {1'h0, accessLaneSelect[7:6] == 2'h2 & ~(notReadSelect[3])}};
  assign accessCountEnq_3 =
    _GEN_75
      ? {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_0) & _slideAddressGen_indexDeq_bits_needRead[0]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_1) & _slideAddressGen_indexDeq_bits_needRead[1]}}
        + {1'h0, {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_2) & _slideAddressGen_indexDeq_bits_needRead[2]} + {1'h0, (&_slideAddressGen_indexDeq_bits_accessLane_3) & _slideAddressGen_indexDeq_bits_needRead[3]}}
      : {1'h0, {1'h0, (&(accessLaneSelect[1:0])) & ~(notReadSelect[0])} + {1'h0, (&(accessLaneSelect[3:2])) & ~(notReadSelect[1])}}
        + {1'h0, {1'h0, (&(accessLaneSelect[5:4])) & ~(notReadSelect[2])} + {1'h0, (&(accessLaneSelect[7:6])) & ~(notReadSelect[3])}};
  assign lastExecuteGroupDeq = requestStageDeq & isLastExecuteGroup;
  wire [3:0]         readMessageQueue_deq_bits_readSource;
  wire               deqAllocate;
  wire               reorderQueueVec_0_deq_valid;
  assign reorderQueueVec_0_deq_valid = ~_reorderQueueVec_fifo_empty;
  wire [31:0]        reorderQueueVec_dataOut_data;
  wire [3:0]         reorderQueueVec_dataOut_write1H;
  wire [31:0]        dataAfterReorderCheck_0 = reorderQueueVec_0_deq_bits_data;
  wire [31:0]        reorderQueueVec_0_enq_bits_data;
  wire [3:0]         reorderQueueVec_0_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn = {reorderQueueVec_0_enq_bits_data, reorderQueueVec_0_enq_bits_write1H};
  assign reorderQueueVec_dataOut_write1H = _reorderQueueVec_fifo_data_out[3:0];
  assign reorderQueueVec_dataOut_data = _reorderQueueVec_fifo_data_out[35:4];
  assign reorderQueueVec_0_deq_bits_data = reorderQueueVec_dataOut_data;
  wire [3:0]         reorderQueueVec_0_deq_bits_write1H = reorderQueueVec_dataOut_write1H;
  wire               reorderQueueVec_0_enq_ready = ~_reorderQueueVec_fifo_full;
  wire               reorderQueueVec_0_deq_ready;
  wire [3:0]         readMessageQueue_1_deq_bits_readSource;
  wire               deqAllocate_1;
  wire               reorderQueueVec_1_deq_valid;
  assign reorderQueueVec_1_deq_valid = ~_reorderQueueVec_fifo_1_empty;
  wire [31:0]        reorderQueueVec_dataOut_1_data;
  wire [3:0]         reorderQueueVec_dataOut_1_write1H;
  wire [31:0]        dataAfterReorderCheck_1 = reorderQueueVec_1_deq_bits_data;
  wire [31:0]        reorderQueueVec_1_enq_bits_data;
  wire [3:0]         reorderQueueVec_1_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn_1 = {reorderQueueVec_1_enq_bits_data, reorderQueueVec_1_enq_bits_write1H};
  assign reorderQueueVec_dataOut_1_write1H = _reorderQueueVec_fifo_1_data_out[3:0];
  assign reorderQueueVec_dataOut_1_data = _reorderQueueVec_fifo_1_data_out[35:4];
  assign reorderQueueVec_1_deq_bits_data = reorderQueueVec_dataOut_1_data;
  wire [3:0]         reorderQueueVec_1_deq_bits_write1H = reorderQueueVec_dataOut_1_write1H;
  wire               reorderQueueVec_1_enq_ready = ~_reorderQueueVec_fifo_1_full;
  wire               reorderQueueVec_1_deq_ready;
  wire [3:0]         readMessageQueue_2_deq_bits_readSource;
  wire               deqAllocate_2;
  wire               reorderQueueVec_2_deq_valid;
  assign reorderQueueVec_2_deq_valid = ~_reorderQueueVec_fifo_2_empty;
  wire [31:0]        reorderQueueVec_dataOut_2_data;
  wire [3:0]         reorderQueueVec_dataOut_2_write1H;
  wire [31:0]        dataAfterReorderCheck_2 = reorderQueueVec_2_deq_bits_data;
  wire [31:0]        reorderQueueVec_2_enq_bits_data;
  wire [3:0]         reorderQueueVec_2_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn_2 = {reorderQueueVec_2_enq_bits_data, reorderQueueVec_2_enq_bits_write1H};
  assign reorderQueueVec_dataOut_2_write1H = _reorderQueueVec_fifo_2_data_out[3:0];
  assign reorderQueueVec_dataOut_2_data = _reorderQueueVec_fifo_2_data_out[35:4];
  assign reorderQueueVec_2_deq_bits_data = reorderQueueVec_dataOut_2_data;
  wire [3:0]         reorderQueueVec_2_deq_bits_write1H = reorderQueueVec_dataOut_2_write1H;
  wire               reorderQueueVec_2_enq_ready = ~_reorderQueueVec_fifo_2_full;
  wire               reorderQueueVec_2_deq_ready;
  wire [3:0]         readMessageQueue_3_deq_bits_readSource;
  wire               deqAllocate_3;
  wire               reorderQueueVec_3_deq_valid;
  assign reorderQueueVec_3_deq_valid = ~_reorderQueueVec_fifo_3_empty;
  wire [31:0]        reorderQueueVec_dataOut_3_data;
  wire [3:0]         reorderQueueVec_dataOut_3_write1H;
  wire [31:0]        dataAfterReorderCheck_3 = reorderQueueVec_3_deq_bits_data;
  wire [31:0]        reorderQueueVec_3_enq_bits_data;
  wire [3:0]         reorderQueueVec_3_enq_bits_write1H;
  wire [35:0]        reorderQueueVec_dataIn_3 = {reorderQueueVec_3_enq_bits_data, reorderQueueVec_3_enq_bits_write1H};
  assign reorderQueueVec_dataOut_3_write1H = _reorderQueueVec_fifo_3_data_out[3:0];
  assign reorderQueueVec_dataOut_3_data = _reorderQueueVec_fifo_3_data_out[35:4];
  assign reorderQueueVec_3_deq_bits_data = reorderQueueVec_dataOut_3_data;
  wire [3:0]         reorderQueueVec_3_deq_bits_write1H = reorderQueueVec_dataOut_3_write1H;
  wire               reorderQueueVec_3_enq_ready = ~_reorderQueueVec_fifo_3_full;
  wire               reorderQueueVec_3_deq_ready;
  reg  [3:0]         reorderQueueAllocate_counter;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate;
  wire               _write1HPipe_0_T = reorderQueueVec_0_deq_ready & reorderQueueVec_0_deq_valid;
  wire               reorderQueueAllocate_release = _write1HPipe_0_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate = readIssueStageEnq ? accessCountEnq_0 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate = reorderQueueAllocate_counter + {1'h0, reorderQueueAllocate_allocate} - {3'h0, reorderQueueAllocate_release};
  reg  [3:0]         reorderQueueAllocate_counter_1;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate_1;
  wire               _write1HPipe_1_T = reorderQueueVec_1_deq_ready & reorderQueueVec_1_deq_valid;
  wire               reorderQueueAllocate_release_1 = _write1HPipe_1_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate_1 = readIssueStageEnq ? accessCountEnq_1 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate_1 = reorderQueueAllocate_counter_1 + {1'h0, reorderQueueAllocate_allocate_1} - {3'h0, reorderQueueAllocate_release_1};
  reg  [3:0]         reorderQueueAllocate_counter_2;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate_2;
  wire               _write1HPipe_2_T = reorderQueueVec_2_deq_ready & reorderQueueVec_2_deq_valid;
  wire               reorderQueueAllocate_release_2 = _write1HPipe_2_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate_2 = readIssueStageEnq ? accessCountEnq_2 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate_2 = reorderQueueAllocate_counter_2 + {1'h0, reorderQueueAllocate_allocate_2} - {3'h0, reorderQueueAllocate_release_2};
  reg  [3:0]         reorderQueueAllocate_counter_3;
  reg  [3:0]         reorderQueueAllocate_counterWillUpdate_3;
  wire               _write1HPipe_3_T = reorderQueueVec_3_deq_ready & reorderQueueVec_3_deq_valid;
  wire               reorderQueueAllocate_release_3 = _write1HPipe_3_T & readValid;
  wire [2:0]         reorderQueueAllocate_allocate_3 = readIssueStageEnq ? accessCountEnq_3 : 3'h0;
  wire [3:0]         reorderQueueAllocate_counterUpdate_3 = reorderQueueAllocate_counter_3 + {1'h0, reorderQueueAllocate_allocate_3} - {3'h0, reorderQueueAllocate_release_3};
  assign reorderQueueAllocate = ~(reorderQueueAllocate_counterWillUpdate[3]) & ~(reorderQueueAllocate_counterWillUpdate_1[3]) & ~(reorderQueueAllocate_counterWillUpdate_2[3]) & ~(reorderQueueAllocate_counterWillUpdate_3[3]);
  reg                reorderStageValid;
  reg  [2:0]         reorderStageState_0;
  reg  [2:0]         reorderStageState_1;
  reg  [2:0]         reorderStageState_2;
  reg  [2:0]         reorderStageState_3;
  reg  [2:0]         reorderStageNeed_0;
  reg  [2:0]         reorderStageNeed_1;
  reg  [2:0]         reorderStageNeed_2;
  reg  [2:0]         reorderStageNeed_3;
  wire               stateCheck = reorderStageState_0 == reorderStageNeed_0 & reorderStageState_1 == reorderStageNeed_1 & reorderStageState_2 == reorderStageNeed_2 & reorderStageState_3 == reorderStageNeed_3;
  assign accessCountQueue_deq_ready = ~reorderStageValid | stateCheck;
  wire               reorderStageEnqFire = accessCountQueue_deq_ready & accessCountQueue_deq_valid;
  wire               reorderStageDeqFire = stateCheck & reorderStageValid;
  wire [3:0]         sourceLane;
  wire               readMessageQueue_deq_valid;
  assign readMessageQueue_deq_valid = ~_readMessageQueue_fifo_empty;
  wire [3:0]         readMessageQueue_dataOut_readSource;
  assign reorderQueueVec_0_enq_bits_write1H = readMessageQueue_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_dataOffset;
  wire [3:0]         readMessageQueue_enq_bits_readSource;
  wire [1:0]         readMessageQueue_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn = {readMessageQueue_enq_bits_readSource, readMessageQueue_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_dataOffset = _readMessageQueue_fifo_data_out[1:0];
  assign readMessageQueue_dataOut_readSource = _readMessageQueue_fifo_data_out[5:2];
  assign readMessageQueue_deq_bits_readSource = readMessageQueue_dataOut_readSource;
  wire [1:0]         readMessageQueue_deq_bits_dataOffset = readMessageQueue_dataOut_dataOffset;
  wire               readMessageQueue_enq_ready = ~_readMessageQueue_fifo_full;
  wire               readMessageQueue_enq_valid;
  assign deqAllocate = ~readValid | reorderStageValid & reorderStageState_0 != reorderStageNeed_0;
  assign reorderQueueVec_0_deq_ready = deqAllocate;
  assign sourceLane = 4'h1 << _readCrossBar_output_0_bits_writeIndex;
  assign readMessageQueue_enq_bits_readSource = sourceLane;
  wire               readChannel_0_valid_0 = maskDestinationType ? _maskedWrite_readChannel_0_valid : _readCrossBar_output_0_valid & readMessageQueue_enq_ready;
  wire [4:0]         readChannel_0_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_vs : _readCrossBar_output_0_bits_vs;
  wire [3:0]         readChannel_0_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_0_bits_offset : _readCrossBar_output_0_bits_offset;
  assign readMessageQueue_enq_valid = readChannel_0_ready_0 & readChannel_0_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_0_enq_bits_data = readResult_0_bits >> {27'h0, readMessageQueue_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_0 = _write1HPipe_0_T & ~maskDestinationType ? reorderQueueVec_0_deq_bits_write1H : 4'h0;
  wire [3:0]         sourceLane_1;
  wire               readMessageQueue_1_deq_valid;
  assign readMessageQueue_1_deq_valid = ~_readMessageQueue_fifo_1_empty;
  wire [3:0]         readMessageQueue_dataOut_1_readSource;
  assign reorderQueueVec_1_enq_bits_write1H = readMessageQueue_1_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_1_dataOffset;
  wire [3:0]         readMessageQueue_1_enq_bits_readSource;
  wire [1:0]         readMessageQueue_1_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn_1 = {readMessageQueue_1_enq_bits_readSource, readMessageQueue_1_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_1_dataOffset = _readMessageQueue_fifo_1_data_out[1:0];
  assign readMessageQueue_dataOut_1_readSource = _readMessageQueue_fifo_1_data_out[5:2];
  assign readMessageQueue_1_deq_bits_readSource = readMessageQueue_dataOut_1_readSource;
  wire [1:0]         readMessageQueue_1_deq_bits_dataOffset = readMessageQueue_dataOut_1_dataOffset;
  wire               readMessageQueue_1_enq_ready = ~_readMessageQueue_fifo_1_full;
  wire               readMessageQueue_1_enq_valid;
  assign deqAllocate_1 = ~readValid | reorderStageValid & reorderStageState_1 != reorderStageNeed_1;
  assign reorderQueueVec_1_deq_ready = deqAllocate_1;
  assign sourceLane_1 = 4'h1 << _readCrossBar_output_1_bits_writeIndex;
  assign readMessageQueue_1_enq_bits_readSource = sourceLane_1;
  wire               readChannel_1_valid_0 = maskDestinationType ? _maskedWrite_readChannel_1_valid : _readCrossBar_output_1_valid & readMessageQueue_1_enq_ready;
  wire [4:0]         readChannel_1_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_vs : _readCrossBar_output_1_bits_vs;
  wire [3:0]         readChannel_1_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_1_bits_offset : _readCrossBar_output_1_bits_offset;
  assign readMessageQueue_1_enq_valid = readChannel_1_ready_0 & readChannel_1_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_1_enq_bits_data = readResult_1_bits >> {27'h0, readMessageQueue_1_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_1 = _write1HPipe_1_T & ~maskDestinationType ? reorderQueueVec_1_deq_bits_write1H : 4'h0;
  wire [3:0]         sourceLane_2;
  wire               readMessageQueue_2_deq_valid;
  assign readMessageQueue_2_deq_valid = ~_readMessageQueue_fifo_2_empty;
  wire [3:0]         readMessageQueue_dataOut_2_readSource;
  assign reorderQueueVec_2_enq_bits_write1H = readMessageQueue_2_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_2_dataOffset;
  wire [3:0]         readMessageQueue_2_enq_bits_readSource;
  wire [1:0]         readMessageQueue_2_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn_2 = {readMessageQueue_2_enq_bits_readSource, readMessageQueue_2_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_2_dataOffset = _readMessageQueue_fifo_2_data_out[1:0];
  assign readMessageQueue_dataOut_2_readSource = _readMessageQueue_fifo_2_data_out[5:2];
  assign readMessageQueue_2_deq_bits_readSource = readMessageQueue_dataOut_2_readSource;
  wire [1:0]         readMessageQueue_2_deq_bits_dataOffset = readMessageQueue_dataOut_2_dataOffset;
  wire               readMessageQueue_2_enq_ready = ~_readMessageQueue_fifo_2_full;
  wire               readMessageQueue_2_enq_valid;
  assign deqAllocate_2 = ~readValid | reorderStageValid & reorderStageState_2 != reorderStageNeed_2;
  assign reorderQueueVec_2_deq_ready = deqAllocate_2;
  assign sourceLane_2 = 4'h1 << _readCrossBar_output_2_bits_writeIndex;
  assign readMessageQueue_2_enq_bits_readSource = sourceLane_2;
  wire               readChannel_2_valid_0 = maskDestinationType ? _maskedWrite_readChannel_2_valid : _readCrossBar_output_2_valid & readMessageQueue_2_enq_ready;
  wire [4:0]         readChannel_2_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_vs : _readCrossBar_output_2_bits_vs;
  wire [3:0]         readChannel_2_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_2_bits_offset : _readCrossBar_output_2_bits_offset;
  assign readMessageQueue_2_enq_valid = readChannel_2_ready_0 & readChannel_2_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_2_enq_bits_data = readResult_2_bits >> {27'h0, readMessageQueue_2_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_2 = _write1HPipe_2_T & ~maskDestinationType ? reorderQueueVec_2_deq_bits_write1H : 4'h0;
  wire [3:0]         sourceLane_3;
  wire               readMessageQueue_3_deq_valid;
  assign readMessageQueue_3_deq_valid = ~_readMessageQueue_fifo_3_empty;
  wire [3:0]         readMessageQueue_dataOut_3_readSource;
  assign reorderQueueVec_3_enq_bits_write1H = readMessageQueue_3_deq_bits_readSource;
  wire [1:0]         readMessageQueue_dataOut_3_dataOffset;
  wire [3:0]         readMessageQueue_3_enq_bits_readSource;
  wire [1:0]         readMessageQueue_3_enq_bits_dataOffset;
  wire [5:0]         readMessageQueue_dataIn_3 = {readMessageQueue_3_enq_bits_readSource, readMessageQueue_3_enq_bits_dataOffset};
  assign readMessageQueue_dataOut_3_dataOffset = _readMessageQueue_fifo_3_data_out[1:0];
  assign readMessageQueue_dataOut_3_readSource = _readMessageQueue_fifo_3_data_out[5:2];
  assign readMessageQueue_3_deq_bits_readSource = readMessageQueue_dataOut_3_readSource;
  wire [1:0]         readMessageQueue_3_deq_bits_dataOffset = readMessageQueue_dataOut_3_dataOffset;
  wire               readMessageQueue_3_enq_ready = ~_readMessageQueue_fifo_3_full;
  wire               readMessageQueue_3_enq_valid;
  assign deqAllocate_3 = ~readValid | reorderStageValid & reorderStageState_3 != reorderStageNeed_3;
  assign reorderQueueVec_3_deq_ready = deqAllocate_3;
  assign sourceLane_3 = 4'h1 << _readCrossBar_output_3_bits_writeIndex;
  assign readMessageQueue_3_enq_bits_readSource = sourceLane_3;
  wire               readChannel_3_valid_0 = maskDestinationType ? _maskedWrite_readChannel_3_valid : _readCrossBar_output_3_valid & readMessageQueue_3_enq_ready;
  wire [4:0]         readChannel_3_bits_vs_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_vs : _readCrossBar_output_3_bits_vs;
  wire [3:0]         readChannel_3_bits_offset_0 = maskDestinationType ? _maskedWrite_readChannel_3_bits_offset : _readCrossBar_output_3_bits_offset;
  assign readMessageQueue_3_enq_valid = readChannel_3_ready_0 & readChannel_3_valid_0 & ~maskDestinationType;
  assign reorderQueueVec_3_enq_bits_data = readResult_3_bits >> {27'h0, readMessageQueue_3_deq_bits_dataOffset, 3'h0};
  wire [3:0]         write1HPipe_3 = _write1HPipe_3_T & ~maskDestinationType ? reorderQueueVec_3_deq_bits_write1H : 4'h0;
  wire [31:0]        readData_data;
  wire               readData_readDataQueue_enq_ready = ~_readData_readDataQueue_fifo_full;
  wire               readData_readDataQueue_deq_ready;
  wire               readData_readDataQueue_enq_valid;
  wire               readData_readDataQueue_deq_valid = ~_readData_readDataQueue_fifo_empty | readData_readDataQueue_enq_valid;
  wire [31:0]        readData_readDataQueue_enq_bits;
  wire [31:0]        readData_readDataQueue_deq_bits = _readData_readDataQueue_fifo_empty ? readData_readDataQueue_enq_bits : _readData_readDataQueue_fifo_data_out;
  wire [1:0]         readData_readResultSelect_lo = {write1HPipe_1[0], write1HPipe_0[0]};
  wire [1:0]         readData_readResultSelect_hi = {write1HPipe_3[0], write1HPipe_2[0]};
  wire [3:0]         readData_readResultSelect = {readData_readResultSelect_hi, readData_readResultSelect_lo};
  assign readData_data =
    (readData_readResultSelect[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_enq_bits = readData_data;
  wire               readTokenRelease_0 = readData_readDataQueue_deq_ready & readData_readDataQueue_deq_valid;
  assign readData_readDataQueue_enq_valid = |readData_readResultSelect;
  wire [31:0]        readData_data_1;
  wire               isWaiteForThisData_1;
  wire               readData_readDataQueue_1_enq_ready = ~_readData_readDataQueue_fifo_1_full;
  wire               readData_readDataQueue_1_deq_ready;
  wire               readData_readDataQueue_1_enq_valid;
  wire               readData_readDataQueue_1_deq_valid = ~_readData_readDataQueue_fifo_1_empty | readData_readDataQueue_1_enq_valid;
  wire [31:0]        readData_readDataQueue_1_enq_bits;
  wire [31:0]        readData_readDataQueue_1_deq_bits = _readData_readDataQueue_fifo_1_empty ? readData_readDataQueue_1_enq_bits : _readData_readDataQueue_fifo_1_data_out;
  wire [1:0]         readData_readResultSelect_lo_1 = {write1HPipe_1[1], write1HPipe_0[1]};
  wire [1:0]         readData_readResultSelect_hi_1 = {write1HPipe_3[1], write1HPipe_2[1]};
  wire [3:0]         readData_readResultSelect_1 = {readData_readResultSelect_hi_1, readData_readResultSelect_lo_1};
  assign readData_data_1 =
    (readData_readResultSelect_1[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_1[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_1[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_1[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_1_enq_bits = readData_data_1;
  wire               readTokenRelease_1 = readData_readDataQueue_1_deq_ready & readData_readDataQueue_1_deq_valid;
  assign readData_readDataQueue_1_enq_valid = |readData_readResultSelect_1;
  wire [31:0]        readData_data_2;
  wire               isWaiteForThisData_2;
  wire               readData_readDataQueue_2_enq_ready = ~_readData_readDataQueue_fifo_2_full;
  wire               readData_readDataQueue_2_deq_ready;
  wire               readData_readDataQueue_2_enq_valid;
  wire               readData_readDataQueue_2_deq_valid = ~_readData_readDataQueue_fifo_2_empty | readData_readDataQueue_2_enq_valid;
  wire [31:0]        readData_readDataQueue_2_enq_bits;
  wire [31:0]        readData_readDataQueue_2_deq_bits = _readData_readDataQueue_fifo_2_empty ? readData_readDataQueue_2_enq_bits : _readData_readDataQueue_fifo_2_data_out;
  wire [1:0]         readData_readResultSelect_lo_2 = {write1HPipe_1[2], write1HPipe_0[2]};
  wire [1:0]         readData_readResultSelect_hi_2 = {write1HPipe_3[2], write1HPipe_2[2]};
  wire [3:0]         readData_readResultSelect_2 = {readData_readResultSelect_hi_2, readData_readResultSelect_lo_2};
  assign readData_data_2 =
    (readData_readResultSelect_2[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_2[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_2[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_2[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_2_enq_bits = readData_data_2;
  wire               readTokenRelease_2 = readData_readDataQueue_2_deq_ready & readData_readDataQueue_2_deq_valid;
  assign readData_readDataQueue_2_enq_valid = |readData_readResultSelect_2;
  wire [31:0]        readData_data_3;
  wire               isWaiteForThisData_3;
  wire               readData_readDataQueue_3_enq_ready = ~_readData_readDataQueue_fifo_3_full;
  wire               readData_readDataQueue_3_deq_ready;
  wire               readData_readDataQueue_3_enq_valid;
  wire               readData_readDataQueue_3_deq_valid = ~_readData_readDataQueue_fifo_3_empty | readData_readDataQueue_3_enq_valid;
  wire [31:0]        readData_readDataQueue_3_enq_bits;
  wire [31:0]        readData_readDataQueue_3_deq_bits = _readData_readDataQueue_fifo_3_empty ? readData_readDataQueue_3_enq_bits : _readData_readDataQueue_fifo_3_data_out;
  wire [1:0]         readData_readResultSelect_lo_3 = {write1HPipe_1[3], write1HPipe_0[3]};
  wire [1:0]         readData_readResultSelect_hi_3 = {write1HPipe_3[3], write1HPipe_2[3]};
  wire [3:0]         readData_readResultSelect_3 = {readData_readResultSelect_hi_3, readData_readResultSelect_lo_3};
  assign readData_data_3 =
    (readData_readResultSelect_3[0] ? dataAfterReorderCheck_0 : 32'h0) | (readData_readResultSelect_3[1] ? dataAfterReorderCheck_1 : 32'h0) | (readData_readResultSelect_3[2] ? dataAfterReorderCheck_2 : 32'h0)
    | (readData_readResultSelect_3[3] ? dataAfterReorderCheck_3 : 32'h0);
  assign readData_readDataQueue_3_enq_bits = readData_data_3;
  wire               readTokenRelease_3 = readData_readDataQueue_3_deq_ready & readData_readDataQueue_3_deq_valid;
  assign readData_readDataQueue_3_enq_valid = |readData_readResultSelect_3;
  reg  [9:0]         waiteReadDataPipeReg_executeGroup;
  reg  [3:0]         waiteReadDataPipeReg_sourceValid;
  reg  [3:0]         waiteReadDataPipeReg_replaceVs1;
  reg  [3:0]         waiteReadDataPipeReg_needRead;
  reg                waiteReadDataPipeReg_last;
  reg  [31:0]        waiteReadData_0;
  reg  [31:0]        waiteReadData_1;
  reg  [31:0]        waiteReadData_2;
  reg  [31:0]        waiteReadData_3;
  reg  [3:0]         waiteReadSate;
  reg                waiteReadStageValid;
  wire [1:0]         executeIndexVec_0 = waiteReadDataPipeReg_executeGroup[1:0];
  wire [1:0]         executeIndexVec_1 = {waiteReadDataPipeReg_executeGroup[0], 1'h0};
  wire               writeDataVec_data_dataIsRead = waiteReadDataPipeReg_needRead[0];
  wire               writeDataVec_data_dataIsRead_4 = waiteReadDataPipeReg_needRead[0];
  wire               writeDataVec_data_dataIsRead_8 = waiteReadDataPipeReg_needRead[0];
  wire [31:0]        _GEN_76 = waiteReadDataPipeReg_replaceVs1[0] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData;
  assign writeDataVec_data_unreadData = _GEN_76;
  wire [31:0]        writeDataVec_data_unreadData_4;
  assign writeDataVec_data_unreadData_4 = _GEN_76;
  wire [31:0]        writeDataVec_data_unreadData_8;
  assign writeDataVec_data_unreadData_8 = _GEN_76;
  wire [7:0]         writeDataVec_data_dataElement = writeDataVec_data_dataIsRead ? waiteReadData_0[7:0] : writeDataVec_data_unreadData[7:0];
  wire               writeDataVec_data_dataIsRead_1 = waiteReadDataPipeReg_needRead[1];
  wire               writeDataVec_data_dataIsRead_5 = waiteReadDataPipeReg_needRead[1];
  wire               writeDataVec_data_dataIsRead_9 = waiteReadDataPipeReg_needRead[1];
  wire [31:0]        _GEN_77 = waiteReadDataPipeReg_replaceVs1[1] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_1;
  assign writeDataVec_data_unreadData_1 = _GEN_77;
  wire [31:0]        writeDataVec_data_unreadData_5;
  assign writeDataVec_data_unreadData_5 = _GEN_77;
  wire [31:0]        writeDataVec_data_unreadData_9;
  assign writeDataVec_data_unreadData_9 = _GEN_77;
  wire [7:0]         writeDataVec_data_dataElement_1 = writeDataVec_data_dataIsRead_1 ? waiteReadData_1[7:0] : writeDataVec_data_unreadData_1[7:0];
  wire               writeDataVec_data_dataIsRead_2 = waiteReadDataPipeReg_needRead[2];
  wire               writeDataVec_data_dataIsRead_6 = waiteReadDataPipeReg_needRead[2];
  wire               writeDataVec_data_dataIsRead_10 = waiteReadDataPipeReg_needRead[2];
  wire [31:0]        _GEN_78 = waiteReadDataPipeReg_replaceVs1[2] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_2;
  assign writeDataVec_data_unreadData_2 = _GEN_78;
  wire [31:0]        writeDataVec_data_unreadData_6;
  assign writeDataVec_data_unreadData_6 = _GEN_78;
  wire [31:0]        writeDataVec_data_unreadData_10;
  assign writeDataVec_data_unreadData_10 = _GEN_78;
  wire [7:0]         writeDataVec_data_dataElement_2 = writeDataVec_data_dataIsRead_2 ? waiteReadData_2[7:0] : writeDataVec_data_unreadData_2[7:0];
  wire               writeDataVec_data_dataIsRead_3 = waiteReadDataPipeReg_needRead[3];
  wire               writeDataVec_data_dataIsRead_7 = waiteReadDataPipeReg_needRead[3];
  wire               writeDataVec_data_dataIsRead_11 = waiteReadDataPipeReg_needRead[3];
  wire [31:0]        _GEN_79 = waiteReadDataPipeReg_replaceVs1[3] ? instReg_readFromScala : 32'h0;
  wire [31:0]        writeDataVec_data_unreadData_3;
  assign writeDataVec_data_unreadData_3 = _GEN_79;
  wire [31:0]        writeDataVec_data_unreadData_7;
  assign writeDataVec_data_unreadData_7 = _GEN_79;
  wire [31:0]        writeDataVec_data_unreadData_11;
  assign writeDataVec_data_unreadData_11 = _GEN_79;
  wire [7:0]         writeDataVec_data_dataElement_3 = writeDataVec_data_dataIsRead_3 ? waiteReadData_3[7:0] : writeDataVec_data_unreadData_3[7:0];
  wire [15:0]        writeDataVec_data_lo = {writeDataVec_data_dataElement_1, writeDataVec_data_dataElement};
  wire [15:0]        writeDataVec_data_hi = {writeDataVec_data_dataElement_3, writeDataVec_data_dataElement_2};
  wire [31:0]        writeDataVec_data = {writeDataVec_data_hi, writeDataVec_data_lo};
  wire [158:0]       writeDataVec_shifterData = {127'h0, writeDataVec_data} << {152'h0, executeIndexVec_0, 5'h0};
  wire [127:0]       writeDataVec_0 = writeDataVec_shifterData[127:0];
  wire [15:0]        writeDataVec_data_dataElement_4 = writeDataVec_data_dataIsRead_4 ? waiteReadData_0[15:0] : writeDataVec_data_unreadData_4[15:0];
  wire [15:0]        writeDataVec_data_dataElement_5 = writeDataVec_data_dataIsRead_5 ? waiteReadData_1[15:0] : writeDataVec_data_unreadData_5[15:0];
  wire [15:0]        writeDataVec_data_dataElement_6 = writeDataVec_data_dataIsRead_6 ? waiteReadData_2[15:0] : writeDataVec_data_unreadData_6[15:0];
  wire [15:0]        writeDataVec_data_dataElement_7 = writeDataVec_data_dataIsRead_7 ? waiteReadData_3[15:0] : writeDataVec_data_unreadData_7[15:0];
  wire [31:0]        writeDataVec_data_lo_1 = {writeDataVec_data_dataElement_5, writeDataVec_data_dataElement_4};
  wire [31:0]        writeDataVec_data_hi_1 = {writeDataVec_data_dataElement_7, writeDataVec_data_dataElement_6};
  wire [63:0]        writeDataVec_data_1 = {writeDataVec_data_hi_1, writeDataVec_data_lo_1};
  wire [190:0]       writeDataVec_shifterData_1 = {127'h0, writeDataVec_data_1} << {184'h0, executeIndexVec_1, 5'h0};
  wire [127:0]       writeDataVec_1 = writeDataVec_shifterData_1[127:0];
  wire [31:0]        writeDataVec_data_dataElement_8 = writeDataVec_data_dataIsRead_8 ? waiteReadData_0 : writeDataVec_data_unreadData_8;
  wire [31:0]        writeDataVec_data_dataElement_9 = writeDataVec_data_dataIsRead_9 ? waiteReadData_1 : writeDataVec_data_unreadData_9;
  wire [31:0]        writeDataVec_data_dataElement_10 = writeDataVec_data_dataIsRead_10 ? waiteReadData_2 : writeDataVec_data_unreadData_10;
  wire [31:0]        writeDataVec_data_dataElement_11 = writeDataVec_data_dataIsRead_11 ? waiteReadData_3 : writeDataVec_data_unreadData_11;
  wire [63:0]        writeDataVec_data_lo_2 = {writeDataVec_data_dataElement_9, writeDataVec_data_dataElement_8};
  wire [63:0]        writeDataVec_data_hi_2 = {writeDataVec_data_dataElement_11, writeDataVec_data_dataElement_10};
  wire [127:0]       writeDataVec_data_2 = {writeDataVec_data_hi_2, writeDataVec_data_lo_2};
  wire [190:0]       writeDataVec_shifterData_2 = {63'h0, writeDataVec_data_2};
  wire [127:0]       writeDataVec_2 = writeDataVec_shifterData_2[127:0];
  wire [127:0]       writeData = (sew1H[0] ? writeDataVec_0 : 128'h0) | (sew1H[1] ? writeDataVec_1 : 128'h0) | (sew1H[2] ? writeDataVec_2 : 128'h0);
  wire [1:0]         writeMaskVec_mask_lo = waiteReadDataPipeReg_sourceValid[1:0];
  wire [1:0]         writeMaskVec_mask_hi = waiteReadDataPipeReg_sourceValid[3:2];
  wire [3:0]         writeMaskVec_mask = {writeMaskVec_mask_hi, writeMaskVec_mask_lo};
  wire [18:0]        writeMaskVec_shifterMask = {15'h0, writeMaskVec_mask} << {15'h0, executeIndexVec_0, 2'h0};
  wire [15:0]        writeMaskVec_0 = writeMaskVec_shifterMask[15:0];
  wire [3:0]         writeMaskVec_mask_lo_1 = {{2{waiteReadDataPipeReg_sourceValid[1]}}, {2{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [3:0]         writeMaskVec_mask_hi_1 = {{2{waiteReadDataPipeReg_sourceValid[3]}}, {2{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [7:0]         writeMaskVec_mask_1 = {writeMaskVec_mask_hi_1, writeMaskVec_mask_lo_1};
  wire [22:0]        writeMaskVec_shifterMask_1 = {15'h0, writeMaskVec_mask_1} << {19'h0, executeIndexVec_1, 2'h0};
  wire [15:0]        writeMaskVec_1 = writeMaskVec_shifterMask_1[15:0];
  wire [7:0]         writeMaskVec_mask_lo_2 = {{4{waiteReadDataPipeReg_sourceValid[1]}}, {4{waiteReadDataPipeReg_sourceValid[0]}}};
  wire [7:0]         writeMaskVec_mask_hi_2 = {{4{waiteReadDataPipeReg_sourceValid[3]}}, {4{waiteReadDataPipeReg_sourceValid[2]}}};
  wire [15:0]        writeMaskVec_mask_2 = {writeMaskVec_mask_hi_2, writeMaskVec_mask_lo_2};
  wire [22:0]        writeMaskVec_shifterMask_2 = {7'h0, writeMaskVec_mask_2};
  wire [15:0]        writeMaskVec_2 = writeMaskVec_shifterMask_2[15:0];
  wire [15:0]        writeMask = (sew1H[0] ? writeMaskVec_0 : 16'h0) | (sew1H[1] ? writeMaskVec_1 : 16'h0) | (sew1H[2] ? writeMaskVec_2 : 16'h0);
  wire [12:0]        _writeRequest_res_writeData_groupCounter_T_6 = {3'h0, waiteReadDataPipeReg_executeGroup} << instReg_sew;
  wire [7:0]         writeRequest_0_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[9:2];
  wire [7:0]         writeRequest_1_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[9:2];
  wire [7:0]         writeRequest_2_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[9:2];
  wire [7:0]         writeRequest_3_writeData_groupCounter = _writeRequest_res_writeData_groupCounter_T_6[9:2];
  wire [31:0]        writeRequest_0_writeData_data = writeData[31:0];
  wire [31:0]        writeRequest_1_writeData_data = writeData[63:32];
  wire [31:0]        writeRequest_2_writeData_data = writeData[95:64];
  wire [31:0]        writeRequest_3_writeData_data = writeData[127:96];
  wire [3:0]         writeRequest_0_writeData_mask = writeMask[3:0];
  wire [3:0]         writeRequest_1_writeData_mask = writeMask[7:4];
  wire [3:0]         writeRequest_2_writeData_mask = writeMask[11:8];
  wire [3:0]         writeRequest_3_writeData_mask = writeMask[15:12];
  wire [1:0]         WillWriteLane_lo = {|writeRequest_1_writeData_mask, |writeRequest_0_writeData_mask};
  wire [1:0]         WillWriteLane_hi = {|writeRequest_3_writeData_mask, |writeRequest_2_writeData_mask};
  wire [3:0]         WillWriteLane = {WillWriteLane_hi, WillWriteLane_lo};
  wire               waiteStageDeqValid = waiteReadStageValid & (waiteReadSate == waiteReadDataPipeReg_needRead | waiteReadDataPipeReg_needRead == 4'h0);
  wire               waiteStageDeqReady;
  wire               waiteStageDeqFire = waiteStageDeqValid & waiteStageDeqReady;
  assign waiteStageEnqReady = ~waiteReadStageValid | waiteStageDeqFire;
  assign readWaitQueue_deq_ready = waiteStageEnqReady;
  wire               waiteStageEnqFire = readWaitQueue_deq_valid & waiteStageEnqReady;
  wire               isWaiteForThisData = waiteReadDataPipeReg_needRead[0] & ~(waiteReadSate[0]) & waiteReadStageValid;
  assign readData_readDataQueue_deq_ready = isWaiteForThisData | unitType[2] | compress | gatherWaiteRead | mvRd;
  assign isWaiteForThisData_1 = waiteReadDataPipeReg_needRead[1] & ~(waiteReadSate[1]) & waiteReadStageValid;
  assign readData_readDataQueue_1_deq_ready = isWaiteForThisData_1;
  assign isWaiteForThisData_2 = waiteReadDataPipeReg_needRead[2] & ~(waiteReadSate[2]) & waiteReadStageValid;
  assign readData_readDataQueue_2_deq_ready = isWaiteForThisData_2;
  assign isWaiteForThisData_3 = waiteReadDataPipeReg_needRead[3] & ~(waiteReadSate[3]) & waiteReadStageValid;
  assign readData_readDataQueue_3_deq_ready = isWaiteForThisData_3;
  wire [1:0]         readResultValid_lo = {readTokenRelease_1, readTokenRelease_0};
  wire [1:0]         readResultValid_hi = {readTokenRelease_3, readTokenRelease_2};
  wire [3:0]         readResultValid = {readResultValid_hi, readResultValid_lo};
  wire               executeEnqValid = otherTypeRequestDeq & ~readType;
  wire [63:0]        source2_lo = {exeReqReg_1_bits_source2, exeReqReg_0_bits_source2};
  wire [63:0]        source2_hi = {exeReqReg_3_bits_source2, exeReqReg_2_bits_source2};
  wire [127:0]       source2 = {source2_hi, source2_lo};
  wire [127:0]       source1 = {source1_hi, source1_lo};
  wire               vs1Split_vs1SetIndex = requestCounter[0];
  wire               vs1Split_0_2 = vs1Split_vs1SetIndex;
  wire [1:0]         vs1Split_vs1SetIndex_1 = requestCounter[1:0];
  wire               vs1Split_1_2 = &vs1Split_vs1SetIndex_1;
  wire [2:0]         vs1Split_vs1SetIndex_2 = requestCounter[2:0];
  wire               vs1Split_2_2 = &vs1Split_vs1SetIndex_2;
  wire [15:0]        _compressSource1_T_3 = sew1H[0] ? (vs1Split_vs1SetIndex ? readVS1Reg_data[31:16] : readVS1Reg_data[15:0]) : 16'h0;
  wire [3:0][7:0]    _GEN_80 = {{readVS1Reg_data[31:24]}, {readVS1Reg_data[23:16]}, {readVS1Reg_data[15:8]}, {readVS1Reg_data[7:0]}};
  wire [7:0][3:0]    _GEN_84 = {{readVS1Reg_data[31:28]}, {readVS1Reg_data[27:24]}, {readVS1Reg_data[23:20]}, {readVS1Reg_data[19:16]}, {readVS1Reg_data[15:12]}, {readVS1Reg_data[11:8]}, {readVS1Reg_data[7:4]}, {readVS1Reg_data[3:0]}};
  wire [7:0]         _GEN_85 = _compressSource1_T_3[7:0] | (sew1H[1] ? _GEN_80[vs1Split_vs1SetIndex_1] : 8'h0);
  wire [15:0]        compressSource1 = {_compressSource1_T_3[15:8], _GEN_85[7:4], _GEN_85[3:0] | (sew1H[2] ? _GEN_84[vs1Split_vs1SetIndex_2] : 4'h0)};
  wire [31:0]        source1Select = mv ? readVS1Reg_data : {16'h0, compressSource1};
  wire               source1Change = sew1H[0] & vs1Split_0_2 | sew1H[1] & vs1Split_1_2 | sew1H[2] & vs1Split_2_2;
  assign viotaCounterAdd = executeEnqValid & unitType[1];
  wire [1:0]         view__in_bits_ffoInput_lo = {exeReqReg_1_bits_ffo, exeReqReg_0_bits_ffo};
  wire [1:0]         view__in_bits_ffoInput_hi = {exeReqReg_3_bits_ffo, exeReqReg_2_bits_ffo};
  wire               reduceUnit_in_valid = executeEnqValid & unitType[2];
  wire               _view__firstGroup_T_1 = _reduceUnit_in_ready & reduceUnit_in_valid;
  wire [9:0]         extendGroupCount = extendType ? (subType[2] ? _extendGroupCount_T_1 : {1'h0, requestCounter, executeIndex[1]}) : {2'h0, requestCounter};
  wire [127:0]       _executeResult_T_4 = unitType[1] ? compressUnitResultQueue_deq_bits_data : 128'h0;
  wire [127:0]       executeResult = {_executeResult_T_4[127:32], _executeResult_T_4[31:0] | (unitType[2] ? _reduceUnit_out_bits_data : 32'h0)} | (unitType[3] ? _extendUnit_out : 128'h0);
  assign executeReady = readType | unitType[1] | unitType[2] & _reduceUnit_in_ready & readVS1Reg_dataValid | unitType[3] & executeEnqValid;
  assign compressUnitResultQueue_deq_ready = &{compressUnitResultQueue_deq_ready_hi, compressUnitResultQueue_deq_ready_lo};
  wire               compressDeq = compressUnitResultQueue_deq_ready & compressUnitResultQueue_deq_valid;
  wire               executeValid = unitType[1] & compressDeq | unitType[3] & executeEnqValid;
  assign executeGroupCounter = (unitType[1] | unitType[2] ? requestCounter : 8'h0) | (unitType[3] ? extendGroupCount[7:0] : 8'h0);
  wire [9:0]         executeDeqGroupCounter = {2'h0, (unitType[1] ? compressUnitResultQueue_deq_bits_groupCounter : 8'h0) | (unitType[2] ? requestCounter : 8'h0)} | (unitType[3] ? extendGroupCount : 10'h0);
  wire [15:0]        executeWriteByteMask = compress | ffo | mvVd ? compressUnitResultQueue_deq_bits_mask : executeByteMask;
  wire               maskFilter = |{~maskDestinationType, currentMaskGroupForDestination[31:0]};
  wire               maskFilter_1 = |{~maskDestinationType, currentMaskGroupForDestination[63:32]};
  wire               maskFilter_2 = |{~maskDestinationType, currentMaskGroupForDestination[95:64]};
  wire               maskFilter_3 = |{~maskDestinationType, currentMaskGroupForDestination[127:96]};
  assign writeQueue_0_deq_valid = ~_writeQueue_fifo_empty;
  wire               exeResp_0_valid_0 = writeQueue_0_deq_valid;
  wire               writeQueue_dataOut_ffoByOther;
  wire [31:0]        writeQueue_dataOut_writeData_data;
  wire [31:0]        exeResp_0_bits_data_0 = writeQueue_0_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_writeData_mask;
  wire [3:0]         exeResp_0_bits_mask_0 = writeQueue_0_deq_bits_writeData_mask;
  wire [7:0]         writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_writeData_vd;
  wire [2:0]         writeQueue_dataOut_index;
  wire [7:0]         writeQueue_0_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_0_enq_bits_writeData_vd;
  wire [12:0]        writeQueue_dataIn_lo = {writeQueue_0_enq_bits_writeData_groupCounter, writeQueue_0_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_0_enq_bits_writeData_data;
  wire [3:0]         writeQueue_0_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi = {writeQueue_0_enq_bits_writeData_data, writeQueue_0_enq_bits_writeData_mask};
  wire               writeQueue_0_enq_bits_ffoByOther;
  wire [49:0]        writeQueue_dataIn_hi_1 = {writeQueue_0_enq_bits_ffoByOther, writeQueue_dataIn_hi, writeQueue_dataIn_lo};
  wire [52:0]        writeQueue_dataIn = {writeQueue_dataIn_hi_1, writeQueue_0_enq_bits_index};
  assign writeQueue_dataOut_index = _writeQueue_fifo_data_out[2:0];
  assign writeQueue_dataOut_writeData_vd = _writeQueue_fifo_data_out[7:3];
  assign writeQueue_dataOut_writeData_groupCounter = _writeQueue_fifo_data_out[15:8];
  assign writeQueue_dataOut_writeData_mask = _writeQueue_fifo_data_out[19:16];
  assign writeQueue_dataOut_writeData_data = _writeQueue_fifo_data_out[51:20];
  assign writeQueue_dataOut_ffoByOther = _writeQueue_fifo_data_out[52];
  wire               writeQueue_0_deq_bits_ffoByOther = writeQueue_dataOut_ffoByOther;
  assign writeQueue_0_deq_bits_writeData_data = writeQueue_dataOut_writeData_data;
  assign writeQueue_0_deq_bits_writeData_mask = writeQueue_dataOut_writeData_mask;
  wire [7:0]         writeQueue_0_deq_bits_writeData_groupCounter = writeQueue_dataOut_writeData_groupCounter;
  wire [4:0]         writeQueue_0_deq_bits_writeData_vd = writeQueue_dataOut_writeData_vd;
  wire [2:0]         writeQueue_0_deq_bits_index = writeQueue_dataOut_index;
  wire               writeQueue_0_enq_ready = ~_writeQueue_fifo_full;
  wire               writeQueue_0_enq_valid;
  assign writeQueue_1_deq_valid = ~_writeQueue_fifo_1_empty;
  wire               exeResp_1_valid_0 = writeQueue_1_deq_valid;
  wire               writeQueue_dataOut_1_ffoByOther;
  wire [31:0]        writeQueue_dataOut_1_writeData_data;
  wire [31:0]        exeResp_1_bits_data_0 = writeQueue_1_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_1_writeData_mask;
  wire [3:0]         exeResp_1_bits_mask_0 = writeQueue_1_deq_bits_writeData_mask;
  wire [7:0]         writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_1_writeData_vd;
  wire [2:0]         writeQueue_dataOut_1_index;
  wire [7:0]         writeQueue_1_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_1_enq_bits_writeData_vd;
  wire [12:0]        writeQueue_dataIn_lo_1 = {writeQueue_1_enq_bits_writeData_groupCounter, writeQueue_1_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_1_enq_bits_writeData_data;
  wire [3:0]         writeQueue_1_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_2 = {writeQueue_1_enq_bits_writeData_data, writeQueue_1_enq_bits_writeData_mask};
  wire               writeQueue_1_enq_bits_ffoByOther;
  wire [49:0]        writeQueue_dataIn_hi_3 = {writeQueue_1_enq_bits_ffoByOther, writeQueue_dataIn_hi_2, writeQueue_dataIn_lo_1};
  wire [52:0]        writeQueue_dataIn_1 = {writeQueue_dataIn_hi_3, writeQueue_1_enq_bits_index};
  assign writeQueue_dataOut_1_index = _writeQueue_fifo_1_data_out[2:0];
  assign writeQueue_dataOut_1_writeData_vd = _writeQueue_fifo_1_data_out[7:3];
  assign writeQueue_dataOut_1_writeData_groupCounter = _writeQueue_fifo_1_data_out[15:8];
  assign writeQueue_dataOut_1_writeData_mask = _writeQueue_fifo_1_data_out[19:16];
  assign writeQueue_dataOut_1_writeData_data = _writeQueue_fifo_1_data_out[51:20];
  assign writeQueue_dataOut_1_ffoByOther = _writeQueue_fifo_1_data_out[52];
  wire               writeQueue_1_deq_bits_ffoByOther = writeQueue_dataOut_1_ffoByOther;
  assign writeQueue_1_deq_bits_writeData_data = writeQueue_dataOut_1_writeData_data;
  assign writeQueue_1_deq_bits_writeData_mask = writeQueue_dataOut_1_writeData_mask;
  wire [7:0]         writeQueue_1_deq_bits_writeData_groupCounter = writeQueue_dataOut_1_writeData_groupCounter;
  wire [4:0]         writeQueue_1_deq_bits_writeData_vd = writeQueue_dataOut_1_writeData_vd;
  wire [2:0]         writeQueue_1_deq_bits_index = writeQueue_dataOut_1_index;
  wire               writeQueue_1_enq_ready = ~_writeQueue_fifo_1_full;
  wire               writeQueue_1_enq_valid;
  assign writeQueue_2_deq_valid = ~_writeQueue_fifo_2_empty;
  wire               exeResp_2_valid_0 = writeQueue_2_deq_valid;
  wire               writeQueue_dataOut_2_ffoByOther;
  wire [31:0]        writeQueue_dataOut_2_writeData_data;
  wire [31:0]        exeResp_2_bits_data_0 = writeQueue_2_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_2_writeData_mask;
  wire [3:0]         exeResp_2_bits_mask_0 = writeQueue_2_deq_bits_writeData_mask;
  wire [7:0]         writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_2_writeData_vd;
  wire [2:0]         writeQueue_dataOut_2_index;
  wire [7:0]         writeQueue_2_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_2_enq_bits_writeData_vd;
  wire [12:0]        writeQueue_dataIn_lo_2 = {writeQueue_2_enq_bits_writeData_groupCounter, writeQueue_2_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_2_enq_bits_writeData_data;
  wire [3:0]         writeQueue_2_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_4 = {writeQueue_2_enq_bits_writeData_data, writeQueue_2_enq_bits_writeData_mask};
  wire               writeQueue_2_enq_bits_ffoByOther;
  wire [49:0]        writeQueue_dataIn_hi_5 = {writeQueue_2_enq_bits_ffoByOther, writeQueue_dataIn_hi_4, writeQueue_dataIn_lo_2};
  wire [52:0]        writeQueue_dataIn_2 = {writeQueue_dataIn_hi_5, writeQueue_2_enq_bits_index};
  assign writeQueue_dataOut_2_index = _writeQueue_fifo_2_data_out[2:0];
  assign writeQueue_dataOut_2_writeData_vd = _writeQueue_fifo_2_data_out[7:3];
  assign writeQueue_dataOut_2_writeData_groupCounter = _writeQueue_fifo_2_data_out[15:8];
  assign writeQueue_dataOut_2_writeData_mask = _writeQueue_fifo_2_data_out[19:16];
  assign writeQueue_dataOut_2_writeData_data = _writeQueue_fifo_2_data_out[51:20];
  assign writeQueue_dataOut_2_ffoByOther = _writeQueue_fifo_2_data_out[52];
  wire               writeQueue_2_deq_bits_ffoByOther = writeQueue_dataOut_2_ffoByOther;
  assign writeQueue_2_deq_bits_writeData_data = writeQueue_dataOut_2_writeData_data;
  assign writeQueue_2_deq_bits_writeData_mask = writeQueue_dataOut_2_writeData_mask;
  wire [7:0]         writeQueue_2_deq_bits_writeData_groupCounter = writeQueue_dataOut_2_writeData_groupCounter;
  wire [4:0]         writeQueue_2_deq_bits_writeData_vd = writeQueue_dataOut_2_writeData_vd;
  wire [2:0]         writeQueue_2_deq_bits_index = writeQueue_dataOut_2_index;
  wire               writeQueue_2_enq_ready = ~_writeQueue_fifo_2_full;
  wire               writeQueue_2_enq_valid;
  assign writeQueue_3_deq_valid = ~_writeQueue_fifo_3_empty;
  wire               exeResp_3_valid_0 = writeQueue_3_deq_valid;
  wire               writeQueue_dataOut_3_ffoByOther;
  wire [31:0]        writeQueue_dataOut_3_writeData_data;
  wire [31:0]        exeResp_3_bits_data_0 = writeQueue_3_deq_bits_writeData_data;
  wire [3:0]         writeQueue_dataOut_3_writeData_mask;
  wire [3:0]         exeResp_3_bits_mask_0 = writeQueue_3_deq_bits_writeData_mask;
  wire [7:0]         writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]         writeQueue_dataOut_3_writeData_vd;
  wire [2:0]         writeQueue_dataOut_3_index;
  wire [7:0]         writeQueue_3_enq_bits_writeData_groupCounter;
  wire [4:0]         writeQueue_3_enq_bits_writeData_vd;
  wire [12:0]        writeQueue_dataIn_lo_3 = {writeQueue_3_enq_bits_writeData_groupCounter, writeQueue_3_enq_bits_writeData_vd};
  wire [31:0]        writeQueue_3_enq_bits_writeData_data;
  wire [3:0]         writeQueue_3_enq_bits_writeData_mask;
  wire [35:0]        writeQueue_dataIn_hi_6 = {writeQueue_3_enq_bits_writeData_data, writeQueue_3_enq_bits_writeData_mask};
  wire               writeQueue_3_enq_bits_ffoByOther;
  wire [49:0]        writeQueue_dataIn_hi_7 = {writeQueue_3_enq_bits_ffoByOther, writeQueue_dataIn_hi_6, writeQueue_dataIn_lo_3};
  wire [52:0]        writeQueue_dataIn_3 = {writeQueue_dataIn_hi_7, writeQueue_3_enq_bits_index};
  assign writeQueue_dataOut_3_index = _writeQueue_fifo_3_data_out[2:0];
  assign writeQueue_dataOut_3_writeData_vd = _writeQueue_fifo_3_data_out[7:3];
  assign writeQueue_dataOut_3_writeData_groupCounter = _writeQueue_fifo_3_data_out[15:8];
  assign writeQueue_dataOut_3_writeData_mask = _writeQueue_fifo_3_data_out[19:16];
  assign writeQueue_dataOut_3_writeData_data = _writeQueue_fifo_3_data_out[51:20];
  assign writeQueue_dataOut_3_ffoByOther = _writeQueue_fifo_3_data_out[52];
  wire               writeQueue_3_deq_bits_ffoByOther = writeQueue_dataOut_3_ffoByOther;
  assign writeQueue_3_deq_bits_writeData_data = writeQueue_dataOut_3_writeData_data;
  assign writeQueue_3_deq_bits_writeData_mask = writeQueue_dataOut_3_writeData_mask;
  wire [7:0]         writeQueue_3_deq_bits_writeData_groupCounter = writeQueue_dataOut_3_writeData_groupCounter;
  wire [4:0]         writeQueue_3_deq_bits_writeData_vd = writeQueue_dataOut_3_writeData_vd;
  wire [2:0]         writeQueue_3_deq_bits_index = writeQueue_dataOut_3_index;
  wire               writeQueue_3_enq_ready = ~_writeQueue_fifo_3_full;
  wire               writeQueue_3_enq_valid;
  wire               dataNotInShifter_readTypeWriteVrf = waiteStageDeqFire & WillWriteLane[0];
  assign writeQueue_0_enq_valid = _maskedWrite_out_0_valid | dataNotInShifter_readTypeWriteVrf;
  assign writeQueue_0_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_vd : 5'h0;
  assign writeQueue_0_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_groupCounter : _maskedWrite_out_0_bits_writeData_groupCounter;
  assign writeQueue_0_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_mask : _maskedWrite_out_0_bits_writeData_mask;
  assign writeQueue_0_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf ? writeRequest_0_writeData_data : _maskedWrite_out_0_bits_writeData_data;
  assign writeQueue_0_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf & _maskedWrite_out_0_bits_ffoByOther;
  wire [4:0]         exeResp_0_bits_vd_0 = instReg_vd + {1'h0, writeQueue_0_deq_bits_writeData_groupCounter[7:4]};
  wire [3:0]         exeResp_0_bits_offset_0 = writeQueue_0_deq_bits_writeData_groupCounter[3:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter;
  wire               _dataNotInShifter_T = exeResp_0_ready_0 & exeResp_0_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange = _dataNotInShifter_T ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_1 = waiteStageDeqFire & WillWriteLane[1];
  assign writeQueue_1_enq_valid = _maskedWrite_out_1_valid | dataNotInShifter_readTypeWriteVrf_1;
  assign writeQueue_1_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_vd : 5'h0;
  assign writeQueue_1_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_groupCounter : _maskedWrite_out_1_bits_writeData_groupCounter;
  assign writeQueue_1_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_mask : _maskedWrite_out_1_bits_writeData_mask;
  assign writeQueue_1_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_1 ? writeRequest_1_writeData_data : _maskedWrite_out_1_bits_writeData_data;
  assign writeQueue_1_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_1 & _maskedWrite_out_1_bits_ffoByOther;
  wire [4:0]         exeResp_1_bits_vd_0 = instReg_vd + {1'h0, writeQueue_1_deq_bits_writeData_groupCounter[7:4]};
  wire [3:0]         exeResp_1_bits_offset_0 = writeQueue_1_deq_bits_writeData_groupCounter[3:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_1;
  wire               _dataNotInShifter_T_3 = exeResp_1_ready_0 & exeResp_1_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_1 = _dataNotInShifter_T_3 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_2 = waiteStageDeqFire & WillWriteLane[2];
  assign writeQueue_2_enq_valid = _maskedWrite_out_2_valid | dataNotInShifter_readTypeWriteVrf_2;
  assign writeQueue_2_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_vd : 5'h0;
  assign writeQueue_2_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_groupCounter : _maskedWrite_out_2_bits_writeData_groupCounter;
  assign writeQueue_2_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_mask : _maskedWrite_out_2_bits_writeData_mask;
  assign writeQueue_2_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_2 ? writeRequest_2_writeData_data : _maskedWrite_out_2_bits_writeData_data;
  assign writeQueue_2_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_2 & _maskedWrite_out_2_bits_ffoByOther;
  wire [4:0]         exeResp_2_bits_vd_0 = instReg_vd + {1'h0, writeQueue_2_deq_bits_writeData_groupCounter[7:4]};
  wire [3:0]         exeResp_2_bits_offset_0 = writeQueue_2_deq_bits_writeData_groupCounter[3:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_2;
  wire               _dataNotInShifter_T_6 = exeResp_2_ready_0 & exeResp_2_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_2 = _dataNotInShifter_T_6 ? 3'h1 : 3'h7;
  wire               dataNotInShifter_readTypeWriteVrf_3 = waiteStageDeqFire & WillWriteLane[3];
  assign writeQueue_3_enq_valid = _maskedWrite_out_3_valid | dataNotInShifter_readTypeWriteVrf_3;
  assign writeQueue_3_enq_bits_writeData_vd = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_vd : 5'h0;
  assign writeQueue_3_enq_bits_writeData_groupCounter = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_groupCounter : _maskedWrite_out_3_bits_writeData_groupCounter;
  assign writeQueue_3_enq_bits_writeData_mask = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_mask : _maskedWrite_out_3_bits_writeData_mask;
  assign writeQueue_3_enq_bits_writeData_data = dataNotInShifter_readTypeWriteVrf_3 ? writeRequest_3_writeData_data : _maskedWrite_out_3_bits_writeData_data;
  assign writeQueue_3_enq_bits_ffoByOther = ~dataNotInShifter_readTypeWriteVrf_3 & _maskedWrite_out_3_bits_ffoByOther;
  wire [4:0]         exeResp_3_bits_vd_0 = instReg_vd + {1'h0, writeQueue_3_deq_bits_writeData_groupCounter[7:4]};
  wire [3:0]         exeResp_3_bits_offset_0 = writeQueue_3_deq_bits_writeData_groupCounter[3:0];
  reg  [2:0]         dataNotInShifter_writeTokenCounter_3;
  wire               _dataNotInShifter_T_9 = exeResp_3_ready_0 & exeResp_3_valid_0;
  wire [2:0]         dataNotInShifter_writeTokenChange_3 = _dataNotInShifter_T_9 ? 3'h1 : 3'h7;
  wire               dataNotInShifter = dataNotInShifter_writeTokenCounter == 3'h0 & dataNotInShifter_writeTokenCounter_1 == 3'h0 & dataNotInShifter_writeTokenCounter_2 == 3'h0 & dataNotInShifter_writeTokenCounter_3 == 3'h0;
  assign waiteStageDeqReady = (~(WillWriteLane[0]) | writeQueue_0_enq_ready) & (~(WillWriteLane[1]) | writeQueue_1_enq_ready) & (~(WillWriteLane[2]) | writeQueue_2_enq_ready) & (~(WillWriteLane[3]) | writeQueue_3_enq_ready);
  reg                waiteLastRequest;
  reg                waitQueueClear;
  wire               lastReportValid = waitQueueClear & ~(writeQueue_0_deq_valid | writeQueue_1_deq_valid | writeQueue_2_deq_valid | writeQueue_3_deq_valid) & dataNotInShifter;
  wire               executeStageInvalid = unitType[1] & ~compressUnitResultQueue_deq_valid & ~_compressUnit_stageValid | unitType[2] & _reduceUnit_in_ready | unitType[3];
  wire               executeStageClean = readType ? waiteStageDeqFire & waiteReadDataPipeReg_last : waiteLastRequest & _maskedWrite_stageClear & executeStageInvalid;
  wire               invalidEnq = instReq_valid & instReq_bits_vl == 12'h0 & ~enqMvRD;
  wire [7:0]         _lastReport_output = lastReportValid ? 8'h1 << instReg_instructionIndex : 8'h0;
  wire [31:0]        gatherData_bits_0 = readVS1Reg_dataValid ? readVS1Reg_data : 32'h0;
  always @(posedge clock) begin
    if (reset) begin
      v0_0 <= 32'h0;
      v0_1 <= 32'h0;
      v0_2 <= 32'h0;
      v0_3 <= 32'h0;
      v0_4 <= 32'h0;
      v0_5 <= 32'h0;
      v0_6 <= 32'h0;
      v0_7 <= 32'h0;
      v0_8 <= 32'h0;
      v0_9 <= 32'h0;
      v0_10 <= 32'h0;
      v0_11 <= 32'h0;
      v0_12 <= 32'h0;
      v0_13 <= 32'h0;
      v0_14 <= 32'h0;
      v0_15 <= 32'h0;
      v0_16 <= 32'h0;
      v0_17 <= 32'h0;
      v0_18 <= 32'h0;
      v0_19 <= 32'h0;
      v0_20 <= 32'h0;
      v0_21 <= 32'h0;
      v0_22 <= 32'h0;
      v0_23 <= 32'h0;
      v0_24 <= 32'h0;
      v0_25 <= 32'h0;
      v0_26 <= 32'h0;
      v0_27 <= 32'h0;
      v0_28 <= 32'h0;
      v0_29 <= 32'h0;
      v0_30 <= 32'h0;
      v0_31 <= 32'h0;
      v0_32 <= 32'h0;
      v0_33 <= 32'h0;
      v0_34 <= 32'h0;
      v0_35 <= 32'h0;
      v0_36 <= 32'h0;
      v0_37 <= 32'h0;
      v0_38 <= 32'h0;
      v0_39 <= 32'h0;
      v0_40 <= 32'h0;
      v0_41 <= 32'h0;
      v0_42 <= 32'h0;
      v0_43 <= 32'h0;
      v0_44 <= 32'h0;
      v0_45 <= 32'h0;
      v0_46 <= 32'h0;
      v0_47 <= 32'h0;
      v0_48 <= 32'h0;
      v0_49 <= 32'h0;
      v0_50 <= 32'h0;
      v0_51 <= 32'h0;
      v0_52 <= 32'h0;
      v0_53 <= 32'h0;
      v0_54 <= 32'h0;
      v0_55 <= 32'h0;
      v0_56 <= 32'h0;
      v0_57 <= 32'h0;
      v0_58 <= 32'h0;
      v0_59 <= 32'h0;
      v0_60 <= 32'h0;
      v0_61 <= 32'h0;
      v0_62 <= 32'h0;
      v0_63 <= 32'h0;
      gatherReadState <= 2'h0;
      gatherDatOffset <= 2'h0;
      gatherLane <= 2'h0;
      gatherOffset <= 4'h0;
      gatherGrowth <= 3'h0;
      instReg_instructionIndex <= 3'h0;
      instReg_decodeResult_specialSlot <= 1'h0;
      instReg_decodeResult_topUop <= 5'h0;
      instReg_decodeResult_popCount <= 1'h0;
      instReg_decodeResult_ffo <= 1'h0;
      instReg_decodeResult_average <= 1'h0;
      instReg_decodeResult_reverse <= 1'h0;
      instReg_decodeResult_dontNeedExecuteInLane <= 1'h0;
      instReg_decodeResult_scheduler <= 1'h0;
      instReg_decodeResult_sReadVD <= 1'h0;
      instReg_decodeResult_vtype <= 1'h0;
      instReg_decodeResult_sWrite <= 1'h0;
      instReg_decodeResult_crossRead <= 1'h0;
      instReg_decodeResult_crossWrite <= 1'h0;
      instReg_decodeResult_maskUnit <= 1'h0;
      instReg_decodeResult_special <= 1'h0;
      instReg_decodeResult_saturate <= 1'h0;
      instReg_decodeResult_vwmacc <= 1'h0;
      instReg_decodeResult_readOnly <= 1'h0;
      instReg_decodeResult_maskSource <= 1'h0;
      instReg_decodeResult_maskDestination <= 1'h0;
      instReg_decodeResult_maskLogic <= 1'h0;
      instReg_decodeResult_uop <= 4'h0;
      instReg_decodeResult_iota <= 1'h0;
      instReg_decodeResult_mv <= 1'h0;
      instReg_decodeResult_extend <= 1'h0;
      instReg_decodeResult_unOrderWrite <= 1'h0;
      instReg_decodeResult_compress <= 1'h0;
      instReg_decodeResult_gather16 <= 1'h0;
      instReg_decodeResult_gather <= 1'h0;
      instReg_decodeResult_slid <= 1'h0;
      instReg_decodeResult_targetRd <= 1'h0;
      instReg_decodeResult_widenReduce <= 1'h0;
      instReg_decodeResult_red <= 1'h0;
      instReg_decodeResult_nr <= 1'h0;
      instReg_decodeResult_itype <= 1'h0;
      instReg_decodeResult_unsigned1 <= 1'h0;
      instReg_decodeResult_unsigned0 <= 1'h0;
      instReg_decodeResult_other <= 1'h0;
      instReg_decodeResult_multiCycle <= 1'h0;
      instReg_decodeResult_divider <= 1'h0;
      instReg_decodeResult_multiplier <= 1'h0;
      instReg_decodeResult_shift <= 1'h0;
      instReg_decodeResult_adder <= 1'h0;
      instReg_decodeResult_logic <= 1'h0;
      instReg_readFromScala <= 32'h0;
      instReg_sew <= 2'h0;
      instReg_vlmul <= 3'h0;
      instReg_maskType <= 1'h0;
      instReg_vxrm <= 3'h0;
      instReg_vs2 <= 5'h0;
      instReg_vs1 <= 5'h0;
      instReg_vd <= 5'h0;
      instReg_vl <= 12'h0;
      instVlValid <= 1'h0;
      readVS1Reg_dataValid <= 1'h0;
      readVS1Reg_requestSend <= 1'h0;
      readVS1Reg_sendToExecution <= 1'h0;
      readVS1Reg_data <= 32'h0;
      readVS1Reg_readIndex <= 7'h0;
      exeReqReg_0_valid <= 1'h0;
      exeReqReg_0_bits_source1 <= 32'h0;
      exeReqReg_0_bits_source2 <= 32'h0;
      exeReqReg_0_bits_index <= 3'h0;
      exeReqReg_0_bits_ffo <= 1'h0;
      exeReqReg_1_valid <= 1'h0;
      exeReqReg_1_bits_source1 <= 32'h0;
      exeReqReg_1_bits_source2 <= 32'h0;
      exeReqReg_1_bits_index <= 3'h0;
      exeReqReg_1_bits_ffo <= 1'h0;
      exeReqReg_2_valid <= 1'h0;
      exeReqReg_2_bits_source1 <= 32'h0;
      exeReqReg_2_bits_source2 <= 32'h0;
      exeReqReg_2_bits_index <= 3'h0;
      exeReqReg_2_bits_ffo <= 1'h0;
      exeReqReg_3_valid <= 1'h0;
      exeReqReg_3_bits_source1 <= 32'h0;
      exeReqReg_3_bits_source2 <= 32'h0;
      exeReqReg_3_bits_index <= 3'h0;
      exeReqReg_3_bits_ffo <= 1'h0;
      requestCounter <= 8'h0;
      executeIndex <= 2'h0;
      readIssueStageState_groupReadState <= 4'h0;
      readIssueStageState_needRead <= 4'h0;
      readIssueStageState_elementValid <= 4'h0;
      readIssueStageState_replaceVs1 <= 4'h0;
      readIssueStageState_readOffset <= 16'h0;
      readIssueStageState_accessLane_0 <= 2'h0;
      readIssueStageState_accessLane_1 <= 2'h0;
      readIssueStageState_accessLane_2 <= 2'h0;
      readIssueStageState_accessLane_3 <= 2'h0;
      readIssueStageState_vsGrowth_0 <= 3'h0;
      readIssueStageState_vsGrowth_1 <= 3'h0;
      readIssueStageState_vsGrowth_2 <= 3'h0;
      readIssueStageState_vsGrowth_3 <= 3'h0;
      readIssueStageState_executeGroup <= 10'h0;
      readIssueStageState_readDataOffset <= 8'h0;
      readIssueStageState_last <= 1'h0;
      readIssueStageValid <= 1'h0;
      tokenCheck_counter <= 4'h0;
      tokenCheck_counter_1 <= 4'h0;
      tokenCheck_counter_2 <= 4'h0;
      tokenCheck_counter_3 <= 4'h0;
      reorderQueueAllocate_counter <= 4'h0;
      reorderQueueAllocate_counterWillUpdate <= 4'h0;
      reorderQueueAllocate_counter_1 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_1 <= 4'h0;
      reorderQueueAllocate_counter_2 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_2 <= 4'h0;
      reorderQueueAllocate_counter_3 <= 4'h0;
      reorderQueueAllocate_counterWillUpdate_3 <= 4'h0;
      reorderStageValid <= 1'h0;
      reorderStageState_0 <= 3'h0;
      reorderStageState_1 <= 3'h0;
      reorderStageState_2 <= 3'h0;
      reorderStageState_3 <= 3'h0;
      reorderStageNeed_0 <= 3'h0;
      reorderStageNeed_1 <= 3'h0;
      reorderStageNeed_2 <= 3'h0;
      reorderStageNeed_3 <= 3'h0;
      waiteReadDataPipeReg_executeGroup <= 10'h0;
      waiteReadDataPipeReg_sourceValid <= 4'h0;
      waiteReadDataPipeReg_replaceVs1 <= 4'h0;
      waiteReadDataPipeReg_needRead <= 4'h0;
      waiteReadDataPipeReg_last <= 1'h0;
      waiteReadData_0 <= 32'h0;
      waiteReadData_1 <= 32'h0;
      waiteReadData_2 <= 32'h0;
      waiteReadData_3 <= 32'h0;
      waiteReadSate <= 4'h0;
      waiteReadStageValid <= 1'h0;
      dataNotInShifter_writeTokenCounter <= 3'h0;
      dataNotInShifter_writeTokenCounter_1 <= 3'h0;
      dataNotInShifter_writeTokenCounter_2 <= 3'h0;
      dataNotInShifter_writeTokenCounter_3 <= 3'h0;
      waiteLastRequest <= 1'h0;
      waitQueueClear <= 1'h0;
    end
    else begin
      automatic logic _GEN_81 = instReq_valid & (viotaReq | enqMvRD) | gatherRequestFire;
      automatic logic _GEN_82;
      automatic logic _GEN_83 = source1Change & viotaCounterAdd;
      _GEN_82 = instReq_valid | gatherRequestFire;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h0)
        v0_0 <= v0_0 & ~maskExt | maskExt & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h0)
        v0_1 <= v0_1 & ~maskExt_1 | maskExt_1 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h0)
        v0_2 <= v0_2 & ~maskExt_2 | maskExt_2 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h0)
        v0_3 <= v0_3 & ~maskExt_3 | maskExt_3 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h1)
        v0_4 <= v0_4 & ~maskExt_4 | maskExt_4 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h1)
        v0_5 <= v0_5 & ~maskExt_5 | maskExt_5 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h1)
        v0_6 <= v0_6 & ~maskExt_6 | maskExt_6 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h1)
        v0_7 <= v0_7 & ~maskExt_7 | maskExt_7 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h2)
        v0_8 <= v0_8 & ~maskExt_8 | maskExt_8 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h2)
        v0_9 <= v0_9 & ~maskExt_9 | maskExt_9 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h2)
        v0_10 <= v0_10 & ~maskExt_10 | maskExt_10 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h2)
        v0_11 <= v0_11 & ~maskExt_11 | maskExt_11 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h3)
        v0_12 <= v0_12 & ~maskExt_12 | maskExt_12 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h3)
        v0_13 <= v0_13 & ~maskExt_13 | maskExt_13 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h3)
        v0_14 <= v0_14 & ~maskExt_14 | maskExt_14 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h3)
        v0_15 <= v0_15 & ~maskExt_15 | maskExt_15 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h4)
        v0_16 <= v0_16 & ~maskExt_16 | maskExt_16 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h4)
        v0_17 <= v0_17 & ~maskExt_17 | maskExt_17 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h4)
        v0_18 <= v0_18 & ~maskExt_18 | maskExt_18 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h4)
        v0_19 <= v0_19 & ~maskExt_19 | maskExt_19 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h5)
        v0_20 <= v0_20 & ~maskExt_20 | maskExt_20 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h5)
        v0_21 <= v0_21 & ~maskExt_21 | maskExt_21 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h5)
        v0_22 <= v0_22 & ~maskExt_22 | maskExt_22 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h5)
        v0_23 <= v0_23 & ~maskExt_23 | maskExt_23 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h6)
        v0_24 <= v0_24 & ~maskExt_24 | maskExt_24 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h6)
        v0_25 <= v0_25 & ~maskExt_25 | maskExt_25 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h6)
        v0_26 <= v0_26 & ~maskExt_26 | maskExt_26 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h6)
        v0_27 <= v0_27 & ~maskExt_27 | maskExt_27 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h7)
        v0_28 <= v0_28 & ~maskExt_28 | maskExt_28 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h7)
        v0_29 <= v0_29 & ~maskExt_29 | maskExt_29 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h7)
        v0_30 <= v0_30 & ~maskExt_30 | maskExt_30 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h7)
        v0_31 <= v0_31 & ~maskExt_31 | maskExt_31 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h8)
        v0_32 <= v0_32 & ~maskExt_32 | maskExt_32 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h8)
        v0_33 <= v0_33 & ~maskExt_33 | maskExt_33 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h8)
        v0_34 <= v0_34 & ~maskExt_34 | maskExt_34 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h8)
        v0_35 <= v0_35 & ~maskExt_35 | maskExt_35 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'h9)
        v0_36 <= v0_36 & ~maskExt_36 | maskExt_36 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'h9)
        v0_37 <= v0_37 & ~maskExt_37 | maskExt_37 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'h9)
        v0_38 <= v0_38 & ~maskExt_38 | maskExt_38 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'h9)
        v0_39 <= v0_39 & ~maskExt_39 | maskExt_39 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'hA)
        v0_40 <= v0_40 & ~maskExt_40 | maskExt_40 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'hA)
        v0_41 <= v0_41 & ~maskExt_41 | maskExt_41 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'hA)
        v0_42 <= v0_42 & ~maskExt_42 | maskExt_42 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'hA)
        v0_43 <= v0_43 & ~maskExt_43 | maskExt_43 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'hB)
        v0_44 <= v0_44 & ~maskExt_44 | maskExt_44 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'hB)
        v0_45 <= v0_45 & ~maskExt_45 | maskExt_45 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'hB)
        v0_46 <= v0_46 & ~maskExt_46 | maskExt_46 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'hB)
        v0_47 <= v0_47 & ~maskExt_47 | maskExt_47 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'hC)
        v0_48 <= v0_48 & ~maskExt_48 | maskExt_48 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'hC)
        v0_49 <= v0_49 & ~maskExt_49 | maskExt_49 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'hC)
        v0_50 <= v0_50 & ~maskExt_50 | maskExt_50 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'hC)
        v0_51 <= v0_51 & ~maskExt_51 | maskExt_51 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'hD)
        v0_52 <= v0_52 & ~maskExt_52 | maskExt_52 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'hD)
        v0_53 <= v0_53 & ~maskExt_53 | maskExt_53 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'hD)
        v0_54 <= v0_54 & ~maskExt_54 | maskExt_54 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'hD)
        v0_55 <= v0_55 & ~maskExt_55 | maskExt_55 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & v0UpdateVec_0_bits_offset == 4'hE)
        v0_56 <= v0_56 & ~maskExt_56 | maskExt_56 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & v0UpdateVec_1_bits_offset == 4'hE)
        v0_57 <= v0_57 & ~maskExt_57 | maskExt_57 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & v0UpdateVec_2_bits_offset == 4'hE)
        v0_58 <= v0_58 & ~maskExt_58 | maskExt_58 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & v0UpdateVec_3_bits_offset == 4'hE)
        v0_59 <= v0_59 & ~maskExt_59 | maskExt_59 & v0UpdateVec_3_bits_data;
      if (v0UpdateVec_0_valid & (&v0UpdateVec_0_bits_offset))
        v0_60 <= v0_60 & ~maskExt_60 | maskExt_60 & v0UpdateVec_0_bits_data;
      if (v0UpdateVec_1_valid & (&v0UpdateVec_1_bits_offset))
        v0_61 <= v0_61 & ~maskExt_61 | maskExt_61 & v0UpdateVec_1_bits_data;
      if (v0UpdateVec_2_valid & (&v0UpdateVec_2_bits_offset))
        v0_62 <= v0_62 & ~maskExt_62 | maskExt_62 & v0UpdateVec_2_bits_data;
      if (v0UpdateVec_3_valid & (&v0UpdateVec_3_bits_offset))
        v0_63 <= v0_63 & ~maskExt_63 | maskExt_63 & v0UpdateVec_3_bits_data;
      if (gatherData_ready_0 & gatherData_valid_0)
        gatherReadState <= 2'h0;
      else if (_tokenCheck_T & gatherSRead)
        gatherReadState <= 2'h2;
      else if (gatherRequestFire)
        gatherReadState <= {notNeedRead, 1'h1};
      else if (readTokenRelease_0 & gatherWaiteRead)
        gatherReadState <= 2'h3;
      if (gatherRequestFire) begin
        gatherDatOffset <= dataOffset;
        gatherLane <= accessLane;
        gatherOffset <= offset;
        gatherGrowth <= reallyGrowth;
      end
      if (_GEN_81 | instReq_valid)
        instReg_instructionIndex <= instReq_bits_instructionIndex;
      if (instReq_valid) begin
        instReg_decodeResult_specialSlot <= instReq_bits_decodeResult_specialSlot;
        instReg_decodeResult_topUop <= instReq_bits_decodeResult_topUop;
        instReg_decodeResult_popCount <= instReq_bits_decodeResult_popCount;
        instReg_decodeResult_ffo <= instReq_bits_decodeResult_ffo;
        instReg_decodeResult_average <= instReq_bits_decodeResult_average;
        instReg_decodeResult_reverse <= instReq_bits_decodeResult_reverse;
        instReg_decodeResult_dontNeedExecuteInLane <= instReq_bits_decodeResult_dontNeedExecuteInLane;
        instReg_decodeResult_scheduler <= instReq_bits_decodeResult_scheduler;
        instReg_decodeResult_sReadVD <= instReq_bits_decodeResult_sReadVD;
        instReg_decodeResult_vtype <= instReq_bits_decodeResult_vtype;
        instReg_decodeResult_sWrite <= instReq_bits_decodeResult_sWrite;
        instReg_decodeResult_crossRead <= instReq_bits_decodeResult_crossRead;
        instReg_decodeResult_crossWrite <= instReq_bits_decodeResult_crossWrite;
        instReg_decodeResult_maskUnit <= instReq_bits_decodeResult_maskUnit;
        instReg_decodeResult_special <= instReq_bits_decodeResult_special;
        instReg_decodeResult_saturate <= instReq_bits_decodeResult_saturate;
        instReg_decodeResult_vwmacc <= instReq_bits_decodeResult_vwmacc;
        instReg_decodeResult_readOnly <= instReq_bits_decodeResult_readOnly;
        instReg_decodeResult_maskSource <= instReq_bits_decodeResult_maskSource;
        instReg_decodeResult_maskDestination <= instReq_bits_decodeResult_maskDestination;
        instReg_decodeResult_maskLogic <= instReq_bits_decodeResult_maskLogic;
        instReg_decodeResult_uop <= instReq_bits_decodeResult_uop;
        instReg_decodeResult_iota <= instReq_bits_decodeResult_iota;
        instReg_decodeResult_mv <= instReq_bits_decodeResult_mv;
        instReg_decodeResult_extend <= instReq_bits_decodeResult_extend;
        instReg_decodeResult_unOrderWrite <= instReq_bits_decodeResult_unOrderWrite;
        instReg_decodeResult_compress <= instReq_bits_decodeResult_compress;
        instReg_decodeResult_gather16 <= instReq_bits_decodeResult_gather16;
        instReg_decodeResult_gather <= instReq_bits_decodeResult_gather;
        instReg_decodeResult_slid <= instReq_bits_decodeResult_slid;
        instReg_decodeResult_targetRd <= instReq_bits_decodeResult_targetRd;
        instReg_decodeResult_widenReduce <= instReq_bits_decodeResult_widenReduce;
        instReg_decodeResult_red <= instReq_bits_decodeResult_red;
        instReg_decodeResult_nr <= instReq_bits_decodeResult_nr;
        instReg_decodeResult_itype <= instReq_bits_decodeResult_itype;
        instReg_decodeResult_unsigned1 <= instReq_bits_decodeResult_unsigned1;
        instReg_decodeResult_unsigned0 <= instReq_bits_decodeResult_unsigned0;
        instReg_decodeResult_other <= instReq_bits_decodeResult_other;
        instReg_decodeResult_multiCycle <= instReq_bits_decodeResult_multiCycle;
        instReg_decodeResult_divider <= instReq_bits_decodeResult_divider;
        instReg_decodeResult_multiplier <= instReq_bits_decodeResult_multiplier;
        instReg_decodeResult_shift <= instReq_bits_decodeResult_shift;
        instReg_decodeResult_adder <= instReq_bits_decodeResult_adder;
        instReg_decodeResult_logic <= instReq_bits_decodeResult_logic;
        instReg_readFromScala <= instReq_bits_readFromScala;
        instReg_sew <= instReq_bits_sew;
        instReg_vlmul <= instReq_bits_vlmul;
        instReg_maskType <= instReq_bits_maskType;
        instReg_vxrm <= instReq_bits_vxrm;
        instReg_vs2 <= instReq_bits_vs2;
        instReg_vd <= instReq_bits_vd;
        instReg_vl <= instReq_bits_vl;
      end
      if (_GEN_81)
        instReg_vs1 <= instReq_bits_vs2;
      else if (instReq_valid)
        instReg_vs1 <= instReq_bits_vs1;
      if (|{instReq_valid, _lastReport_output})
        instVlValid <= ((|instReq_bits_vl) | enqMvRD) & instReq_valid;
      readVS1Reg_dataValid <= ~_GEN_83 & (readTokenRelease_0 | ~_GEN_82 & readVS1Reg_dataValid);
      readVS1Reg_requestSend <= ~_GEN_83 & (_tokenCheck_T | ~_GEN_82 & readVS1Reg_requestSend);
      readVS1Reg_sendToExecution <= _view__firstGroup_T_1 | viotaCounterAdd | ~_GEN_82 & readVS1Reg_sendToExecution;
      if (readTokenRelease_0) begin
        readVS1Reg_data <= readData_readDataQueue_deq_bits;
        waiteReadData_0 <= readData_readDataQueue_deq_bits;
      end
      if (_GEN_83)
        readVS1Reg_readIndex <= readVS1Reg_readIndex + 7'h1;
      else if (_GEN_82)
        readVS1Reg_readIndex <= 7'h0;
      if (tokenIO_0_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_0_valid <= tokenIO_0_maskRequestRelease_0 & ~viota;
      if (tokenIO_0_maskRequestRelease_0) begin
        exeReqReg_0_bits_source1 <= exeRequestQueue_0_deq_bits_source1;
        exeReqReg_0_bits_source2 <= exeRequestQueue_0_deq_bits_source2;
        exeReqReg_0_bits_index <= exeRequestQueue_0_deq_bits_index;
        exeReqReg_0_bits_ffo <= exeRequestQueue_0_deq_bits_ffo;
      end
      if (tokenIO_1_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_1_valid <= tokenIO_1_maskRequestRelease_0 & ~viota;
      if (tokenIO_1_maskRequestRelease_0) begin
        exeReqReg_1_bits_source1 <= exeRequestQueue_1_deq_bits_source1;
        exeReqReg_1_bits_source2 <= exeRequestQueue_1_deq_bits_source2;
        exeReqReg_1_bits_index <= exeRequestQueue_1_deq_bits_index;
        exeReqReg_1_bits_ffo <= exeRequestQueue_1_deq_bits_ffo;
      end
      if (tokenIO_2_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_2_valid <= tokenIO_2_maskRequestRelease_0 & ~viota;
      if (tokenIO_2_maskRequestRelease_0) begin
        exeReqReg_2_bits_source1 <= exeRequestQueue_2_deq_bits_source1;
        exeReqReg_2_bits_source2 <= exeRequestQueue_2_deq_bits_source2;
        exeReqReg_2_bits_index <= exeRequestQueue_2_deq_bits_index;
        exeReqReg_2_bits_ffo <= exeRequestQueue_2_deq_bits_ffo;
      end
      if (tokenIO_3_maskRequestRelease_0 ^ lastExecuteGroupDeq)
        exeReqReg_3_valid <= tokenIO_3_maskRequestRelease_0 & ~viota;
      if (tokenIO_3_maskRequestRelease_0) begin
        exeReqReg_3_bits_source1 <= exeRequestQueue_3_deq_bits_source1;
        exeReqReg_3_bits_source2 <= exeRequestQueue_3_deq_bits_source2;
        exeReqReg_3_bits_index <= exeRequestQueue_3_deq_bits_index;
        exeReqReg_3_bits_ffo <= exeRequestQueue_3_deq_bits_ffo;
      end
      if (instReq_valid | groupCounterAdd)
        requestCounter <= instReq_valid ? 8'h0 : requestCounter + 8'h1;
      if (requestStageDeq & anyDataValid)
        executeIndex <= executeIndex + executeIndexGrowth[1:0];
      if (readIssueStageEnq) begin
        readIssueStageState_groupReadState <= 4'h0;
        readIssueStageState_needRead <= _GEN_74 ? _slideAddressGen_indexDeq_bits_needRead : ~notReadSelect;
        readIssueStageState_elementValid <= _GEN_74 ? _slideAddressGen_indexDeq_bits_elementValid : elementValidSelect;
        readIssueStageState_replaceVs1 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_replaceVs1 : 4'h0;
        readIssueStageState_readOffset <= _GEN_74 ? _slideAddressGen_indexDeq_bits_readOffset : offsetSelect;
        readIssueStageState_accessLane_0 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_accessLane_0 : accessLaneSelect[1:0];
        readIssueStageState_accessLane_1 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_accessLane_1 : accessLaneSelect[3:2];
        readIssueStageState_accessLane_2 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_accessLane_2 : accessLaneSelect[5:4];
        readIssueStageState_accessLane_3 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_accessLane_3 : accessLaneSelect[7:6];
        readIssueStageState_vsGrowth_0 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_vsGrowth_0 : growthSelect[2:0];
        readIssueStageState_vsGrowth_1 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_vsGrowth_1 : growthSelect[5:3];
        readIssueStageState_vsGrowth_2 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_vsGrowth_2 : growthSelect[8:6];
        readIssueStageState_vsGrowth_3 <= _GEN_74 ? _slideAddressGen_indexDeq_bits_vsGrowth_3 : growthSelect[11:9];
        readIssueStageState_executeGroup <= _GEN_74 ? _slideAddressGen_indexDeq_bits_executeGroup : executeGroup;
        readIssueStageState_readDataOffset <= _GEN_74 ? _slideAddressGen_indexDeq_bits_readDataOffset : dataOffsetSelect;
        readIssueStageState_last <= _GEN_74 ? _slideAddressGen_indexDeq_bits_last : isVlBoundary;
      end
      else if (anyReadFire)
        readIssueStageState_groupReadState <= readStateUpdate;
      if (readTypeRequestDeq ^ readIssueStageEnq)
        readIssueStageValid <= readIssueStageEnq;
      if (_tokenCheck_T ^ readTokenRelease_0)
        tokenCheck_counter <= tokenCheck_counter + tokenCheck_counterChange;
      if (pipeReadFire_1 ^ readTokenRelease_1)
        tokenCheck_counter_1 <= tokenCheck_counter_1 + tokenCheck_counterChange_1;
      if (pipeReadFire_2 ^ readTokenRelease_2)
        tokenCheck_counter_2 <= tokenCheck_counter_2 + tokenCheck_counterChange_2;
      if (pipeReadFire_3 ^ readTokenRelease_3)
        tokenCheck_counter_3 <= tokenCheck_counter_3 + tokenCheck_counterChange_3;
      if (reorderQueueAllocate_release | readIssueStageEnq) begin
        reorderQueueAllocate_counter <= reorderQueueAllocate_counterUpdate;
        reorderQueueAllocate_counterWillUpdate <= reorderQueueAllocate_counterUpdate + 4'h4;
      end
      if (reorderQueueAllocate_release_1 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_1 <= reorderQueueAllocate_counterUpdate_1;
        reorderQueueAllocate_counterWillUpdate_1 <= reorderQueueAllocate_counterUpdate_1 + 4'h4;
      end
      if (reorderQueueAllocate_release_2 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_2 <= reorderQueueAllocate_counterUpdate_2;
        reorderQueueAllocate_counterWillUpdate_2 <= reorderQueueAllocate_counterUpdate_2 + 4'h4;
      end
      if (reorderQueueAllocate_release_3 | readIssueStageEnq) begin
        reorderQueueAllocate_counter_3 <= reorderQueueAllocate_counterUpdate_3;
        reorderQueueAllocate_counterWillUpdate_3 <= reorderQueueAllocate_counterUpdate_3 + 4'h4;
      end
      if (reorderStageEnqFire ^ reorderStageDeqFire)
        reorderStageValid <= reorderStageEnqFire;
      if (_write1HPipe_0_T & readType)
        reorderStageState_0 <= reorderStageState_0 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_0 <= 3'h0;
      if (_write1HPipe_1_T & readType)
        reorderStageState_1 <= reorderStageState_1 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_1 <= 3'h0;
      if (_write1HPipe_2_T & readType)
        reorderStageState_2 <= reorderStageState_2 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_2 <= 3'h0;
      if (_write1HPipe_3_T & readType)
        reorderStageState_3 <= reorderStageState_3 + 3'h1;
      else if (reorderStageEnqFire)
        reorderStageState_3 <= 3'h0;
      if (reorderStageEnqFire) begin
        reorderStageNeed_0 <= accessCountQueue_deq_bits_0;
        reorderStageNeed_1 <= accessCountQueue_deq_bits_1;
        reorderStageNeed_2 <= accessCountQueue_deq_bits_2;
        reorderStageNeed_3 <= accessCountQueue_deq_bits_3;
      end
      if (waiteStageEnqFire) begin
        waiteReadDataPipeReg_executeGroup <= readWaitQueue_deq_bits_executeGroup;
        waiteReadDataPipeReg_sourceValid <= readWaitQueue_deq_bits_sourceValid;
        waiteReadDataPipeReg_replaceVs1 <= readWaitQueue_deq_bits_replaceVs1;
        waiteReadDataPipeReg_needRead <= readWaitQueue_deq_bits_needRead;
        waiteReadDataPipeReg_last <= readWaitQueue_deq_bits_last;
      end
      if (readTokenRelease_1)
        waiteReadData_1 <= readData_readDataQueue_1_deq_bits;
      if (readTokenRelease_2)
        waiteReadData_2 <= readData_readDataQueue_2_deq_bits;
      if (readTokenRelease_3)
        waiteReadData_3 <= readData_readDataQueue_3_deq_bits;
      if (waiteStageEnqFire & (|readResultValid))
        waiteReadSate <= readResultValid;
      else if (|readResultValid)
        waiteReadSate <= waiteReadSate | readResultValid;
      else if (waiteStageEnqFire)
        waiteReadSate <= 4'h0;
      if (waiteStageDeqFire ^ waiteStageEnqFire)
        waiteReadStageValid <= waiteStageEnqFire;
      if (_dataNotInShifter_T ^ writeRelease_0)
        dataNotInShifter_writeTokenCounter <= dataNotInShifter_writeTokenCounter + dataNotInShifter_writeTokenChange;
      if (_dataNotInShifter_T_3 ^ writeRelease_1)
        dataNotInShifter_writeTokenCounter_1 <= dataNotInShifter_writeTokenCounter_1 + dataNotInShifter_writeTokenChange_1;
      if (_dataNotInShifter_T_6 ^ writeRelease_2)
        dataNotInShifter_writeTokenCounter_2 <= dataNotInShifter_writeTokenCounter_2 + dataNotInShifter_writeTokenChange_2;
      if (_dataNotInShifter_T_9 ^ writeRelease_3)
        dataNotInShifter_writeTokenCounter_3 <= dataNotInShifter_writeTokenCounter_3 + dataNotInShifter_writeTokenChange_3;
      waiteLastRequest <= ~readType & requestStageDeq & lastGroup | ~lastReportValid & waiteLastRequest;
      waitQueueClear <= executeStageClean | invalidEnq | ~lastReportValid & waitQueueClear;
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:88];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [6:0] i = 7'h0; i < 7'h59; i += 7'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        v0_0 = _RANDOM[7'h0];
        v0_1 = _RANDOM[7'h1];
        v0_2 = _RANDOM[7'h2];
        v0_3 = _RANDOM[7'h3];
        v0_4 = _RANDOM[7'h4];
        v0_5 = _RANDOM[7'h5];
        v0_6 = _RANDOM[7'h6];
        v0_7 = _RANDOM[7'h7];
        v0_8 = _RANDOM[7'h8];
        v0_9 = _RANDOM[7'h9];
        v0_10 = _RANDOM[7'hA];
        v0_11 = _RANDOM[7'hB];
        v0_12 = _RANDOM[7'hC];
        v0_13 = _RANDOM[7'hD];
        v0_14 = _RANDOM[7'hE];
        v0_15 = _RANDOM[7'hF];
        v0_16 = _RANDOM[7'h10];
        v0_17 = _RANDOM[7'h11];
        v0_18 = _RANDOM[7'h12];
        v0_19 = _RANDOM[7'h13];
        v0_20 = _RANDOM[7'h14];
        v0_21 = _RANDOM[7'h15];
        v0_22 = _RANDOM[7'h16];
        v0_23 = _RANDOM[7'h17];
        v0_24 = _RANDOM[7'h18];
        v0_25 = _RANDOM[7'h19];
        v0_26 = _RANDOM[7'h1A];
        v0_27 = _RANDOM[7'h1B];
        v0_28 = _RANDOM[7'h1C];
        v0_29 = _RANDOM[7'h1D];
        v0_30 = _RANDOM[7'h1E];
        v0_31 = _RANDOM[7'h1F];
        v0_32 = _RANDOM[7'h20];
        v0_33 = _RANDOM[7'h21];
        v0_34 = _RANDOM[7'h22];
        v0_35 = _RANDOM[7'h23];
        v0_36 = _RANDOM[7'h24];
        v0_37 = _RANDOM[7'h25];
        v0_38 = _RANDOM[7'h26];
        v0_39 = _RANDOM[7'h27];
        v0_40 = _RANDOM[7'h28];
        v0_41 = _RANDOM[7'h29];
        v0_42 = _RANDOM[7'h2A];
        v0_43 = _RANDOM[7'h2B];
        v0_44 = _RANDOM[7'h2C];
        v0_45 = _RANDOM[7'h2D];
        v0_46 = _RANDOM[7'h2E];
        v0_47 = _RANDOM[7'h2F];
        v0_48 = _RANDOM[7'h30];
        v0_49 = _RANDOM[7'h31];
        v0_50 = _RANDOM[7'h32];
        v0_51 = _RANDOM[7'h33];
        v0_52 = _RANDOM[7'h34];
        v0_53 = _RANDOM[7'h35];
        v0_54 = _RANDOM[7'h36];
        v0_55 = _RANDOM[7'h37];
        v0_56 = _RANDOM[7'h38];
        v0_57 = _RANDOM[7'h39];
        v0_58 = _RANDOM[7'h3A];
        v0_59 = _RANDOM[7'h3B];
        v0_60 = _RANDOM[7'h3C];
        v0_61 = _RANDOM[7'h3D];
        v0_62 = _RANDOM[7'h3E];
        v0_63 = _RANDOM[7'h3F];
        gatherReadState = _RANDOM[7'h40][1:0];
        gatherDatOffset = _RANDOM[7'h40][3:2];
        gatherLane = _RANDOM[7'h40][5:4];
        gatherOffset = _RANDOM[7'h40][9:6];
        gatherGrowth = _RANDOM[7'h40][12:10];
        instReg_instructionIndex = _RANDOM[7'h40][15:13];
        instReg_decodeResult_specialSlot = _RANDOM[7'h40][16];
        instReg_decodeResult_topUop = _RANDOM[7'h40][21:17];
        instReg_decodeResult_popCount = _RANDOM[7'h40][22];
        instReg_decodeResult_ffo = _RANDOM[7'h40][23];
        instReg_decodeResult_average = _RANDOM[7'h40][24];
        instReg_decodeResult_reverse = _RANDOM[7'h40][25];
        instReg_decodeResult_dontNeedExecuteInLane = _RANDOM[7'h40][26];
        instReg_decodeResult_scheduler = _RANDOM[7'h40][27];
        instReg_decodeResult_sReadVD = _RANDOM[7'h40][28];
        instReg_decodeResult_vtype = _RANDOM[7'h40][29];
        instReg_decodeResult_sWrite = _RANDOM[7'h40][30];
        instReg_decodeResult_crossRead = _RANDOM[7'h40][31];
        instReg_decodeResult_crossWrite = _RANDOM[7'h41][0];
        instReg_decodeResult_maskUnit = _RANDOM[7'h41][1];
        instReg_decodeResult_special = _RANDOM[7'h41][2];
        instReg_decodeResult_saturate = _RANDOM[7'h41][3];
        instReg_decodeResult_vwmacc = _RANDOM[7'h41][4];
        instReg_decodeResult_readOnly = _RANDOM[7'h41][5];
        instReg_decodeResult_maskSource = _RANDOM[7'h41][6];
        instReg_decodeResult_maskDestination = _RANDOM[7'h41][7];
        instReg_decodeResult_maskLogic = _RANDOM[7'h41][8];
        instReg_decodeResult_uop = _RANDOM[7'h41][12:9];
        instReg_decodeResult_iota = _RANDOM[7'h41][13];
        instReg_decodeResult_mv = _RANDOM[7'h41][14];
        instReg_decodeResult_extend = _RANDOM[7'h41][15];
        instReg_decodeResult_unOrderWrite = _RANDOM[7'h41][16];
        instReg_decodeResult_compress = _RANDOM[7'h41][17];
        instReg_decodeResult_gather16 = _RANDOM[7'h41][18];
        instReg_decodeResult_gather = _RANDOM[7'h41][19];
        instReg_decodeResult_slid = _RANDOM[7'h41][20];
        instReg_decodeResult_targetRd = _RANDOM[7'h41][21];
        instReg_decodeResult_widenReduce = _RANDOM[7'h41][22];
        instReg_decodeResult_red = _RANDOM[7'h41][23];
        instReg_decodeResult_nr = _RANDOM[7'h41][24];
        instReg_decodeResult_itype = _RANDOM[7'h41][25];
        instReg_decodeResult_unsigned1 = _RANDOM[7'h41][26];
        instReg_decodeResult_unsigned0 = _RANDOM[7'h41][27];
        instReg_decodeResult_other = _RANDOM[7'h41][28];
        instReg_decodeResult_multiCycle = _RANDOM[7'h41][29];
        instReg_decodeResult_divider = _RANDOM[7'h41][30];
        instReg_decodeResult_multiplier = _RANDOM[7'h41][31];
        instReg_decodeResult_shift = _RANDOM[7'h42][0];
        instReg_decodeResult_adder = _RANDOM[7'h42][1];
        instReg_decodeResult_logic = _RANDOM[7'h42][2];
        instReg_readFromScala = {_RANDOM[7'h42][31:3], _RANDOM[7'h43][2:0]};
        instReg_sew = _RANDOM[7'h43][4:3];
        instReg_vlmul = _RANDOM[7'h43][7:5];
        instReg_maskType = _RANDOM[7'h43][8];
        instReg_vxrm = _RANDOM[7'h43][11:9];
        instReg_vs2 = _RANDOM[7'h43][16:12];
        instReg_vs1 = _RANDOM[7'h43][21:17];
        instReg_vd = _RANDOM[7'h43][26:22];
        instReg_vl = {_RANDOM[7'h43][31:27], _RANDOM[7'h44][6:0]};
        instVlValid = _RANDOM[7'h44][7];
        readVS1Reg_dataValid = _RANDOM[7'h44][8];
        readVS1Reg_requestSend = _RANDOM[7'h44][9];
        readVS1Reg_sendToExecution = _RANDOM[7'h44][10];
        readVS1Reg_data = {_RANDOM[7'h44][31:11], _RANDOM[7'h45][10:0]};
        readVS1Reg_readIndex = _RANDOM[7'h45][17:11];
        exeReqReg_0_valid = _RANDOM[7'h45][22];
        exeReqReg_0_bits_source1 = {_RANDOM[7'h45][31:23], _RANDOM[7'h46][22:0]};
        exeReqReg_0_bits_source2 = {_RANDOM[7'h46][31:23], _RANDOM[7'h47][22:0]};
        exeReqReg_0_bits_index = _RANDOM[7'h47][25:23];
        exeReqReg_0_bits_ffo = _RANDOM[7'h47][26];
        exeReqReg_1_valid = _RANDOM[7'h47][27];
        exeReqReg_1_bits_source1 = {_RANDOM[7'h47][31:28], _RANDOM[7'h48][27:0]};
        exeReqReg_1_bits_source2 = {_RANDOM[7'h48][31:28], _RANDOM[7'h49][27:0]};
        exeReqReg_1_bits_index = _RANDOM[7'h49][30:28];
        exeReqReg_1_bits_ffo = _RANDOM[7'h49][31];
        exeReqReg_2_valid = _RANDOM[7'h4A][0];
        exeReqReg_2_bits_source1 = {_RANDOM[7'h4A][31:1], _RANDOM[7'h4B][0]};
        exeReqReg_2_bits_source2 = {_RANDOM[7'h4B][31:1], _RANDOM[7'h4C][0]};
        exeReqReg_2_bits_index = _RANDOM[7'h4C][3:1];
        exeReqReg_2_bits_ffo = _RANDOM[7'h4C][4];
        exeReqReg_3_valid = _RANDOM[7'h4C][5];
        exeReqReg_3_bits_source1 = {_RANDOM[7'h4C][31:6], _RANDOM[7'h4D][5:0]};
        exeReqReg_3_bits_source2 = {_RANDOM[7'h4D][31:6], _RANDOM[7'h4E][5:0]};
        exeReqReg_3_bits_index = _RANDOM[7'h4E][8:6];
        exeReqReg_3_bits_ffo = _RANDOM[7'h4E][9];
        requestCounter = _RANDOM[7'h4E][17:10];
        executeIndex = _RANDOM[7'h4E][19:18];
        readIssueStageState_groupReadState = _RANDOM[7'h4E][23:20];
        readIssueStageState_needRead = _RANDOM[7'h4E][27:24];
        readIssueStageState_elementValid = _RANDOM[7'h4E][31:28];
        readIssueStageState_replaceVs1 = _RANDOM[7'h4F][3:0];
        readIssueStageState_readOffset = _RANDOM[7'h4F][19:4];
        readIssueStageState_accessLane_0 = _RANDOM[7'h4F][21:20];
        readIssueStageState_accessLane_1 = _RANDOM[7'h4F][23:22];
        readIssueStageState_accessLane_2 = _RANDOM[7'h4F][25:24];
        readIssueStageState_accessLane_3 = _RANDOM[7'h4F][27:26];
        readIssueStageState_vsGrowth_0 = _RANDOM[7'h4F][30:28];
        readIssueStageState_vsGrowth_1 = {_RANDOM[7'h4F][31], _RANDOM[7'h50][1:0]};
        readIssueStageState_vsGrowth_2 = _RANDOM[7'h50][4:2];
        readIssueStageState_vsGrowth_3 = _RANDOM[7'h50][7:5];
        readIssueStageState_executeGroup = _RANDOM[7'h50][17:8];
        readIssueStageState_readDataOffset = _RANDOM[7'h50][25:18];
        readIssueStageState_last = _RANDOM[7'h50][26];
        readIssueStageValid = _RANDOM[7'h50][27];
        tokenCheck_counter = _RANDOM[7'h50][31:28];
        tokenCheck_counter_1 = _RANDOM[7'h51][3:0];
        tokenCheck_counter_2 = _RANDOM[7'h51][7:4];
        tokenCheck_counter_3 = _RANDOM[7'h51][11:8];
        reorderQueueAllocate_counter = _RANDOM[7'h51][15:12];
        reorderQueueAllocate_counterWillUpdate = _RANDOM[7'h51][19:16];
        reorderQueueAllocate_counter_1 = _RANDOM[7'h51][23:20];
        reorderQueueAllocate_counterWillUpdate_1 = _RANDOM[7'h51][27:24];
        reorderQueueAllocate_counter_2 = _RANDOM[7'h51][31:28];
        reorderQueueAllocate_counterWillUpdate_2 = _RANDOM[7'h52][3:0];
        reorderQueueAllocate_counter_3 = _RANDOM[7'h52][7:4];
        reorderQueueAllocate_counterWillUpdate_3 = _RANDOM[7'h52][11:8];
        reorderStageValid = _RANDOM[7'h52][12];
        reorderStageState_0 = _RANDOM[7'h52][15:13];
        reorderStageState_1 = _RANDOM[7'h52][18:16];
        reorderStageState_2 = _RANDOM[7'h52][21:19];
        reorderStageState_3 = _RANDOM[7'h52][24:22];
        reorderStageNeed_0 = _RANDOM[7'h52][27:25];
        reorderStageNeed_1 = _RANDOM[7'h52][30:28];
        reorderStageNeed_2 = {_RANDOM[7'h52][31], _RANDOM[7'h53][1:0]};
        reorderStageNeed_3 = _RANDOM[7'h53][4:2];
        waiteReadDataPipeReg_executeGroup = _RANDOM[7'h53][14:5];
        waiteReadDataPipeReg_sourceValid = _RANDOM[7'h53][18:15];
        waiteReadDataPipeReg_replaceVs1 = _RANDOM[7'h53][22:19];
        waiteReadDataPipeReg_needRead = _RANDOM[7'h53][26:23];
        waiteReadDataPipeReg_last = _RANDOM[7'h53][27];
        waiteReadData_0 = {_RANDOM[7'h53][31:28], _RANDOM[7'h54][27:0]};
        waiteReadData_1 = {_RANDOM[7'h54][31:28], _RANDOM[7'h55][27:0]};
        waiteReadData_2 = {_RANDOM[7'h55][31:28], _RANDOM[7'h56][27:0]};
        waiteReadData_3 = {_RANDOM[7'h56][31:28], _RANDOM[7'h57][27:0]};
        waiteReadSate = _RANDOM[7'h57][31:28];
        waiteReadStageValid = _RANDOM[7'h58][0];
        dataNotInShifter_writeTokenCounter = _RANDOM[7'h58][3:1];
        dataNotInShifter_writeTokenCounter_1 = _RANDOM[7'h58][6:4];
        dataNotInShifter_writeTokenCounter_2 = _RANDOM[7'h58][9:7];
        dataNotInShifter_writeTokenCounter_3 = _RANDOM[7'h58][12:10];
        waiteLastRequest = _RANDOM[7'h58][13];
        waitQueueClear = _RANDOM[7'h58][14];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire               exeRequestQueue_0_empty;
  assign exeRequestQueue_0_empty = _exeRequestQueue_queue_fifo_empty;
  wire               exeRequestQueue_0_full;
  assign exeRequestQueue_0_full = _exeRequestQueue_queue_fifo_full;
  wire               exeRequestQueue_1_empty;
  assign exeRequestQueue_1_empty = _exeRequestQueue_queue_fifo_1_empty;
  wire               exeRequestQueue_1_full;
  assign exeRequestQueue_1_full = _exeRequestQueue_queue_fifo_1_full;
  wire               exeRequestQueue_2_empty;
  assign exeRequestQueue_2_empty = _exeRequestQueue_queue_fifo_2_empty;
  wire               exeRequestQueue_2_full;
  assign exeRequestQueue_2_full = _exeRequestQueue_queue_fifo_2_full;
  wire               exeRequestQueue_3_empty;
  assign exeRequestQueue_3_empty = _exeRequestQueue_queue_fifo_3_empty;
  wire               exeRequestQueue_3_full;
  assign exeRequestQueue_3_full = _exeRequestQueue_queue_fifo_3_full;
  wire               accessCountQueue_empty;
  assign accessCountQueue_empty = _accessCountQueue_fifo_empty;
  wire               accessCountQueue_full;
  assign accessCountQueue_full = _accessCountQueue_fifo_full;
  wire               readWaitQueue_empty;
  assign readWaitQueue_empty = _readWaitQueue_fifo_empty;
  wire               readWaitQueue_full;
  assign readWaitQueue_full = _readWaitQueue_fifo_full;
  assign compressUnitResultQueue_empty = _compressUnitResultQueue_fifo_empty;
  wire               compressUnitResultQueue_full;
  assign compressUnitResultQueue_full = _compressUnitResultQueue_fifo_full;
  wire               reorderQueueVec_0_empty;
  assign reorderQueueVec_0_empty = _reorderQueueVec_fifo_empty;
  wire               reorderQueueVec_0_full;
  assign reorderQueueVec_0_full = _reorderQueueVec_fifo_full;
  wire               reorderQueueVec_1_empty;
  assign reorderQueueVec_1_empty = _reorderQueueVec_fifo_1_empty;
  wire               reorderQueueVec_1_full;
  assign reorderQueueVec_1_full = _reorderQueueVec_fifo_1_full;
  wire               reorderQueueVec_2_empty;
  assign reorderQueueVec_2_empty = _reorderQueueVec_fifo_2_empty;
  wire               reorderQueueVec_2_full;
  assign reorderQueueVec_2_full = _reorderQueueVec_fifo_2_full;
  wire               reorderQueueVec_3_empty;
  assign reorderQueueVec_3_empty = _reorderQueueVec_fifo_3_empty;
  wire               reorderQueueVec_3_full;
  assign reorderQueueVec_3_full = _reorderQueueVec_fifo_3_full;
  wire               readMessageQueue_empty;
  assign readMessageQueue_empty = _readMessageQueue_fifo_empty;
  wire               readMessageQueue_full;
  assign readMessageQueue_full = _readMessageQueue_fifo_full;
  wire               readMessageQueue_1_empty;
  assign readMessageQueue_1_empty = _readMessageQueue_fifo_1_empty;
  wire               readMessageQueue_1_full;
  assign readMessageQueue_1_full = _readMessageQueue_fifo_1_full;
  wire               readMessageQueue_2_empty;
  assign readMessageQueue_2_empty = _readMessageQueue_fifo_2_empty;
  wire               readMessageQueue_2_full;
  assign readMessageQueue_2_full = _readMessageQueue_fifo_2_full;
  wire               readMessageQueue_3_empty;
  assign readMessageQueue_3_empty = _readMessageQueue_fifo_3_empty;
  wire               readMessageQueue_3_full;
  assign readMessageQueue_3_full = _readMessageQueue_fifo_3_full;
  wire               readData_readDataQueue_empty;
  assign readData_readDataQueue_empty = _readData_readDataQueue_fifo_empty;
  wire               readData_readDataQueue_full;
  assign readData_readDataQueue_full = _readData_readDataQueue_fifo_full;
  wire               readData_readDataQueue_1_empty;
  assign readData_readDataQueue_1_empty = _readData_readDataQueue_fifo_1_empty;
  wire               readData_readDataQueue_1_full;
  assign readData_readDataQueue_1_full = _readData_readDataQueue_fifo_1_full;
  wire               readData_readDataQueue_2_empty;
  assign readData_readDataQueue_2_empty = _readData_readDataQueue_fifo_2_empty;
  wire               readData_readDataQueue_2_full;
  assign readData_readDataQueue_2_full = _readData_readDataQueue_fifo_2_full;
  wire               readData_readDataQueue_3_empty;
  assign readData_readDataQueue_3_empty = _readData_readDataQueue_fifo_3_empty;
  wire               readData_readDataQueue_3_full;
  assign readData_readDataQueue_3_full = _readData_readDataQueue_fifo_3_full;
  assign compressUnitResultQueue_enq_valid = _compressUnit_out_compressValid;
  assign compressUnitResultQueue_enq_bits_compressValid = _compressUnit_out_compressValid;
  wire               writeQueue_0_empty;
  assign writeQueue_0_empty = _writeQueue_fifo_empty;
  wire               writeQueue_0_full;
  assign writeQueue_0_full = _writeQueue_fifo_full;
  wire               writeQueue_1_empty;
  assign writeQueue_1_empty = _writeQueue_fifo_1_empty;
  wire               writeQueue_1_full;
  assign writeQueue_1_full = _writeQueue_fifo_1_full;
  wire               writeQueue_2_empty;
  assign writeQueue_2_empty = _writeQueue_fifo_2_empty;
  wire               writeQueue_2_full;
  assign writeQueue_2_full = _writeQueue_fifo_2_full;
  wire               writeQueue_3_empty;
  assign writeQueue_3_empty = _writeQueue_fifo_3_empty;
  wire               writeQueue_3_full;
  assign writeQueue_3_full = _writeQueue_fifo_3_full;
  BitLevelMaskWrite maskedWrite (
    .clock                             (clock),
    .reset                             (reset),
    .needWAR                           (maskDestinationType),
    .vd                                (instReg_vd),
    .in_0_ready                        (_maskedWrite_in_0_ready),
    .in_0_valid                        (unitType[2] ? _reduceUnit_out_valid : executeValid & maskFilter),
    .in_0_bits_data                    (unitType[2] ? _reduceUnit_out_bits_data : executeResult[31:0]),
    .in_0_bits_bitMask                 (currentMaskGroupForDestination[31:0]),
    .in_0_bits_mask                    (unitType[2] ? _reduceUnit_out_bits_mask : executeWriteByteMask[3:0]),
    .in_0_bits_groupCounter            (unitType[2] ? 8'h0 : executeDeqGroupCounter[7:0]),
    .in_0_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[0] & ffo),
    .in_1_ready                        (_maskedWrite_in_1_ready),
    .in_1_valid                        (executeValid & maskFilter_1),
    .in_1_bits_data                    (executeResult[63:32]),
    .in_1_bits_bitMask                 (currentMaskGroupForDestination[63:32]),
    .in_1_bits_mask                    (executeWriteByteMask[7:4]),
    .in_1_bits_groupCounter            (executeDeqGroupCounter[7:0]),
    .in_1_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[1] & ffo),
    .in_2_ready                        (_maskedWrite_in_2_ready),
    .in_2_valid                        (executeValid & maskFilter_2),
    .in_2_bits_data                    (executeResult[95:64]),
    .in_2_bits_bitMask                 (currentMaskGroupForDestination[95:64]),
    .in_2_bits_mask                    (executeWriteByteMask[11:8]),
    .in_2_bits_groupCounter            (executeDeqGroupCounter[7:0]),
    .in_2_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[2] & ffo),
    .in_3_ready                        (_maskedWrite_in_3_ready),
    .in_3_valid                        (executeValid & maskFilter_3),
    .in_3_bits_data                    (executeResult[127:96]),
    .in_3_bits_bitMask                 (currentMaskGroupForDestination[127:96]),
    .in_3_bits_mask                    (executeWriteByteMask[15:12]),
    .in_3_bits_groupCounter            (executeDeqGroupCounter[7:0]),
    .in_3_bits_ffoByOther              (compressUnitResultQueue_deq_bits_ffoOutput[3] & ffo),
    .out_0_ready                       (writeQueue_0_enq_ready),
    .out_0_valid                       (_maskedWrite_out_0_valid),
    .out_0_bits_ffoByOther             (_maskedWrite_out_0_bits_ffoByOther),
    .out_0_bits_writeData_data         (_maskedWrite_out_0_bits_writeData_data),
    .out_0_bits_writeData_mask         (_maskedWrite_out_0_bits_writeData_mask),
    .out_0_bits_writeData_groupCounter (_maskedWrite_out_0_bits_writeData_groupCounter),
    .out_1_ready                       (writeQueue_1_enq_ready),
    .out_1_valid                       (_maskedWrite_out_1_valid),
    .out_1_bits_ffoByOther             (_maskedWrite_out_1_bits_ffoByOther),
    .out_1_bits_writeData_data         (_maskedWrite_out_1_bits_writeData_data),
    .out_1_bits_writeData_mask         (_maskedWrite_out_1_bits_writeData_mask),
    .out_1_bits_writeData_groupCounter (_maskedWrite_out_1_bits_writeData_groupCounter),
    .out_2_ready                       (writeQueue_2_enq_ready),
    .out_2_valid                       (_maskedWrite_out_2_valid),
    .out_2_bits_ffoByOther             (_maskedWrite_out_2_bits_ffoByOther),
    .out_2_bits_writeData_data         (_maskedWrite_out_2_bits_writeData_data),
    .out_2_bits_writeData_mask         (_maskedWrite_out_2_bits_writeData_mask),
    .out_2_bits_writeData_groupCounter (_maskedWrite_out_2_bits_writeData_groupCounter),
    .out_3_ready                       (writeQueue_3_enq_ready),
    .out_3_valid                       (_maskedWrite_out_3_valid),
    .out_3_bits_ffoByOther             (_maskedWrite_out_3_bits_ffoByOther),
    .out_3_bits_writeData_data         (_maskedWrite_out_3_bits_writeData_data),
    .out_3_bits_writeData_mask         (_maskedWrite_out_3_bits_writeData_mask),
    .out_3_bits_writeData_groupCounter (_maskedWrite_out_3_bits_writeData_groupCounter),
    .readChannel_0_ready               (readChannel_0_ready_0),
    .readChannel_0_valid               (_maskedWrite_readChannel_0_valid),
    .readChannel_0_bits_vs             (_maskedWrite_readChannel_0_bits_vs),
    .readChannel_0_bits_offset         (_maskedWrite_readChannel_0_bits_offset),
    .readChannel_1_ready               (readChannel_1_ready_0),
    .readChannel_1_valid               (_maskedWrite_readChannel_1_valid),
    .readChannel_1_bits_vs             (_maskedWrite_readChannel_1_bits_vs),
    .readChannel_1_bits_offset         (_maskedWrite_readChannel_1_bits_offset),
    .readChannel_2_ready               (readChannel_2_ready_0),
    .readChannel_2_valid               (_maskedWrite_readChannel_2_valid),
    .readChannel_2_bits_vs             (_maskedWrite_readChannel_2_bits_vs),
    .readChannel_2_bits_offset         (_maskedWrite_readChannel_2_bits_offset),
    .readChannel_3_ready               (readChannel_3_ready_0),
    .readChannel_3_valid               (_maskedWrite_readChannel_3_valid),
    .readChannel_3_bits_vs             (_maskedWrite_readChannel_3_bits_vs),
    .readChannel_3_bits_offset         (_maskedWrite_readChannel_3_bits_offset),
    .readResult_0_valid                (readResult_0_valid),
    .readResult_0_bits                 (readResult_0_bits),
    .readResult_1_valid                (readResult_1_valid),
    .readResult_1_bits                 (readResult_1_bits),
    .readResult_2_valid                (readResult_2_valid),
    .readResult_2_bits                 (readResult_2_bits),
    .readResult_3_valid                (readResult_3_valid),
    .readResult_3_bits                 (readResult_3_bits),
    .stageClear                        (_maskedWrite_stageClear)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_0_enq_ready & exeRequestQueue_0_enq_valid & ~(_exeRequestQueue_queue_fifo_empty & exeRequestQueue_0_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_0_deq_ready & ~_exeRequestQueue_queue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn),
    .empty        (_exeRequestQueue_queue_fifo_empty),
    .almost_empty (exeRequestQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_0_almostFull),
    .full         (_exeRequestQueue_queue_fifo_full),
    .error        (_exeRequestQueue_queue_fifo_error),
    .data_out     (_exeRequestQueue_queue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_1_enq_ready & exeRequestQueue_1_enq_valid & ~(_exeRequestQueue_queue_fifo_1_empty & exeRequestQueue_1_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_1_deq_ready & ~_exeRequestQueue_queue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_1),
    .empty        (_exeRequestQueue_queue_fifo_1_empty),
    .almost_empty (exeRequestQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_1_almostFull),
    .full         (_exeRequestQueue_queue_fifo_1_full),
    .error        (_exeRequestQueue_queue_fifo_1_error),
    .data_out     (_exeRequestQueue_queue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_2_enq_ready & exeRequestQueue_2_enq_valid & ~(_exeRequestQueue_queue_fifo_2_empty & exeRequestQueue_2_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_2_deq_ready & ~_exeRequestQueue_queue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_2),
    .empty        (_exeRequestQueue_queue_fifo_2_empty),
    .almost_empty (exeRequestQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_2_almostFull),
    .full         (_exeRequestQueue_queue_fifo_2_full),
    .error        (_exeRequestQueue_queue_fifo_2_error),
    .data_out     (_exeRequestQueue_queue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(68)
  ) exeRequestQueue_queue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(exeRequestQueue_3_enq_ready & exeRequestQueue_3_enq_valid & ~(_exeRequestQueue_queue_fifo_3_empty & exeRequestQueue_3_deq_ready))),
    .pop_req_n    (~(exeRequestQueue_3_deq_ready & ~_exeRequestQueue_queue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (exeRequestQueue_queue_dataIn_3),
    .empty        (_exeRequestQueue_queue_fifo_3_empty),
    .almost_empty (exeRequestQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (exeRequestQueue_3_almostFull),
    .full         (_exeRequestQueue_queue_fifo_3_full),
    .error        (_exeRequestQueue_queue_fifo_3_error),
    .data_out     (_exeRequestQueue_queue_fifo_3_data_out)
  );
  SlideIndexGen slideAddressGen (
    .clock                              (clock),
    .reset                              (reset),
    .newInstruction                     (instReq_valid & (|instReq_bits_vl)),
    .instructionReq_decodeResult_topUop (instReg_decodeResult_topUop),
    .instructionReq_readFromScala       (instReg_readFromScala),
    .instructionReq_sew                 (instReg_sew),
    .instructionReq_vlmul               (instReg_vlmul),
    .instructionReq_maskType            (instReg_maskType),
    .instructionReq_vl                  (instReg_vl),
    .indexDeq_ready                     (slideAddressGen_indexDeq_ready),
    .indexDeq_valid                     (_slideAddressGen_indexDeq_valid),
    .indexDeq_bits_needRead             (_slideAddressGen_indexDeq_bits_needRead),
    .indexDeq_bits_elementValid         (_slideAddressGen_indexDeq_bits_elementValid),
    .indexDeq_bits_replaceVs1           (_slideAddressGen_indexDeq_bits_replaceVs1),
    .indexDeq_bits_readOffset           (_slideAddressGen_indexDeq_bits_readOffset),
    .indexDeq_bits_accessLane_0         (_slideAddressGen_indexDeq_bits_accessLane_0),
    .indexDeq_bits_accessLane_1         (_slideAddressGen_indexDeq_bits_accessLane_1),
    .indexDeq_bits_accessLane_2         (_slideAddressGen_indexDeq_bits_accessLane_2),
    .indexDeq_bits_accessLane_3         (_slideAddressGen_indexDeq_bits_accessLane_3),
    .indexDeq_bits_vsGrowth_0           (_slideAddressGen_indexDeq_bits_vsGrowth_0),
    .indexDeq_bits_vsGrowth_1           (_slideAddressGen_indexDeq_bits_vsGrowth_1),
    .indexDeq_bits_vsGrowth_2           (_slideAddressGen_indexDeq_bits_vsGrowth_2),
    .indexDeq_bits_vsGrowth_3           (_slideAddressGen_indexDeq_bits_vsGrowth_3),
    .indexDeq_bits_executeGroup         (_slideAddressGen_indexDeq_bits_executeGroup),
    .indexDeq_bits_readDataOffset       (_slideAddressGen_indexDeq_bits_readDataOffset),
    .indexDeq_bits_last                 (_slideAddressGen_indexDeq_bits_last),
    .slideGroupOut                      (_slideAddressGen_slideGroupOut),
    .slideMaskInput                     (_GEN_44[_slideAddressGen_slideGroupOut[8:0]])
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(12)
  ) accessCountQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(accessCountQueue_enq_ready & accessCountQueue_enq_valid)),
    .pop_req_n    (~(accessCountQueue_deq_ready & ~_accessCountQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (accessCountQueue_dataIn),
    .empty        (_accessCountQueue_fifo_empty),
    .almost_empty (accessCountQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (accessCountQueue_almostFull),
    .full         (_accessCountQueue_fifo_full),
    .error        (_accessCountQueue_fifo_error),
    .data_out     (_accessCountQueue_fifo_data_out)
  );
  MaskUnitReadCrossBar readCrossBar (
    .input_0_ready            (_readCrossBar_input_0_ready),
    .input_0_valid            (readCrossBar_input_0_valid),
    .input_0_bits_vs          (selectExecuteReq_0_bits_vs),
    .input_0_bits_offset      (selectExecuteReq_0_bits_offset),
    .input_0_bits_readLane    (selectExecuteReq_0_bits_readLane),
    .input_0_bits_dataOffset  (selectExecuteReq_0_bits_dataOffset),
    .input_1_ready            (_readCrossBar_input_1_ready),
    .input_1_valid            (readCrossBar_input_1_valid),
    .input_1_bits_vs          (selectExecuteReq_1_bits_vs),
    .input_1_bits_offset      (selectExecuteReq_1_bits_offset),
    .input_1_bits_readLane    (selectExecuteReq_1_bits_readLane),
    .input_1_bits_dataOffset  (selectExecuteReq_1_bits_dataOffset),
    .input_2_ready            (_readCrossBar_input_2_ready),
    .input_2_valid            (readCrossBar_input_2_valid),
    .input_2_bits_vs          (selectExecuteReq_2_bits_vs),
    .input_2_bits_offset      (selectExecuteReq_2_bits_offset),
    .input_2_bits_readLane    (selectExecuteReq_2_bits_readLane),
    .input_2_bits_dataOffset  (selectExecuteReq_2_bits_dataOffset),
    .input_3_ready            (_readCrossBar_input_3_ready),
    .input_3_valid            (readCrossBar_input_3_valid),
    .input_3_bits_vs          (selectExecuteReq_3_bits_vs),
    .input_3_bits_offset      (selectExecuteReq_3_bits_offset),
    .input_3_bits_readLane    (selectExecuteReq_3_bits_readLane),
    .input_3_bits_dataOffset  (selectExecuteReq_3_bits_dataOffset),
    .output_0_ready           (readChannel_0_ready_0 & readMessageQueue_enq_ready),
    .output_0_valid           (_readCrossBar_output_0_valid),
    .output_0_bits_vs         (_readCrossBar_output_0_bits_vs),
    .output_0_bits_offset     (_readCrossBar_output_0_bits_offset),
    .output_0_bits_writeIndex (_readCrossBar_output_0_bits_writeIndex),
    .output_0_bits_dataOffset (readMessageQueue_enq_bits_dataOffset),
    .output_1_ready           (readChannel_1_ready_0 & readMessageQueue_1_enq_ready),
    .output_1_valid           (_readCrossBar_output_1_valid),
    .output_1_bits_vs         (_readCrossBar_output_1_bits_vs),
    .output_1_bits_offset     (_readCrossBar_output_1_bits_offset),
    .output_1_bits_writeIndex (_readCrossBar_output_1_bits_writeIndex),
    .output_1_bits_dataOffset (readMessageQueue_1_enq_bits_dataOffset),
    .output_2_ready           (readChannel_2_ready_0 & readMessageQueue_2_enq_ready),
    .output_2_valid           (_readCrossBar_output_2_valid),
    .output_2_bits_vs         (_readCrossBar_output_2_bits_vs),
    .output_2_bits_offset     (_readCrossBar_output_2_bits_offset),
    .output_2_bits_writeIndex (_readCrossBar_output_2_bits_writeIndex),
    .output_2_bits_dataOffset (readMessageQueue_2_enq_bits_dataOffset),
    .output_3_ready           (readChannel_3_ready_0 & readMessageQueue_3_enq_ready),
    .output_3_valid           (_readCrossBar_output_3_valid),
    .output_3_bits_vs         (_readCrossBar_output_3_bits_vs),
    .output_3_bits_offset     (_readCrossBar_output_3_bits_offset),
    .output_3_bits_writeIndex (_readCrossBar_output_3_bits_writeIndex),
    .output_3_bits_dataOffset (readMessageQueue_3_enq_bits_dataOffset)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(64),
    .err_mode(2),
    .rst_mode(3),
    .width(23)
  ) readWaitQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readWaitQueue_enq_ready & readWaitQueue_enq_valid)),
    .pop_req_n    (~(readWaitQueue_deq_ready & ~_readWaitQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readWaitQueue_dataIn),
    .empty        (_readWaitQueue_fifo_empty),
    .almost_empty (readWaitQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readWaitQueue_almostFull),
    .full         (_readWaitQueue_fifo_full),
    .error        (_readWaitQueue_fifo_error),
    .data_out     (_readWaitQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(4),
    .err_mode(2),
    .rst_mode(3),
    .width(157)
  ) compressUnitResultQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(compressUnitResultQueue_enq_ready & compressUnitResultQueue_enq_valid & ~(_compressUnitResultQueue_fifo_empty & compressUnitResultQueue_deq_ready))),
    .pop_req_n    (~(compressUnitResultQueue_deq_ready & ~_compressUnitResultQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (compressUnitResultQueue_dataIn),
    .empty        (_compressUnitResultQueue_fifo_empty),
    .almost_empty (compressUnitResultQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (compressUnitResultQueue_almostFull),
    .full         (_compressUnitResultQueue_fifo_full),
    .error        (_compressUnitResultQueue_fifo_error),
    .data_out     (_compressUnitResultQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_0_enq_ready & reorderQueueVec_0_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_0_deq_ready & ~_reorderQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn),
    .empty        (_reorderQueueVec_fifo_empty),
    .almost_empty (reorderQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_0_almostFull),
    .full         (_reorderQueueVec_fifo_full),
    .error        (_reorderQueueVec_fifo_error),
    .data_out     (_reorderQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_1_enq_ready & reorderQueueVec_1_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_1_deq_ready & ~_reorderQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_1),
    .empty        (_reorderQueueVec_fifo_1_empty),
    .almost_empty (reorderQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_1_almostFull),
    .full         (_reorderQueueVec_fifo_1_full),
    .error        (_reorderQueueVec_fifo_1_error),
    .data_out     (_reorderQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_2_enq_ready & reorderQueueVec_2_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_2_deq_ready & ~_reorderQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_2),
    .empty        (_reorderQueueVec_fifo_2_empty),
    .almost_empty (reorderQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_2_almostFull),
    .full         (_reorderQueueVec_fifo_2_full),
    .error        (_reorderQueueVec_fifo_2_error),
    .data_out     (_reorderQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(36)
  ) reorderQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(reorderQueueVec_3_enq_ready & reorderQueueVec_3_enq_valid)),
    .pop_req_n    (~(reorderQueueVec_3_deq_ready & ~_reorderQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (reorderQueueVec_dataIn_3),
    .empty        (_reorderQueueVec_fifo_3_empty),
    .almost_empty (reorderQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (reorderQueueVec_3_almostFull),
    .full         (_reorderQueueVec_fifo_3_full),
    .error        (_reorderQueueVec_fifo_3_error),
    .data_out     (_reorderQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_enq_ready & readMessageQueue_enq_valid)),
    .pop_req_n    (~(readMessageQueue_deq_ready & ~_readMessageQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn),
    .empty        (_readMessageQueue_fifo_empty),
    .almost_empty (readMessageQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_almostFull),
    .full         (_readMessageQueue_fifo_full),
    .error        (_readMessageQueue_fifo_error),
    .data_out     (_readMessageQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_1_enq_ready & readMessageQueue_1_enq_valid)),
    .pop_req_n    (~(readMessageQueue_1_deq_ready & ~_readMessageQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_1),
    .empty        (_readMessageQueue_fifo_1_empty),
    .almost_empty (readMessageQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_1_almostFull),
    .full         (_readMessageQueue_fifo_1_full),
    .error        (_readMessageQueue_fifo_1_error),
    .data_out     (_readMessageQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_2_enq_ready & readMessageQueue_2_enq_valid)),
    .pop_req_n    (~(readMessageQueue_2_deq_ready & ~_readMessageQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_2),
    .empty        (_readMessageQueue_fifo_2_empty),
    .almost_empty (readMessageQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_2_almostFull),
    .full         (_readMessageQueue_fifo_2_full),
    .error        (_readMessageQueue_fifo_2_error),
    .data_out     (_readMessageQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(7),
    .err_mode(2),
    .rst_mode(3),
    .width(6)
  ) readMessageQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readMessageQueue_3_enq_ready & readMessageQueue_3_enq_valid)),
    .pop_req_n    (~(readMessageQueue_3_deq_ready & ~_readMessageQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readMessageQueue_dataIn_3),
    .empty        (_readMessageQueue_fifo_3_empty),
    .almost_empty (readMessageQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readMessageQueue_3_almostFull),
    .full         (_readMessageQueue_fifo_3_full),
    .error        (_readMessageQueue_fifo_3_error),
    .data_out     (_readMessageQueue_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_enq_ready & readData_readDataQueue_enq_valid & ~(_readData_readDataQueue_fifo_empty & readData_readDataQueue_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_deq_ready & ~_readData_readDataQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_enq_bits),
    .empty        (_readData_readDataQueue_fifo_empty),
    .almost_empty (readData_readDataQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_almostFull),
    .full         (_readData_readDataQueue_fifo_full),
    .error        (_readData_readDataQueue_fifo_error),
    .data_out     (_readData_readDataQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_1_enq_ready & readData_readDataQueue_1_enq_valid & ~(_readData_readDataQueue_fifo_1_empty & readData_readDataQueue_1_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_1_deq_ready & ~_readData_readDataQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_1_enq_bits),
    .empty        (_readData_readDataQueue_fifo_1_empty),
    .almost_empty (readData_readDataQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_1_almostFull),
    .full         (_readData_readDataQueue_fifo_1_full),
    .error        (_readData_readDataQueue_fifo_1_error),
    .data_out     (_readData_readDataQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_2_enq_ready & readData_readDataQueue_2_enq_valid & ~(_readData_readDataQueue_fifo_2_empty & readData_readDataQueue_2_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_2_deq_ready & ~_readData_readDataQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_2_enq_bits),
    .empty        (_readData_readDataQueue_fifo_2_empty),
    .almost_empty (readData_readDataQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_2_almostFull),
    .full         (_readData_readDataQueue_fifo_2_full),
    .error        (_readData_readDataQueue_fifo_2_error),
    .data_out     (_readData_readDataQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) readData_readDataQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(readData_readDataQueue_3_enq_ready & readData_readDataQueue_3_enq_valid & ~(_readData_readDataQueue_fifo_3_empty & readData_readDataQueue_3_deq_ready))),
    .pop_req_n    (~(readData_readDataQueue_3_deq_ready & ~_readData_readDataQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (readData_readDataQueue_3_enq_bits),
    .empty        (_readData_readDataQueue_fifo_3_empty),
    .almost_empty (readData_readDataQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (readData_readDataQueue_3_almostFull),
    .full         (_readData_readDataQueue_fifo_3_full),
    .error        (_readData_readDataQueue_fifo_3_error),
    .data_out     (_readData_readDataQueue_fifo_3_data_out)
  );
  MaskCompress compressUnit (
    .clock                  (clock),
    .reset                  (reset),
    .in_valid               (viotaCounterAdd),
    .in_bits_maskType       (instReg_maskType),
    .in_bits_eew            (instReg_sew),
    .in_bits_uop            (instReg_decodeResult_topUop[2:0]),
    .in_bits_readFromScalar (instReg_readFromScala),
    .in_bits_source1        (source1Select),
    .in_bits_mask           ({16'h0, executeElementMask}),
    .in_bits_source2        (source2),
    .in_bits_pipeData       (source1),
    .in_bits_groupCounter   (requestCounter),
    .in_bits_ffoInput       ({view__in_bits_ffoInput_hi, view__in_bits_ffoInput_lo}),
    .in_bits_validInput     ({view__in_bits_validInput_hi, view__in_bits_validInput_lo}),
    .in_bits_lastCompress   (lastGroup),
    .out_data               (compressUnitResultQueue_enq_bits_data),
    .out_mask               (compressUnitResultQueue_enq_bits_mask),
    .out_groupCounter       (compressUnitResultQueue_enq_bits_groupCounter),
    .out_ffoOutput          (compressUnitResultQueue_enq_bits_ffoOutput),
    .out_compressValid      (_compressUnit_out_compressValid),
    .newInstruction         (instReq_valid),
    .ffoInstruction         (&(instReq_bits_decodeResult_topUop[2:1])),
    .writeData              (_compressUnit_writeData),
    .stageValid             (_compressUnit_stageValid)
  );
  MaskReduce reduceUnit (
    .clock               (clock),
    .reset               (reset),
    .in_ready            (_reduceUnit_in_ready),
    .in_valid            (reduceUnit_in_valid),
    .in_bits_maskType    (instReg_maskType),
    .in_bits_eew         (instReg_sew),
    .in_bits_uop         (instReg_decodeResult_topUop[2:0]),
    .in_bits_readVS1     (readVS1Reg_data),
    .in_bits_source2     (source2),
    .in_bits_sourceValid ({view__in_bits_sourceValid_hi, view__in_bits_sourceValid_lo}),
    .in_bits_lastGroup   (lastGroup),
    .in_bits_vxrm        (instReg_vxrm),
    .in_bits_aluUop      (instReg_decodeResult_uop),
    .in_bits_sign        (~instReg_decodeResult_unsigned1),
    .out_valid           (_reduceUnit_out_valid),
    .out_bits_data       (_reduceUnit_out_bits_data),
    .out_bits_mask       (_reduceUnit_out_bits_mask),
    .firstGroup          (~readVS1Reg_sendToExecution & _view__firstGroup_T_1),
    .newInstruction      (instReq_valid),
    .validInst           (|instReg_vl),
    .pop                 (instReg_decodeResult_popCount)
  );
  MaskExtend extendUnit (
    .in_eew          (instReg_sew),
    .in_uop          (instReg_decodeResult_topUop[2:0]),
    .in_source2      (source2),
    .in_groupCounter (extendGroupCount[7:0]),
    .out             (_extendUnit_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(53)
  ) writeQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_0_enq_ready & writeQueue_0_enq_valid)),
    .pop_req_n    (~(writeQueue_0_deq_ready & ~_writeQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn),
    .empty        (_writeQueue_fifo_empty),
    .almost_empty (writeQueue_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_0_almostFull),
    .full         (_writeQueue_fifo_full),
    .error        (_writeQueue_fifo_error),
    .data_out     (_writeQueue_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(53)
  ) writeQueue_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_1_enq_ready & writeQueue_1_enq_valid)),
    .pop_req_n    (~(writeQueue_1_deq_ready & ~_writeQueue_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_1),
    .empty        (_writeQueue_fifo_1_empty),
    .almost_empty (writeQueue_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_1_almostFull),
    .full         (_writeQueue_fifo_1_full),
    .error        (_writeQueue_fifo_1_error),
    .data_out     (_writeQueue_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(53)
  ) writeQueue_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_2_enq_ready & writeQueue_2_enq_valid)),
    .pop_req_n    (~(writeQueue_2_deq_ready & ~_writeQueue_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_2),
    .empty        (_writeQueue_fifo_2_empty),
    .almost_empty (writeQueue_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_2_almostFull),
    .full         (_writeQueue_fifo_2_full),
    .error        (_writeQueue_fifo_2_error),
    .data_out     (_writeQueue_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(53)
  ) writeQueue_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(writeQueue_3_enq_ready & writeQueue_3_enq_valid)),
    .pop_req_n    (~(writeQueue_3_deq_ready & ~_writeQueue_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (writeQueue_dataIn_3),
    .empty        (_writeQueue_fifo_3_empty),
    .almost_empty (writeQueue_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (writeQueue_3_almostFull),
    .full         (_writeQueue_fifo_3_full),
    .error        (_writeQueue_fifo_3_error),
    .data_out     (_writeQueue_fifo_3_data_out)
  );
  assign exeResp_0_valid = exeResp_0_valid_0;
  assign exeResp_0_bits_vd = exeResp_0_bits_vd_0;
  assign exeResp_0_bits_offset = exeResp_0_bits_offset_0;
  assign exeResp_0_bits_mask = exeResp_0_bits_mask_0;
  assign exeResp_0_bits_data = exeResp_0_bits_data_0;
  assign exeResp_0_bits_instructionIndex = exeResp_0_bits_instructionIndex_0;
  assign exeResp_1_valid = exeResp_1_valid_0;
  assign exeResp_1_bits_vd = exeResp_1_bits_vd_0;
  assign exeResp_1_bits_offset = exeResp_1_bits_offset_0;
  assign exeResp_1_bits_mask = exeResp_1_bits_mask_0;
  assign exeResp_1_bits_data = exeResp_1_bits_data_0;
  assign exeResp_1_bits_instructionIndex = exeResp_1_bits_instructionIndex_0;
  assign exeResp_2_valid = exeResp_2_valid_0;
  assign exeResp_2_bits_vd = exeResp_2_bits_vd_0;
  assign exeResp_2_bits_offset = exeResp_2_bits_offset_0;
  assign exeResp_2_bits_mask = exeResp_2_bits_mask_0;
  assign exeResp_2_bits_data = exeResp_2_bits_data_0;
  assign exeResp_2_bits_instructionIndex = exeResp_2_bits_instructionIndex_0;
  assign exeResp_3_valid = exeResp_3_valid_0;
  assign exeResp_3_bits_vd = exeResp_3_bits_vd_0;
  assign exeResp_3_bits_offset = exeResp_3_bits_offset_0;
  assign exeResp_3_bits_mask = exeResp_3_bits_mask_0;
  assign exeResp_3_bits_data = exeResp_3_bits_data_0;
  assign exeResp_3_bits_instructionIndex = exeResp_3_bits_instructionIndex_0;
  assign tokenIO_0_maskRequestRelease = tokenIO_0_maskRequestRelease_0;
  assign tokenIO_1_maskRequestRelease = tokenIO_1_maskRequestRelease_0;
  assign tokenIO_2_maskRequestRelease = tokenIO_2_maskRequestRelease_0;
  assign tokenIO_3_maskRequestRelease = tokenIO_3_maskRequestRelease_0;
  assign readChannel_0_valid = readChannel_0_valid_0;
  assign readChannel_0_bits_vs = readChannel_0_bits_vs_0;
  assign readChannel_0_bits_offset = readChannel_0_bits_offset_0;
  assign readChannel_0_bits_instructionIndex = readChannel_0_bits_instructionIndex_0;
  assign readChannel_1_valid = readChannel_1_valid_0;
  assign readChannel_1_bits_vs = readChannel_1_bits_vs_0;
  assign readChannel_1_bits_offset = readChannel_1_bits_offset_0;
  assign readChannel_1_bits_instructionIndex = readChannel_1_bits_instructionIndex_0;
  assign readChannel_2_valid = readChannel_2_valid_0;
  assign readChannel_2_bits_vs = readChannel_2_bits_vs_0;
  assign readChannel_2_bits_offset = readChannel_2_bits_offset_0;
  assign readChannel_2_bits_instructionIndex = readChannel_2_bits_instructionIndex_0;
  assign readChannel_3_valid = readChannel_3_valid_0;
  assign readChannel_3_bits_vs = readChannel_3_bits_vs_0;
  assign readChannel_3_bits_offset = readChannel_3_bits_offset_0;
  assign readChannel_3_bits_instructionIndex = readChannel_3_bits_instructionIndex_0;
  assign lastReport = _lastReport_output;
  assign laneMaskInput_0 = _GEN_31[laneMaskSelect_0[3:0]];
  assign laneMaskInput_1 = _GEN_32[laneMaskSelect_1[3:0]];
  assign laneMaskInput_2 = _GEN_33[laneMaskSelect_2[3:0]];
  assign laneMaskInput_3 = _GEN_34[laneMaskSelect_3[3:0]];
  assign writeRDData = instReg_decodeResult_popCount ? _reduceUnit_out_bits_data : _compressUnit_writeData;
  assign gatherData_valid = gatherData_valid_0;
  assign gatherData_bits = gatherData_bits_0;
endmodule

