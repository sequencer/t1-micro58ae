
// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module StoreUnit(
  input           clock,
                  reset,
                  lsuRequest_valid,
  input  [2:0]    lsuRequest_bits_instructionInformation_nf,
  input           lsuRequest_bits_instructionInformation_mew,
  input  [1:0]    lsuRequest_bits_instructionInformation_mop,
  input  [4:0]    lsuRequest_bits_instructionInformation_lumop,
  input  [1:0]    lsuRequest_bits_instructionInformation_eew,
  input  [4:0]    lsuRequest_bits_instructionInformation_vs3,
  input           lsuRequest_bits_instructionInformation_isStore,
                  lsuRequest_bits_instructionInformation_maskedLoadStore,
  input  [31:0]   lsuRequest_bits_rs1Data,
                  lsuRequest_bits_rs2Data,
  input  [2:0]    lsuRequest_bits_instructionIndex,
  input  [10:0]   csrInterface_vl,
                  csrInterface_vStart,
  input  [2:0]    csrInterface_vlmul,
  input  [1:0]    csrInterface_vSew,
                  csrInterface_vxrm,
  input           csrInterface_vta,
                  csrInterface_vma,
  input  [127:0]  maskInput,
  output          maskSelect_valid,
  output [2:0]    maskSelect_bits,
  input           memRequest_ready,
  output          memRequest_valid,
  output [1023:0] memRequest_bits_data,
  output [127:0]  memRequest_bits_mask,
  output [3:0]    memRequest_bits_index,
  output [31:0]   memRequest_bits_address,
  output          status_idle,
                  status_last,
  output [2:0]    status_instructionIndex,
  output          status_changeMaskGroup,
  output [31:0]   status_startAddress,
                  status_endAddress,
  input           vrfReadDataPorts_0_ready,
  output          vrfReadDataPorts_0_valid,
  output [4:0]    vrfReadDataPorts_0_bits_vs,
  output [2:0]    vrfReadDataPorts_0_bits_instructionIndex,
  input           vrfReadDataPorts_1_ready,
  output          vrfReadDataPorts_1_valid,
  output [4:0]    vrfReadDataPorts_1_bits_vs,
  output [2:0]    vrfReadDataPorts_1_bits_instructionIndex,
  input           vrfReadDataPorts_2_ready,
  output          vrfReadDataPorts_2_valid,
  output [4:0]    vrfReadDataPorts_2_bits_vs,
  output [2:0]    vrfReadDataPorts_2_bits_instructionIndex,
  input           vrfReadDataPorts_3_ready,
  output          vrfReadDataPorts_3_valid,
  output [4:0]    vrfReadDataPorts_3_bits_vs,
  output [2:0]    vrfReadDataPorts_3_bits_instructionIndex,
  input           vrfReadDataPorts_4_ready,
  output          vrfReadDataPorts_4_valid,
  output [4:0]    vrfReadDataPorts_4_bits_vs,
  output [2:0]    vrfReadDataPorts_4_bits_instructionIndex,
  input           vrfReadDataPorts_5_ready,
  output          vrfReadDataPorts_5_valid,
  output [4:0]    vrfReadDataPorts_5_bits_vs,
  output [2:0]    vrfReadDataPorts_5_bits_instructionIndex,
  input           vrfReadDataPorts_6_ready,
  output          vrfReadDataPorts_6_valid,
  output [4:0]    vrfReadDataPorts_6_bits_vs,
  output [2:0]    vrfReadDataPorts_6_bits_instructionIndex,
  input           vrfReadDataPorts_7_ready,
  output          vrfReadDataPorts_7_valid,
  output [4:0]    vrfReadDataPorts_7_bits_vs,
  output [2:0]    vrfReadDataPorts_7_bits_instructionIndex,
  input           vrfReadDataPorts_8_ready,
  output          vrfReadDataPorts_8_valid,
  output [4:0]    vrfReadDataPorts_8_bits_vs,
  output [2:0]    vrfReadDataPorts_8_bits_instructionIndex,
  input           vrfReadDataPorts_9_ready,
  output          vrfReadDataPorts_9_valid,
  output [4:0]    vrfReadDataPorts_9_bits_vs,
  output [2:0]    vrfReadDataPorts_9_bits_instructionIndex,
  input           vrfReadDataPorts_10_ready,
  output          vrfReadDataPorts_10_valid,
  output [4:0]    vrfReadDataPorts_10_bits_vs,
  output [2:0]    vrfReadDataPorts_10_bits_instructionIndex,
  input           vrfReadDataPorts_11_ready,
  output          vrfReadDataPorts_11_valid,
  output [4:0]    vrfReadDataPorts_11_bits_vs,
  output [2:0]    vrfReadDataPorts_11_bits_instructionIndex,
  input           vrfReadDataPorts_12_ready,
  output          vrfReadDataPorts_12_valid,
  output [4:0]    vrfReadDataPorts_12_bits_vs,
  output [2:0]    vrfReadDataPorts_12_bits_instructionIndex,
  input           vrfReadDataPorts_13_ready,
  output          vrfReadDataPorts_13_valid,
  output [4:0]    vrfReadDataPorts_13_bits_vs,
  output [2:0]    vrfReadDataPorts_13_bits_instructionIndex,
  input           vrfReadDataPorts_14_ready,
  output          vrfReadDataPorts_14_valid,
  output [4:0]    vrfReadDataPorts_14_bits_vs,
  output [2:0]    vrfReadDataPorts_14_bits_instructionIndex,
  input           vrfReadDataPorts_15_ready,
  output          vrfReadDataPorts_15_valid,
  output [4:0]    vrfReadDataPorts_15_bits_vs,
  output [2:0]    vrfReadDataPorts_15_bits_instructionIndex,
  input           vrfReadDataPorts_16_ready,
  output          vrfReadDataPorts_16_valid,
  output [4:0]    vrfReadDataPorts_16_bits_vs,
  output [2:0]    vrfReadDataPorts_16_bits_instructionIndex,
  input           vrfReadDataPorts_17_ready,
  output          vrfReadDataPorts_17_valid,
  output [4:0]    vrfReadDataPorts_17_bits_vs,
  output [2:0]    vrfReadDataPorts_17_bits_instructionIndex,
  input           vrfReadDataPorts_18_ready,
  output          vrfReadDataPorts_18_valid,
  output [4:0]    vrfReadDataPorts_18_bits_vs,
  output [2:0]    vrfReadDataPorts_18_bits_instructionIndex,
  input           vrfReadDataPorts_19_ready,
  output          vrfReadDataPorts_19_valid,
  output [4:0]    vrfReadDataPorts_19_bits_vs,
  output [2:0]    vrfReadDataPorts_19_bits_instructionIndex,
  input           vrfReadDataPorts_20_ready,
  output          vrfReadDataPorts_20_valid,
  output [4:0]    vrfReadDataPorts_20_bits_vs,
  output [2:0]    vrfReadDataPorts_20_bits_instructionIndex,
  input           vrfReadDataPorts_21_ready,
  output          vrfReadDataPorts_21_valid,
  output [4:0]    vrfReadDataPorts_21_bits_vs,
  output [2:0]    vrfReadDataPorts_21_bits_instructionIndex,
  input           vrfReadDataPorts_22_ready,
  output          vrfReadDataPorts_22_valid,
  output [4:0]    vrfReadDataPorts_22_bits_vs,
  output [2:0]    vrfReadDataPorts_22_bits_instructionIndex,
  input           vrfReadDataPorts_23_ready,
  output          vrfReadDataPorts_23_valid,
  output [4:0]    vrfReadDataPorts_23_bits_vs,
  output [2:0]    vrfReadDataPorts_23_bits_instructionIndex,
  input           vrfReadDataPorts_24_ready,
  output          vrfReadDataPorts_24_valid,
  output [4:0]    vrfReadDataPorts_24_bits_vs,
  output [2:0]    vrfReadDataPorts_24_bits_instructionIndex,
  input           vrfReadDataPorts_25_ready,
  output          vrfReadDataPorts_25_valid,
  output [4:0]    vrfReadDataPorts_25_bits_vs,
  output [2:0]    vrfReadDataPorts_25_bits_instructionIndex,
  input           vrfReadDataPorts_26_ready,
  output          vrfReadDataPorts_26_valid,
  output [4:0]    vrfReadDataPorts_26_bits_vs,
  output [2:0]    vrfReadDataPorts_26_bits_instructionIndex,
  input           vrfReadDataPorts_27_ready,
  output          vrfReadDataPorts_27_valid,
  output [4:0]    vrfReadDataPorts_27_bits_vs,
  output [2:0]    vrfReadDataPorts_27_bits_instructionIndex,
  input           vrfReadDataPorts_28_ready,
  output          vrfReadDataPorts_28_valid,
  output [4:0]    vrfReadDataPorts_28_bits_vs,
  output [2:0]    vrfReadDataPorts_28_bits_instructionIndex,
  input           vrfReadDataPorts_29_ready,
  output          vrfReadDataPorts_29_valid,
  output [4:0]    vrfReadDataPorts_29_bits_vs,
  output [2:0]    vrfReadDataPorts_29_bits_instructionIndex,
  input           vrfReadDataPorts_30_ready,
  output          vrfReadDataPorts_30_valid,
  output [4:0]    vrfReadDataPorts_30_bits_vs,
  output [2:0]    vrfReadDataPorts_30_bits_instructionIndex,
  input           vrfReadDataPorts_31_ready,
  output          vrfReadDataPorts_31_valid,
  output [4:0]    vrfReadDataPorts_31_bits_vs,
  output [2:0]    vrfReadDataPorts_31_bits_instructionIndex,
  input           vrfReadResults_0_valid,
  input  [31:0]   vrfReadResults_0_bits,
  input           vrfReadResults_1_valid,
  input  [31:0]   vrfReadResults_1_bits,
  input           vrfReadResults_2_valid,
  input  [31:0]   vrfReadResults_2_bits,
  input           vrfReadResults_3_valid,
  input  [31:0]   vrfReadResults_3_bits,
  input           vrfReadResults_4_valid,
  input  [31:0]   vrfReadResults_4_bits,
  input           vrfReadResults_5_valid,
  input  [31:0]   vrfReadResults_5_bits,
  input           vrfReadResults_6_valid,
  input  [31:0]   vrfReadResults_6_bits,
  input           vrfReadResults_7_valid,
  input  [31:0]   vrfReadResults_7_bits,
  input           vrfReadResults_8_valid,
  input  [31:0]   vrfReadResults_8_bits,
  input           vrfReadResults_9_valid,
  input  [31:0]   vrfReadResults_9_bits,
  input           vrfReadResults_10_valid,
  input  [31:0]   vrfReadResults_10_bits,
  input           vrfReadResults_11_valid,
  input  [31:0]   vrfReadResults_11_bits,
  input           vrfReadResults_12_valid,
  input  [31:0]   vrfReadResults_12_bits,
  input           vrfReadResults_13_valid,
  input  [31:0]   vrfReadResults_13_bits,
  input           vrfReadResults_14_valid,
  input  [31:0]   vrfReadResults_14_bits,
  input           vrfReadResults_15_valid,
  input  [31:0]   vrfReadResults_15_bits,
  input           vrfReadResults_16_valid,
  input  [31:0]   vrfReadResults_16_bits,
  input           vrfReadResults_17_valid,
  input  [31:0]   vrfReadResults_17_bits,
  input           vrfReadResults_18_valid,
  input  [31:0]   vrfReadResults_18_bits,
  input           vrfReadResults_19_valid,
  input  [31:0]   vrfReadResults_19_bits,
  input           vrfReadResults_20_valid,
  input  [31:0]   vrfReadResults_20_bits,
  input           vrfReadResults_21_valid,
  input  [31:0]   vrfReadResults_21_bits,
  input           vrfReadResults_22_valid,
  input  [31:0]   vrfReadResults_22_bits,
  input           vrfReadResults_23_valid,
  input  [31:0]   vrfReadResults_23_bits,
  input           vrfReadResults_24_valid,
  input  [31:0]   vrfReadResults_24_bits,
  input           vrfReadResults_25_valid,
  input  [31:0]   vrfReadResults_25_bits,
  input           vrfReadResults_26_valid,
  input  [31:0]   vrfReadResults_26_bits,
  input           vrfReadResults_27_valid,
  input  [31:0]   vrfReadResults_27_bits,
  input           vrfReadResults_28_valid,
  input  [31:0]   vrfReadResults_28_bits,
  input           vrfReadResults_29_valid,
  input  [31:0]   vrfReadResults_29_bits,
  input           vrfReadResults_30_valid,
  input  [31:0]   vrfReadResults_30_bits,
  input           vrfReadResults_31_valid,
  input  [31:0]   vrfReadResults_31_bits,
  input           storeResponse
);

  wire              _addressQueue_fifo_empty;
  wire              _addressQueue_fifo_full;
  wire              _addressQueue_fifo_error;
  wire              _vrfReadQueueVec_fifo_31_empty;
  wire              _vrfReadQueueVec_fifo_31_full;
  wire              _vrfReadQueueVec_fifo_31_error;
  wire [31:0]       _vrfReadQueueVec_fifo_31_data_out;
  wire              _vrfReadQueueVec_fifo_30_empty;
  wire              _vrfReadQueueVec_fifo_30_full;
  wire              _vrfReadQueueVec_fifo_30_error;
  wire [31:0]       _vrfReadQueueVec_fifo_30_data_out;
  wire              _vrfReadQueueVec_fifo_29_empty;
  wire              _vrfReadQueueVec_fifo_29_full;
  wire              _vrfReadQueueVec_fifo_29_error;
  wire [31:0]       _vrfReadQueueVec_fifo_29_data_out;
  wire              _vrfReadQueueVec_fifo_28_empty;
  wire              _vrfReadQueueVec_fifo_28_full;
  wire              _vrfReadQueueVec_fifo_28_error;
  wire [31:0]       _vrfReadQueueVec_fifo_28_data_out;
  wire              _vrfReadQueueVec_fifo_27_empty;
  wire              _vrfReadQueueVec_fifo_27_full;
  wire              _vrfReadQueueVec_fifo_27_error;
  wire [31:0]       _vrfReadQueueVec_fifo_27_data_out;
  wire              _vrfReadQueueVec_fifo_26_empty;
  wire              _vrfReadQueueVec_fifo_26_full;
  wire              _vrfReadQueueVec_fifo_26_error;
  wire [31:0]       _vrfReadQueueVec_fifo_26_data_out;
  wire              _vrfReadQueueVec_fifo_25_empty;
  wire              _vrfReadQueueVec_fifo_25_full;
  wire              _vrfReadQueueVec_fifo_25_error;
  wire [31:0]       _vrfReadQueueVec_fifo_25_data_out;
  wire              _vrfReadQueueVec_fifo_24_empty;
  wire              _vrfReadQueueVec_fifo_24_full;
  wire              _vrfReadQueueVec_fifo_24_error;
  wire [31:0]       _vrfReadQueueVec_fifo_24_data_out;
  wire              _vrfReadQueueVec_fifo_23_empty;
  wire              _vrfReadQueueVec_fifo_23_full;
  wire              _vrfReadQueueVec_fifo_23_error;
  wire [31:0]       _vrfReadQueueVec_fifo_23_data_out;
  wire              _vrfReadQueueVec_fifo_22_empty;
  wire              _vrfReadQueueVec_fifo_22_full;
  wire              _vrfReadQueueVec_fifo_22_error;
  wire [31:0]       _vrfReadQueueVec_fifo_22_data_out;
  wire              _vrfReadQueueVec_fifo_21_empty;
  wire              _vrfReadQueueVec_fifo_21_full;
  wire              _vrfReadQueueVec_fifo_21_error;
  wire [31:0]       _vrfReadQueueVec_fifo_21_data_out;
  wire              _vrfReadQueueVec_fifo_20_empty;
  wire              _vrfReadQueueVec_fifo_20_full;
  wire              _vrfReadQueueVec_fifo_20_error;
  wire [31:0]       _vrfReadQueueVec_fifo_20_data_out;
  wire              _vrfReadQueueVec_fifo_19_empty;
  wire              _vrfReadQueueVec_fifo_19_full;
  wire              _vrfReadQueueVec_fifo_19_error;
  wire [31:0]       _vrfReadQueueVec_fifo_19_data_out;
  wire              _vrfReadQueueVec_fifo_18_empty;
  wire              _vrfReadQueueVec_fifo_18_full;
  wire              _vrfReadQueueVec_fifo_18_error;
  wire [31:0]       _vrfReadQueueVec_fifo_18_data_out;
  wire              _vrfReadQueueVec_fifo_17_empty;
  wire              _vrfReadQueueVec_fifo_17_full;
  wire              _vrfReadQueueVec_fifo_17_error;
  wire [31:0]       _vrfReadQueueVec_fifo_17_data_out;
  wire              _vrfReadQueueVec_fifo_16_empty;
  wire              _vrfReadQueueVec_fifo_16_full;
  wire              _vrfReadQueueVec_fifo_16_error;
  wire [31:0]       _vrfReadQueueVec_fifo_16_data_out;
  wire              _vrfReadQueueVec_fifo_15_empty;
  wire              _vrfReadQueueVec_fifo_15_full;
  wire              _vrfReadQueueVec_fifo_15_error;
  wire [31:0]       _vrfReadQueueVec_fifo_15_data_out;
  wire              _vrfReadQueueVec_fifo_14_empty;
  wire              _vrfReadQueueVec_fifo_14_full;
  wire              _vrfReadQueueVec_fifo_14_error;
  wire [31:0]       _vrfReadQueueVec_fifo_14_data_out;
  wire              _vrfReadQueueVec_fifo_13_empty;
  wire              _vrfReadQueueVec_fifo_13_full;
  wire              _vrfReadQueueVec_fifo_13_error;
  wire [31:0]       _vrfReadQueueVec_fifo_13_data_out;
  wire              _vrfReadQueueVec_fifo_12_empty;
  wire              _vrfReadQueueVec_fifo_12_full;
  wire              _vrfReadQueueVec_fifo_12_error;
  wire [31:0]       _vrfReadQueueVec_fifo_12_data_out;
  wire              _vrfReadQueueVec_fifo_11_empty;
  wire              _vrfReadQueueVec_fifo_11_full;
  wire              _vrfReadQueueVec_fifo_11_error;
  wire [31:0]       _vrfReadQueueVec_fifo_11_data_out;
  wire              _vrfReadQueueVec_fifo_10_empty;
  wire              _vrfReadQueueVec_fifo_10_full;
  wire              _vrfReadQueueVec_fifo_10_error;
  wire [31:0]       _vrfReadQueueVec_fifo_10_data_out;
  wire              _vrfReadQueueVec_fifo_9_empty;
  wire              _vrfReadQueueVec_fifo_9_full;
  wire              _vrfReadQueueVec_fifo_9_error;
  wire [31:0]       _vrfReadQueueVec_fifo_9_data_out;
  wire              _vrfReadQueueVec_fifo_8_empty;
  wire              _vrfReadQueueVec_fifo_8_full;
  wire              _vrfReadQueueVec_fifo_8_error;
  wire [31:0]       _vrfReadQueueVec_fifo_8_data_out;
  wire              _vrfReadQueueVec_fifo_7_empty;
  wire              _vrfReadQueueVec_fifo_7_full;
  wire              _vrfReadQueueVec_fifo_7_error;
  wire [31:0]       _vrfReadQueueVec_fifo_7_data_out;
  wire              _vrfReadQueueVec_fifo_6_empty;
  wire              _vrfReadQueueVec_fifo_6_full;
  wire              _vrfReadQueueVec_fifo_6_error;
  wire [31:0]       _vrfReadQueueVec_fifo_6_data_out;
  wire              _vrfReadQueueVec_fifo_5_empty;
  wire              _vrfReadQueueVec_fifo_5_full;
  wire              _vrfReadQueueVec_fifo_5_error;
  wire [31:0]       _vrfReadQueueVec_fifo_5_data_out;
  wire              _vrfReadQueueVec_fifo_4_empty;
  wire              _vrfReadQueueVec_fifo_4_full;
  wire              _vrfReadQueueVec_fifo_4_error;
  wire [31:0]       _vrfReadQueueVec_fifo_4_data_out;
  wire              _vrfReadQueueVec_fifo_3_empty;
  wire              _vrfReadQueueVec_fifo_3_full;
  wire              _vrfReadQueueVec_fifo_3_error;
  wire [31:0]       _vrfReadQueueVec_fifo_3_data_out;
  wire              _vrfReadQueueVec_fifo_2_empty;
  wire              _vrfReadQueueVec_fifo_2_full;
  wire              _vrfReadQueueVec_fifo_2_error;
  wire [31:0]       _vrfReadQueueVec_fifo_2_data_out;
  wire              _vrfReadQueueVec_fifo_1_empty;
  wire              _vrfReadQueueVec_fifo_1_full;
  wire              _vrfReadQueueVec_fifo_1_error;
  wire [31:0]       _vrfReadQueueVec_fifo_1_data_out;
  wire              _vrfReadQueueVec_fifo_empty;
  wire              _vrfReadQueueVec_fifo_full;
  wire              _vrfReadQueueVec_fifo_error;
  wire [31:0]       _vrfReadQueueVec_fifo_data_out;
  wire              addressQueue_almostFull;
  wire              addressQueue_almostEmpty;
  wire              vrfReadQueueVec_31_almostFull;
  wire              vrfReadQueueVec_31_almostEmpty;
  wire              vrfReadQueueVec_30_almostFull;
  wire              vrfReadQueueVec_30_almostEmpty;
  wire              vrfReadQueueVec_29_almostFull;
  wire              vrfReadQueueVec_29_almostEmpty;
  wire              vrfReadQueueVec_28_almostFull;
  wire              vrfReadQueueVec_28_almostEmpty;
  wire              vrfReadQueueVec_27_almostFull;
  wire              vrfReadQueueVec_27_almostEmpty;
  wire              vrfReadQueueVec_26_almostFull;
  wire              vrfReadQueueVec_26_almostEmpty;
  wire              vrfReadQueueVec_25_almostFull;
  wire              vrfReadQueueVec_25_almostEmpty;
  wire              vrfReadQueueVec_24_almostFull;
  wire              vrfReadQueueVec_24_almostEmpty;
  wire              vrfReadQueueVec_23_almostFull;
  wire              vrfReadQueueVec_23_almostEmpty;
  wire              vrfReadQueueVec_22_almostFull;
  wire              vrfReadQueueVec_22_almostEmpty;
  wire              vrfReadQueueVec_21_almostFull;
  wire              vrfReadQueueVec_21_almostEmpty;
  wire              vrfReadQueueVec_20_almostFull;
  wire              vrfReadQueueVec_20_almostEmpty;
  wire              vrfReadQueueVec_19_almostFull;
  wire              vrfReadQueueVec_19_almostEmpty;
  wire              vrfReadQueueVec_18_almostFull;
  wire              vrfReadQueueVec_18_almostEmpty;
  wire              vrfReadQueueVec_17_almostFull;
  wire              vrfReadQueueVec_17_almostEmpty;
  wire              vrfReadQueueVec_16_almostFull;
  wire              vrfReadQueueVec_16_almostEmpty;
  wire              vrfReadQueueVec_15_almostFull;
  wire              vrfReadQueueVec_15_almostEmpty;
  wire              vrfReadQueueVec_14_almostFull;
  wire              vrfReadQueueVec_14_almostEmpty;
  wire              vrfReadQueueVec_13_almostFull;
  wire              vrfReadQueueVec_13_almostEmpty;
  wire              vrfReadQueueVec_12_almostFull;
  wire              vrfReadQueueVec_12_almostEmpty;
  wire              vrfReadQueueVec_11_almostFull;
  wire              vrfReadQueueVec_11_almostEmpty;
  wire              vrfReadQueueVec_10_almostFull;
  wire              vrfReadQueueVec_10_almostEmpty;
  wire              vrfReadQueueVec_9_almostFull;
  wire              vrfReadQueueVec_9_almostEmpty;
  wire              vrfReadQueueVec_8_almostFull;
  wire              vrfReadQueueVec_8_almostEmpty;
  wire              vrfReadQueueVec_7_almostFull;
  wire              vrfReadQueueVec_7_almostEmpty;
  wire              vrfReadQueueVec_6_almostFull;
  wire              vrfReadQueueVec_6_almostEmpty;
  wire              vrfReadQueueVec_5_almostFull;
  wire              vrfReadQueueVec_5_almostEmpty;
  wire              vrfReadQueueVec_4_almostFull;
  wire              vrfReadQueueVec_4_almostEmpty;
  wire              vrfReadQueueVec_3_almostFull;
  wire              vrfReadQueueVec_3_almostEmpty;
  wire              vrfReadQueueVec_2_almostFull;
  wire              vrfReadQueueVec_2_almostEmpty;
  wire              vrfReadQueueVec_1_almostFull;
  wire              vrfReadQueueVec_1_almostEmpty;
  wire              vrfReadQueueVec_0_almostFull;
  wire              vrfReadQueueVec_0_almostEmpty;
  wire              memRequest_ready_0 = memRequest_ready;
  wire              vrfReadDataPorts_0_ready_0 = vrfReadDataPorts_0_ready;
  wire              vrfReadDataPorts_1_ready_0 = vrfReadDataPorts_1_ready;
  wire              vrfReadDataPorts_2_ready_0 = vrfReadDataPorts_2_ready;
  wire              vrfReadDataPorts_3_ready_0 = vrfReadDataPorts_3_ready;
  wire              vrfReadDataPorts_4_ready_0 = vrfReadDataPorts_4_ready;
  wire              vrfReadDataPorts_5_ready_0 = vrfReadDataPorts_5_ready;
  wire              vrfReadDataPorts_6_ready_0 = vrfReadDataPorts_6_ready;
  wire              vrfReadDataPorts_7_ready_0 = vrfReadDataPorts_7_ready;
  wire              vrfReadDataPorts_8_ready_0 = vrfReadDataPorts_8_ready;
  wire              vrfReadDataPorts_9_ready_0 = vrfReadDataPorts_9_ready;
  wire              vrfReadDataPorts_10_ready_0 = vrfReadDataPorts_10_ready;
  wire              vrfReadDataPorts_11_ready_0 = vrfReadDataPorts_11_ready;
  wire              vrfReadDataPorts_12_ready_0 = vrfReadDataPorts_12_ready;
  wire              vrfReadDataPorts_13_ready_0 = vrfReadDataPorts_13_ready;
  wire              vrfReadDataPorts_14_ready_0 = vrfReadDataPorts_14_ready;
  wire              vrfReadDataPorts_15_ready_0 = vrfReadDataPorts_15_ready;
  wire              vrfReadDataPorts_16_ready_0 = vrfReadDataPorts_16_ready;
  wire              vrfReadDataPorts_17_ready_0 = vrfReadDataPorts_17_ready;
  wire              vrfReadDataPorts_18_ready_0 = vrfReadDataPorts_18_ready;
  wire              vrfReadDataPorts_19_ready_0 = vrfReadDataPorts_19_ready;
  wire              vrfReadDataPorts_20_ready_0 = vrfReadDataPorts_20_ready;
  wire              vrfReadDataPorts_21_ready_0 = vrfReadDataPorts_21_ready;
  wire              vrfReadDataPorts_22_ready_0 = vrfReadDataPorts_22_ready;
  wire              vrfReadDataPorts_23_ready_0 = vrfReadDataPorts_23_ready;
  wire              vrfReadDataPorts_24_ready_0 = vrfReadDataPorts_24_ready;
  wire              vrfReadDataPorts_25_ready_0 = vrfReadDataPorts_25_ready;
  wire              vrfReadDataPorts_26_ready_0 = vrfReadDataPorts_26_ready;
  wire              vrfReadDataPorts_27_ready_0 = vrfReadDataPorts_27_ready;
  wire              vrfReadDataPorts_28_ready_0 = vrfReadDataPorts_28_ready;
  wire              vrfReadDataPorts_29_ready_0 = vrfReadDataPorts_29_ready;
  wire              vrfReadDataPorts_30_ready_0 = vrfReadDataPorts_30_ready;
  wire              vrfReadDataPorts_31_ready_0 = vrfReadDataPorts_31_ready;
  wire              vrfReadQueueVec_0_enq_valid = vrfReadResults_0_valid;
  wire [31:0]       vrfReadQueueVec_0_enq_bits = vrfReadResults_0_bits;
  wire              vrfReadQueueVec_1_enq_valid = vrfReadResults_1_valid;
  wire [31:0]       vrfReadQueueVec_1_enq_bits = vrfReadResults_1_bits;
  wire              vrfReadQueueVec_2_enq_valid = vrfReadResults_2_valid;
  wire [31:0]       vrfReadQueueVec_2_enq_bits = vrfReadResults_2_bits;
  wire              vrfReadQueueVec_3_enq_valid = vrfReadResults_3_valid;
  wire [31:0]       vrfReadQueueVec_3_enq_bits = vrfReadResults_3_bits;
  wire              vrfReadQueueVec_4_enq_valid = vrfReadResults_4_valid;
  wire [31:0]       vrfReadQueueVec_4_enq_bits = vrfReadResults_4_bits;
  wire              vrfReadQueueVec_5_enq_valid = vrfReadResults_5_valid;
  wire [31:0]       vrfReadQueueVec_5_enq_bits = vrfReadResults_5_bits;
  wire              vrfReadQueueVec_6_enq_valid = vrfReadResults_6_valid;
  wire [31:0]       vrfReadQueueVec_6_enq_bits = vrfReadResults_6_bits;
  wire              vrfReadQueueVec_7_enq_valid = vrfReadResults_7_valid;
  wire [31:0]       vrfReadQueueVec_7_enq_bits = vrfReadResults_7_bits;
  wire              vrfReadQueueVec_8_enq_valid = vrfReadResults_8_valid;
  wire [31:0]       vrfReadQueueVec_8_enq_bits = vrfReadResults_8_bits;
  wire              vrfReadQueueVec_9_enq_valid = vrfReadResults_9_valid;
  wire [31:0]       vrfReadQueueVec_9_enq_bits = vrfReadResults_9_bits;
  wire              vrfReadQueueVec_10_enq_valid = vrfReadResults_10_valid;
  wire [31:0]       vrfReadQueueVec_10_enq_bits = vrfReadResults_10_bits;
  wire              vrfReadQueueVec_11_enq_valid = vrfReadResults_11_valid;
  wire [31:0]       vrfReadQueueVec_11_enq_bits = vrfReadResults_11_bits;
  wire              vrfReadQueueVec_12_enq_valid = vrfReadResults_12_valid;
  wire [31:0]       vrfReadQueueVec_12_enq_bits = vrfReadResults_12_bits;
  wire              vrfReadQueueVec_13_enq_valid = vrfReadResults_13_valid;
  wire [31:0]       vrfReadQueueVec_13_enq_bits = vrfReadResults_13_bits;
  wire              vrfReadQueueVec_14_enq_valid = vrfReadResults_14_valid;
  wire [31:0]       vrfReadQueueVec_14_enq_bits = vrfReadResults_14_bits;
  wire              vrfReadQueueVec_15_enq_valid = vrfReadResults_15_valid;
  wire [31:0]       vrfReadQueueVec_15_enq_bits = vrfReadResults_15_bits;
  wire              vrfReadQueueVec_16_enq_valid = vrfReadResults_16_valid;
  wire [31:0]       vrfReadQueueVec_16_enq_bits = vrfReadResults_16_bits;
  wire              vrfReadQueueVec_17_enq_valid = vrfReadResults_17_valid;
  wire [31:0]       vrfReadQueueVec_17_enq_bits = vrfReadResults_17_bits;
  wire              vrfReadQueueVec_18_enq_valid = vrfReadResults_18_valid;
  wire [31:0]       vrfReadQueueVec_18_enq_bits = vrfReadResults_18_bits;
  wire              vrfReadQueueVec_19_enq_valid = vrfReadResults_19_valid;
  wire [31:0]       vrfReadQueueVec_19_enq_bits = vrfReadResults_19_bits;
  wire              vrfReadQueueVec_20_enq_valid = vrfReadResults_20_valid;
  wire [31:0]       vrfReadQueueVec_20_enq_bits = vrfReadResults_20_bits;
  wire              vrfReadQueueVec_21_enq_valid = vrfReadResults_21_valid;
  wire [31:0]       vrfReadQueueVec_21_enq_bits = vrfReadResults_21_bits;
  wire              vrfReadQueueVec_22_enq_valid = vrfReadResults_22_valid;
  wire [31:0]       vrfReadQueueVec_22_enq_bits = vrfReadResults_22_bits;
  wire              vrfReadQueueVec_23_enq_valid = vrfReadResults_23_valid;
  wire [31:0]       vrfReadQueueVec_23_enq_bits = vrfReadResults_23_bits;
  wire              vrfReadQueueVec_24_enq_valid = vrfReadResults_24_valid;
  wire [31:0]       vrfReadQueueVec_24_enq_bits = vrfReadResults_24_bits;
  wire              vrfReadQueueVec_25_enq_valid = vrfReadResults_25_valid;
  wire [31:0]       vrfReadQueueVec_25_enq_bits = vrfReadResults_25_bits;
  wire              vrfReadQueueVec_26_enq_valid = vrfReadResults_26_valid;
  wire [31:0]       vrfReadQueueVec_26_enq_bits = vrfReadResults_26_bits;
  wire              vrfReadQueueVec_27_enq_valid = vrfReadResults_27_valid;
  wire [31:0]       vrfReadQueueVec_27_enq_bits = vrfReadResults_27_bits;
  wire              vrfReadQueueVec_28_enq_valid = vrfReadResults_28_valid;
  wire [31:0]       vrfReadQueueVec_28_enq_bits = vrfReadResults_28_bits;
  wire              vrfReadQueueVec_29_enq_valid = vrfReadResults_29_valid;
  wire [31:0]       vrfReadQueueVec_29_enq_bits = vrfReadResults_29_bits;
  wire              vrfReadQueueVec_30_enq_valid = vrfReadResults_30_valid;
  wire [31:0]       vrfReadQueueVec_30_enq_bits = vrfReadResults_30_bits;
  wire              vrfReadQueueVec_31_enq_valid = vrfReadResults_31_valid;
  wire [31:0]       vrfReadQueueVec_31_enq_bits = vrfReadResults_31_bits;
  wire              addressQueue_deq_ready = storeResponse;
  wire [1:0]        accessStateCheck_lo_lo_lo_lo = 2'h0;
  wire [1:0]        accessStateCheck_lo_lo_lo_hi = 2'h0;
  wire [1:0]        accessStateCheck_lo_lo_hi_lo = 2'h0;
  wire [1:0]        accessStateCheck_lo_lo_hi_hi = 2'h0;
  wire [1:0]        accessStateCheck_lo_hi_lo_lo = 2'h0;
  wire [1:0]        accessStateCheck_lo_hi_lo_hi = 2'h0;
  wire [1:0]        accessStateCheck_lo_hi_hi_lo = 2'h0;
  wire [1:0]        accessStateCheck_lo_hi_hi_hi = 2'h0;
  wire [1:0]        accessStateCheck_hi_lo_lo_lo = 2'h0;
  wire [1:0]        accessStateCheck_hi_lo_lo_hi = 2'h0;
  wire [1:0]        accessStateCheck_hi_lo_hi_lo = 2'h0;
  wire [1:0]        accessStateCheck_hi_lo_hi_hi = 2'h0;
  wire [1:0]        accessStateCheck_hi_hi_lo_lo = 2'h0;
  wire [1:0]        accessStateCheck_hi_hi_lo_hi = 2'h0;
  wire [1:0]        accessStateCheck_hi_hi_hi_lo = 2'h0;
  wire [1:0]        accessStateCheck_hi_hi_hi_hi = 2'h0;
  wire [3:0]        accessStateCheck_lo_lo_lo = 4'h0;
  wire [3:0]        accessStateCheck_lo_lo_hi = 4'h0;
  wire [3:0]        accessStateCheck_lo_hi_lo = 4'h0;
  wire [3:0]        accessStateCheck_lo_hi_hi = 4'h0;
  wire [3:0]        accessStateCheck_hi_lo_lo = 4'h0;
  wire [3:0]        accessStateCheck_hi_lo_hi = 4'h0;
  wire [3:0]        accessStateCheck_hi_hi_lo = 4'h0;
  wire [3:0]        accessStateCheck_hi_hi_hi = 4'h0;
  wire [7:0]        accessStateCheck_lo_lo = 8'h0;
  wire [7:0]        accessStateCheck_lo_hi = 8'h0;
  wire [7:0]        accessStateCheck_hi_lo = 8'h0;
  wire [7:0]        accessStateCheck_hi_hi = 8'h0;
  wire [15:0]       accessStateCheck_lo = 16'h0;
  wire [15:0]       accessStateCheck_hi = 16'h0;
  wire              accessStateCheck = 1'h1;
  wire              accessStateUpdate_0 = 1'h0;
  wire              accessStateUpdate_1 = 1'h0;
  wire              accessStateUpdate_2 = 1'h0;
  wire              accessStateUpdate_3 = 1'h0;
  wire              accessStateUpdate_4 = 1'h0;
  wire              accessStateUpdate_5 = 1'h0;
  wire              accessStateUpdate_6 = 1'h0;
  wire              accessStateUpdate_7 = 1'h0;
  wire              accessStateUpdate_8 = 1'h0;
  wire              accessStateUpdate_9 = 1'h0;
  wire              accessStateUpdate_10 = 1'h0;
  wire              accessStateUpdate_11 = 1'h0;
  wire              accessStateUpdate_12 = 1'h0;
  wire              accessStateUpdate_13 = 1'h0;
  wire              accessStateUpdate_14 = 1'h0;
  wire              accessStateUpdate_15 = 1'h0;
  wire              accessStateUpdate_16 = 1'h0;
  wire              accessStateUpdate_17 = 1'h0;
  wire              accessStateUpdate_18 = 1'h0;
  wire              accessStateUpdate_19 = 1'h0;
  wire              accessStateUpdate_20 = 1'h0;
  wire              accessStateUpdate_21 = 1'h0;
  wire              accessStateUpdate_22 = 1'h0;
  wire              accessStateUpdate_23 = 1'h0;
  wire              accessStateUpdate_24 = 1'h0;
  wire              accessStateUpdate_25 = 1'h0;
  wire              accessStateUpdate_26 = 1'h0;
  wire              accessStateUpdate_27 = 1'h0;
  wire              accessStateUpdate_28 = 1'h0;
  wire              accessStateUpdate_29 = 1'h0;
  wire              accessStateUpdate_30 = 1'h0;
  wire              accessStateUpdate_31 = 1'h0;
  wire [4095:0]     hi = 4096'h0;
  wire [4095:0]     hi_1 = 4096'h0;
  wire [4095:0]     hi_2 = 4096'h0;
  wire [4095:0]     hi_3 = 4096'h0;
  wire [4095:0]     hi_8 = 4096'h0;
  wire [4095:0]     hi_9 = 4096'h0;
  wire [4095:0]     hi_10 = 4096'h0;
  wire [4095:0]     hi_11 = 4096'h0;
  wire [4095:0]     hi_16 = 4096'h0;
  wire [4095:0]     hi_17 = 4096'h0;
  wire [4095:0]     hi_18 = 4096'h0;
  wire [4095:0]     hi_19 = 4096'h0;
  wire [2047:0]     lo_hi = 2048'h0;
  wire [2047:0]     hi_lo = 2048'h0;
  wire [2047:0]     hi_hi = 2048'h0;
  wire [2047:0]     lo_hi_1 = 2048'h0;
  wire [2047:0]     hi_lo_1 = 2048'h0;
  wire [2047:0]     hi_hi_1 = 2048'h0;
  wire [2047:0]     hi_lo_2 = 2048'h0;
  wire [2047:0]     hi_hi_2 = 2048'h0;
  wire [2047:0]     hi_lo_3 = 2048'h0;
  wire [2047:0]     hi_hi_3 = 2048'h0;
  wire [2047:0]     hi_hi_4 = 2048'h0;
  wire [2047:0]     hi_hi_5 = 2048'h0;
  wire [2047:0]     lo_hi_8 = 2048'h0;
  wire [2047:0]     hi_lo_8 = 2048'h0;
  wire [2047:0]     hi_hi_8 = 2048'h0;
  wire [2047:0]     lo_hi_9 = 2048'h0;
  wire [2047:0]     hi_lo_9 = 2048'h0;
  wire [2047:0]     hi_hi_9 = 2048'h0;
  wire [2047:0]     hi_lo_10 = 2048'h0;
  wire [2047:0]     hi_hi_10 = 2048'h0;
  wire [2047:0]     hi_lo_11 = 2048'h0;
  wire [2047:0]     hi_hi_11 = 2048'h0;
  wire [2047:0]     hi_hi_12 = 2048'h0;
  wire [2047:0]     hi_hi_13 = 2048'h0;
  wire [2047:0]     lo_hi_16 = 2048'h0;
  wire [2047:0]     hi_lo_16 = 2048'h0;
  wire [2047:0]     hi_hi_16 = 2048'h0;
  wire [2047:0]     lo_hi_17 = 2048'h0;
  wire [2047:0]     hi_lo_17 = 2048'h0;
  wire [2047:0]     hi_hi_17 = 2048'h0;
  wire [2047:0]     hi_lo_18 = 2048'h0;
  wire [2047:0]     hi_hi_18 = 2048'h0;
  wire [2047:0]     hi_lo_19 = 2048'h0;
  wire [2047:0]     hi_hi_19 = 2048'h0;
  wire [2047:0]     hi_hi_20 = 2048'h0;
  wire [2047:0]     hi_hi_21 = 2048'h0;
  wire [1023:0]     res_1 = 1024'h0;
  wire [1023:0]     res_2 = 1024'h0;
  wire [1023:0]     res_3 = 1024'h0;
  wire [1023:0]     res_4 = 1024'h0;
  wire [1023:0]     res_5 = 1024'h0;
  wire [1023:0]     res_6 = 1024'h0;
  wire [1023:0]     res_7 = 1024'h0;
  wire [1023:0]     res_10 = 1024'h0;
  wire [1023:0]     res_11 = 1024'h0;
  wire [1023:0]     res_12 = 1024'h0;
  wire [1023:0]     res_13 = 1024'h0;
  wire [1023:0]     res_14 = 1024'h0;
  wire [1023:0]     res_15 = 1024'h0;
  wire [1023:0]     res_19 = 1024'h0;
  wire [1023:0]     res_20 = 1024'h0;
  wire [1023:0]     res_21 = 1024'h0;
  wire [1023:0]     res_22 = 1024'h0;
  wire [1023:0]     res_23 = 1024'h0;
  wire [1023:0]     res_28 = 1024'h0;
  wire [1023:0]     res_29 = 1024'h0;
  wire [1023:0]     res_30 = 1024'h0;
  wire [1023:0]     res_31 = 1024'h0;
  wire [1023:0]     res_37 = 1024'h0;
  wire [1023:0]     res_38 = 1024'h0;
  wire [1023:0]     res_39 = 1024'h0;
  wire [1023:0]     res_46 = 1024'h0;
  wire [1023:0]     res_47 = 1024'h0;
  wire [1023:0]     res_55 = 1024'h0;
  wire [1023:0]     res_65 = 1024'h0;
  wire [1023:0]     res_66 = 1024'h0;
  wire [1023:0]     res_67 = 1024'h0;
  wire [1023:0]     res_68 = 1024'h0;
  wire [1023:0]     res_69 = 1024'h0;
  wire [1023:0]     res_70 = 1024'h0;
  wire [1023:0]     res_71 = 1024'h0;
  wire [1023:0]     res_74 = 1024'h0;
  wire [1023:0]     res_75 = 1024'h0;
  wire [1023:0]     res_76 = 1024'h0;
  wire [1023:0]     res_77 = 1024'h0;
  wire [1023:0]     res_78 = 1024'h0;
  wire [1023:0]     res_79 = 1024'h0;
  wire [1023:0]     res_83 = 1024'h0;
  wire [1023:0]     res_84 = 1024'h0;
  wire [1023:0]     res_85 = 1024'h0;
  wire [1023:0]     res_86 = 1024'h0;
  wire [1023:0]     res_87 = 1024'h0;
  wire [1023:0]     res_92 = 1024'h0;
  wire [1023:0]     res_93 = 1024'h0;
  wire [1023:0]     res_94 = 1024'h0;
  wire [1023:0]     res_95 = 1024'h0;
  wire [1023:0]     res_101 = 1024'h0;
  wire [1023:0]     res_102 = 1024'h0;
  wire [1023:0]     res_103 = 1024'h0;
  wire [1023:0]     res_110 = 1024'h0;
  wire [1023:0]     res_111 = 1024'h0;
  wire [1023:0]     res_119 = 1024'h0;
  wire [1023:0]     res_129 = 1024'h0;
  wire [1023:0]     res_130 = 1024'h0;
  wire [1023:0]     res_131 = 1024'h0;
  wire [1023:0]     res_132 = 1024'h0;
  wire [1023:0]     res_133 = 1024'h0;
  wire [1023:0]     res_134 = 1024'h0;
  wire [1023:0]     res_135 = 1024'h0;
  wire [1023:0]     res_138 = 1024'h0;
  wire [1023:0]     res_139 = 1024'h0;
  wire [1023:0]     res_140 = 1024'h0;
  wire [1023:0]     res_141 = 1024'h0;
  wire [1023:0]     res_142 = 1024'h0;
  wire [1023:0]     res_143 = 1024'h0;
  wire [1023:0]     res_147 = 1024'h0;
  wire [1023:0]     res_148 = 1024'h0;
  wire [1023:0]     res_149 = 1024'h0;
  wire [1023:0]     res_150 = 1024'h0;
  wire [1023:0]     res_151 = 1024'h0;
  wire [1023:0]     res_156 = 1024'h0;
  wire [1023:0]     res_157 = 1024'h0;
  wire [1023:0]     res_158 = 1024'h0;
  wire [1023:0]     res_159 = 1024'h0;
  wire [1023:0]     res_165 = 1024'h0;
  wire [1023:0]     res_166 = 1024'h0;
  wire [1023:0]     res_167 = 1024'h0;
  wire [1023:0]     res_174 = 1024'h0;
  wire [1023:0]     res_175 = 1024'h0;
  wire [1023:0]     res_183 = 1024'h0;
  wire [1:0]        vrfReadDataPorts_0_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_1_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_2_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_3_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_4_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_5_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_6_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_7_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_8_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_9_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_10_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_11_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_12_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_13_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_14_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_15_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_16_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_17_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_18_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_19_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_20_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_21_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_22_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_23_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_24_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_25_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_26_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_27_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_28_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_29_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_30_bits_readSource = 2'h2;
  wire [1:0]        vrfReadDataPorts_31_bits_readSource = 2'h2;
  wire [31:0]       alignedDequeueAddress;
  reg  [2:0]        lsuRequestReg_instructionInformation_nf;
  reg               lsuRequestReg_instructionInformation_mew;
  reg  [1:0]        lsuRequestReg_instructionInformation_mop;
  reg  [4:0]        lsuRequestReg_instructionInformation_lumop;
  reg  [1:0]        lsuRequestReg_instructionInformation_eew;
  reg  [4:0]        lsuRequestReg_instructionInformation_vs3;
  reg               lsuRequestReg_instructionInformation_isStore;
  reg               lsuRequestReg_instructionInformation_maskedLoadStore;
  reg  [31:0]       lsuRequestReg_rs1Data;
  reg  [31:0]       lsuRequestReg_rs2Data;
  reg  [2:0]        lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_0_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_1_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_2_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_3_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_4_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_5_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_6_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_7_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_8_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_9_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_10_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_11_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_12_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_13_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_14_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_15_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_16_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_17_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_18_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_19_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_20_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_21_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_22_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_23_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_24_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_25_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_26_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_27_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_28_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_29_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_30_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  wire [2:0]        vrfReadDataPorts_31_bits_instructionIndex_0 = lsuRequestReg_instructionIndex;
  reg  [10:0]       csrInterfaceReg_vl;
  reg  [10:0]       csrInterfaceReg_vStart;
  reg  [2:0]        csrInterfaceReg_vlmul;
  reg  [1:0]        csrInterfaceReg_vSew;
  reg  [1:0]        csrInterfaceReg_vxrm;
  reg               csrInterfaceReg_vta;
  reg               csrInterfaceReg_vma;
  reg               requestFireNext;
  reg  [1:0]        dataEEW;
  wire [3:0]        _dataEEWOH_T = 4'h1 << dataEEW;
  wire [2:0]        dataEEWOH = _dataEEWOH_T[2:0];
  wire              isMaskType = lsuRequest_valid ? lsuRequest_bits_instructionInformation_maskedLoadStore : lsuRequestReg_instructionInformation_maskedLoadStore;
  wire [127:0]      maskAmend = isMaskType ? maskInput : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
  reg  [127:0]      maskReg;
  wire [127:0]      _lastMaskAmend_T_1 = 128'h1 << csrInterface_vl[6:0];
  wire [125:0]      _GEN = _lastMaskAmend_T_1[126:1] | _lastMaskAmend_T_1[127:2];
  wire [124:0]      _GEN_0 = _GEN[124:0] | {_lastMaskAmend_T_1[127], _GEN[125:2]};
  wire [122:0]      _GEN_1 = _GEN_0[122:0] | {_lastMaskAmend_T_1[127], _GEN[125], _GEN_0[124:4]};
  wire [118:0]      _GEN_2 = _GEN_1[118:0] | {_lastMaskAmend_T_1[127], _GEN[125], _GEN_0[124:123], _GEN_1[122:8]};
  wire [110:0]      _GEN_3 = _GEN_2[110:0] | {_lastMaskAmend_T_1[127], _GEN[125], _GEN_0[124:123], _GEN_1[122:119], _GEN_2[118:16]};
  wire [94:0]       _GEN_4 = _GEN_3[94:0] | {_lastMaskAmend_T_1[127], _GEN[125], _GEN_0[124:123], _GEN_1[122:119], _GEN_2[118:111], _GEN_3[110:32]};
  wire [126:0]      lastMaskAmend =
    {_lastMaskAmend_T_1[127],
     _GEN[125],
     _GEN_0[124:123],
     _GEN_1[122:119],
     _GEN_2[118:111],
     _GEN_3[110:95],
     _GEN_4[94:63],
     _GEN_4[62:0] | {_lastMaskAmend_T_1[127], _GEN[125], _GEN_0[124:123], _GEN_1[122:119], _GEN_2[118:111], _GEN_3[110:95], _GEN_4[94:64]}};
  reg               needAmend;
  reg  [126:0]      lastMaskAmendReg;
  wire [1:0]        countEndForGroup = {1'h0, dataEEWOH[1]} | {2{dataEEWOH[2]}};
  reg  [2:0]        maskGroupCounter;
  wire [2:0]        nextMaskGroup = maskGroupCounter + 3'h1;
  reg  [1:0]        maskCounterInGroup;
  wire [1:0]        nextMaskCount = maskCounterInGroup + 2'h1;
  wire              isLastDataGroup = maskCounterInGroup == countEndForGroup;
  wire [2:0]        _maskSelect_bits_output = lsuRequest_valid ? 3'h0 : nextMaskGroup;
  reg               isLastMaskGroup;
  wire [127:0]      maskWire = maskReg & (needAmend & isLastMaskGroup ? {1'h0, lastMaskAmendReg} : 128'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF);
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_lo_lo = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_lo_hi = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo = {maskForGroupWire_lo_lo_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_hi_lo = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_hi_hi = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi = {maskForGroupWire_lo_lo_lo_lo_hi_hi, maskForGroupWire_lo_lo_lo_lo_hi_lo};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo = {maskForGroupWire_lo_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_lo_lo = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_lo_hi = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo = {maskForGroupWire_lo_lo_lo_hi_lo_hi, maskForGroupWire_lo_lo_lo_hi_lo_lo};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_hi_lo = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_hi_hi = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi = {maskForGroupWire_lo_lo_lo_hi_hi_hi, maskForGroupWire_lo_lo_lo_hi_hi_lo};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi = {maskForGroupWire_lo_lo_lo_hi_hi, maskForGroupWire_lo_lo_lo_hi_lo};
  wire [31:0]       maskForGroupWire_lo_lo_lo = {maskForGroupWire_lo_lo_lo_hi, maskForGroupWire_lo_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_lo_lo = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_lo_hi = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo = {maskForGroupWire_lo_lo_hi_lo_lo_hi, maskForGroupWire_lo_lo_hi_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_hi_lo = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_hi_hi = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi = {maskForGroupWire_lo_lo_hi_lo_hi_hi, maskForGroupWire_lo_lo_hi_lo_hi_lo};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo = {maskForGroupWire_lo_lo_hi_lo_hi, maskForGroupWire_lo_lo_hi_lo_lo};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_lo_lo = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_lo_hi = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo = {maskForGroupWire_lo_lo_hi_hi_lo_hi, maskForGroupWire_lo_lo_hi_hi_lo_lo};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_hi_lo = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_hi_hi = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi = {maskForGroupWire_lo_lo_hi_hi_hi_hi, maskForGroupWire_lo_lo_hi_hi_hi_lo};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi = {maskForGroupWire_lo_lo_hi_hi_hi, maskForGroupWire_lo_lo_hi_hi_lo};
  wire [31:0]       maskForGroupWire_lo_lo_hi = {maskForGroupWire_lo_lo_hi_hi, maskForGroupWire_lo_lo_hi_lo};
  wire [63:0]       maskForGroupWire_lo_lo = {maskForGroupWire_lo_lo_hi, maskForGroupWire_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_lo_lo = {{2{maskWire[33]}}, {2{maskWire[32]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_lo_hi = {{2{maskWire[35]}}, {2{maskWire[34]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo = {maskForGroupWire_lo_hi_lo_lo_lo_hi, maskForGroupWire_lo_hi_lo_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_hi_lo = {{2{maskWire[37]}}, {2{maskWire[36]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_hi_hi = {{2{maskWire[39]}}, {2{maskWire[38]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi = {maskForGroupWire_lo_hi_lo_lo_hi_hi, maskForGroupWire_lo_hi_lo_lo_hi_lo};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo = {maskForGroupWire_lo_hi_lo_lo_hi, maskForGroupWire_lo_hi_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_lo_lo = {{2{maskWire[41]}}, {2{maskWire[40]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_lo_hi = {{2{maskWire[43]}}, {2{maskWire[42]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo = {maskForGroupWire_lo_hi_lo_hi_lo_hi, maskForGroupWire_lo_hi_lo_hi_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_hi_lo = {{2{maskWire[45]}}, {2{maskWire[44]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_hi_hi = {{2{maskWire[47]}}, {2{maskWire[46]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi = {maskForGroupWire_lo_hi_lo_hi_hi_hi, maskForGroupWire_lo_hi_lo_hi_hi_lo};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi = {maskForGroupWire_lo_hi_lo_hi_hi, maskForGroupWire_lo_hi_lo_hi_lo};
  wire [31:0]       maskForGroupWire_lo_hi_lo = {maskForGroupWire_lo_hi_lo_hi, maskForGroupWire_lo_hi_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_lo_lo = {{2{maskWire[49]}}, {2{maskWire[48]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_lo_hi = {{2{maskWire[51]}}, {2{maskWire[50]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo = {maskForGroupWire_lo_hi_hi_lo_lo_hi, maskForGroupWire_lo_hi_hi_lo_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_hi_lo = {{2{maskWire[53]}}, {2{maskWire[52]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_hi_hi = {{2{maskWire[55]}}, {2{maskWire[54]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi = {maskForGroupWire_lo_hi_hi_lo_hi_hi, maskForGroupWire_lo_hi_hi_lo_hi_lo};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo = {maskForGroupWire_lo_hi_hi_lo_hi, maskForGroupWire_lo_hi_hi_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_lo_lo = {{2{maskWire[57]}}, {2{maskWire[56]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_lo_hi = {{2{maskWire[59]}}, {2{maskWire[58]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo = {maskForGroupWire_lo_hi_hi_hi_lo_hi, maskForGroupWire_lo_hi_hi_hi_lo_lo};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_hi_lo = {{2{maskWire[61]}}, {2{maskWire[60]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_hi_hi = {{2{maskWire[63]}}, {2{maskWire[62]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi = {maskForGroupWire_lo_hi_hi_hi_hi_hi, maskForGroupWire_lo_hi_hi_hi_hi_lo};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi = {maskForGroupWire_lo_hi_hi_hi_hi, maskForGroupWire_lo_hi_hi_hi_lo};
  wire [31:0]       maskForGroupWire_lo_hi_hi = {maskForGroupWire_lo_hi_hi_hi, maskForGroupWire_lo_hi_hi_lo};
  wire [63:0]       maskForGroupWire_lo_hi = {maskForGroupWire_lo_hi_hi, maskForGroupWire_lo_hi_lo};
  wire [127:0]      maskForGroupWire_lo = {maskForGroupWire_lo_hi, maskForGroupWire_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_lo_lo = {{2{maskWire[65]}}, {2{maskWire[64]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_lo_hi = {{2{maskWire[67]}}, {2{maskWire[66]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo = {maskForGroupWire_hi_lo_lo_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_hi_lo = {{2{maskWire[69]}}, {2{maskWire[68]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_hi_hi = {{2{maskWire[71]}}, {2{maskWire[70]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi = {maskForGroupWire_hi_lo_lo_lo_hi_hi, maskForGroupWire_hi_lo_lo_lo_hi_lo};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo = {maskForGroupWire_hi_lo_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_lo_lo = {{2{maskWire[73]}}, {2{maskWire[72]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_lo_hi = {{2{maskWire[75]}}, {2{maskWire[74]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo = {maskForGroupWire_hi_lo_lo_hi_lo_hi, maskForGroupWire_hi_lo_lo_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_hi_lo = {{2{maskWire[77]}}, {2{maskWire[76]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_hi_hi = {{2{maskWire[79]}}, {2{maskWire[78]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi = {maskForGroupWire_hi_lo_lo_hi_hi_hi, maskForGroupWire_hi_lo_lo_hi_hi_lo};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi = {maskForGroupWire_hi_lo_lo_hi_hi, maskForGroupWire_hi_lo_lo_hi_lo};
  wire [31:0]       maskForGroupWire_hi_lo_lo = {maskForGroupWire_hi_lo_lo_hi, maskForGroupWire_hi_lo_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_lo_lo = {{2{maskWire[81]}}, {2{maskWire[80]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_lo_hi = {{2{maskWire[83]}}, {2{maskWire[82]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo = {maskForGroupWire_hi_lo_hi_lo_lo_hi, maskForGroupWire_hi_lo_hi_lo_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_hi_lo = {{2{maskWire[85]}}, {2{maskWire[84]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_hi_hi = {{2{maskWire[87]}}, {2{maskWire[86]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi = {maskForGroupWire_hi_lo_hi_lo_hi_hi, maskForGroupWire_hi_lo_hi_lo_hi_lo};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo = {maskForGroupWire_hi_lo_hi_lo_hi, maskForGroupWire_hi_lo_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_lo_lo = {{2{maskWire[89]}}, {2{maskWire[88]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_lo_hi = {{2{maskWire[91]}}, {2{maskWire[90]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo = {maskForGroupWire_hi_lo_hi_hi_lo_hi, maskForGroupWire_hi_lo_hi_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_hi_lo = {{2{maskWire[93]}}, {2{maskWire[92]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_hi_hi = {{2{maskWire[95]}}, {2{maskWire[94]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi = {maskForGroupWire_hi_lo_hi_hi_hi_hi, maskForGroupWire_hi_lo_hi_hi_hi_lo};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi = {maskForGroupWire_hi_lo_hi_hi_hi, maskForGroupWire_hi_lo_hi_hi_lo};
  wire [31:0]       maskForGroupWire_hi_lo_hi = {maskForGroupWire_hi_lo_hi_hi, maskForGroupWire_hi_lo_hi_lo};
  wire [63:0]       maskForGroupWire_hi_lo = {maskForGroupWire_hi_lo_hi, maskForGroupWire_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_lo_lo = {{2{maskWire[97]}}, {2{maskWire[96]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_lo_hi = {{2{maskWire[99]}}, {2{maskWire[98]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo = {maskForGroupWire_hi_hi_lo_lo_lo_hi, maskForGroupWire_hi_hi_lo_lo_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_hi_lo = {{2{maskWire[101]}}, {2{maskWire[100]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_hi_hi = {{2{maskWire[103]}}, {2{maskWire[102]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi = {maskForGroupWire_hi_hi_lo_lo_hi_hi, maskForGroupWire_hi_hi_lo_lo_hi_lo};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo = {maskForGroupWire_hi_hi_lo_lo_hi, maskForGroupWire_hi_hi_lo_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_lo_lo = {{2{maskWire[105]}}, {2{maskWire[104]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_lo_hi = {{2{maskWire[107]}}, {2{maskWire[106]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo = {maskForGroupWire_hi_hi_lo_hi_lo_hi, maskForGroupWire_hi_hi_lo_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_hi_lo = {{2{maskWire[109]}}, {2{maskWire[108]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_hi_hi = {{2{maskWire[111]}}, {2{maskWire[110]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi = {maskForGroupWire_hi_hi_lo_hi_hi_hi, maskForGroupWire_hi_hi_lo_hi_hi_lo};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi = {maskForGroupWire_hi_hi_lo_hi_hi, maskForGroupWire_hi_hi_lo_hi_lo};
  wire [31:0]       maskForGroupWire_hi_hi_lo = {maskForGroupWire_hi_hi_lo_hi, maskForGroupWire_hi_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_lo_lo = {{2{maskWire[113]}}, {2{maskWire[112]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_lo_hi = {{2{maskWire[115]}}, {2{maskWire[114]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo = {maskForGroupWire_hi_hi_hi_lo_lo_hi, maskForGroupWire_hi_hi_hi_lo_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_hi_lo = {{2{maskWire[117]}}, {2{maskWire[116]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_hi_hi = {{2{maskWire[119]}}, {2{maskWire[118]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi = {maskForGroupWire_hi_hi_hi_lo_hi_hi, maskForGroupWire_hi_hi_hi_lo_hi_lo};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo = {maskForGroupWire_hi_hi_hi_lo_hi, maskForGroupWire_hi_hi_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_lo_lo = {{2{maskWire[121]}}, {2{maskWire[120]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_lo_hi = {{2{maskWire[123]}}, {2{maskWire[122]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo = {maskForGroupWire_hi_hi_hi_hi_lo_hi, maskForGroupWire_hi_hi_hi_hi_lo_lo};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_hi_lo = {{2{maskWire[125]}}, {2{maskWire[124]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_hi_hi = {{2{maskWire[127]}}, {2{maskWire[126]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_hi_hi_lo};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_hi_lo};
  wire [31:0]       maskForGroupWire_hi_hi_hi = {maskForGroupWire_hi_hi_hi_hi, maskForGroupWire_hi_hi_hi_lo};
  wire [63:0]       maskForGroupWire_hi_hi = {maskForGroupWire_hi_hi_hi, maskForGroupWire_hi_hi_lo};
  wire [127:0]      maskForGroupWire_hi = {maskForGroupWire_hi_hi, maskForGroupWire_hi_lo};
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_lo_lo_1 = {{2{maskWire[1]}}, {2{maskWire[0]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_lo_hi_1 = {{2{maskWire[3]}}, {2{maskWire[2]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_hi_lo_1 = {{2{maskWire[5]}}, {2{maskWire[4]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_lo_hi_hi_1 = {{2{maskWire[7]}}, {2{maskWire[6]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_1 = {maskForGroupWire_lo_lo_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_lo_lo_1 = {{2{maskWire[9]}}, {2{maskWire[8]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_lo_hi_1 = {{2{maskWire[11]}}, {2{maskWire[10]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_1 = {maskForGroupWire_lo_lo_lo_hi_lo_hi_1, maskForGroupWire_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_hi_lo_1 = {{2{maskWire[13]}}, {2{maskWire[12]}}};
  wire [3:0]        maskForGroupWire_lo_lo_lo_hi_hi_hi_1 = {{2{maskWire[15]}}, {2{maskWire[14]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_1 = {maskForGroupWire_lo_lo_lo_hi_hi_hi_1, maskForGroupWire_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_1 = {maskForGroupWire_lo_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_lo_hi_lo_1};
  wire [31:0]       maskForGroupWire_lo_lo_lo_1 = {maskForGroupWire_lo_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_lo_lo_1 = {{2{maskWire[17]}}, {2{maskWire[16]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_lo_hi_1 = {{2{maskWire[19]}}, {2{maskWire[18]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_1 = {maskForGroupWire_lo_lo_hi_lo_lo_hi_1, maskForGroupWire_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_hi_lo_1 = {{2{maskWire[21]}}, {2{maskWire[20]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_lo_hi_hi_1 = {{2{maskWire[23]}}, {2{maskWire[22]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_1 = {maskForGroupWire_lo_lo_hi_lo_hi_hi_1, maskForGroupWire_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_1 = {maskForGroupWire_lo_lo_hi_lo_hi_1, maskForGroupWire_lo_lo_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_lo_lo_1 = {{2{maskWire[25]}}, {2{maskWire[24]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_lo_hi_1 = {{2{maskWire[27]}}, {2{maskWire[26]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_1 = {maskForGroupWire_lo_lo_hi_hi_lo_hi_1, maskForGroupWire_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_hi_lo_1 = {{2{maskWire[29]}}, {2{maskWire[28]}}};
  wire [3:0]        maskForGroupWire_lo_lo_hi_hi_hi_hi_1 = {{2{maskWire[31]}}, {2{maskWire[30]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_1 = {maskForGroupWire_lo_lo_hi_hi_hi_hi_1, maskForGroupWire_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_1 = {maskForGroupWire_lo_lo_hi_hi_hi_1, maskForGroupWire_lo_lo_hi_hi_lo_1};
  wire [31:0]       maskForGroupWire_lo_lo_hi_1 = {maskForGroupWire_lo_lo_hi_hi_1, maskForGroupWire_lo_lo_hi_lo_1};
  wire [63:0]       maskForGroupWire_lo_lo_1 = {maskForGroupWire_lo_lo_hi_1, maskForGroupWire_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_lo_lo_1 = {{2{maskWire[33]}}, {2{maskWire[32]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_lo_hi_1 = {{2{maskWire[35]}}, {2{maskWire[34]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_1 = {maskForGroupWire_lo_hi_lo_lo_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_hi_lo_1 = {{2{maskWire[37]}}, {2{maskWire[36]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_lo_hi_hi_1 = {{2{maskWire[39]}}, {2{maskWire[38]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_1 = {maskForGroupWire_lo_hi_lo_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_1 = {maskForGroupWire_lo_hi_lo_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_lo_lo_1 = {{2{maskWire[41]}}, {2{maskWire[40]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_lo_hi_1 = {{2{maskWire[43]}}, {2{maskWire[42]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_1 = {maskForGroupWire_lo_hi_lo_hi_lo_hi_1, maskForGroupWire_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_hi_lo_1 = {{2{maskWire[45]}}, {2{maskWire[44]}}};
  wire [3:0]        maskForGroupWire_lo_hi_lo_hi_hi_hi_1 = {{2{maskWire[47]}}, {2{maskWire[46]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_1 = {maskForGroupWire_lo_hi_lo_hi_hi_hi_1, maskForGroupWire_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_1 = {maskForGroupWire_lo_hi_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_hi_lo_1};
  wire [31:0]       maskForGroupWire_lo_hi_lo_1 = {maskForGroupWire_lo_hi_lo_hi_1, maskForGroupWire_lo_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_lo_lo_1 = {{2{maskWire[49]}}, {2{maskWire[48]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_lo_hi_1 = {{2{maskWire[51]}}, {2{maskWire[50]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_1 = {maskForGroupWire_lo_hi_hi_lo_lo_hi_1, maskForGroupWire_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_hi_lo_1 = {{2{maskWire[53]}}, {2{maskWire[52]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_lo_hi_hi_1 = {{2{maskWire[55]}}, {2{maskWire[54]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_1 = {maskForGroupWire_lo_hi_hi_lo_hi_hi_1, maskForGroupWire_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_1 = {maskForGroupWire_lo_hi_hi_lo_hi_1, maskForGroupWire_lo_hi_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_lo_lo_1 = {{2{maskWire[57]}}, {2{maskWire[56]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_lo_hi_1 = {{2{maskWire[59]}}, {2{maskWire[58]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_1 = {maskForGroupWire_lo_hi_hi_hi_lo_hi_1, maskForGroupWire_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_hi_lo_1 = {{2{maskWire[61]}}, {2{maskWire[60]}}};
  wire [3:0]        maskForGroupWire_lo_hi_hi_hi_hi_hi_1 = {{2{maskWire[63]}}, {2{maskWire[62]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_hi_lo_1};
  wire [31:0]       maskForGroupWire_lo_hi_hi_1 = {maskForGroupWire_lo_hi_hi_hi_1, maskForGroupWire_lo_hi_hi_lo_1};
  wire [63:0]       maskForGroupWire_lo_hi_1 = {maskForGroupWire_lo_hi_hi_1, maskForGroupWire_lo_hi_lo_1};
  wire [127:0]      maskForGroupWire_lo_1 = {maskForGroupWire_lo_hi_1, maskForGroupWire_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_lo_lo_1 = {{2{maskWire[65]}}, {2{maskWire[64]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_lo_hi_1 = {{2{maskWire[67]}}, {2{maskWire[66]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_1 = {maskForGroupWire_hi_lo_lo_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_hi_lo_1 = {{2{maskWire[69]}}, {2{maskWire[68]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_lo_hi_hi_1 = {{2{maskWire[71]}}, {2{maskWire[70]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_1 = {maskForGroupWire_hi_lo_lo_lo_hi_hi_1, maskForGroupWire_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_1 = {maskForGroupWire_hi_lo_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_lo_lo_1 = {{2{maskWire[73]}}, {2{maskWire[72]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_lo_hi_1 = {{2{maskWire[75]}}, {2{maskWire[74]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_1 = {maskForGroupWire_hi_lo_lo_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_hi_lo_1 = {{2{maskWire[77]}}, {2{maskWire[76]}}};
  wire [3:0]        maskForGroupWire_hi_lo_lo_hi_hi_hi_1 = {{2{maskWire[79]}}, {2{maskWire[78]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_1 = {maskForGroupWire_hi_lo_lo_hi_hi_hi_1, maskForGroupWire_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_1 = {maskForGroupWire_hi_lo_lo_hi_hi_1, maskForGroupWire_hi_lo_lo_hi_lo_1};
  wire [31:0]       maskForGroupWire_hi_lo_lo_1 = {maskForGroupWire_hi_lo_lo_hi_1, maskForGroupWire_hi_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_lo_lo_1 = {{2{maskWire[81]}}, {2{maskWire[80]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_lo_hi_1 = {{2{maskWire[83]}}, {2{maskWire[82]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_1 = {maskForGroupWire_hi_lo_hi_lo_lo_hi_1, maskForGroupWire_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_hi_lo_1 = {{2{maskWire[85]}}, {2{maskWire[84]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_lo_hi_hi_1 = {{2{maskWire[87]}}, {2{maskWire[86]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_1 = {maskForGroupWire_hi_lo_hi_lo_hi_hi_1, maskForGroupWire_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_1 = {maskForGroupWire_hi_lo_hi_lo_hi_1, maskForGroupWire_hi_lo_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_lo_lo_1 = {{2{maskWire[89]}}, {2{maskWire[88]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_lo_hi_1 = {{2{maskWire[91]}}, {2{maskWire[90]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_1 = {maskForGroupWire_hi_lo_hi_hi_lo_hi_1, maskForGroupWire_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_hi_lo_1 = {{2{maskWire[93]}}, {2{maskWire[92]}}};
  wire [3:0]        maskForGroupWire_hi_lo_hi_hi_hi_hi_1 = {{2{maskWire[95]}}, {2{maskWire[94]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_1 = {maskForGroupWire_hi_lo_hi_hi_hi_hi_1, maskForGroupWire_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_1 = {maskForGroupWire_hi_lo_hi_hi_hi_1, maskForGroupWire_hi_lo_hi_hi_lo_1};
  wire [31:0]       maskForGroupWire_hi_lo_hi_1 = {maskForGroupWire_hi_lo_hi_hi_1, maskForGroupWire_hi_lo_hi_lo_1};
  wire [63:0]       maskForGroupWire_hi_lo_1 = {maskForGroupWire_hi_lo_hi_1, maskForGroupWire_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_lo_lo_1 = {{2{maskWire[97]}}, {2{maskWire[96]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_lo_hi_1 = {{2{maskWire[99]}}, {2{maskWire[98]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_1 = {maskForGroupWire_hi_hi_lo_lo_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_hi_lo_1 = {{2{maskWire[101]}}, {2{maskWire[100]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_lo_hi_hi_1 = {{2{maskWire[103]}}, {2{maskWire[102]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_1 = {maskForGroupWire_hi_hi_lo_lo_hi_hi_1, maskForGroupWire_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_1 = {maskForGroupWire_hi_hi_lo_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_lo_lo_1 = {{2{maskWire[105]}}, {2{maskWire[104]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_lo_hi_1 = {{2{maskWire[107]}}, {2{maskWire[106]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_1 = {maskForGroupWire_hi_hi_lo_hi_lo_hi_1, maskForGroupWire_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_hi_lo_1 = {{2{maskWire[109]}}, {2{maskWire[108]}}};
  wire [3:0]        maskForGroupWire_hi_hi_lo_hi_hi_hi_1 = {{2{maskWire[111]}}, {2{maskWire[110]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_1 = {maskForGroupWire_hi_hi_lo_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_1 = {maskForGroupWire_hi_hi_lo_hi_hi_1, maskForGroupWire_hi_hi_lo_hi_lo_1};
  wire [31:0]       maskForGroupWire_hi_hi_lo_1 = {maskForGroupWire_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_lo_lo_1 = {{2{maskWire[113]}}, {2{maskWire[112]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_lo_hi_1 = {{2{maskWire[115]}}, {2{maskWire[114]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_1 = {maskForGroupWire_hi_hi_hi_lo_lo_hi_1, maskForGroupWire_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_hi_lo_1 = {{2{maskWire[117]}}, {2{maskWire[116]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_lo_hi_hi_1 = {{2{maskWire[119]}}, {2{maskWire[118]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_1 = {maskForGroupWire_hi_hi_hi_lo_hi_hi_1, maskForGroupWire_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_1 = {maskForGroupWire_hi_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_lo_lo_1 = {{2{maskWire[121]}}, {2{maskWire[120]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_lo_hi_1 = {{2{maskWire[123]}}, {2{maskWire[122]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_1 = {maskForGroupWire_hi_hi_hi_hi_lo_hi_1, maskForGroupWire_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_hi_lo_1 = {{2{maskWire[125]}}, {2{maskWire[124]}}};
  wire [3:0]        maskForGroupWire_hi_hi_hi_hi_hi_hi_1 = {{2{maskWire[127]}}, {2{maskWire[126]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_hi_lo_1};
  wire [31:0]       maskForGroupWire_hi_hi_hi_1 = {maskForGroupWire_hi_hi_hi_hi_1, maskForGroupWire_hi_hi_hi_lo_1};
  wire [63:0]       maskForGroupWire_hi_hi_1 = {maskForGroupWire_hi_hi_hi_1, maskForGroupWire_hi_hi_lo_1};
  wire [127:0]      maskForGroupWire_hi_1 = {maskForGroupWire_hi_hi_1, maskForGroupWire_hi_lo_1};
  wire [3:0]        _maskForGroupWire_T_517 = 4'h1 << maskCounterInGroup;
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_lo_2 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_hi_2 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_lo_2 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_hi_2 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_hi_2 = {maskForGroupWire_lo_lo_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_lo_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_lo_2 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_hi_2 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_lo_2 = {maskForGroupWire_lo_lo_lo_hi_lo_hi_2, maskForGroupWire_lo_lo_lo_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_lo_2 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_hi_2 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_hi_2 = {maskForGroupWire_lo_lo_lo_hi_hi_hi_2, maskForGroupWire_lo_lo_lo_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_lo_lo_hi_2 = {maskForGroupWire_lo_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_lo_hi_lo_2};
  wire [63:0]       maskForGroupWire_lo_lo_lo_2 = {maskForGroupWire_lo_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_lo_2 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_hi_2 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_lo_2 = {maskForGroupWire_lo_lo_hi_lo_lo_hi_2, maskForGroupWire_lo_lo_hi_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_lo_2 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_hi_2 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_hi_2 = {maskForGroupWire_lo_lo_hi_lo_hi_hi_2, maskForGroupWire_lo_lo_hi_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_lo_hi_lo_2 = {maskForGroupWire_lo_lo_hi_lo_hi_2, maskForGroupWire_lo_lo_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_lo_2 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_hi_2 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_lo_2 = {maskForGroupWire_lo_lo_hi_hi_lo_hi_2, maskForGroupWire_lo_lo_hi_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_lo_2 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_hi_2 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_hi_2 = {maskForGroupWire_lo_lo_hi_hi_hi_hi_2, maskForGroupWire_lo_lo_hi_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_lo_hi_hi_2 = {maskForGroupWire_lo_lo_hi_hi_hi_2, maskForGroupWire_lo_lo_hi_hi_lo_2};
  wire [63:0]       maskForGroupWire_lo_lo_hi_2 = {maskForGroupWire_lo_lo_hi_hi_2, maskForGroupWire_lo_lo_hi_lo_2};
  wire [127:0]      maskForGroupWire_lo_lo_2 = {maskForGroupWire_lo_lo_hi_2, maskForGroupWire_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_lo_2 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_hi_2 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_lo_2 = {maskForGroupWire_lo_hi_lo_lo_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_lo_2 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_hi_2 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_hi_2 = {maskForGroupWire_lo_hi_lo_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_hi_lo_lo_2 = {maskForGroupWire_lo_hi_lo_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_lo_2 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_hi_2 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_lo_2 = {maskForGroupWire_lo_hi_lo_hi_lo_hi_2, maskForGroupWire_lo_hi_lo_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_lo_2 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_hi_2 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_hi_2 = {maskForGroupWire_lo_hi_lo_hi_hi_hi_2, maskForGroupWire_lo_hi_lo_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_hi_lo_hi_2 = {maskForGroupWire_lo_hi_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_hi_lo_2};
  wire [63:0]       maskForGroupWire_lo_hi_lo_2 = {maskForGroupWire_lo_hi_lo_hi_2, maskForGroupWire_lo_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_lo_2 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_hi_2 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_lo_2 = {maskForGroupWire_lo_hi_hi_lo_lo_hi_2, maskForGroupWire_lo_hi_hi_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_lo_2 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_hi_2 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_hi_2 = {maskForGroupWire_lo_hi_hi_lo_hi_hi_2, maskForGroupWire_lo_hi_hi_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_hi_hi_lo_2 = {maskForGroupWire_lo_hi_hi_lo_hi_2, maskForGroupWire_lo_hi_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_lo_2 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_hi_2 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_lo_2 = {maskForGroupWire_lo_hi_hi_hi_lo_hi_2, maskForGroupWire_lo_hi_hi_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_lo_2 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_hi_2 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_lo_hi_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_hi_lo_2};
  wire [63:0]       maskForGroupWire_lo_hi_hi_2 = {maskForGroupWire_lo_hi_hi_hi_2, maskForGroupWire_lo_hi_hi_lo_2};
  wire [127:0]      maskForGroupWire_lo_hi_2 = {maskForGroupWire_lo_hi_hi_2, maskForGroupWire_lo_hi_lo_2};
  wire [255:0]      maskForGroupWire_lo_2 = {maskForGroupWire_lo_hi_2, maskForGroupWire_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_lo_2 = {{4{maskWire[65]}}, {4{maskWire[64]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_hi_2 = {{4{maskWire[67]}}, {4{maskWire[66]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_lo_2 = {maskForGroupWire_hi_lo_lo_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_lo_2 = {{4{maskWire[69]}}, {4{maskWire[68]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_hi_2 = {{4{maskWire[71]}}, {4{maskWire[70]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_hi_2 = {maskForGroupWire_hi_lo_lo_lo_hi_hi_2, maskForGroupWire_hi_lo_lo_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_lo_lo_lo_2 = {maskForGroupWire_hi_lo_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_lo_2 = {{4{maskWire[73]}}, {4{maskWire[72]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_hi_2 = {{4{maskWire[75]}}, {4{maskWire[74]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_lo_2 = {maskForGroupWire_hi_lo_lo_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_lo_2 = {{4{maskWire[77]}}, {4{maskWire[76]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_hi_2 = {{4{maskWire[79]}}, {4{maskWire[78]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_hi_2 = {maskForGroupWire_hi_lo_lo_hi_hi_hi_2, maskForGroupWire_hi_lo_lo_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_lo_lo_hi_2 = {maskForGroupWire_hi_lo_lo_hi_hi_2, maskForGroupWire_hi_lo_lo_hi_lo_2};
  wire [63:0]       maskForGroupWire_hi_lo_lo_2 = {maskForGroupWire_hi_lo_lo_hi_2, maskForGroupWire_hi_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_lo_2 = {{4{maskWire[81]}}, {4{maskWire[80]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_hi_2 = {{4{maskWire[83]}}, {4{maskWire[82]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_lo_2 = {maskForGroupWire_hi_lo_hi_lo_lo_hi_2, maskForGroupWire_hi_lo_hi_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_lo_2 = {{4{maskWire[85]}}, {4{maskWire[84]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_hi_2 = {{4{maskWire[87]}}, {4{maskWire[86]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_hi_2 = {maskForGroupWire_hi_lo_hi_lo_hi_hi_2, maskForGroupWire_hi_lo_hi_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_lo_hi_lo_2 = {maskForGroupWire_hi_lo_hi_lo_hi_2, maskForGroupWire_hi_lo_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_lo_2 = {{4{maskWire[89]}}, {4{maskWire[88]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_hi_2 = {{4{maskWire[91]}}, {4{maskWire[90]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_lo_2 = {maskForGroupWire_hi_lo_hi_hi_lo_hi_2, maskForGroupWire_hi_lo_hi_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_lo_2 = {{4{maskWire[93]}}, {4{maskWire[92]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_hi_2 = {{4{maskWire[95]}}, {4{maskWire[94]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_hi_2 = {maskForGroupWire_hi_lo_hi_hi_hi_hi_2, maskForGroupWire_hi_lo_hi_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_lo_hi_hi_2 = {maskForGroupWire_hi_lo_hi_hi_hi_2, maskForGroupWire_hi_lo_hi_hi_lo_2};
  wire [63:0]       maskForGroupWire_hi_lo_hi_2 = {maskForGroupWire_hi_lo_hi_hi_2, maskForGroupWire_hi_lo_hi_lo_2};
  wire [127:0]      maskForGroupWire_hi_lo_2 = {maskForGroupWire_hi_lo_hi_2, maskForGroupWire_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_lo_2 = {{4{maskWire[97]}}, {4{maskWire[96]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_hi_2 = {{4{maskWire[99]}}, {4{maskWire[98]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_lo_2 = {maskForGroupWire_hi_hi_lo_lo_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_lo_2 = {{4{maskWire[101]}}, {4{maskWire[100]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_hi_2 = {{4{maskWire[103]}}, {4{maskWire[102]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_hi_2 = {maskForGroupWire_hi_hi_lo_lo_hi_hi_2, maskForGroupWire_hi_hi_lo_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_hi_lo_lo_2 = {maskForGroupWire_hi_hi_lo_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_lo_2 = {{4{maskWire[105]}}, {4{maskWire[104]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_hi_2 = {{4{maskWire[107]}}, {4{maskWire[106]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_lo_2 = {maskForGroupWire_hi_hi_lo_hi_lo_hi_2, maskForGroupWire_hi_hi_lo_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_lo_2 = {{4{maskWire[109]}}, {4{maskWire[108]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_hi_2 = {{4{maskWire[111]}}, {4{maskWire[110]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_hi_2 = {maskForGroupWire_hi_hi_lo_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_hi_lo_hi_2 = {maskForGroupWire_hi_hi_lo_hi_hi_2, maskForGroupWire_hi_hi_lo_hi_lo_2};
  wire [63:0]       maskForGroupWire_hi_hi_lo_2 = {maskForGroupWire_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_lo_2 = {{4{maskWire[113]}}, {4{maskWire[112]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_hi_2 = {{4{maskWire[115]}}, {4{maskWire[114]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_lo_2 = {maskForGroupWire_hi_hi_hi_lo_lo_hi_2, maskForGroupWire_hi_hi_hi_lo_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_lo_2 = {{4{maskWire[117]}}, {4{maskWire[116]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_hi_2 = {{4{maskWire[119]}}, {4{maskWire[118]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_hi_2 = {maskForGroupWire_hi_hi_hi_lo_hi_hi_2, maskForGroupWire_hi_hi_hi_lo_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_hi_hi_lo_2 = {maskForGroupWire_hi_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_lo_2 = {{4{maskWire[121]}}, {4{maskWire[120]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_hi_2 = {{4{maskWire[123]}}, {4{maskWire[122]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_lo_2 = {maskForGroupWire_hi_hi_hi_hi_lo_hi_2, maskForGroupWire_hi_hi_hi_hi_lo_lo_2};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_lo_2 = {{4{maskWire[125]}}, {4{maskWire[124]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_hi_2 = {{4{maskWire[127]}}, {4{maskWire[126]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_hi_hi_lo_2};
  wire [31:0]       maskForGroupWire_hi_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_hi_lo_2};
  wire [63:0]       maskForGroupWire_hi_hi_hi_2 = {maskForGroupWire_hi_hi_hi_hi_2, maskForGroupWire_hi_hi_hi_lo_2};
  wire [127:0]      maskForGroupWire_hi_hi_2 = {maskForGroupWire_hi_hi_hi_2, maskForGroupWire_hi_hi_lo_2};
  wire [255:0]      maskForGroupWire_hi_2 = {maskForGroupWire_hi_hi_2, maskForGroupWire_hi_lo_2};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_lo_3 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_hi_3 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_lo_3 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_hi_3 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_hi_3 = {maskForGroupWire_lo_lo_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_lo_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_lo_3 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_hi_3 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_lo_3 = {maskForGroupWire_lo_lo_lo_hi_lo_hi_3, maskForGroupWire_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_lo_3 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_hi_3 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_hi_3 = {maskForGroupWire_lo_lo_lo_hi_hi_hi_3, maskForGroupWire_lo_lo_lo_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_lo_lo_hi_3 = {maskForGroupWire_lo_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_lo_hi_lo_3};
  wire [63:0]       maskForGroupWire_lo_lo_lo_3 = {maskForGroupWire_lo_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_lo_3 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_hi_3 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_lo_3 = {maskForGroupWire_lo_lo_hi_lo_lo_hi_3, maskForGroupWire_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_lo_3 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_hi_3 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_hi_3 = {maskForGroupWire_lo_lo_hi_lo_hi_hi_3, maskForGroupWire_lo_lo_hi_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_lo_hi_lo_3 = {maskForGroupWire_lo_lo_hi_lo_hi_3, maskForGroupWire_lo_lo_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_lo_3 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_hi_3 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_lo_3 = {maskForGroupWire_lo_lo_hi_hi_lo_hi_3, maskForGroupWire_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_lo_3 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_hi_3 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_hi_3 = {maskForGroupWire_lo_lo_hi_hi_hi_hi_3, maskForGroupWire_lo_lo_hi_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_lo_hi_hi_3 = {maskForGroupWire_lo_lo_hi_hi_hi_3, maskForGroupWire_lo_lo_hi_hi_lo_3};
  wire [63:0]       maskForGroupWire_lo_lo_hi_3 = {maskForGroupWire_lo_lo_hi_hi_3, maskForGroupWire_lo_lo_hi_lo_3};
  wire [127:0]      maskForGroupWire_lo_lo_3 = {maskForGroupWire_lo_lo_hi_3, maskForGroupWire_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_lo_3 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_hi_3 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_lo_3 = {maskForGroupWire_lo_hi_lo_lo_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_lo_3 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_hi_3 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_hi_3 = {maskForGroupWire_lo_hi_lo_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_hi_lo_lo_3 = {maskForGroupWire_lo_hi_lo_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_lo_3 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_hi_3 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_lo_3 = {maskForGroupWire_lo_hi_lo_hi_lo_hi_3, maskForGroupWire_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_lo_3 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_hi_3 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_hi_3 = {maskForGroupWire_lo_hi_lo_hi_hi_hi_3, maskForGroupWire_lo_hi_lo_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_hi_lo_hi_3 = {maskForGroupWire_lo_hi_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_hi_lo_3};
  wire [63:0]       maskForGroupWire_lo_hi_lo_3 = {maskForGroupWire_lo_hi_lo_hi_3, maskForGroupWire_lo_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_lo_3 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_hi_3 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_lo_3 = {maskForGroupWire_lo_hi_hi_lo_lo_hi_3, maskForGroupWire_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_lo_3 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_hi_3 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_hi_3 = {maskForGroupWire_lo_hi_hi_lo_hi_hi_3, maskForGroupWire_lo_hi_hi_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_hi_hi_lo_3 = {maskForGroupWire_lo_hi_hi_lo_hi_3, maskForGroupWire_lo_hi_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_lo_3 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_hi_3 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_lo_3 = {maskForGroupWire_lo_hi_hi_hi_lo_hi_3, maskForGroupWire_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_lo_3 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_hi_3 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_lo_hi_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_hi_lo_3};
  wire [63:0]       maskForGroupWire_lo_hi_hi_3 = {maskForGroupWire_lo_hi_hi_hi_3, maskForGroupWire_lo_hi_hi_lo_3};
  wire [127:0]      maskForGroupWire_lo_hi_3 = {maskForGroupWire_lo_hi_hi_3, maskForGroupWire_lo_hi_lo_3};
  wire [255:0]      maskForGroupWire_lo_3 = {maskForGroupWire_lo_hi_3, maskForGroupWire_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_lo_3 = {{4{maskWire[65]}}, {4{maskWire[64]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_hi_3 = {{4{maskWire[67]}}, {4{maskWire[66]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_lo_3 = {maskForGroupWire_hi_lo_lo_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_lo_3 = {{4{maskWire[69]}}, {4{maskWire[68]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_hi_3 = {{4{maskWire[71]}}, {4{maskWire[70]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_hi_3 = {maskForGroupWire_hi_lo_lo_lo_hi_hi_3, maskForGroupWire_hi_lo_lo_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_lo_lo_lo_3 = {maskForGroupWire_hi_lo_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_lo_3 = {{4{maskWire[73]}}, {4{maskWire[72]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_hi_3 = {{4{maskWire[75]}}, {4{maskWire[74]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_lo_3 = {maskForGroupWire_hi_lo_lo_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_lo_3 = {{4{maskWire[77]}}, {4{maskWire[76]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_hi_3 = {{4{maskWire[79]}}, {4{maskWire[78]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_hi_3 = {maskForGroupWire_hi_lo_lo_hi_hi_hi_3, maskForGroupWire_hi_lo_lo_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_lo_lo_hi_3 = {maskForGroupWire_hi_lo_lo_hi_hi_3, maskForGroupWire_hi_lo_lo_hi_lo_3};
  wire [63:0]       maskForGroupWire_hi_lo_lo_3 = {maskForGroupWire_hi_lo_lo_hi_3, maskForGroupWire_hi_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_lo_3 = {{4{maskWire[81]}}, {4{maskWire[80]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_hi_3 = {{4{maskWire[83]}}, {4{maskWire[82]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_lo_3 = {maskForGroupWire_hi_lo_hi_lo_lo_hi_3, maskForGroupWire_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_lo_3 = {{4{maskWire[85]}}, {4{maskWire[84]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_hi_3 = {{4{maskWire[87]}}, {4{maskWire[86]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_hi_3 = {maskForGroupWire_hi_lo_hi_lo_hi_hi_3, maskForGroupWire_hi_lo_hi_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_lo_hi_lo_3 = {maskForGroupWire_hi_lo_hi_lo_hi_3, maskForGroupWire_hi_lo_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_lo_3 = {{4{maskWire[89]}}, {4{maskWire[88]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_hi_3 = {{4{maskWire[91]}}, {4{maskWire[90]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_lo_3 = {maskForGroupWire_hi_lo_hi_hi_lo_hi_3, maskForGroupWire_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_lo_3 = {{4{maskWire[93]}}, {4{maskWire[92]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_hi_3 = {{4{maskWire[95]}}, {4{maskWire[94]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_hi_3 = {maskForGroupWire_hi_lo_hi_hi_hi_hi_3, maskForGroupWire_hi_lo_hi_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_lo_hi_hi_3 = {maskForGroupWire_hi_lo_hi_hi_hi_3, maskForGroupWire_hi_lo_hi_hi_lo_3};
  wire [63:0]       maskForGroupWire_hi_lo_hi_3 = {maskForGroupWire_hi_lo_hi_hi_3, maskForGroupWire_hi_lo_hi_lo_3};
  wire [127:0]      maskForGroupWire_hi_lo_3 = {maskForGroupWire_hi_lo_hi_3, maskForGroupWire_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_lo_3 = {{4{maskWire[97]}}, {4{maskWire[96]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_hi_3 = {{4{maskWire[99]}}, {4{maskWire[98]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_lo_3 = {maskForGroupWire_hi_hi_lo_lo_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_lo_3 = {{4{maskWire[101]}}, {4{maskWire[100]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_hi_3 = {{4{maskWire[103]}}, {4{maskWire[102]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_hi_3 = {maskForGroupWire_hi_hi_lo_lo_hi_hi_3, maskForGroupWire_hi_hi_lo_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_hi_lo_lo_3 = {maskForGroupWire_hi_hi_lo_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_lo_3 = {{4{maskWire[105]}}, {4{maskWire[104]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_hi_3 = {{4{maskWire[107]}}, {4{maskWire[106]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_lo_3 = {maskForGroupWire_hi_hi_lo_hi_lo_hi_3, maskForGroupWire_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_lo_3 = {{4{maskWire[109]}}, {4{maskWire[108]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_hi_3 = {{4{maskWire[111]}}, {4{maskWire[110]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_hi_3 = {maskForGroupWire_hi_hi_lo_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_hi_lo_hi_3 = {maskForGroupWire_hi_hi_lo_hi_hi_3, maskForGroupWire_hi_hi_lo_hi_lo_3};
  wire [63:0]       maskForGroupWire_hi_hi_lo_3 = {maskForGroupWire_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_lo_3 = {{4{maskWire[113]}}, {4{maskWire[112]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_hi_3 = {{4{maskWire[115]}}, {4{maskWire[114]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_lo_3 = {maskForGroupWire_hi_hi_hi_lo_lo_hi_3, maskForGroupWire_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_lo_3 = {{4{maskWire[117]}}, {4{maskWire[116]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_hi_3 = {{4{maskWire[119]}}, {4{maskWire[118]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_hi_3 = {maskForGroupWire_hi_hi_hi_lo_hi_hi_3, maskForGroupWire_hi_hi_hi_lo_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_hi_hi_lo_3 = {maskForGroupWire_hi_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_lo_3 = {{4{maskWire[121]}}, {4{maskWire[120]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_hi_3 = {{4{maskWire[123]}}, {4{maskWire[122]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_lo_3 = {maskForGroupWire_hi_hi_hi_hi_lo_hi_3, maskForGroupWire_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_lo_3 = {{4{maskWire[125]}}, {4{maskWire[124]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_hi_3 = {{4{maskWire[127]}}, {4{maskWire[126]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_hi_hi_lo_3};
  wire [31:0]       maskForGroupWire_hi_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_hi_lo_3};
  wire [63:0]       maskForGroupWire_hi_hi_hi_3 = {maskForGroupWire_hi_hi_hi_hi_3, maskForGroupWire_hi_hi_hi_lo_3};
  wire [127:0]      maskForGroupWire_hi_hi_3 = {maskForGroupWire_hi_hi_hi_3, maskForGroupWire_hi_hi_lo_3};
  wire [255:0]      maskForGroupWire_hi_3 = {maskForGroupWire_hi_hi_3, maskForGroupWire_hi_lo_3};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_lo_4 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_hi_4 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_lo_4 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_hi_4 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_hi_4 = {maskForGroupWire_lo_lo_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_lo_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_lo_4 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_hi_4 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_lo_4 = {maskForGroupWire_lo_lo_lo_hi_lo_hi_4, maskForGroupWire_lo_lo_lo_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_lo_4 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_hi_4 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_hi_4 = {maskForGroupWire_lo_lo_lo_hi_hi_hi_4, maskForGroupWire_lo_lo_lo_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_lo_lo_hi_4 = {maskForGroupWire_lo_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_lo_hi_lo_4};
  wire [63:0]       maskForGroupWire_lo_lo_lo_4 = {maskForGroupWire_lo_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_lo_4 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_hi_4 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_lo_4 = {maskForGroupWire_lo_lo_hi_lo_lo_hi_4, maskForGroupWire_lo_lo_hi_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_lo_4 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_hi_4 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_hi_4 = {maskForGroupWire_lo_lo_hi_lo_hi_hi_4, maskForGroupWire_lo_lo_hi_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_lo_hi_lo_4 = {maskForGroupWire_lo_lo_hi_lo_hi_4, maskForGroupWire_lo_lo_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_lo_4 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_hi_4 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_lo_4 = {maskForGroupWire_lo_lo_hi_hi_lo_hi_4, maskForGroupWire_lo_lo_hi_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_lo_4 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_hi_4 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_hi_4 = {maskForGroupWire_lo_lo_hi_hi_hi_hi_4, maskForGroupWire_lo_lo_hi_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_lo_hi_hi_4 = {maskForGroupWire_lo_lo_hi_hi_hi_4, maskForGroupWire_lo_lo_hi_hi_lo_4};
  wire [63:0]       maskForGroupWire_lo_lo_hi_4 = {maskForGroupWire_lo_lo_hi_hi_4, maskForGroupWire_lo_lo_hi_lo_4};
  wire [127:0]      maskForGroupWire_lo_lo_4 = {maskForGroupWire_lo_lo_hi_4, maskForGroupWire_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_lo_4 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_hi_4 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_lo_4 = {maskForGroupWire_lo_hi_lo_lo_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_lo_4 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_hi_4 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_hi_4 = {maskForGroupWire_lo_hi_lo_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_hi_lo_lo_4 = {maskForGroupWire_lo_hi_lo_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_lo_4 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_hi_4 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_lo_4 = {maskForGroupWire_lo_hi_lo_hi_lo_hi_4, maskForGroupWire_lo_hi_lo_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_lo_4 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_hi_4 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_hi_4 = {maskForGroupWire_lo_hi_lo_hi_hi_hi_4, maskForGroupWire_lo_hi_lo_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_hi_lo_hi_4 = {maskForGroupWire_lo_hi_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_hi_lo_4};
  wire [63:0]       maskForGroupWire_lo_hi_lo_4 = {maskForGroupWire_lo_hi_lo_hi_4, maskForGroupWire_lo_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_lo_4 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_hi_4 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_lo_4 = {maskForGroupWire_lo_hi_hi_lo_lo_hi_4, maskForGroupWire_lo_hi_hi_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_lo_4 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_hi_4 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_hi_4 = {maskForGroupWire_lo_hi_hi_lo_hi_hi_4, maskForGroupWire_lo_hi_hi_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_hi_hi_lo_4 = {maskForGroupWire_lo_hi_hi_lo_hi_4, maskForGroupWire_lo_hi_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_lo_4 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_hi_4 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_lo_4 = {maskForGroupWire_lo_hi_hi_hi_lo_hi_4, maskForGroupWire_lo_hi_hi_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_lo_4 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_hi_4 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_lo_hi_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_hi_lo_4};
  wire [63:0]       maskForGroupWire_lo_hi_hi_4 = {maskForGroupWire_lo_hi_hi_hi_4, maskForGroupWire_lo_hi_hi_lo_4};
  wire [127:0]      maskForGroupWire_lo_hi_4 = {maskForGroupWire_lo_hi_hi_4, maskForGroupWire_lo_hi_lo_4};
  wire [255:0]      maskForGroupWire_lo_4 = {maskForGroupWire_lo_hi_4, maskForGroupWire_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_lo_4 = {{4{maskWire[65]}}, {4{maskWire[64]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_hi_4 = {{4{maskWire[67]}}, {4{maskWire[66]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_lo_4 = {maskForGroupWire_hi_lo_lo_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_lo_4 = {{4{maskWire[69]}}, {4{maskWire[68]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_hi_4 = {{4{maskWire[71]}}, {4{maskWire[70]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_hi_4 = {maskForGroupWire_hi_lo_lo_lo_hi_hi_4, maskForGroupWire_hi_lo_lo_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_lo_lo_lo_4 = {maskForGroupWire_hi_lo_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_lo_4 = {{4{maskWire[73]}}, {4{maskWire[72]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_hi_4 = {{4{maskWire[75]}}, {4{maskWire[74]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_lo_4 = {maskForGroupWire_hi_lo_lo_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_lo_4 = {{4{maskWire[77]}}, {4{maskWire[76]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_hi_4 = {{4{maskWire[79]}}, {4{maskWire[78]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_hi_4 = {maskForGroupWire_hi_lo_lo_hi_hi_hi_4, maskForGroupWire_hi_lo_lo_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_lo_lo_hi_4 = {maskForGroupWire_hi_lo_lo_hi_hi_4, maskForGroupWire_hi_lo_lo_hi_lo_4};
  wire [63:0]       maskForGroupWire_hi_lo_lo_4 = {maskForGroupWire_hi_lo_lo_hi_4, maskForGroupWire_hi_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_lo_4 = {{4{maskWire[81]}}, {4{maskWire[80]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_hi_4 = {{4{maskWire[83]}}, {4{maskWire[82]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_lo_4 = {maskForGroupWire_hi_lo_hi_lo_lo_hi_4, maskForGroupWire_hi_lo_hi_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_lo_4 = {{4{maskWire[85]}}, {4{maskWire[84]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_hi_4 = {{4{maskWire[87]}}, {4{maskWire[86]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_hi_4 = {maskForGroupWire_hi_lo_hi_lo_hi_hi_4, maskForGroupWire_hi_lo_hi_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_lo_hi_lo_4 = {maskForGroupWire_hi_lo_hi_lo_hi_4, maskForGroupWire_hi_lo_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_lo_4 = {{4{maskWire[89]}}, {4{maskWire[88]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_hi_4 = {{4{maskWire[91]}}, {4{maskWire[90]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_lo_4 = {maskForGroupWire_hi_lo_hi_hi_lo_hi_4, maskForGroupWire_hi_lo_hi_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_lo_4 = {{4{maskWire[93]}}, {4{maskWire[92]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_hi_4 = {{4{maskWire[95]}}, {4{maskWire[94]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_hi_4 = {maskForGroupWire_hi_lo_hi_hi_hi_hi_4, maskForGroupWire_hi_lo_hi_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_lo_hi_hi_4 = {maskForGroupWire_hi_lo_hi_hi_hi_4, maskForGroupWire_hi_lo_hi_hi_lo_4};
  wire [63:0]       maskForGroupWire_hi_lo_hi_4 = {maskForGroupWire_hi_lo_hi_hi_4, maskForGroupWire_hi_lo_hi_lo_4};
  wire [127:0]      maskForGroupWire_hi_lo_4 = {maskForGroupWire_hi_lo_hi_4, maskForGroupWire_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_lo_4 = {{4{maskWire[97]}}, {4{maskWire[96]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_hi_4 = {{4{maskWire[99]}}, {4{maskWire[98]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_lo_4 = {maskForGroupWire_hi_hi_lo_lo_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_lo_4 = {{4{maskWire[101]}}, {4{maskWire[100]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_hi_4 = {{4{maskWire[103]}}, {4{maskWire[102]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_hi_4 = {maskForGroupWire_hi_hi_lo_lo_hi_hi_4, maskForGroupWire_hi_hi_lo_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_hi_lo_lo_4 = {maskForGroupWire_hi_hi_lo_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_lo_4 = {{4{maskWire[105]}}, {4{maskWire[104]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_hi_4 = {{4{maskWire[107]}}, {4{maskWire[106]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_lo_4 = {maskForGroupWire_hi_hi_lo_hi_lo_hi_4, maskForGroupWire_hi_hi_lo_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_lo_4 = {{4{maskWire[109]}}, {4{maskWire[108]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_hi_4 = {{4{maskWire[111]}}, {4{maskWire[110]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_hi_4 = {maskForGroupWire_hi_hi_lo_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_hi_lo_hi_4 = {maskForGroupWire_hi_hi_lo_hi_hi_4, maskForGroupWire_hi_hi_lo_hi_lo_4};
  wire [63:0]       maskForGroupWire_hi_hi_lo_4 = {maskForGroupWire_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_lo_4 = {{4{maskWire[113]}}, {4{maskWire[112]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_hi_4 = {{4{maskWire[115]}}, {4{maskWire[114]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_lo_4 = {maskForGroupWire_hi_hi_hi_lo_lo_hi_4, maskForGroupWire_hi_hi_hi_lo_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_lo_4 = {{4{maskWire[117]}}, {4{maskWire[116]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_hi_4 = {{4{maskWire[119]}}, {4{maskWire[118]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_hi_4 = {maskForGroupWire_hi_hi_hi_lo_hi_hi_4, maskForGroupWire_hi_hi_hi_lo_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_hi_hi_lo_4 = {maskForGroupWire_hi_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_lo_4 = {{4{maskWire[121]}}, {4{maskWire[120]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_hi_4 = {{4{maskWire[123]}}, {4{maskWire[122]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_lo_4 = {maskForGroupWire_hi_hi_hi_hi_lo_hi_4, maskForGroupWire_hi_hi_hi_hi_lo_lo_4};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_lo_4 = {{4{maskWire[125]}}, {4{maskWire[124]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_hi_4 = {{4{maskWire[127]}}, {4{maskWire[126]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_hi_hi_lo_4};
  wire [31:0]       maskForGroupWire_hi_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_hi_lo_4};
  wire [63:0]       maskForGroupWire_hi_hi_hi_4 = {maskForGroupWire_hi_hi_hi_hi_4, maskForGroupWire_hi_hi_hi_lo_4};
  wire [127:0]      maskForGroupWire_hi_hi_4 = {maskForGroupWire_hi_hi_hi_4, maskForGroupWire_hi_hi_lo_4};
  wire [255:0]      maskForGroupWire_hi_4 = {maskForGroupWire_hi_hi_4, maskForGroupWire_hi_lo_4};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_lo_5 = {{4{maskWire[1]}}, {4{maskWire[0]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_lo_hi_5 = {{4{maskWire[3]}}, {4{maskWire[2]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_lo_5 = {{4{maskWire[5]}}, {4{maskWire[4]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_lo_hi_hi_5 = {{4{maskWire[7]}}, {4{maskWire[6]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_lo_hi_5 = {maskForGroupWire_lo_lo_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_lo_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_lo_5 = {{4{maskWire[9]}}, {4{maskWire[8]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_lo_hi_5 = {{4{maskWire[11]}}, {4{maskWire[10]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_lo_5 = {maskForGroupWire_lo_lo_lo_hi_lo_hi_5, maskForGroupWire_lo_lo_lo_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_lo_5 = {{4{maskWire[13]}}, {4{maskWire[12]}}};
  wire [7:0]        maskForGroupWire_lo_lo_lo_hi_hi_hi_5 = {{4{maskWire[15]}}, {4{maskWire[14]}}};
  wire [15:0]       maskForGroupWire_lo_lo_lo_hi_hi_5 = {maskForGroupWire_lo_lo_lo_hi_hi_hi_5, maskForGroupWire_lo_lo_lo_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_lo_lo_hi_5 = {maskForGroupWire_lo_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_lo_hi_lo_5};
  wire [63:0]       maskForGroupWire_lo_lo_lo_5 = {maskForGroupWire_lo_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_lo_5 = {{4{maskWire[17]}}, {4{maskWire[16]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_lo_hi_5 = {{4{maskWire[19]}}, {4{maskWire[18]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_lo_5 = {maskForGroupWire_lo_lo_hi_lo_lo_hi_5, maskForGroupWire_lo_lo_hi_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_lo_5 = {{4{maskWire[21]}}, {4{maskWire[20]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_lo_hi_hi_5 = {{4{maskWire[23]}}, {4{maskWire[22]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_lo_hi_5 = {maskForGroupWire_lo_lo_hi_lo_hi_hi_5, maskForGroupWire_lo_lo_hi_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_lo_hi_lo_5 = {maskForGroupWire_lo_lo_hi_lo_hi_5, maskForGroupWire_lo_lo_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_lo_5 = {{4{maskWire[25]}}, {4{maskWire[24]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_lo_hi_5 = {{4{maskWire[27]}}, {4{maskWire[26]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_lo_5 = {maskForGroupWire_lo_lo_hi_hi_lo_hi_5, maskForGroupWire_lo_lo_hi_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_lo_5 = {{4{maskWire[29]}}, {4{maskWire[28]}}};
  wire [7:0]        maskForGroupWire_lo_lo_hi_hi_hi_hi_5 = {{4{maskWire[31]}}, {4{maskWire[30]}}};
  wire [15:0]       maskForGroupWire_lo_lo_hi_hi_hi_5 = {maskForGroupWire_lo_lo_hi_hi_hi_hi_5, maskForGroupWire_lo_lo_hi_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_lo_hi_hi_5 = {maskForGroupWire_lo_lo_hi_hi_hi_5, maskForGroupWire_lo_lo_hi_hi_lo_5};
  wire [63:0]       maskForGroupWire_lo_lo_hi_5 = {maskForGroupWire_lo_lo_hi_hi_5, maskForGroupWire_lo_lo_hi_lo_5};
  wire [127:0]      maskForGroupWire_lo_lo_5 = {maskForGroupWire_lo_lo_hi_5, maskForGroupWire_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_lo_5 = {{4{maskWire[33]}}, {4{maskWire[32]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_lo_hi_5 = {{4{maskWire[35]}}, {4{maskWire[34]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_lo_5 = {maskForGroupWire_lo_hi_lo_lo_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_lo_5 = {{4{maskWire[37]}}, {4{maskWire[36]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_lo_hi_hi_5 = {{4{maskWire[39]}}, {4{maskWire[38]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_lo_hi_5 = {maskForGroupWire_lo_hi_lo_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_hi_lo_lo_5 = {maskForGroupWire_lo_hi_lo_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_lo_5 = {{4{maskWire[41]}}, {4{maskWire[40]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_lo_hi_5 = {{4{maskWire[43]}}, {4{maskWire[42]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_lo_5 = {maskForGroupWire_lo_hi_lo_hi_lo_hi_5, maskForGroupWire_lo_hi_lo_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_lo_5 = {{4{maskWire[45]}}, {4{maskWire[44]}}};
  wire [7:0]        maskForGroupWire_lo_hi_lo_hi_hi_hi_5 = {{4{maskWire[47]}}, {4{maskWire[46]}}};
  wire [15:0]       maskForGroupWire_lo_hi_lo_hi_hi_5 = {maskForGroupWire_lo_hi_lo_hi_hi_hi_5, maskForGroupWire_lo_hi_lo_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_hi_lo_hi_5 = {maskForGroupWire_lo_hi_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_hi_lo_5};
  wire [63:0]       maskForGroupWire_lo_hi_lo_5 = {maskForGroupWire_lo_hi_lo_hi_5, maskForGroupWire_lo_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_lo_5 = {{4{maskWire[49]}}, {4{maskWire[48]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_lo_hi_5 = {{4{maskWire[51]}}, {4{maskWire[50]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_lo_5 = {maskForGroupWire_lo_hi_hi_lo_lo_hi_5, maskForGroupWire_lo_hi_hi_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_lo_5 = {{4{maskWire[53]}}, {4{maskWire[52]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_lo_hi_hi_5 = {{4{maskWire[55]}}, {4{maskWire[54]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_lo_hi_5 = {maskForGroupWire_lo_hi_hi_lo_hi_hi_5, maskForGroupWire_lo_hi_hi_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_hi_hi_lo_5 = {maskForGroupWire_lo_hi_hi_lo_hi_5, maskForGroupWire_lo_hi_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_lo_5 = {{4{maskWire[57]}}, {4{maskWire[56]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_lo_hi_5 = {{4{maskWire[59]}}, {4{maskWire[58]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_lo_5 = {maskForGroupWire_lo_hi_hi_hi_lo_hi_5, maskForGroupWire_lo_hi_hi_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_lo_5 = {{4{maskWire[61]}}, {4{maskWire[60]}}};
  wire [7:0]        maskForGroupWire_lo_hi_hi_hi_hi_hi_5 = {{4{maskWire[63]}}, {4{maskWire[62]}}};
  wire [15:0]       maskForGroupWire_lo_hi_hi_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_lo_hi_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_hi_lo_5};
  wire [63:0]       maskForGroupWire_lo_hi_hi_5 = {maskForGroupWire_lo_hi_hi_hi_5, maskForGroupWire_lo_hi_hi_lo_5};
  wire [127:0]      maskForGroupWire_lo_hi_5 = {maskForGroupWire_lo_hi_hi_5, maskForGroupWire_lo_hi_lo_5};
  wire [255:0]      maskForGroupWire_lo_5 = {maskForGroupWire_lo_hi_5, maskForGroupWire_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_lo_5 = {{4{maskWire[65]}}, {4{maskWire[64]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_lo_hi_5 = {{4{maskWire[67]}}, {4{maskWire[66]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_lo_5 = {maskForGroupWire_hi_lo_lo_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_lo_5 = {{4{maskWire[69]}}, {4{maskWire[68]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_lo_hi_hi_5 = {{4{maskWire[71]}}, {4{maskWire[70]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_lo_hi_5 = {maskForGroupWire_hi_lo_lo_lo_hi_hi_5, maskForGroupWire_hi_lo_lo_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_lo_lo_lo_5 = {maskForGroupWire_hi_lo_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_lo_5 = {{4{maskWire[73]}}, {4{maskWire[72]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_lo_hi_5 = {{4{maskWire[75]}}, {4{maskWire[74]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_lo_5 = {maskForGroupWire_hi_lo_lo_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_lo_5 = {{4{maskWire[77]}}, {4{maskWire[76]}}};
  wire [7:0]        maskForGroupWire_hi_lo_lo_hi_hi_hi_5 = {{4{maskWire[79]}}, {4{maskWire[78]}}};
  wire [15:0]       maskForGroupWire_hi_lo_lo_hi_hi_5 = {maskForGroupWire_hi_lo_lo_hi_hi_hi_5, maskForGroupWire_hi_lo_lo_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_lo_lo_hi_5 = {maskForGroupWire_hi_lo_lo_hi_hi_5, maskForGroupWire_hi_lo_lo_hi_lo_5};
  wire [63:0]       maskForGroupWire_hi_lo_lo_5 = {maskForGroupWire_hi_lo_lo_hi_5, maskForGroupWire_hi_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_lo_5 = {{4{maskWire[81]}}, {4{maskWire[80]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_lo_hi_5 = {{4{maskWire[83]}}, {4{maskWire[82]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_lo_5 = {maskForGroupWire_hi_lo_hi_lo_lo_hi_5, maskForGroupWire_hi_lo_hi_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_lo_5 = {{4{maskWire[85]}}, {4{maskWire[84]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_lo_hi_hi_5 = {{4{maskWire[87]}}, {4{maskWire[86]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_lo_hi_5 = {maskForGroupWire_hi_lo_hi_lo_hi_hi_5, maskForGroupWire_hi_lo_hi_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_lo_hi_lo_5 = {maskForGroupWire_hi_lo_hi_lo_hi_5, maskForGroupWire_hi_lo_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_lo_5 = {{4{maskWire[89]}}, {4{maskWire[88]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_lo_hi_5 = {{4{maskWire[91]}}, {4{maskWire[90]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_lo_5 = {maskForGroupWire_hi_lo_hi_hi_lo_hi_5, maskForGroupWire_hi_lo_hi_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_lo_5 = {{4{maskWire[93]}}, {4{maskWire[92]}}};
  wire [7:0]        maskForGroupWire_hi_lo_hi_hi_hi_hi_5 = {{4{maskWire[95]}}, {4{maskWire[94]}}};
  wire [15:0]       maskForGroupWire_hi_lo_hi_hi_hi_5 = {maskForGroupWire_hi_lo_hi_hi_hi_hi_5, maskForGroupWire_hi_lo_hi_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_lo_hi_hi_5 = {maskForGroupWire_hi_lo_hi_hi_hi_5, maskForGroupWire_hi_lo_hi_hi_lo_5};
  wire [63:0]       maskForGroupWire_hi_lo_hi_5 = {maskForGroupWire_hi_lo_hi_hi_5, maskForGroupWire_hi_lo_hi_lo_5};
  wire [127:0]      maskForGroupWire_hi_lo_5 = {maskForGroupWire_hi_lo_hi_5, maskForGroupWire_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_lo_5 = {{4{maskWire[97]}}, {4{maskWire[96]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_lo_hi_5 = {{4{maskWire[99]}}, {4{maskWire[98]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_lo_5 = {maskForGroupWire_hi_hi_lo_lo_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_lo_5 = {{4{maskWire[101]}}, {4{maskWire[100]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_lo_hi_hi_5 = {{4{maskWire[103]}}, {4{maskWire[102]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_lo_hi_5 = {maskForGroupWire_hi_hi_lo_lo_hi_hi_5, maskForGroupWire_hi_hi_lo_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_hi_lo_lo_5 = {maskForGroupWire_hi_hi_lo_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_lo_5 = {{4{maskWire[105]}}, {4{maskWire[104]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_lo_hi_5 = {{4{maskWire[107]}}, {4{maskWire[106]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_lo_5 = {maskForGroupWire_hi_hi_lo_hi_lo_hi_5, maskForGroupWire_hi_hi_lo_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_lo_5 = {{4{maskWire[109]}}, {4{maskWire[108]}}};
  wire [7:0]        maskForGroupWire_hi_hi_lo_hi_hi_hi_5 = {{4{maskWire[111]}}, {4{maskWire[110]}}};
  wire [15:0]       maskForGroupWire_hi_hi_lo_hi_hi_5 = {maskForGroupWire_hi_hi_lo_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_hi_lo_hi_5 = {maskForGroupWire_hi_hi_lo_hi_hi_5, maskForGroupWire_hi_hi_lo_hi_lo_5};
  wire [63:0]       maskForGroupWire_hi_hi_lo_5 = {maskForGroupWire_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_lo_5 = {{4{maskWire[113]}}, {4{maskWire[112]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_lo_hi_5 = {{4{maskWire[115]}}, {4{maskWire[114]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_lo_5 = {maskForGroupWire_hi_hi_hi_lo_lo_hi_5, maskForGroupWire_hi_hi_hi_lo_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_lo_5 = {{4{maskWire[117]}}, {4{maskWire[116]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_lo_hi_hi_5 = {{4{maskWire[119]}}, {4{maskWire[118]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_lo_hi_5 = {maskForGroupWire_hi_hi_hi_lo_hi_hi_5, maskForGroupWire_hi_hi_hi_lo_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_hi_hi_lo_5 = {maskForGroupWire_hi_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_lo_5 = {{4{maskWire[121]}}, {4{maskWire[120]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_lo_hi_5 = {{4{maskWire[123]}}, {4{maskWire[122]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_lo_5 = {maskForGroupWire_hi_hi_hi_hi_lo_hi_5, maskForGroupWire_hi_hi_hi_hi_lo_lo_5};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_lo_5 = {{4{maskWire[125]}}, {4{maskWire[124]}}};
  wire [7:0]        maskForGroupWire_hi_hi_hi_hi_hi_hi_5 = {{4{maskWire[127]}}, {4{maskWire[126]}}};
  wire [15:0]       maskForGroupWire_hi_hi_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_hi_hi_lo_5};
  wire [31:0]       maskForGroupWire_hi_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_hi_lo_5};
  wire [63:0]       maskForGroupWire_hi_hi_hi_5 = {maskForGroupWire_hi_hi_hi_hi_5, maskForGroupWire_hi_hi_hi_lo_5};
  wire [127:0]      maskForGroupWire_hi_hi_5 = {maskForGroupWire_hi_hi_hi_5, maskForGroupWire_hi_hi_lo_5};
  wire [255:0]      maskForGroupWire_hi_5 = {maskForGroupWire_hi_hi_5, maskForGroupWire_hi_lo_5};
  wire [127:0]      maskForGroupWire =
    (dataEEWOH[0] ? maskWire : 128'h0) | (dataEEWOH[1] ? (maskCounterInGroup[0] ? maskForGroupWire_hi : maskForGroupWire_lo_1) : 128'h0)
    | (dataEEWOH[2]
         ? (_maskForGroupWire_T_517[0] ? maskForGroupWire_lo_2[127:0] : 128'h0) | (_maskForGroupWire_T_517[1] ? maskForGroupWire_lo_3[255:128] : 128'h0) | (_maskForGroupWire_T_517[2] ? maskForGroupWire_hi_4[127:0] : 128'h0)
           | (_maskForGroupWire_T_517[3] ? maskForGroupWire_hi_5[255:128] : 128'h0)
         : 128'h0);
  wire [1:0]        initSendState_lo = maskForGroupWire[1:0];
  wire [1:0]        fillBySeg_lo_lo_lo_lo_lo_lo = maskForGroupWire[1:0];
  wire [1:0]        initSendState_hi = maskForGroupWire[3:2];
  wire [1:0]        fillBySeg_lo_lo_lo_lo_lo_hi = maskForGroupWire[3:2];
  wire              initSendState_0 = |{initSendState_hi, initSendState_lo};
  wire [1:0]        initSendState_lo_1 = maskForGroupWire[5:4];
  wire [1:0]        fillBySeg_lo_lo_lo_lo_hi_lo = maskForGroupWire[5:4];
  wire [1:0]        initSendState_hi_1 = maskForGroupWire[7:6];
  wire [1:0]        fillBySeg_lo_lo_lo_lo_hi_hi = maskForGroupWire[7:6];
  wire              initSendState_1 = |{initSendState_hi_1, initSendState_lo_1};
  wire [1:0]        initSendState_lo_2 = maskForGroupWire[9:8];
  wire [1:0]        fillBySeg_lo_lo_lo_hi_lo_lo = maskForGroupWire[9:8];
  wire [1:0]        initSendState_hi_2 = maskForGroupWire[11:10];
  wire [1:0]        fillBySeg_lo_lo_lo_hi_lo_hi = maskForGroupWire[11:10];
  wire              initSendState_2 = |{initSendState_hi_2, initSendState_lo_2};
  wire [1:0]        initSendState_lo_3 = maskForGroupWire[13:12];
  wire [1:0]        fillBySeg_lo_lo_lo_hi_hi_lo = maskForGroupWire[13:12];
  wire [1:0]        initSendState_hi_3 = maskForGroupWire[15:14];
  wire [1:0]        fillBySeg_lo_lo_lo_hi_hi_hi = maskForGroupWire[15:14];
  wire              initSendState_3 = |{initSendState_hi_3, initSendState_lo_3};
  wire [1:0]        initSendState_lo_4 = maskForGroupWire[17:16];
  wire [1:0]        fillBySeg_lo_lo_hi_lo_lo_lo = maskForGroupWire[17:16];
  wire [1:0]        initSendState_hi_4 = maskForGroupWire[19:18];
  wire [1:0]        fillBySeg_lo_lo_hi_lo_lo_hi = maskForGroupWire[19:18];
  wire              initSendState_4 = |{initSendState_hi_4, initSendState_lo_4};
  wire [1:0]        initSendState_lo_5 = maskForGroupWire[21:20];
  wire [1:0]        fillBySeg_lo_lo_hi_lo_hi_lo = maskForGroupWire[21:20];
  wire [1:0]        initSendState_hi_5 = maskForGroupWire[23:22];
  wire [1:0]        fillBySeg_lo_lo_hi_lo_hi_hi = maskForGroupWire[23:22];
  wire              initSendState_5 = |{initSendState_hi_5, initSendState_lo_5};
  wire [1:0]        initSendState_lo_6 = maskForGroupWire[25:24];
  wire [1:0]        fillBySeg_lo_lo_hi_hi_lo_lo = maskForGroupWire[25:24];
  wire [1:0]        initSendState_hi_6 = maskForGroupWire[27:26];
  wire [1:0]        fillBySeg_lo_lo_hi_hi_lo_hi = maskForGroupWire[27:26];
  wire              initSendState_6 = |{initSendState_hi_6, initSendState_lo_6};
  wire [1:0]        initSendState_lo_7 = maskForGroupWire[29:28];
  wire [1:0]        fillBySeg_lo_lo_hi_hi_hi_lo = maskForGroupWire[29:28];
  wire [1:0]        initSendState_hi_7 = maskForGroupWire[31:30];
  wire [1:0]        fillBySeg_lo_lo_hi_hi_hi_hi = maskForGroupWire[31:30];
  wire              initSendState_7 = |{initSendState_hi_7, initSendState_lo_7};
  wire [1:0]        initSendState_lo_8 = maskForGroupWire[33:32];
  wire [1:0]        fillBySeg_lo_hi_lo_lo_lo_lo = maskForGroupWire[33:32];
  wire [1:0]        initSendState_hi_8 = maskForGroupWire[35:34];
  wire [1:0]        fillBySeg_lo_hi_lo_lo_lo_hi = maskForGroupWire[35:34];
  wire              initSendState_8 = |{initSendState_hi_8, initSendState_lo_8};
  wire [1:0]        initSendState_lo_9 = maskForGroupWire[37:36];
  wire [1:0]        fillBySeg_lo_hi_lo_lo_hi_lo = maskForGroupWire[37:36];
  wire [1:0]        initSendState_hi_9 = maskForGroupWire[39:38];
  wire [1:0]        fillBySeg_lo_hi_lo_lo_hi_hi = maskForGroupWire[39:38];
  wire              initSendState_9 = |{initSendState_hi_9, initSendState_lo_9};
  wire [1:0]        initSendState_lo_10 = maskForGroupWire[41:40];
  wire [1:0]        fillBySeg_lo_hi_lo_hi_lo_lo = maskForGroupWire[41:40];
  wire [1:0]        initSendState_hi_10 = maskForGroupWire[43:42];
  wire [1:0]        fillBySeg_lo_hi_lo_hi_lo_hi = maskForGroupWire[43:42];
  wire              initSendState_10 = |{initSendState_hi_10, initSendState_lo_10};
  wire [1:0]        initSendState_lo_11 = maskForGroupWire[45:44];
  wire [1:0]        fillBySeg_lo_hi_lo_hi_hi_lo = maskForGroupWire[45:44];
  wire [1:0]        initSendState_hi_11 = maskForGroupWire[47:46];
  wire [1:0]        fillBySeg_lo_hi_lo_hi_hi_hi = maskForGroupWire[47:46];
  wire              initSendState_11 = |{initSendState_hi_11, initSendState_lo_11};
  wire [1:0]        initSendState_lo_12 = maskForGroupWire[49:48];
  wire [1:0]        fillBySeg_lo_hi_hi_lo_lo_lo = maskForGroupWire[49:48];
  wire [1:0]        initSendState_hi_12 = maskForGroupWire[51:50];
  wire [1:0]        fillBySeg_lo_hi_hi_lo_lo_hi = maskForGroupWire[51:50];
  wire              initSendState_12 = |{initSendState_hi_12, initSendState_lo_12};
  wire [1:0]        initSendState_lo_13 = maskForGroupWire[53:52];
  wire [1:0]        fillBySeg_lo_hi_hi_lo_hi_lo = maskForGroupWire[53:52];
  wire [1:0]        initSendState_hi_13 = maskForGroupWire[55:54];
  wire [1:0]        fillBySeg_lo_hi_hi_lo_hi_hi = maskForGroupWire[55:54];
  wire              initSendState_13 = |{initSendState_hi_13, initSendState_lo_13};
  wire [1:0]        initSendState_lo_14 = maskForGroupWire[57:56];
  wire [1:0]        fillBySeg_lo_hi_hi_hi_lo_lo = maskForGroupWire[57:56];
  wire [1:0]        initSendState_hi_14 = maskForGroupWire[59:58];
  wire [1:0]        fillBySeg_lo_hi_hi_hi_lo_hi = maskForGroupWire[59:58];
  wire              initSendState_14 = |{initSendState_hi_14, initSendState_lo_14};
  wire [1:0]        initSendState_lo_15 = maskForGroupWire[61:60];
  wire [1:0]        fillBySeg_lo_hi_hi_hi_hi_lo = maskForGroupWire[61:60];
  wire [1:0]        initSendState_hi_15 = maskForGroupWire[63:62];
  wire [1:0]        fillBySeg_lo_hi_hi_hi_hi_hi = maskForGroupWire[63:62];
  wire              initSendState_15 = |{initSendState_hi_15, initSendState_lo_15};
  wire [1:0]        initSendState_lo_16 = maskForGroupWire[65:64];
  wire [1:0]        fillBySeg_hi_lo_lo_lo_lo_lo = maskForGroupWire[65:64];
  wire [1:0]        initSendState_hi_16 = maskForGroupWire[67:66];
  wire [1:0]        fillBySeg_hi_lo_lo_lo_lo_hi = maskForGroupWire[67:66];
  wire              initSendState_16 = |{initSendState_hi_16, initSendState_lo_16};
  wire [1:0]        initSendState_lo_17 = maskForGroupWire[69:68];
  wire [1:0]        fillBySeg_hi_lo_lo_lo_hi_lo = maskForGroupWire[69:68];
  wire [1:0]        initSendState_hi_17 = maskForGroupWire[71:70];
  wire [1:0]        fillBySeg_hi_lo_lo_lo_hi_hi = maskForGroupWire[71:70];
  wire              initSendState_17 = |{initSendState_hi_17, initSendState_lo_17};
  wire [1:0]        initSendState_lo_18 = maskForGroupWire[73:72];
  wire [1:0]        fillBySeg_hi_lo_lo_hi_lo_lo = maskForGroupWire[73:72];
  wire [1:0]        initSendState_hi_18 = maskForGroupWire[75:74];
  wire [1:0]        fillBySeg_hi_lo_lo_hi_lo_hi = maskForGroupWire[75:74];
  wire              initSendState_18 = |{initSendState_hi_18, initSendState_lo_18};
  wire [1:0]        initSendState_lo_19 = maskForGroupWire[77:76];
  wire [1:0]        fillBySeg_hi_lo_lo_hi_hi_lo = maskForGroupWire[77:76];
  wire [1:0]        initSendState_hi_19 = maskForGroupWire[79:78];
  wire [1:0]        fillBySeg_hi_lo_lo_hi_hi_hi = maskForGroupWire[79:78];
  wire              initSendState_19 = |{initSendState_hi_19, initSendState_lo_19};
  wire [1:0]        initSendState_lo_20 = maskForGroupWire[81:80];
  wire [1:0]        fillBySeg_hi_lo_hi_lo_lo_lo = maskForGroupWire[81:80];
  wire [1:0]        initSendState_hi_20 = maskForGroupWire[83:82];
  wire [1:0]        fillBySeg_hi_lo_hi_lo_lo_hi = maskForGroupWire[83:82];
  wire              initSendState_20 = |{initSendState_hi_20, initSendState_lo_20};
  wire [1:0]        initSendState_lo_21 = maskForGroupWire[85:84];
  wire [1:0]        fillBySeg_hi_lo_hi_lo_hi_lo = maskForGroupWire[85:84];
  wire [1:0]        initSendState_hi_21 = maskForGroupWire[87:86];
  wire [1:0]        fillBySeg_hi_lo_hi_lo_hi_hi = maskForGroupWire[87:86];
  wire              initSendState_21 = |{initSendState_hi_21, initSendState_lo_21};
  wire [1:0]        initSendState_lo_22 = maskForGroupWire[89:88];
  wire [1:0]        fillBySeg_hi_lo_hi_hi_lo_lo = maskForGroupWire[89:88];
  wire [1:0]        initSendState_hi_22 = maskForGroupWire[91:90];
  wire [1:0]        fillBySeg_hi_lo_hi_hi_lo_hi = maskForGroupWire[91:90];
  wire              initSendState_22 = |{initSendState_hi_22, initSendState_lo_22};
  wire [1:0]        initSendState_lo_23 = maskForGroupWire[93:92];
  wire [1:0]        fillBySeg_hi_lo_hi_hi_hi_lo = maskForGroupWire[93:92];
  wire [1:0]        initSendState_hi_23 = maskForGroupWire[95:94];
  wire [1:0]        fillBySeg_hi_lo_hi_hi_hi_hi = maskForGroupWire[95:94];
  wire              initSendState_23 = |{initSendState_hi_23, initSendState_lo_23};
  wire [1:0]        initSendState_lo_24 = maskForGroupWire[97:96];
  wire [1:0]        fillBySeg_hi_hi_lo_lo_lo_lo = maskForGroupWire[97:96];
  wire [1:0]        initSendState_hi_24 = maskForGroupWire[99:98];
  wire [1:0]        fillBySeg_hi_hi_lo_lo_lo_hi = maskForGroupWire[99:98];
  wire              initSendState_24 = |{initSendState_hi_24, initSendState_lo_24};
  wire [1:0]        initSendState_lo_25 = maskForGroupWire[101:100];
  wire [1:0]        fillBySeg_hi_hi_lo_lo_hi_lo = maskForGroupWire[101:100];
  wire [1:0]        initSendState_hi_25 = maskForGroupWire[103:102];
  wire [1:0]        fillBySeg_hi_hi_lo_lo_hi_hi = maskForGroupWire[103:102];
  wire              initSendState_25 = |{initSendState_hi_25, initSendState_lo_25};
  wire [1:0]        initSendState_lo_26 = maskForGroupWire[105:104];
  wire [1:0]        fillBySeg_hi_hi_lo_hi_lo_lo = maskForGroupWire[105:104];
  wire [1:0]        initSendState_hi_26 = maskForGroupWire[107:106];
  wire [1:0]        fillBySeg_hi_hi_lo_hi_lo_hi = maskForGroupWire[107:106];
  wire              initSendState_26 = |{initSendState_hi_26, initSendState_lo_26};
  wire [1:0]        initSendState_lo_27 = maskForGroupWire[109:108];
  wire [1:0]        fillBySeg_hi_hi_lo_hi_hi_lo = maskForGroupWire[109:108];
  wire [1:0]        initSendState_hi_27 = maskForGroupWire[111:110];
  wire [1:0]        fillBySeg_hi_hi_lo_hi_hi_hi = maskForGroupWire[111:110];
  wire              initSendState_27 = |{initSendState_hi_27, initSendState_lo_27};
  wire [1:0]        initSendState_lo_28 = maskForGroupWire[113:112];
  wire [1:0]        fillBySeg_hi_hi_hi_lo_lo_lo = maskForGroupWire[113:112];
  wire [1:0]        initSendState_hi_28 = maskForGroupWire[115:114];
  wire [1:0]        fillBySeg_hi_hi_hi_lo_lo_hi = maskForGroupWire[115:114];
  wire              initSendState_28 = |{initSendState_hi_28, initSendState_lo_28};
  wire [1:0]        initSendState_lo_29 = maskForGroupWire[117:116];
  wire [1:0]        fillBySeg_hi_hi_hi_lo_hi_lo = maskForGroupWire[117:116];
  wire [1:0]        initSendState_hi_29 = maskForGroupWire[119:118];
  wire [1:0]        fillBySeg_hi_hi_hi_lo_hi_hi = maskForGroupWire[119:118];
  wire              initSendState_29 = |{initSendState_hi_29, initSendState_lo_29};
  wire [1:0]        initSendState_lo_30 = maskForGroupWire[121:120];
  wire [1:0]        fillBySeg_hi_hi_hi_hi_lo_lo = maskForGroupWire[121:120];
  wire [1:0]        initSendState_hi_30 = maskForGroupWire[123:122];
  wire [1:0]        fillBySeg_hi_hi_hi_hi_lo_hi = maskForGroupWire[123:122];
  wire              initSendState_30 = |{initSendState_hi_30, initSendState_lo_30};
  wire [1:0]        initSendState_lo_31 = maskForGroupWire[125:124];
  wire [1:0]        fillBySeg_hi_hi_hi_hi_hi_lo = maskForGroupWire[125:124];
  wire [1:0]        initSendState_hi_31 = maskForGroupWire[127:126];
  wire [1:0]        fillBySeg_hi_hi_hi_hi_hi_hi = maskForGroupWire[127:126];
  wire              initSendState_31 = |{initSendState_hi_31, initSendState_lo_31};
  reg  [1023:0]     accessData_0;
  wire [1023:0]     accessDataUpdate_1 = accessData_0;
  reg  [1023:0]     accessData_1;
  wire [1023:0]     accessDataUpdate_2 = accessData_1;
  reg  [1023:0]     accessData_2;
  wire [1023:0]     accessDataUpdate_3 = accessData_2;
  reg  [1023:0]     accessData_3;
  wire [1023:0]     accessDataUpdate_4 = accessData_3;
  reg  [1023:0]     accessData_4;
  wire [1023:0]     accessDataUpdate_5 = accessData_4;
  reg  [1023:0]     accessData_5;
  wire [1023:0]     accessDataUpdate_6 = accessData_5;
  reg  [1023:0]     accessData_6;
  wire [1023:0]     accessDataUpdate_7 = accessData_6;
  reg  [1023:0]     accessData_7;
  reg  [2:0]        accessPtr;
  reg  [2:0]        dataGroup;
  reg  [1023:0]     dataBuffer_0;
  reg  [1023:0]     dataBuffer_1;
  reg  [1023:0]     dataBuffer_2;
  reg  [1023:0]     dataBuffer_3;
  reg  [1023:0]     dataBuffer_4;
  reg  [1023:0]     dataBuffer_5;
  reg  [1023:0]     dataBuffer_6;
  reg  [1023:0]     dataBuffer_7;
  reg  [3:0]        bufferBaseCacheLineIndex;
  wire [3:0]        memRequest_bits_index_0 = bufferBaseCacheLineIndex;
  reg  [2:0]        cacheLineIndexInBuffer;
  wire [6:0]        initOffset = lsuRequestReg_rs1Data[6:0];
  wire              invalidInstruction = csrInterface_vl == 11'h0;
  reg               invalidInstructionNext;
  wire              wholeType = lsuRequest_bits_instructionInformation_lumop[3];
  wire [2:0]        nfCorrection = wholeType ? 3'h0 : lsuRequest_bits_instructionInformation_nf;
  reg  [3:0]        segmentInstructionIndexInterval;
  wire [17:0]       bytePerInstruction = {3'h0, {11'h0, {1'h0, nfCorrection} + 4'h1} * {4'h0, csrInterface_vl}} << lsuRequest_bits_instructionInformation_eew;
  wire [17:0]       accessMemSize = bytePerInstruction + {11'h0, lsuRequest_bits_rs1Data[6:0]};
  wire [10:0]       lastCacheLineIndex = accessMemSize[17:7] - {10'h0, accessMemSize[6:0] == 7'h0};
  wire [10:0]       lastWriteVrfIndex = bytePerInstruction[17:7] - {10'h0, bytePerInstruction[6:0] == 7'h0};
  reg  [10:0]       lastWriteVrfIndexReg;
  reg               lastCacheNeedPush;
  reg  [10:0]       cacheLineNumberReg;
  wire [13:0]       dataByteSize = {3'h0, csrInterface_vl} << lsuRequest_bits_instructionInformation_eew;
  wire [6:0]        lastDataGroupForInstruction = dataByteSize[13:7] - {6'h0, dataByteSize[6:0] == 7'h0};
  reg  [6:0]        lastDataGroupReg;
  wire [2:0]        nextDataGroup = lsuRequest_valid ? 3'h0 : dataGroup + 3'h1;
  wire              isLastRead = {4'h0, dataGroup} == lastDataGroupReg;
  reg               hazardCheck;
  wire              accessBufferEnqueueFire;
  wire              vrfReadQueueVec_0_deq_ready;
  wire              vrfReadQueueVec_0_enq_ready = ~_vrfReadQueueVec_fifo_full | vrfReadQueueVec_0_deq_ready;
  wire              vrfReadQueueVec_0_deq_valid = ~_vrfReadQueueVec_fifo_empty | vrfReadQueueVec_0_enq_valid;
  wire [31:0]       vrfReadQueueVec_0_deq_bits = _vrfReadQueueVec_fifo_empty ? vrfReadQueueVec_0_enq_bits : _vrfReadQueueVec_fifo_data_out;
  wire              vrfReadQueueVec_1_deq_ready;
  wire              vrfReadQueueVec_1_enq_ready = ~_vrfReadQueueVec_fifo_1_full | vrfReadQueueVec_1_deq_ready;
  wire              vrfReadQueueVec_1_deq_valid = ~_vrfReadQueueVec_fifo_1_empty | vrfReadQueueVec_1_enq_valid;
  wire [31:0]       vrfReadQueueVec_1_deq_bits = _vrfReadQueueVec_fifo_1_empty ? vrfReadQueueVec_1_enq_bits : _vrfReadQueueVec_fifo_1_data_out;
  wire              vrfReadQueueVec_2_deq_ready;
  wire              vrfReadQueueVec_2_enq_ready = ~_vrfReadQueueVec_fifo_2_full | vrfReadQueueVec_2_deq_ready;
  wire              vrfReadQueueVec_2_deq_valid = ~_vrfReadQueueVec_fifo_2_empty | vrfReadQueueVec_2_enq_valid;
  wire [31:0]       vrfReadQueueVec_2_deq_bits = _vrfReadQueueVec_fifo_2_empty ? vrfReadQueueVec_2_enq_bits : _vrfReadQueueVec_fifo_2_data_out;
  wire              vrfReadQueueVec_3_deq_ready;
  wire              vrfReadQueueVec_3_enq_ready = ~_vrfReadQueueVec_fifo_3_full | vrfReadQueueVec_3_deq_ready;
  wire              vrfReadQueueVec_3_deq_valid = ~_vrfReadQueueVec_fifo_3_empty | vrfReadQueueVec_3_enq_valid;
  wire [31:0]       vrfReadQueueVec_3_deq_bits = _vrfReadQueueVec_fifo_3_empty ? vrfReadQueueVec_3_enq_bits : _vrfReadQueueVec_fifo_3_data_out;
  wire              vrfReadQueueVec_4_deq_ready;
  wire              vrfReadQueueVec_4_enq_ready = ~_vrfReadQueueVec_fifo_4_full | vrfReadQueueVec_4_deq_ready;
  wire              vrfReadQueueVec_4_deq_valid = ~_vrfReadQueueVec_fifo_4_empty | vrfReadQueueVec_4_enq_valid;
  wire [31:0]       vrfReadQueueVec_4_deq_bits = _vrfReadQueueVec_fifo_4_empty ? vrfReadQueueVec_4_enq_bits : _vrfReadQueueVec_fifo_4_data_out;
  wire              vrfReadQueueVec_5_deq_ready;
  wire              vrfReadQueueVec_5_enq_ready = ~_vrfReadQueueVec_fifo_5_full | vrfReadQueueVec_5_deq_ready;
  wire              vrfReadQueueVec_5_deq_valid = ~_vrfReadQueueVec_fifo_5_empty | vrfReadQueueVec_5_enq_valid;
  wire [31:0]       vrfReadQueueVec_5_deq_bits = _vrfReadQueueVec_fifo_5_empty ? vrfReadQueueVec_5_enq_bits : _vrfReadQueueVec_fifo_5_data_out;
  wire              vrfReadQueueVec_6_deq_ready;
  wire              vrfReadQueueVec_6_enq_ready = ~_vrfReadQueueVec_fifo_6_full | vrfReadQueueVec_6_deq_ready;
  wire              vrfReadQueueVec_6_deq_valid = ~_vrfReadQueueVec_fifo_6_empty | vrfReadQueueVec_6_enq_valid;
  wire [31:0]       vrfReadQueueVec_6_deq_bits = _vrfReadQueueVec_fifo_6_empty ? vrfReadQueueVec_6_enq_bits : _vrfReadQueueVec_fifo_6_data_out;
  wire              vrfReadQueueVec_7_deq_ready;
  wire              vrfReadQueueVec_7_enq_ready = ~_vrfReadQueueVec_fifo_7_full | vrfReadQueueVec_7_deq_ready;
  wire              vrfReadQueueVec_7_deq_valid = ~_vrfReadQueueVec_fifo_7_empty | vrfReadQueueVec_7_enq_valid;
  wire [31:0]       vrfReadQueueVec_7_deq_bits = _vrfReadQueueVec_fifo_7_empty ? vrfReadQueueVec_7_enq_bits : _vrfReadQueueVec_fifo_7_data_out;
  wire              vrfReadQueueVec_8_deq_ready;
  wire              vrfReadQueueVec_8_enq_ready = ~_vrfReadQueueVec_fifo_8_full | vrfReadQueueVec_8_deq_ready;
  wire              vrfReadQueueVec_8_deq_valid = ~_vrfReadQueueVec_fifo_8_empty | vrfReadQueueVec_8_enq_valid;
  wire [31:0]       vrfReadQueueVec_8_deq_bits = _vrfReadQueueVec_fifo_8_empty ? vrfReadQueueVec_8_enq_bits : _vrfReadQueueVec_fifo_8_data_out;
  wire              vrfReadQueueVec_9_deq_ready;
  wire              vrfReadQueueVec_9_enq_ready = ~_vrfReadQueueVec_fifo_9_full | vrfReadQueueVec_9_deq_ready;
  wire              vrfReadQueueVec_9_deq_valid = ~_vrfReadQueueVec_fifo_9_empty | vrfReadQueueVec_9_enq_valid;
  wire [31:0]       vrfReadQueueVec_9_deq_bits = _vrfReadQueueVec_fifo_9_empty ? vrfReadQueueVec_9_enq_bits : _vrfReadQueueVec_fifo_9_data_out;
  wire              vrfReadQueueVec_10_deq_ready;
  wire              vrfReadQueueVec_10_enq_ready = ~_vrfReadQueueVec_fifo_10_full | vrfReadQueueVec_10_deq_ready;
  wire              vrfReadQueueVec_10_deq_valid = ~_vrfReadQueueVec_fifo_10_empty | vrfReadQueueVec_10_enq_valid;
  wire [31:0]       vrfReadQueueVec_10_deq_bits = _vrfReadQueueVec_fifo_10_empty ? vrfReadQueueVec_10_enq_bits : _vrfReadQueueVec_fifo_10_data_out;
  wire              vrfReadQueueVec_11_deq_ready;
  wire              vrfReadQueueVec_11_enq_ready = ~_vrfReadQueueVec_fifo_11_full | vrfReadQueueVec_11_deq_ready;
  wire              vrfReadQueueVec_11_deq_valid = ~_vrfReadQueueVec_fifo_11_empty | vrfReadQueueVec_11_enq_valid;
  wire [31:0]       vrfReadQueueVec_11_deq_bits = _vrfReadQueueVec_fifo_11_empty ? vrfReadQueueVec_11_enq_bits : _vrfReadQueueVec_fifo_11_data_out;
  wire              vrfReadQueueVec_12_deq_ready;
  wire              vrfReadQueueVec_12_enq_ready = ~_vrfReadQueueVec_fifo_12_full | vrfReadQueueVec_12_deq_ready;
  wire              vrfReadQueueVec_12_deq_valid = ~_vrfReadQueueVec_fifo_12_empty | vrfReadQueueVec_12_enq_valid;
  wire [31:0]       vrfReadQueueVec_12_deq_bits = _vrfReadQueueVec_fifo_12_empty ? vrfReadQueueVec_12_enq_bits : _vrfReadQueueVec_fifo_12_data_out;
  wire              vrfReadQueueVec_13_deq_ready;
  wire              vrfReadQueueVec_13_enq_ready = ~_vrfReadQueueVec_fifo_13_full | vrfReadQueueVec_13_deq_ready;
  wire              vrfReadQueueVec_13_deq_valid = ~_vrfReadQueueVec_fifo_13_empty | vrfReadQueueVec_13_enq_valid;
  wire [31:0]       vrfReadQueueVec_13_deq_bits = _vrfReadQueueVec_fifo_13_empty ? vrfReadQueueVec_13_enq_bits : _vrfReadQueueVec_fifo_13_data_out;
  wire              vrfReadQueueVec_14_deq_ready;
  wire              vrfReadQueueVec_14_enq_ready = ~_vrfReadQueueVec_fifo_14_full | vrfReadQueueVec_14_deq_ready;
  wire              vrfReadQueueVec_14_deq_valid = ~_vrfReadQueueVec_fifo_14_empty | vrfReadQueueVec_14_enq_valid;
  wire [31:0]       vrfReadQueueVec_14_deq_bits = _vrfReadQueueVec_fifo_14_empty ? vrfReadQueueVec_14_enq_bits : _vrfReadQueueVec_fifo_14_data_out;
  wire              vrfReadQueueVec_15_deq_ready;
  wire              vrfReadQueueVec_15_enq_ready = ~_vrfReadQueueVec_fifo_15_full | vrfReadQueueVec_15_deq_ready;
  wire              vrfReadQueueVec_15_deq_valid = ~_vrfReadQueueVec_fifo_15_empty | vrfReadQueueVec_15_enq_valid;
  wire [31:0]       vrfReadQueueVec_15_deq_bits = _vrfReadQueueVec_fifo_15_empty ? vrfReadQueueVec_15_enq_bits : _vrfReadQueueVec_fifo_15_data_out;
  wire              vrfReadQueueVec_16_deq_ready;
  wire              vrfReadQueueVec_16_enq_ready = ~_vrfReadQueueVec_fifo_16_full | vrfReadQueueVec_16_deq_ready;
  wire              vrfReadQueueVec_16_deq_valid = ~_vrfReadQueueVec_fifo_16_empty | vrfReadQueueVec_16_enq_valid;
  wire [31:0]       vrfReadQueueVec_16_deq_bits = _vrfReadQueueVec_fifo_16_empty ? vrfReadQueueVec_16_enq_bits : _vrfReadQueueVec_fifo_16_data_out;
  wire              vrfReadQueueVec_17_deq_ready;
  wire              vrfReadQueueVec_17_enq_ready = ~_vrfReadQueueVec_fifo_17_full | vrfReadQueueVec_17_deq_ready;
  wire              vrfReadQueueVec_17_deq_valid = ~_vrfReadQueueVec_fifo_17_empty | vrfReadQueueVec_17_enq_valid;
  wire [31:0]       vrfReadQueueVec_17_deq_bits = _vrfReadQueueVec_fifo_17_empty ? vrfReadQueueVec_17_enq_bits : _vrfReadQueueVec_fifo_17_data_out;
  wire              vrfReadQueueVec_18_deq_ready;
  wire              vrfReadQueueVec_18_enq_ready = ~_vrfReadQueueVec_fifo_18_full | vrfReadQueueVec_18_deq_ready;
  wire              vrfReadQueueVec_18_deq_valid = ~_vrfReadQueueVec_fifo_18_empty | vrfReadQueueVec_18_enq_valid;
  wire [31:0]       vrfReadQueueVec_18_deq_bits = _vrfReadQueueVec_fifo_18_empty ? vrfReadQueueVec_18_enq_bits : _vrfReadQueueVec_fifo_18_data_out;
  wire              vrfReadQueueVec_19_deq_ready;
  wire              vrfReadQueueVec_19_enq_ready = ~_vrfReadQueueVec_fifo_19_full | vrfReadQueueVec_19_deq_ready;
  wire              vrfReadQueueVec_19_deq_valid = ~_vrfReadQueueVec_fifo_19_empty | vrfReadQueueVec_19_enq_valid;
  wire [31:0]       vrfReadQueueVec_19_deq_bits = _vrfReadQueueVec_fifo_19_empty ? vrfReadQueueVec_19_enq_bits : _vrfReadQueueVec_fifo_19_data_out;
  wire              vrfReadQueueVec_20_deq_ready;
  wire              vrfReadQueueVec_20_enq_ready = ~_vrfReadQueueVec_fifo_20_full | vrfReadQueueVec_20_deq_ready;
  wire              vrfReadQueueVec_20_deq_valid = ~_vrfReadQueueVec_fifo_20_empty | vrfReadQueueVec_20_enq_valid;
  wire [31:0]       vrfReadQueueVec_20_deq_bits = _vrfReadQueueVec_fifo_20_empty ? vrfReadQueueVec_20_enq_bits : _vrfReadQueueVec_fifo_20_data_out;
  wire              vrfReadQueueVec_21_deq_ready;
  wire              vrfReadQueueVec_21_enq_ready = ~_vrfReadQueueVec_fifo_21_full | vrfReadQueueVec_21_deq_ready;
  wire              vrfReadQueueVec_21_deq_valid = ~_vrfReadQueueVec_fifo_21_empty | vrfReadQueueVec_21_enq_valid;
  wire [31:0]       vrfReadQueueVec_21_deq_bits = _vrfReadQueueVec_fifo_21_empty ? vrfReadQueueVec_21_enq_bits : _vrfReadQueueVec_fifo_21_data_out;
  wire              vrfReadQueueVec_22_deq_ready;
  wire              vrfReadQueueVec_22_enq_ready = ~_vrfReadQueueVec_fifo_22_full | vrfReadQueueVec_22_deq_ready;
  wire              vrfReadQueueVec_22_deq_valid = ~_vrfReadQueueVec_fifo_22_empty | vrfReadQueueVec_22_enq_valid;
  wire [31:0]       vrfReadQueueVec_22_deq_bits = _vrfReadQueueVec_fifo_22_empty ? vrfReadQueueVec_22_enq_bits : _vrfReadQueueVec_fifo_22_data_out;
  wire              vrfReadQueueVec_23_deq_ready;
  wire              vrfReadQueueVec_23_enq_ready = ~_vrfReadQueueVec_fifo_23_full | vrfReadQueueVec_23_deq_ready;
  wire              vrfReadQueueVec_23_deq_valid = ~_vrfReadQueueVec_fifo_23_empty | vrfReadQueueVec_23_enq_valid;
  wire [31:0]       vrfReadQueueVec_23_deq_bits = _vrfReadQueueVec_fifo_23_empty ? vrfReadQueueVec_23_enq_bits : _vrfReadQueueVec_fifo_23_data_out;
  wire              vrfReadQueueVec_24_deq_ready;
  wire              vrfReadQueueVec_24_enq_ready = ~_vrfReadQueueVec_fifo_24_full | vrfReadQueueVec_24_deq_ready;
  wire              vrfReadQueueVec_24_deq_valid = ~_vrfReadQueueVec_fifo_24_empty | vrfReadQueueVec_24_enq_valid;
  wire [31:0]       vrfReadQueueVec_24_deq_bits = _vrfReadQueueVec_fifo_24_empty ? vrfReadQueueVec_24_enq_bits : _vrfReadQueueVec_fifo_24_data_out;
  wire              vrfReadQueueVec_25_deq_ready;
  wire              vrfReadQueueVec_25_enq_ready = ~_vrfReadQueueVec_fifo_25_full | vrfReadQueueVec_25_deq_ready;
  wire              vrfReadQueueVec_25_deq_valid = ~_vrfReadQueueVec_fifo_25_empty | vrfReadQueueVec_25_enq_valid;
  wire [31:0]       vrfReadQueueVec_25_deq_bits = _vrfReadQueueVec_fifo_25_empty ? vrfReadQueueVec_25_enq_bits : _vrfReadQueueVec_fifo_25_data_out;
  wire              vrfReadQueueVec_26_deq_ready;
  wire              vrfReadQueueVec_26_enq_ready = ~_vrfReadQueueVec_fifo_26_full | vrfReadQueueVec_26_deq_ready;
  wire              vrfReadQueueVec_26_deq_valid = ~_vrfReadQueueVec_fifo_26_empty | vrfReadQueueVec_26_enq_valid;
  wire [31:0]       vrfReadQueueVec_26_deq_bits = _vrfReadQueueVec_fifo_26_empty ? vrfReadQueueVec_26_enq_bits : _vrfReadQueueVec_fifo_26_data_out;
  wire              vrfReadQueueVec_27_deq_ready;
  wire              vrfReadQueueVec_27_enq_ready = ~_vrfReadQueueVec_fifo_27_full | vrfReadQueueVec_27_deq_ready;
  wire              vrfReadQueueVec_27_deq_valid = ~_vrfReadQueueVec_fifo_27_empty | vrfReadQueueVec_27_enq_valid;
  wire [31:0]       vrfReadQueueVec_27_deq_bits = _vrfReadQueueVec_fifo_27_empty ? vrfReadQueueVec_27_enq_bits : _vrfReadQueueVec_fifo_27_data_out;
  wire              vrfReadQueueVec_28_deq_ready;
  wire              vrfReadQueueVec_28_enq_ready = ~_vrfReadQueueVec_fifo_28_full | vrfReadQueueVec_28_deq_ready;
  wire              vrfReadQueueVec_28_deq_valid = ~_vrfReadQueueVec_fifo_28_empty | vrfReadQueueVec_28_enq_valid;
  wire [31:0]       vrfReadQueueVec_28_deq_bits = _vrfReadQueueVec_fifo_28_empty ? vrfReadQueueVec_28_enq_bits : _vrfReadQueueVec_fifo_28_data_out;
  wire              vrfReadQueueVec_29_deq_ready;
  wire              vrfReadQueueVec_29_enq_ready = ~_vrfReadQueueVec_fifo_29_full | vrfReadQueueVec_29_deq_ready;
  wire              vrfReadQueueVec_29_deq_valid = ~_vrfReadQueueVec_fifo_29_empty | vrfReadQueueVec_29_enq_valid;
  wire [31:0]       vrfReadQueueVec_29_deq_bits = _vrfReadQueueVec_fifo_29_empty ? vrfReadQueueVec_29_enq_bits : _vrfReadQueueVec_fifo_29_data_out;
  wire              vrfReadQueueVec_30_deq_ready;
  wire              vrfReadQueueVec_30_enq_ready = ~_vrfReadQueueVec_fifo_30_full | vrfReadQueueVec_30_deq_ready;
  wire              vrfReadQueueVec_30_deq_valid = ~_vrfReadQueueVec_fifo_30_empty | vrfReadQueueVec_30_enq_valid;
  wire [31:0]       vrfReadQueueVec_30_deq_bits = _vrfReadQueueVec_fifo_30_empty ? vrfReadQueueVec_30_enq_bits : _vrfReadQueueVec_fifo_30_data_out;
  wire              vrfReadQueueVec_31_deq_ready;
  wire              vrfReadQueueVec_31_enq_ready = ~_vrfReadQueueVec_fifo_31_full | vrfReadQueueVec_31_deq_ready;
  wire              vrfReadQueueVec_31_deq_valid = ~_vrfReadQueueVec_fifo_31_empty | vrfReadQueueVec_31_enq_valid;
  wire [31:0]       vrfReadQueueVec_31_deq_bits = _vrfReadQueueVec_fifo_31_empty ? vrfReadQueueVec_31_enq_bits : _vrfReadQueueVec_fifo_31_data_out;
  reg  [2:0]        readStageValid_segPtr;
  reg  [2:0]        readStageValid_readCount;
  reg               readStageValid_stageValid;
  wire              readStageValid_lastReadPtr = readStageValid_segPtr == 3'h0;
  wire [2:0]        readStageValid_nextReadCount = lsuRequest_valid ? 3'h0 : readStageValid_readCount + 3'h1;
  wire              readStageValid_lastReadGroup = {4'h0, readStageValid_readCount} == lastDataGroupReg;
  wire              vrfReadDataPorts_0_valid_0;
  wire              _readStageValid_T_11 = vrfReadDataPorts_0_ready_0 & vrfReadDataPorts_0_valid_0;
  reg  [3:0]        readStageValid_readCounter;
  wire [3:0]        readStageValid_counterChange = _readStageValid_T_11 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_0_valid_0 = readStageValid_stageValid & ~(readStageValid_readCounter[3]);
  wire [4:0]        _GEN_5 = {1'h0, segmentInstructionIndexInterval};
  wire [4:0]        vrfReadDataPorts_0_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr} * _GEN_5 + {2'h0, readStageValid_readCount};
  reg  [2:0]        readStageValid_segPtr_1;
  reg  [2:0]        readStageValid_readCount_1;
  reg               readStageValid_stageValid_1;
  wire              readStageValid_lastReadPtr_1 = readStageValid_segPtr_1 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_1 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_1 + 3'h1;
  wire              readStageValid_lastReadGroup_1 = {4'h0, readStageValid_readCount_1} == lastDataGroupReg;
  wire              vrfReadDataPorts_1_valid_0;
  wire              _readStageValid_T_30 = vrfReadDataPorts_1_ready_0 & vrfReadDataPorts_1_valid_0;
  reg  [3:0]        readStageValid_readCounter_1;
  wire [3:0]        readStageValid_counterChange_1 = _readStageValid_T_30 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_1_valid_0 = readStageValid_stageValid_1 & ~(readStageValid_readCounter_1[3]);
  wire [4:0]        vrfReadDataPorts_1_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_1} * _GEN_5 + {2'h0, readStageValid_readCount_1};
  reg  [2:0]        readStageValid_segPtr_2;
  reg  [2:0]        readStageValid_readCount_2;
  reg               readStageValid_stageValid_2;
  wire              readStageValid_lastReadPtr_2 = readStageValid_segPtr_2 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_2 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_2 + 3'h1;
  wire              readStageValid_lastReadGroup_2 = {4'h0, readStageValid_readCount_2} == lastDataGroupReg;
  wire              vrfReadDataPorts_2_valid_0;
  wire              _readStageValid_T_49 = vrfReadDataPorts_2_ready_0 & vrfReadDataPorts_2_valid_0;
  reg  [3:0]        readStageValid_readCounter_2;
  wire [3:0]        readStageValid_counterChange_2 = _readStageValid_T_49 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_2_valid_0 = readStageValid_stageValid_2 & ~(readStageValid_readCounter_2[3]);
  wire [4:0]        vrfReadDataPorts_2_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_2} * _GEN_5 + {2'h0, readStageValid_readCount_2};
  reg  [2:0]        readStageValid_segPtr_3;
  reg  [2:0]        readStageValid_readCount_3;
  reg               readStageValid_stageValid_3;
  wire              readStageValid_lastReadPtr_3 = readStageValid_segPtr_3 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_3 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_3 + 3'h1;
  wire              readStageValid_lastReadGroup_3 = {4'h0, readStageValid_readCount_3} == lastDataGroupReg;
  wire              vrfReadDataPorts_3_valid_0;
  wire              _readStageValid_T_68 = vrfReadDataPorts_3_ready_0 & vrfReadDataPorts_3_valid_0;
  reg  [3:0]        readStageValid_readCounter_3;
  wire [3:0]        readStageValid_counterChange_3 = _readStageValid_T_68 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_3_valid_0 = readStageValid_stageValid_3 & ~(readStageValid_readCounter_3[3]);
  wire [4:0]        vrfReadDataPorts_3_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_3} * _GEN_5 + {2'h0, readStageValid_readCount_3};
  reg  [2:0]        readStageValid_segPtr_4;
  reg  [2:0]        readStageValid_readCount_4;
  reg               readStageValid_stageValid_4;
  wire              readStageValid_lastReadPtr_4 = readStageValid_segPtr_4 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_4 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_4 + 3'h1;
  wire              readStageValid_lastReadGroup_4 = {4'h0, readStageValid_readCount_4} == lastDataGroupReg;
  wire              vrfReadDataPorts_4_valid_0;
  wire              _readStageValid_T_87 = vrfReadDataPorts_4_ready_0 & vrfReadDataPorts_4_valid_0;
  reg  [3:0]        readStageValid_readCounter_4;
  wire [3:0]        readStageValid_counterChange_4 = _readStageValid_T_87 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_4_valid_0 = readStageValid_stageValid_4 & ~(readStageValid_readCounter_4[3]);
  wire [4:0]        vrfReadDataPorts_4_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_4} * _GEN_5 + {2'h0, readStageValid_readCount_4};
  reg  [2:0]        readStageValid_segPtr_5;
  reg  [2:0]        readStageValid_readCount_5;
  reg               readStageValid_stageValid_5;
  wire              readStageValid_lastReadPtr_5 = readStageValid_segPtr_5 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_5 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_5 + 3'h1;
  wire              readStageValid_lastReadGroup_5 = {4'h0, readStageValid_readCount_5} == lastDataGroupReg;
  wire              vrfReadDataPorts_5_valid_0;
  wire              _readStageValid_T_106 = vrfReadDataPorts_5_ready_0 & vrfReadDataPorts_5_valid_0;
  reg  [3:0]        readStageValid_readCounter_5;
  wire [3:0]        readStageValid_counterChange_5 = _readStageValid_T_106 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_5_valid_0 = readStageValid_stageValid_5 & ~(readStageValid_readCounter_5[3]);
  wire [4:0]        vrfReadDataPorts_5_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_5} * _GEN_5 + {2'h0, readStageValid_readCount_5};
  reg  [2:0]        readStageValid_segPtr_6;
  reg  [2:0]        readStageValid_readCount_6;
  reg               readStageValid_stageValid_6;
  wire              readStageValid_lastReadPtr_6 = readStageValid_segPtr_6 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_6 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_6 + 3'h1;
  wire              readStageValid_lastReadGroup_6 = {4'h0, readStageValid_readCount_6} == lastDataGroupReg;
  wire              vrfReadDataPorts_6_valid_0;
  wire              _readStageValid_T_125 = vrfReadDataPorts_6_ready_0 & vrfReadDataPorts_6_valid_0;
  reg  [3:0]        readStageValid_readCounter_6;
  wire [3:0]        readStageValid_counterChange_6 = _readStageValid_T_125 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_6_valid_0 = readStageValid_stageValid_6 & ~(readStageValid_readCounter_6[3]);
  wire [4:0]        vrfReadDataPorts_6_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_6} * _GEN_5 + {2'h0, readStageValid_readCount_6};
  reg  [2:0]        readStageValid_segPtr_7;
  reg  [2:0]        readStageValid_readCount_7;
  reg               readStageValid_stageValid_7;
  wire              readStageValid_lastReadPtr_7 = readStageValid_segPtr_7 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_7 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_7 + 3'h1;
  wire              readStageValid_lastReadGroup_7 = {4'h0, readStageValid_readCount_7} == lastDataGroupReg;
  wire              vrfReadDataPorts_7_valid_0;
  wire              _readStageValid_T_144 = vrfReadDataPorts_7_ready_0 & vrfReadDataPorts_7_valid_0;
  reg  [3:0]        readStageValid_readCounter_7;
  wire [3:0]        readStageValid_counterChange_7 = _readStageValid_T_144 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_7_valid_0 = readStageValid_stageValid_7 & ~(readStageValid_readCounter_7[3]);
  wire [4:0]        vrfReadDataPorts_7_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_7} * _GEN_5 + {2'h0, readStageValid_readCount_7};
  reg  [2:0]        readStageValid_segPtr_8;
  reg  [2:0]        readStageValid_readCount_8;
  reg               readStageValid_stageValid_8;
  wire              readStageValid_lastReadPtr_8 = readStageValid_segPtr_8 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_8 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_8 + 3'h1;
  wire              readStageValid_lastReadGroup_8 = {4'h0, readStageValid_readCount_8} == lastDataGroupReg;
  wire              vrfReadDataPorts_8_valid_0;
  wire              _readStageValid_T_163 = vrfReadDataPorts_8_ready_0 & vrfReadDataPorts_8_valid_0;
  reg  [3:0]        readStageValid_readCounter_8;
  wire [3:0]        readStageValid_counterChange_8 = _readStageValid_T_163 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_8_valid_0 = readStageValid_stageValid_8 & ~(readStageValid_readCounter_8[3]);
  wire [4:0]        vrfReadDataPorts_8_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_8} * _GEN_5 + {2'h0, readStageValid_readCount_8};
  reg  [2:0]        readStageValid_segPtr_9;
  reg  [2:0]        readStageValid_readCount_9;
  reg               readStageValid_stageValid_9;
  wire              readStageValid_lastReadPtr_9 = readStageValid_segPtr_9 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_9 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_9 + 3'h1;
  wire              readStageValid_lastReadGroup_9 = {4'h0, readStageValid_readCount_9} == lastDataGroupReg;
  wire              vrfReadDataPorts_9_valid_0;
  wire              _readStageValid_T_182 = vrfReadDataPorts_9_ready_0 & vrfReadDataPorts_9_valid_0;
  reg  [3:0]        readStageValid_readCounter_9;
  wire [3:0]        readStageValid_counterChange_9 = _readStageValid_T_182 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_9_valid_0 = readStageValid_stageValid_9 & ~(readStageValid_readCounter_9[3]);
  wire [4:0]        vrfReadDataPorts_9_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_9} * _GEN_5 + {2'h0, readStageValid_readCount_9};
  reg  [2:0]        readStageValid_segPtr_10;
  reg  [2:0]        readStageValid_readCount_10;
  reg               readStageValid_stageValid_10;
  wire              readStageValid_lastReadPtr_10 = readStageValid_segPtr_10 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_10 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_10 + 3'h1;
  wire              readStageValid_lastReadGroup_10 = {4'h0, readStageValid_readCount_10} == lastDataGroupReg;
  wire              vrfReadDataPorts_10_valid_0;
  wire              _readStageValid_T_201 = vrfReadDataPorts_10_ready_0 & vrfReadDataPorts_10_valid_0;
  reg  [3:0]        readStageValid_readCounter_10;
  wire [3:0]        readStageValid_counterChange_10 = _readStageValid_T_201 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_10_valid_0 = readStageValid_stageValid_10 & ~(readStageValid_readCounter_10[3]);
  wire [4:0]        vrfReadDataPorts_10_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_10} * _GEN_5 + {2'h0, readStageValid_readCount_10};
  reg  [2:0]        readStageValid_segPtr_11;
  reg  [2:0]        readStageValid_readCount_11;
  reg               readStageValid_stageValid_11;
  wire              readStageValid_lastReadPtr_11 = readStageValid_segPtr_11 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_11 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_11 + 3'h1;
  wire              readStageValid_lastReadGroup_11 = {4'h0, readStageValid_readCount_11} == lastDataGroupReg;
  wire              vrfReadDataPorts_11_valid_0;
  wire              _readStageValid_T_220 = vrfReadDataPorts_11_ready_0 & vrfReadDataPorts_11_valid_0;
  reg  [3:0]        readStageValid_readCounter_11;
  wire [3:0]        readStageValid_counterChange_11 = _readStageValid_T_220 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_11_valid_0 = readStageValid_stageValid_11 & ~(readStageValid_readCounter_11[3]);
  wire [4:0]        vrfReadDataPorts_11_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_11} * _GEN_5 + {2'h0, readStageValid_readCount_11};
  reg  [2:0]        readStageValid_segPtr_12;
  reg  [2:0]        readStageValid_readCount_12;
  reg               readStageValid_stageValid_12;
  wire              readStageValid_lastReadPtr_12 = readStageValid_segPtr_12 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_12 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_12 + 3'h1;
  wire              readStageValid_lastReadGroup_12 = {4'h0, readStageValid_readCount_12} == lastDataGroupReg;
  wire              vrfReadDataPorts_12_valid_0;
  wire              _readStageValid_T_239 = vrfReadDataPorts_12_ready_0 & vrfReadDataPorts_12_valid_0;
  reg  [3:0]        readStageValid_readCounter_12;
  wire [3:0]        readStageValid_counterChange_12 = _readStageValid_T_239 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_12_valid_0 = readStageValid_stageValid_12 & ~(readStageValid_readCounter_12[3]);
  wire [4:0]        vrfReadDataPorts_12_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_12} * _GEN_5 + {2'h0, readStageValid_readCount_12};
  reg  [2:0]        readStageValid_segPtr_13;
  reg  [2:0]        readStageValid_readCount_13;
  reg               readStageValid_stageValid_13;
  wire              readStageValid_lastReadPtr_13 = readStageValid_segPtr_13 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_13 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_13 + 3'h1;
  wire              readStageValid_lastReadGroup_13 = {4'h0, readStageValid_readCount_13} == lastDataGroupReg;
  wire              vrfReadDataPorts_13_valid_0;
  wire              _readStageValid_T_258 = vrfReadDataPorts_13_ready_0 & vrfReadDataPorts_13_valid_0;
  reg  [3:0]        readStageValid_readCounter_13;
  wire [3:0]        readStageValid_counterChange_13 = _readStageValid_T_258 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_13_valid_0 = readStageValid_stageValid_13 & ~(readStageValid_readCounter_13[3]);
  wire [4:0]        vrfReadDataPorts_13_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_13} * _GEN_5 + {2'h0, readStageValid_readCount_13};
  reg  [2:0]        readStageValid_segPtr_14;
  reg  [2:0]        readStageValid_readCount_14;
  reg               readStageValid_stageValid_14;
  wire              readStageValid_lastReadPtr_14 = readStageValid_segPtr_14 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_14 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_14 + 3'h1;
  wire              readStageValid_lastReadGroup_14 = {4'h0, readStageValid_readCount_14} == lastDataGroupReg;
  wire              vrfReadDataPorts_14_valid_0;
  wire              _readStageValid_T_277 = vrfReadDataPorts_14_ready_0 & vrfReadDataPorts_14_valid_0;
  reg  [3:0]        readStageValid_readCounter_14;
  wire [3:0]        readStageValid_counterChange_14 = _readStageValid_T_277 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_14_valid_0 = readStageValid_stageValid_14 & ~(readStageValid_readCounter_14[3]);
  wire [4:0]        vrfReadDataPorts_14_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_14} * _GEN_5 + {2'h0, readStageValid_readCount_14};
  reg  [2:0]        readStageValid_segPtr_15;
  reg  [2:0]        readStageValid_readCount_15;
  reg               readStageValid_stageValid_15;
  wire              readStageValid_lastReadPtr_15 = readStageValid_segPtr_15 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_15 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_15 + 3'h1;
  wire              readStageValid_lastReadGroup_15 = {4'h0, readStageValid_readCount_15} == lastDataGroupReg;
  wire              vrfReadDataPorts_15_valid_0;
  wire              _readStageValid_T_296 = vrfReadDataPorts_15_ready_0 & vrfReadDataPorts_15_valid_0;
  reg  [3:0]        readStageValid_readCounter_15;
  wire [3:0]        readStageValid_counterChange_15 = _readStageValid_T_296 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_15_valid_0 = readStageValid_stageValid_15 & ~(readStageValid_readCounter_15[3]);
  wire [4:0]        vrfReadDataPorts_15_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_15} * _GEN_5 + {2'h0, readStageValid_readCount_15};
  reg  [2:0]        readStageValid_segPtr_16;
  reg  [2:0]        readStageValid_readCount_16;
  reg               readStageValid_stageValid_16;
  wire              readStageValid_lastReadPtr_16 = readStageValid_segPtr_16 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_16 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_16 + 3'h1;
  wire              readStageValid_lastReadGroup_16 = {4'h0, readStageValid_readCount_16} == lastDataGroupReg;
  wire              vrfReadDataPorts_16_valid_0;
  wire              _readStageValid_T_315 = vrfReadDataPorts_16_ready_0 & vrfReadDataPorts_16_valid_0;
  reg  [3:0]        readStageValid_readCounter_16;
  wire [3:0]        readStageValid_counterChange_16 = _readStageValid_T_315 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_16_valid_0 = readStageValid_stageValid_16 & ~(readStageValid_readCounter_16[3]);
  wire [4:0]        vrfReadDataPorts_16_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_16} * _GEN_5 + {2'h0, readStageValid_readCount_16};
  reg  [2:0]        readStageValid_segPtr_17;
  reg  [2:0]        readStageValid_readCount_17;
  reg               readStageValid_stageValid_17;
  wire              readStageValid_lastReadPtr_17 = readStageValid_segPtr_17 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_17 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_17 + 3'h1;
  wire              readStageValid_lastReadGroup_17 = {4'h0, readStageValid_readCount_17} == lastDataGroupReg;
  wire              vrfReadDataPorts_17_valid_0;
  wire              _readStageValid_T_334 = vrfReadDataPorts_17_ready_0 & vrfReadDataPorts_17_valid_0;
  reg  [3:0]        readStageValid_readCounter_17;
  wire [3:0]        readStageValid_counterChange_17 = _readStageValid_T_334 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_17_valid_0 = readStageValid_stageValid_17 & ~(readStageValid_readCounter_17[3]);
  wire [4:0]        vrfReadDataPorts_17_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_17} * _GEN_5 + {2'h0, readStageValid_readCount_17};
  reg  [2:0]        readStageValid_segPtr_18;
  reg  [2:0]        readStageValid_readCount_18;
  reg               readStageValid_stageValid_18;
  wire              readStageValid_lastReadPtr_18 = readStageValid_segPtr_18 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_18 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_18 + 3'h1;
  wire              readStageValid_lastReadGroup_18 = {4'h0, readStageValid_readCount_18} == lastDataGroupReg;
  wire              vrfReadDataPorts_18_valid_0;
  wire              _readStageValid_T_353 = vrfReadDataPorts_18_ready_0 & vrfReadDataPorts_18_valid_0;
  reg  [3:0]        readStageValid_readCounter_18;
  wire [3:0]        readStageValid_counterChange_18 = _readStageValid_T_353 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_18_valid_0 = readStageValid_stageValid_18 & ~(readStageValid_readCounter_18[3]);
  wire [4:0]        vrfReadDataPorts_18_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_18} * _GEN_5 + {2'h0, readStageValid_readCount_18};
  reg  [2:0]        readStageValid_segPtr_19;
  reg  [2:0]        readStageValid_readCount_19;
  reg               readStageValid_stageValid_19;
  wire              readStageValid_lastReadPtr_19 = readStageValid_segPtr_19 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_19 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_19 + 3'h1;
  wire              readStageValid_lastReadGroup_19 = {4'h0, readStageValid_readCount_19} == lastDataGroupReg;
  wire              vrfReadDataPorts_19_valid_0;
  wire              _readStageValid_T_372 = vrfReadDataPorts_19_ready_0 & vrfReadDataPorts_19_valid_0;
  reg  [3:0]        readStageValid_readCounter_19;
  wire [3:0]        readStageValid_counterChange_19 = _readStageValid_T_372 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_19_valid_0 = readStageValid_stageValid_19 & ~(readStageValid_readCounter_19[3]);
  wire [4:0]        vrfReadDataPorts_19_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_19} * _GEN_5 + {2'h0, readStageValid_readCount_19};
  reg  [2:0]        readStageValid_segPtr_20;
  reg  [2:0]        readStageValid_readCount_20;
  reg               readStageValid_stageValid_20;
  wire              readStageValid_lastReadPtr_20 = readStageValid_segPtr_20 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_20 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_20 + 3'h1;
  wire              readStageValid_lastReadGroup_20 = {4'h0, readStageValid_readCount_20} == lastDataGroupReg;
  wire              vrfReadDataPorts_20_valid_0;
  wire              _readStageValid_T_391 = vrfReadDataPorts_20_ready_0 & vrfReadDataPorts_20_valid_0;
  reg  [3:0]        readStageValid_readCounter_20;
  wire [3:0]        readStageValid_counterChange_20 = _readStageValid_T_391 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_20_valid_0 = readStageValid_stageValid_20 & ~(readStageValid_readCounter_20[3]);
  wire [4:0]        vrfReadDataPorts_20_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_20} * _GEN_5 + {2'h0, readStageValid_readCount_20};
  reg  [2:0]        readStageValid_segPtr_21;
  reg  [2:0]        readStageValid_readCount_21;
  reg               readStageValid_stageValid_21;
  wire              readStageValid_lastReadPtr_21 = readStageValid_segPtr_21 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_21 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_21 + 3'h1;
  wire              readStageValid_lastReadGroup_21 = {4'h0, readStageValid_readCount_21} == lastDataGroupReg;
  wire              vrfReadDataPorts_21_valid_0;
  wire              _readStageValid_T_410 = vrfReadDataPorts_21_ready_0 & vrfReadDataPorts_21_valid_0;
  reg  [3:0]        readStageValid_readCounter_21;
  wire [3:0]        readStageValid_counterChange_21 = _readStageValid_T_410 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_21_valid_0 = readStageValid_stageValid_21 & ~(readStageValid_readCounter_21[3]);
  wire [4:0]        vrfReadDataPorts_21_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_21} * _GEN_5 + {2'h0, readStageValid_readCount_21};
  reg  [2:0]        readStageValid_segPtr_22;
  reg  [2:0]        readStageValid_readCount_22;
  reg               readStageValid_stageValid_22;
  wire              readStageValid_lastReadPtr_22 = readStageValid_segPtr_22 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_22 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_22 + 3'h1;
  wire              readStageValid_lastReadGroup_22 = {4'h0, readStageValid_readCount_22} == lastDataGroupReg;
  wire              vrfReadDataPorts_22_valid_0;
  wire              _readStageValid_T_429 = vrfReadDataPorts_22_ready_0 & vrfReadDataPorts_22_valid_0;
  reg  [3:0]        readStageValid_readCounter_22;
  wire [3:0]        readStageValid_counterChange_22 = _readStageValid_T_429 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_22_valid_0 = readStageValid_stageValid_22 & ~(readStageValid_readCounter_22[3]);
  wire [4:0]        vrfReadDataPorts_22_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_22} * _GEN_5 + {2'h0, readStageValid_readCount_22};
  reg  [2:0]        readStageValid_segPtr_23;
  reg  [2:0]        readStageValid_readCount_23;
  reg               readStageValid_stageValid_23;
  wire              readStageValid_lastReadPtr_23 = readStageValid_segPtr_23 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_23 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_23 + 3'h1;
  wire              readStageValid_lastReadGroup_23 = {4'h0, readStageValid_readCount_23} == lastDataGroupReg;
  wire              vrfReadDataPorts_23_valid_0;
  wire              _readStageValid_T_448 = vrfReadDataPorts_23_ready_0 & vrfReadDataPorts_23_valid_0;
  reg  [3:0]        readStageValid_readCounter_23;
  wire [3:0]        readStageValid_counterChange_23 = _readStageValid_T_448 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_23_valid_0 = readStageValid_stageValid_23 & ~(readStageValid_readCounter_23[3]);
  wire [4:0]        vrfReadDataPorts_23_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_23} * _GEN_5 + {2'h0, readStageValid_readCount_23};
  reg  [2:0]        readStageValid_segPtr_24;
  reg  [2:0]        readStageValid_readCount_24;
  reg               readStageValid_stageValid_24;
  wire              readStageValid_lastReadPtr_24 = readStageValid_segPtr_24 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_24 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_24 + 3'h1;
  wire              readStageValid_lastReadGroup_24 = {4'h0, readStageValid_readCount_24} == lastDataGroupReg;
  wire              vrfReadDataPorts_24_valid_0;
  wire              _readStageValid_T_467 = vrfReadDataPorts_24_ready_0 & vrfReadDataPorts_24_valid_0;
  reg  [3:0]        readStageValid_readCounter_24;
  wire [3:0]        readStageValid_counterChange_24 = _readStageValid_T_467 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_24_valid_0 = readStageValid_stageValid_24 & ~(readStageValid_readCounter_24[3]);
  wire [4:0]        vrfReadDataPorts_24_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_24} * _GEN_5 + {2'h0, readStageValid_readCount_24};
  reg  [2:0]        readStageValid_segPtr_25;
  reg  [2:0]        readStageValid_readCount_25;
  reg               readStageValid_stageValid_25;
  wire              readStageValid_lastReadPtr_25 = readStageValid_segPtr_25 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_25 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_25 + 3'h1;
  wire              readStageValid_lastReadGroup_25 = {4'h0, readStageValid_readCount_25} == lastDataGroupReg;
  wire              vrfReadDataPorts_25_valid_0;
  wire              _readStageValid_T_486 = vrfReadDataPorts_25_ready_0 & vrfReadDataPorts_25_valid_0;
  reg  [3:0]        readStageValid_readCounter_25;
  wire [3:0]        readStageValid_counterChange_25 = _readStageValid_T_486 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_25_valid_0 = readStageValid_stageValid_25 & ~(readStageValid_readCounter_25[3]);
  wire [4:0]        vrfReadDataPorts_25_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_25} * _GEN_5 + {2'h0, readStageValid_readCount_25};
  reg  [2:0]        readStageValid_segPtr_26;
  reg  [2:0]        readStageValid_readCount_26;
  reg               readStageValid_stageValid_26;
  wire              readStageValid_lastReadPtr_26 = readStageValid_segPtr_26 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_26 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_26 + 3'h1;
  wire              readStageValid_lastReadGroup_26 = {4'h0, readStageValid_readCount_26} == lastDataGroupReg;
  wire              vrfReadDataPorts_26_valid_0;
  wire              _readStageValid_T_505 = vrfReadDataPorts_26_ready_0 & vrfReadDataPorts_26_valid_0;
  reg  [3:0]        readStageValid_readCounter_26;
  wire [3:0]        readStageValid_counterChange_26 = _readStageValid_T_505 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_26_valid_0 = readStageValid_stageValid_26 & ~(readStageValid_readCounter_26[3]);
  wire [4:0]        vrfReadDataPorts_26_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_26} * _GEN_5 + {2'h0, readStageValid_readCount_26};
  reg  [2:0]        readStageValid_segPtr_27;
  reg  [2:0]        readStageValid_readCount_27;
  reg               readStageValid_stageValid_27;
  wire              readStageValid_lastReadPtr_27 = readStageValid_segPtr_27 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_27 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_27 + 3'h1;
  wire              readStageValid_lastReadGroup_27 = {4'h0, readStageValid_readCount_27} == lastDataGroupReg;
  wire              vrfReadDataPorts_27_valid_0;
  wire              _readStageValid_T_524 = vrfReadDataPorts_27_ready_0 & vrfReadDataPorts_27_valid_0;
  reg  [3:0]        readStageValid_readCounter_27;
  wire [3:0]        readStageValid_counterChange_27 = _readStageValid_T_524 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_27_valid_0 = readStageValid_stageValid_27 & ~(readStageValid_readCounter_27[3]);
  wire [4:0]        vrfReadDataPorts_27_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_27} * _GEN_5 + {2'h0, readStageValid_readCount_27};
  reg  [2:0]        readStageValid_segPtr_28;
  reg  [2:0]        readStageValid_readCount_28;
  reg               readStageValid_stageValid_28;
  wire              readStageValid_lastReadPtr_28 = readStageValid_segPtr_28 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_28 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_28 + 3'h1;
  wire              readStageValid_lastReadGroup_28 = {4'h0, readStageValid_readCount_28} == lastDataGroupReg;
  wire              vrfReadDataPorts_28_valid_0;
  wire              _readStageValid_T_543 = vrfReadDataPorts_28_ready_0 & vrfReadDataPorts_28_valid_0;
  reg  [3:0]        readStageValid_readCounter_28;
  wire [3:0]        readStageValid_counterChange_28 = _readStageValid_T_543 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_28_valid_0 = readStageValid_stageValid_28 & ~(readStageValid_readCounter_28[3]);
  wire [4:0]        vrfReadDataPorts_28_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_28} * _GEN_5 + {2'h0, readStageValid_readCount_28};
  reg  [2:0]        readStageValid_segPtr_29;
  reg  [2:0]        readStageValid_readCount_29;
  reg               readStageValid_stageValid_29;
  wire              readStageValid_lastReadPtr_29 = readStageValid_segPtr_29 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_29 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_29 + 3'h1;
  wire              readStageValid_lastReadGroup_29 = {4'h0, readStageValid_readCount_29} == lastDataGroupReg;
  wire              vrfReadDataPorts_29_valid_0;
  wire              _readStageValid_T_562 = vrfReadDataPorts_29_ready_0 & vrfReadDataPorts_29_valid_0;
  reg  [3:0]        readStageValid_readCounter_29;
  wire [3:0]        readStageValid_counterChange_29 = _readStageValid_T_562 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_29_valid_0 = readStageValid_stageValid_29 & ~(readStageValid_readCounter_29[3]);
  wire [4:0]        vrfReadDataPorts_29_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_29} * _GEN_5 + {2'h0, readStageValid_readCount_29};
  reg  [2:0]        readStageValid_segPtr_30;
  reg  [2:0]        readStageValid_readCount_30;
  reg               readStageValid_stageValid_30;
  wire              readStageValid_lastReadPtr_30 = readStageValid_segPtr_30 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_30 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_30 + 3'h1;
  wire              readStageValid_lastReadGroup_30 = {4'h0, readStageValid_readCount_30} == lastDataGroupReg;
  wire              vrfReadDataPorts_30_valid_0;
  wire              _readStageValid_T_581 = vrfReadDataPorts_30_ready_0 & vrfReadDataPorts_30_valid_0;
  reg  [3:0]        readStageValid_readCounter_30;
  wire [3:0]        readStageValid_counterChange_30 = _readStageValid_T_581 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_30_valid_0 = readStageValid_stageValid_30 & ~(readStageValid_readCounter_30[3]);
  wire [4:0]        vrfReadDataPorts_30_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_30} * _GEN_5 + {2'h0, readStageValid_readCount_30};
  reg  [2:0]        readStageValid_segPtr_31;
  reg  [2:0]        readStageValid_readCount_31;
  reg               readStageValid_stageValid_31;
  wire              readStageValid_lastReadPtr_31 = readStageValid_segPtr_31 == 3'h0;
  wire [2:0]        readStageValid_nextReadCount_31 = lsuRequest_valid ? 3'h0 : readStageValid_readCount_31 + 3'h1;
  wire              readStageValid_lastReadGroup_31 = {4'h0, readStageValid_readCount_31} == lastDataGroupReg;
  wire              vrfReadDataPorts_31_valid_0;
  wire              _readStageValid_T_600 = vrfReadDataPorts_31_ready_0 & vrfReadDataPorts_31_valid_0;
  reg  [3:0]        readStageValid_readCounter_31;
  wire [3:0]        readStageValid_counterChange_31 = _readStageValid_T_600 ? 4'h1 : 4'hF;
  assign vrfReadDataPorts_31_valid_0 = readStageValid_stageValid_31 & ~(readStageValid_readCounter_31[3]);
  wire [4:0]        vrfReadDataPorts_31_bits_vs_0 = lsuRequestReg_instructionInformation_vs3 + {2'h0, readStageValid_segPtr_31} * _GEN_5 + {2'h0, readStageValid_readCount_31};
  wire              readStageValid =
    |{readStageValid_stageValid,
      readStageValid_readCounter,
      readStageValid_stageValid_1,
      readStageValid_readCounter_1,
      readStageValid_stageValid_2,
      readStageValid_readCounter_2,
      readStageValid_stageValid_3,
      readStageValid_readCounter_3,
      readStageValid_stageValid_4,
      readStageValid_readCounter_4,
      readStageValid_stageValid_5,
      readStageValid_readCounter_5,
      readStageValid_stageValid_6,
      readStageValid_readCounter_6,
      readStageValid_stageValid_7,
      readStageValid_readCounter_7,
      readStageValid_stageValid_8,
      readStageValid_readCounter_8,
      readStageValid_stageValid_9,
      readStageValid_readCounter_9,
      readStageValid_stageValid_10,
      readStageValid_readCounter_10,
      readStageValid_stageValid_11,
      readStageValid_readCounter_11,
      readStageValid_stageValid_12,
      readStageValid_readCounter_12,
      readStageValid_stageValid_13,
      readStageValid_readCounter_13,
      readStageValid_stageValid_14,
      readStageValid_readCounter_14,
      readStageValid_stageValid_15,
      readStageValid_readCounter_15,
      readStageValid_stageValid_16,
      readStageValid_readCounter_16,
      readStageValid_stageValid_17,
      readStageValid_readCounter_17,
      readStageValid_stageValid_18,
      readStageValid_readCounter_18,
      readStageValid_stageValid_19,
      readStageValid_readCounter_19,
      readStageValid_stageValid_20,
      readStageValid_readCounter_20,
      readStageValid_stageValid_21,
      readStageValid_readCounter_21,
      readStageValid_stageValid_22,
      readStageValid_readCounter_22,
      readStageValid_stageValid_23,
      readStageValid_readCounter_23,
      readStageValid_stageValid_24,
      readStageValid_readCounter_24,
      readStageValid_stageValid_25,
      readStageValid_readCounter_25,
      readStageValid_stageValid_26,
      readStageValid_readCounter_26,
      readStageValid_stageValid_27,
      readStageValid_readCounter_27,
      readStageValid_stageValid_28,
      readStageValid_readCounter_28,
      readStageValid_stageValid_29,
      readStageValid_readCounter_29,
      readStageValid_stageValid_30,
      readStageValid_readCounter_30,
      readStageValid_stageValid_31,
      readStageValid_readCounter_31};
  reg               bufferFull;
  wire              accessBufferDequeueReady;
  wire              accessBufferEnqueueReady = ~bufferFull | accessBufferDequeueReady;
  wire              accessBufferEnqueueValid =
    vrfReadQueueVec_0_deq_valid & vrfReadQueueVec_1_deq_valid & vrfReadQueueVec_2_deq_valid & vrfReadQueueVec_3_deq_valid & vrfReadQueueVec_4_deq_valid & vrfReadQueueVec_5_deq_valid & vrfReadQueueVec_6_deq_valid
    & vrfReadQueueVec_7_deq_valid & vrfReadQueueVec_8_deq_valid & vrfReadQueueVec_9_deq_valid & vrfReadQueueVec_10_deq_valid & vrfReadQueueVec_11_deq_valid & vrfReadQueueVec_12_deq_valid & vrfReadQueueVec_13_deq_valid
    & vrfReadQueueVec_14_deq_valid & vrfReadQueueVec_15_deq_valid & vrfReadQueueVec_16_deq_valid & vrfReadQueueVec_17_deq_valid & vrfReadQueueVec_18_deq_valid & vrfReadQueueVec_19_deq_valid & vrfReadQueueVec_20_deq_valid
    & vrfReadQueueVec_21_deq_valid & vrfReadQueueVec_22_deq_valid & vrfReadQueueVec_23_deq_valid & vrfReadQueueVec_24_deq_valid & vrfReadQueueVec_25_deq_valid & vrfReadQueueVec_26_deq_valid & vrfReadQueueVec_27_deq_valid
    & vrfReadQueueVec_28_deq_valid & vrfReadQueueVec_29_deq_valid & vrfReadQueueVec_30_deq_valid & vrfReadQueueVec_31_deq_valid;
  wire              readQueueClear =
    ~(vrfReadQueueVec_0_deq_valid | vrfReadQueueVec_1_deq_valid | vrfReadQueueVec_2_deq_valid | vrfReadQueueVec_3_deq_valid | vrfReadQueueVec_4_deq_valid | vrfReadQueueVec_5_deq_valid | vrfReadQueueVec_6_deq_valid
      | vrfReadQueueVec_7_deq_valid | vrfReadQueueVec_8_deq_valid | vrfReadQueueVec_9_deq_valid | vrfReadQueueVec_10_deq_valid | vrfReadQueueVec_11_deq_valid | vrfReadQueueVec_12_deq_valid | vrfReadQueueVec_13_deq_valid
      | vrfReadQueueVec_14_deq_valid | vrfReadQueueVec_15_deq_valid | vrfReadQueueVec_16_deq_valid | vrfReadQueueVec_17_deq_valid | vrfReadQueueVec_18_deq_valid | vrfReadQueueVec_19_deq_valid | vrfReadQueueVec_20_deq_valid
      | vrfReadQueueVec_21_deq_valid | vrfReadQueueVec_22_deq_valid | vrfReadQueueVec_23_deq_valid | vrfReadQueueVec_24_deq_valid | vrfReadQueueVec_25_deq_valid | vrfReadQueueVec_26_deq_valid | vrfReadQueueVec_27_deq_valid
      | vrfReadQueueVec_28_deq_valid | vrfReadQueueVec_29_deq_valid | vrfReadQueueVec_30_deq_valid | vrfReadQueueVec_31_deq_valid);
  assign accessBufferEnqueueFire = accessBufferEnqueueValid & accessBufferEnqueueReady;
  assign vrfReadQueueVec_0_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_1_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_2_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_3_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_4_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_5_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_6_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_7_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_8_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_9_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_10_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_11_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_12_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_13_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_14_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_15_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_16_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_17_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_18_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_19_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_20_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_21_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_22_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_23_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_24_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_25_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_26_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_27_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_28_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_29_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_30_deq_ready = accessBufferEnqueueFire;
  assign vrfReadQueueVec_31_deq_ready = accessBufferEnqueueFire;
  wire              lastPtr = accessPtr == 3'h0;
  wire              lastPtrEnq = lastPtr & accessBufferEnqueueFire;
  wire              accessBufferDequeueValid = bufferFull | lastPtrEnq;
  wire              accessBufferDequeueFire = accessBufferDequeueValid & accessBufferDequeueReady;
  wire [63:0]       accessDataUpdate_lo_lo_lo_lo = {vrfReadQueueVec_1_deq_bits, vrfReadQueueVec_0_deq_bits};
  wire [63:0]       accessDataUpdate_lo_lo_lo_hi = {vrfReadQueueVec_3_deq_bits, vrfReadQueueVec_2_deq_bits};
  wire [127:0]      accessDataUpdate_lo_lo_lo = {accessDataUpdate_lo_lo_lo_hi, accessDataUpdate_lo_lo_lo_lo};
  wire [63:0]       accessDataUpdate_lo_lo_hi_lo = {vrfReadQueueVec_5_deq_bits, vrfReadQueueVec_4_deq_bits};
  wire [63:0]       accessDataUpdate_lo_lo_hi_hi = {vrfReadQueueVec_7_deq_bits, vrfReadQueueVec_6_deq_bits};
  wire [127:0]      accessDataUpdate_lo_lo_hi = {accessDataUpdate_lo_lo_hi_hi, accessDataUpdate_lo_lo_hi_lo};
  wire [255:0]      accessDataUpdate_lo_lo = {accessDataUpdate_lo_lo_hi, accessDataUpdate_lo_lo_lo};
  wire [63:0]       accessDataUpdate_lo_hi_lo_lo = {vrfReadQueueVec_9_deq_bits, vrfReadQueueVec_8_deq_bits};
  wire [63:0]       accessDataUpdate_lo_hi_lo_hi = {vrfReadQueueVec_11_deq_bits, vrfReadQueueVec_10_deq_bits};
  wire [127:0]      accessDataUpdate_lo_hi_lo = {accessDataUpdate_lo_hi_lo_hi, accessDataUpdate_lo_hi_lo_lo};
  wire [63:0]       accessDataUpdate_lo_hi_hi_lo = {vrfReadQueueVec_13_deq_bits, vrfReadQueueVec_12_deq_bits};
  wire [63:0]       accessDataUpdate_lo_hi_hi_hi = {vrfReadQueueVec_15_deq_bits, vrfReadQueueVec_14_deq_bits};
  wire [127:0]      accessDataUpdate_lo_hi_hi = {accessDataUpdate_lo_hi_hi_hi, accessDataUpdate_lo_hi_hi_lo};
  wire [255:0]      accessDataUpdate_lo_hi = {accessDataUpdate_lo_hi_hi, accessDataUpdate_lo_hi_lo};
  wire [511:0]      accessDataUpdate_lo = {accessDataUpdate_lo_hi, accessDataUpdate_lo_lo};
  wire [63:0]       accessDataUpdate_hi_lo_lo_lo = {vrfReadQueueVec_17_deq_bits, vrfReadQueueVec_16_deq_bits};
  wire [63:0]       accessDataUpdate_hi_lo_lo_hi = {vrfReadQueueVec_19_deq_bits, vrfReadQueueVec_18_deq_bits};
  wire [127:0]      accessDataUpdate_hi_lo_lo = {accessDataUpdate_hi_lo_lo_hi, accessDataUpdate_hi_lo_lo_lo};
  wire [63:0]       accessDataUpdate_hi_lo_hi_lo = {vrfReadQueueVec_21_deq_bits, vrfReadQueueVec_20_deq_bits};
  wire [63:0]       accessDataUpdate_hi_lo_hi_hi = {vrfReadQueueVec_23_deq_bits, vrfReadQueueVec_22_deq_bits};
  wire [127:0]      accessDataUpdate_hi_lo_hi = {accessDataUpdate_hi_lo_hi_hi, accessDataUpdate_hi_lo_hi_lo};
  wire [255:0]      accessDataUpdate_hi_lo = {accessDataUpdate_hi_lo_hi, accessDataUpdate_hi_lo_lo};
  wire [63:0]       accessDataUpdate_hi_hi_lo_lo = {vrfReadQueueVec_25_deq_bits, vrfReadQueueVec_24_deq_bits};
  wire [63:0]       accessDataUpdate_hi_hi_lo_hi = {vrfReadQueueVec_27_deq_bits, vrfReadQueueVec_26_deq_bits};
  wire [127:0]      accessDataUpdate_hi_hi_lo = {accessDataUpdate_hi_hi_lo_hi, accessDataUpdate_hi_hi_lo_lo};
  wire [63:0]       accessDataUpdate_hi_hi_hi_lo = {vrfReadQueueVec_29_deq_bits, vrfReadQueueVec_28_deq_bits};
  wire [63:0]       accessDataUpdate_hi_hi_hi_hi = {vrfReadQueueVec_31_deq_bits, vrfReadQueueVec_30_deq_bits};
  wire [127:0]      accessDataUpdate_hi_hi_hi = {accessDataUpdate_hi_hi_hi_hi, accessDataUpdate_hi_hi_hi_lo};
  wire [255:0]      accessDataUpdate_hi_hi = {accessDataUpdate_hi_hi_hi, accessDataUpdate_hi_hi_lo};
  wire [511:0]      accessDataUpdate_hi = {accessDataUpdate_hi_hi, accessDataUpdate_hi_lo};
  wire [1023:0]     accessDataUpdate_0 = {accessDataUpdate_hi, accessDataUpdate_lo};
  reg               bufferValid;
  reg  [127:0]      maskForBufferData_0;
  reg  [127:0]      maskForBufferData_1;
  reg  [127:0]      maskForBufferData_2;
  reg  [127:0]      maskForBufferData_3;
  reg  [127:0]      maskForBufferData_4;
  reg  [127:0]      maskForBufferData_5;
  reg  [127:0]      maskForBufferData_6;
  reg  [127:0]      maskForBufferData_7;
  reg               lastDataGroupInDataBuffer;
  wire              memRequest_valid_0;
  wire              _addressQueue_enq_valid_T = memRequest_ready_0 & memRequest_valid_0;
  wire              alignedDequeueFire;
  assign alignedDequeueFire = _addressQueue_enq_valid_T;
  wire              addressQueue_enq_valid;
  assign addressQueue_enq_valid = _addressQueue_enq_valid_T;
  reg  [1023:0]     cacheLineTemp;
  reg  [127:0]      maskTemp;
  reg               canSendTail;
  wire              isLastCacheLineInBuffer = cacheLineIndexInBuffer == lsuRequestReg_instructionInformation_nf;
  wire              bufferWillClear = alignedDequeueFire & isLastCacheLineInBuffer;
  wire              addressQueue_enq_ready;
  wire              addressQueueFree;
  assign accessBufferDequeueReady = ~bufferValid | memRequest_ready_0 & isLastCacheLineInBuffer & addressQueueFree;
  wire [1023:0]     bufferStageEnqueueData_0 = bufferFull ? accessData_0 : accessDataUpdate_0;
  wire [1023:0]     bufferStageEnqueueData_1 = bufferFull ? accessData_1 : accessDataUpdate_1;
  wire [1023:0]     bufferStageEnqueueData_2 = bufferFull ? accessData_2 : accessDataUpdate_2;
  wire [1023:0]     bufferStageEnqueueData_3 = bufferFull ? accessData_3 : accessDataUpdate_3;
  wire [1023:0]     bufferStageEnqueueData_4 = bufferFull ? accessData_4 : accessDataUpdate_4;
  wire [1023:0]     bufferStageEnqueueData_5 = bufferFull ? accessData_5 : accessDataUpdate_5;
  wire [1023:0]     bufferStageEnqueueData_6 = bufferFull ? accessData_6 : accessDataUpdate_6;
  wire [1023:0]     bufferStageEnqueueData_7 = bufferFull ? accessData_7 : accessDataUpdate_7;
  wire [7:0]        _fillBySeg_T = 8'h1 << lsuRequestReg_instructionInformation_nf;
  wire [3:0]        fillBySeg_lo_lo_lo_lo_lo = {fillBySeg_lo_lo_lo_lo_lo_hi, fillBySeg_lo_lo_lo_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_lo_lo_lo_hi = {fillBySeg_lo_lo_lo_lo_hi_hi, fillBySeg_lo_lo_lo_lo_hi_lo};
  wire [7:0]        fillBySeg_lo_lo_lo_lo = {fillBySeg_lo_lo_lo_lo_hi, fillBySeg_lo_lo_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_lo_lo_hi_lo = {fillBySeg_lo_lo_lo_hi_lo_hi, fillBySeg_lo_lo_lo_hi_lo_lo};
  wire [3:0]        fillBySeg_lo_lo_lo_hi_hi = {fillBySeg_lo_lo_lo_hi_hi_hi, fillBySeg_lo_lo_lo_hi_hi_lo};
  wire [7:0]        fillBySeg_lo_lo_lo_hi = {fillBySeg_lo_lo_lo_hi_hi, fillBySeg_lo_lo_lo_hi_lo};
  wire [15:0]       fillBySeg_lo_lo_lo = {fillBySeg_lo_lo_lo_hi, fillBySeg_lo_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_lo_hi_lo_lo = {fillBySeg_lo_lo_hi_lo_lo_hi, fillBySeg_lo_lo_hi_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_lo_hi_lo_hi = {fillBySeg_lo_lo_hi_lo_hi_hi, fillBySeg_lo_lo_hi_lo_hi_lo};
  wire [7:0]        fillBySeg_lo_lo_hi_lo = {fillBySeg_lo_lo_hi_lo_hi, fillBySeg_lo_lo_hi_lo_lo};
  wire [3:0]        fillBySeg_lo_lo_hi_hi_lo = {fillBySeg_lo_lo_hi_hi_lo_hi, fillBySeg_lo_lo_hi_hi_lo_lo};
  wire [3:0]        fillBySeg_lo_lo_hi_hi_hi = {fillBySeg_lo_lo_hi_hi_hi_hi, fillBySeg_lo_lo_hi_hi_hi_lo};
  wire [7:0]        fillBySeg_lo_lo_hi_hi = {fillBySeg_lo_lo_hi_hi_hi, fillBySeg_lo_lo_hi_hi_lo};
  wire [15:0]       fillBySeg_lo_lo_hi = {fillBySeg_lo_lo_hi_hi, fillBySeg_lo_lo_hi_lo};
  wire [31:0]       fillBySeg_lo_lo = {fillBySeg_lo_lo_hi, fillBySeg_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_lo_lo_lo = {fillBySeg_lo_hi_lo_lo_lo_hi, fillBySeg_lo_hi_lo_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_lo_lo_hi = {fillBySeg_lo_hi_lo_lo_hi_hi, fillBySeg_lo_hi_lo_lo_hi_lo};
  wire [7:0]        fillBySeg_lo_hi_lo_lo = {fillBySeg_lo_hi_lo_lo_hi, fillBySeg_lo_hi_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_lo_hi_lo = {fillBySeg_lo_hi_lo_hi_lo_hi, fillBySeg_lo_hi_lo_hi_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_lo_hi_hi = {fillBySeg_lo_hi_lo_hi_hi_hi, fillBySeg_lo_hi_lo_hi_hi_lo};
  wire [7:0]        fillBySeg_lo_hi_lo_hi = {fillBySeg_lo_hi_lo_hi_hi, fillBySeg_lo_hi_lo_hi_lo};
  wire [15:0]       fillBySeg_lo_hi_lo = {fillBySeg_lo_hi_lo_hi, fillBySeg_lo_hi_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_hi_lo_lo = {fillBySeg_lo_hi_hi_lo_lo_hi, fillBySeg_lo_hi_hi_lo_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_hi_lo_hi = {fillBySeg_lo_hi_hi_lo_hi_hi, fillBySeg_lo_hi_hi_lo_hi_lo};
  wire [7:0]        fillBySeg_lo_hi_hi_lo = {fillBySeg_lo_hi_hi_lo_hi, fillBySeg_lo_hi_hi_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_hi_hi_lo = {fillBySeg_lo_hi_hi_hi_lo_hi, fillBySeg_lo_hi_hi_hi_lo_lo};
  wire [3:0]        fillBySeg_lo_hi_hi_hi_hi = {fillBySeg_lo_hi_hi_hi_hi_hi, fillBySeg_lo_hi_hi_hi_hi_lo};
  wire [7:0]        fillBySeg_lo_hi_hi_hi = {fillBySeg_lo_hi_hi_hi_hi, fillBySeg_lo_hi_hi_hi_lo};
  wire [15:0]       fillBySeg_lo_hi_hi = {fillBySeg_lo_hi_hi_hi, fillBySeg_lo_hi_hi_lo};
  wire [31:0]       fillBySeg_lo_hi = {fillBySeg_lo_hi_hi, fillBySeg_lo_hi_lo};
  wire [63:0]       fillBySeg_lo = {fillBySeg_lo_hi, fillBySeg_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_lo_lo_lo = {fillBySeg_hi_lo_lo_lo_lo_hi, fillBySeg_hi_lo_lo_lo_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_lo_lo_hi = {fillBySeg_hi_lo_lo_lo_hi_hi, fillBySeg_hi_lo_lo_lo_hi_lo};
  wire [7:0]        fillBySeg_hi_lo_lo_lo = {fillBySeg_hi_lo_lo_lo_hi, fillBySeg_hi_lo_lo_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_lo_hi_lo = {fillBySeg_hi_lo_lo_hi_lo_hi, fillBySeg_hi_lo_lo_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_lo_hi_hi = {fillBySeg_hi_lo_lo_hi_hi_hi, fillBySeg_hi_lo_lo_hi_hi_lo};
  wire [7:0]        fillBySeg_hi_lo_lo_hi = {fillBySeg_hi_lo_lo_hi_hi, fillBySeg_hi_lo_lo_hi_lo};
  wire [15:0]       fillBySeg_hi_lo_lo = {fillBySeg_hi_lo_lo_hi, fillBySeg_hi_lo_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_hi_lo_lo = {fillBySeg_hi_lo_hi_lo_lo_hi, fillBySeg_hi_lo_hi_lo_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_hi_lo_hi = {fillBySeg_hi_lo_hi_lo_hi_hi, fillBySeg_hi_lo_hi_lo_hi_lo};
  wire [7:0]        fillBySeg_hi_lo_hi_lo = {fillBySeg_hi_lo_hi_lo_hi, fillBySeg_hi_lo_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_hi_hi_lo = {fillBySeg_hi_lo_hi_hi_lo_hi, fillBySeg_hi_lo_hi_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_lo_hi_hi_hi = {fillBySeg_hi_lo_hi_hi_hi_hi, fillBySeg_hi_lo_hi_hi_hi_lo};
  wire [7:0]        fillBySeg_hi_lo_hi_hi = {fillBySeg_hi_lo_hi_hi_hi, fillBySeg_hi_lo_hi_hi_lo};
  wire [15:0]       fillBySeg_hi_lo_hi = {fillBySeg_hi_lo_hi_hi, fillBySeg_hi_lo_hi_lo};
  wire [31:0]       fillBySeg_hi_lo = {fillBySeg_hi_lo_hi, fillBySeg_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_lo_lo_lo = {fillBySeg_hi_hi_lo_lo_lo_hi, fillBySeg_hi_hi_lo_lo_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_lo_lo_hi = {fillBySeg_hi_hi_lo_lo_hi_hi, fillBySeg_hi_hi_lo_lo_hi_lo};
  wire [7:0]        fillBySeg_hi_hi_lo_lo = {fillBySeg_hi_hi_lo_lo_hi, fillBySeg_hi_hi_lo_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_lo_hi_lo = {fillBySeg_hi_hi_lo_hi_lo_hi, fillBySeg_hi_hi_lo_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_lo_hi_hi = {fillBySeg_hi_hi_lo_hi_hi_hi, fillBySeg_hi_hi_lo_hi_hi_lo};
  wire [7:0]        fillBySeg_hi_hi_lo_hi = {fillBySeg_hi_hi_lo_hi_hi, fillBySeg_hi_hi_lo_hi_lo};
  wire [15:0]       fillBySeg_hi_hi_lo = {fillBySeg_hi_hi_lo_hi, fillBySeg_hi_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_hi_lo_lo = {fillBySeg_hi_hi_hi_lo_lo_hi, fillBySeg_hi_hi_hi_lo_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_hi_lo_hi = {fillBySeg_hi_hi_hi_lo_hi_hi, fillBySeg_hi_hi_hi_lo_hi_lo};
  wire [7:0]        fillBySeg_hi_hi_hi_lo = {fillBySeg_hi_hi_hi_lo_hi, fillBySeg_hi_hi_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_hi_hi_lo = {fillBySeg_hi_hi_hi_hi_lo_hi, fillBySeg_hi_hi_hi_hi_lo_lo};
  wire [3:0]        fillBySeg_hi_hi_hi_hi_hi = {fillBySeg_hi_hi_hi_hi_hi_hi, fillBySeg_hi_hi_hi_hi_hi_lo};
  wire [7:0]        fillBySeg_hi_hi_hi_hi = {fillBySeg_hi_hi_hi_hi_hi, fillBySeg_hi_hi_hi_hi_lo};
  wire [15:0]       fillBySeg_hi_hi_hi = {fillBySeg_hi_hi_hi_hi, fillBySeg_hi_hi_hi_lo};
  wire [31:0]       fillBySeg_hi_hi = {fillBySeg_hi_hi_hi, fillBySeg_hi_hi_lo};
  wire [63:0]       fillBySeg_hi = {fillBySeg_hi_hi, fillBySeg_hi_lo};
  wire [3:0]        fillBySeg_lo_lo_lo_lo_lo_lo_1 = {{2{maskForGroupWire[1]}}, {2{maskForGroupWire[0]}}};
  wire [3:0]        fillBySeg_lo_lo_lo_lo_lo_hi_1 = {{2{maskForGroupWire[3]}}, {2{maskForGroupWire[2]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_lo_lo_1 = {fillBySeg_lo_lo_lo_lo_lo_hi_1, fillBySeg_lo_lo_lo_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_lo_lo_lo_hi_lo_1 = {{2{maskForGroupWire[5]}}, {2{maskForGroupWire[4]}}};
  wire [3:0]        fillBySeg_lo_lo_lo_lo_hi_hi_1 = {{2{maskForGroupWire[7]}}, {2{maskForGroupWire[6]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_lo_hi_1 = {fillBySeg_lo_lo_lo_lo_hi_hi_1, fillBySeg_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]       fillBySeg_lo_lo_lo_lo_1 = {fillBySeg_lo_lo_lo_lo_hi_1, fillBySeg_lo_lo_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_lo_lo_hi_lo_lo_1 = {{2{maskForGroupWire[9]}}, {2{maskForGroupWire[8]}}};
  wire [3:0]        fillBySeg_lo_lo_lo_hi_lo_hi_1 = {{2{maskForGroupWire[11]}}, {2{maskForGroupWire[10]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_hi_lo_1 = {fillBySeg_lo_lo_lo_hi_lo_hi_1, fillBySeg_lo_lo_lo_hi_lo_lo_1};
  wire [3:0]        fillBySeg_lo_lo_lo_hi_hi_lo_1 = {{2{maskForGroupWire[13]}}, {2{maskForGroupWire[12]}}};
  wire [3:0]        fillBySeg_lo_lo_lo_hi_hi_hi_1 = {{2{maskForGroupWire[15]}}, {2{maskForGroupWire[14]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_hi_hi_1 = {fillBySeg_lo_lo_lo_hi_hi_hi_1, fillBySeg_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]       fillBySeg_lo_lo_lo_hi_1 = {fillBySeg_lo_lo_lo_hi_hi_1, fillBySeg_lo_lo_lo_hi_lo_1};
  wire [31:0]       fillBySeg_lo_lo_lo_1 = {fillBySeg_lo_lo_lo_hi_1, fillBySeg_lo_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_lo_hi_lo_lo_lo_1 = {{2{maskForGroupWire[17]}}, {2{maskForGroupWire[16]}}};
  wire [3:0]        fillBySeg_lo_lo_hi_lo_lo_hi_1 = {{2{maskForGroupWire[19]}}, {2{maskForGroupWire[18]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_lo_lo_1 = {fillBySeg_lo_lo_hi_lo_lo_hi_1, fillBySeg_lo_lo_hi_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_lo_hi_lo_hi_lo_1 = {{2{maskForGroupWire[21]}}, {2{maskForGroupWire[20]}}};
  wire [3:0]        fillBySeg_lo_lo_hi_lo_hi_hi_1 = {{2{maskForGroupWire[23]}}, {2{maskForGroupWire[22]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_lo_hi_1 = {fillBySeg_lo_lo_hi_lo_hi_hi_1, fillBySeg_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]       fillBySeg_lo_lo_hi_lo_1 = {fillBySeg_lo_lo_hi_lo_hi_1, fillBySeg_lo_lo_hi_lo_lo_1};
  wire [3:0]        fillBySeg_lo_lo_hi_hi_lo_lo_1 = {{2{maskForGroupWire[25]}}, {2{maskForGroupWire[24]}}};
  wire [3:0]        fillBySeg_lo_lo_hi_hi_lo_hi_1 = {{2{maskForGroupWire[27]}}, {2{maskForGroupWire[26]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_hi_lo_1 = {fillBySeg_lo_lo_hi_hi_lo_hi_1, fillBySeg_lo_lo_hi_hi_lo_lo_1};
  wire [3:0]        fillBySeg_lo_lo_hi_hi_hi_lo_1 = {{2{maskForGroupWire[29]}}, {2{maskForGroupWire[28]}}};
  wire [3:0]        fillBySeg_lo_lo_hi_hi_hi_hi_1 = {{2{maskForGroupWire[31]}}, {2{maskForGroupWire[30]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_hi_hi_1 = {fillBySeg_lo_lo_hi_hi_hi_hi_1, fillBySeg_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]       fillBySeg_lo_lo_hi_hi_1 = {fillBySeg_lo_lo_hi_hi_hi_1, fillBySeg_lo_lo_hi_hi_lo_1};
  wire [31:0]       fillBySeg_lo_lo_hi_1 = {fillBySeg_lo_lo_hi_hi_1, fillBySeg_lo_lo_hi_lo_1};
  wire [63:0]       fillBySeg_lo_lo_1 = {fillBySeg_lo_lo_hi_1, fillBySeg_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_lo_lo_lo_lo_1 = {{2{maskForGroupWire[33]}}, {2{maskForGroupWire[32]}}};
  wire [3:0]        fillBySeg_lo_hi_lo_lo_lo_hi_1 = {{2{maskForGroupWire[35]}}, {2{maskForGroupWire[34]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_lo_lo_1 = {fillBySeg_lo_hi_lo_lo_lo_hi_1, fillBySeg_lo_hi_lo_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_lo_lo_hi_lo_1 = {{2{maskForGroupWire[37]}}, {2{maskForGroupWire[36]}}};
  wire [3:0]        fillBySeg_lo_hi_lo_lo_hi_hi_1 = {{2{maskForGroupWire[39]}}, {2{maskForGroupWire[38]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_lo_hi_1 = {fillBySeg_lo_hi_lo_lo_hi_hi_1, fillBySeg_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]       fillBySeg_lo_hi_lo_lo_1 = {fillBySeg_lo_hi_lo_lo_hi_1, fillBySeg_lo_hi_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_lo_hi_lo_lo_1 = {{2{maskForGroupWire[41]}}, {2{maskForGroupWire[40]}}};
  wire [3:0]        fillBySeg_lo_hi_lo_hi_lo_hi_1 = {{2{maskForGroupWire[43]}}, {2{maskForGroupWire[42]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_hi_lo_1 = {fillBySeg_lo_hi_lo_hi_lo_hi_1, fillBySeg_lo_hi_lo_hi_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_lo_hi_hi_lo_1 = {{2{maskForGroupWire[45]}}, {2{maskForGroupWire[44]}}};
  wire [3:0]        fillBySeg_lo_hi_lo_hi_hi_hi_1 = {{2{maskForGroupWire[47]}}, {2{maskForGroupWire[46]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_hi_hi_1 = {fillBySeg_lo_hi_lo_hi_hi_hi_1, fillBySeg_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]       fillBySeg_lo_hi_lo_hi_1 = {fillBySeg_lo_hi_lo_hi_hi_1, fillBySeg_lo_hi_lo_hi_lo_1};
  wire [31:0]       fillBySeg_lo_hi_lo_1 = {fillBySeg_lo_hi_lo_hi_1, fillBySeg_lo_hi_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_hi_lo_lo_lo_1 = {{2{maskForGroupWire[49]}}, {2{maskForGroupWire[48]}}};
  wire [3:0]        fillBySeg_lo_hi_hi_lo_lo_hi_1 = {{2{maskForGroupWire[51]}}, {2{maskForGroupWire[50]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_lo_lo_1 = {fillBySeg_lo_hi_hi_lo_lo_hi_1, fillBySeg_lo_hi_hi_lo_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_hi_lo_hi_lo_1 = {{2{maskForGroupWire[53]}}, {2{maskForGroupWire[52]}}};
  wire [3:0]        fillBySeg_lo_hi_hi_lo_hi_hi_1 = {{2{maskForGroupWire[55]}}, {2{maskForGroupWire[54]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_lo_hi_1 = {fillBySeg_lo_hi_hi_lo_hi_hi_1, fillBySeg_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]       fillBySeg_lo_hi_hi_lo_1 = {fillBySeg_lo_hi_hi_lo_hi_1, fillBySeg_lo_hi_hi_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_hi_hi_lo_lo_1 = {{2{maskForGroupWire[57]}}, {2{maskForGroupWire[56]}}};
  wire [3:0]        fillBySeg_lo_hi_hi_hi_lo_hi_1 = {{2{maskForGroupWire[59]}}, {2{maskForGroupWire[58]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_hi_lo_1 = {fillBySeg_lo_hi_hi_hi_lo_hi_1, fillBySeg_lo_hi_hi_hi_lo_lo_1};
  wire [3:0]        fillBySeg_lo_hi_hi_hi_hi_lo_1 = {{2{maskForGroupWire[61]}}, {2{maskForGroupWire[60]}}};
  wire [3:0]        fillBySeg_lo_hi_hi_hi_hi_hi_1 = {{2{maskForGroupWire[63]}}, {2{maskForGroupWire[62]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_hi_hi_1 = {fillBySeg_lo_hi_hi_hi_hi_hi_1, fillBySeg_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]       fillBySeg_lo_hi_hi_hi_1 = {fillBySeg_lo_hi_hi_hi_hi_1, fillBySeg_lo_hi_hi_hi_lo_1};
  wire [31:0]       fillBySeg_lo_hi_hi_1 = {fillBySeg_lo_hi_hi_hi_1, fillBySeg_lo_hi_hi_lo_1};
  wire [63:0]       fillBySeg_lo_hi_1 = {fillBySeg_lo_hi_hi_1, fillBySeg_lo_hi_lo_1};
  wire [127:0]      fillBySeg_lo_1 = {fillBySeg_lo_hi_1, fillBySeg_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_lo_lo_lo_lo_1 = {{2{maskForGroupWire[65]}}, {2{maskForGroupWire[64]}}};
  wire [3:0]        fillBySeg_hi_lo_lo_lo_lo_hi_1 = {{2{maskForGroupWire[67]}}, {2{maskForGroupWire[66]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_lo_lo_1 = {fillBySeg_hi_lo_lo_lo_lo_hi_1, fillBySeg_hi_lo_lo_lo_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_lo_lo_hi_lo_1 = {{2{maskForGroupWire[69]}}, {2{maskForGroupWire[68]}}};
  wire [3:0]        fillBySeg_hi_lo_lo_lo_hi_hi_1 = {{2{maskForGroupWire[71]}}, {2{maskForGroupWire[70]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_lo_hi_1 = {fillBySeg_hi_lo_lo_lo_hi_hi_1, fillBySeg_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]       fillBySeg_hi_lo_lo_lo_1 = {fillBySeg_hi_lo_lo_lo_hi_1, fillBySeg_hi_lo_lo_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_lo_hi_lo_lo_1 = {{2{maskForGroupWire[73]}}, {2{maskForGroupWire[72]}}};
  wire [3:0]        fillBySeg_hi_lo_lo_hi_lo_hi_1 = {{2{maskForGroupWire[75]}}, {2{maskForGroupWire[74]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_hi_lo_1 = {fillBySeg_hi_lo_lo_hi_lo_hi_1, fillBySeg_hi_lo_lo_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_lo_hi_hi_lo_1 = {{2{maskForGroupWire[77]}}, {2{maskForGroupWire[76]}}};
  wire [3:0]        fillBySeg_hi_lo_lo_hi_hi_hi_1 = {{2{maskForGroupWire[79]}}, {2{maskForGroupWire[78]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_hi_hi_1 = {fillBySeg_hi_lo_lo_hi_hi_hi_1, fillBySeg_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]       fillBySeg_hi_lo_lo_hi_1 = {fillBySeg_hi_lo_lo_hi_hi_1, fillBySeg_hi_lo_lo_hi_lo_1};
  wire [31:0]       fillBySeg_hi_lo_lo_1 = {fillBySeg_hi_lo_lo_hi_1, fillBySeg_hi_lo_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_hi_lo_lo_lo_1 = {{2{maskForGroupWire[81]}}, {2{maskForGroupWire[80]}}};
  wire [3:0]        fillBySeg_hi_lo_hi_lo_lo_hi_1 = {{2{maskForGroupWire[83]}}, {2{maskForGroupWire[82]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_lo_lo_1 = {fillBySeg_hi_lo_hi_lo_lo_hi_1, fillBySeg_hi_lo_hi_lo_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_hi_lo_hi_lo_1 = {{2{maskForGroupWire[85]}}, {2{maskForGroupWire[84]}}};
  wire [3:0]        fillBySeg_hi_lo_hi_lo_hi_hi_1 = {{2{maskForGroupWire[87]}}, {2{maskForGroupWire[86]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_lo_hi_1 = {fillBySeg_hi_lo_hi_lo_hi_hi_1, fillBySeg_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]       fillBySeg_hi_lo_hi_lo_1 = {fillBySeg_hi_lo_hi_lo_hi_1, fillBySeg_hi_lo_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_hi_hi_lo_lo_1 = {{2{maskForGroupWire[89]}}, {2{maskForGroupWire[88]}}};
  wire [3:0]        fillBySeg_hi_lo_hi_hi_lo_hi_1 = {{2{maskForGroupWire[91]}}, {2{maskForGroupWire[90]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_hi_lo_1 = {fillBySeg_hi_lo_hi_hi_lo_hi_1, fillBySeg_hi_lo_hi_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_lo_hi_hi_hi_lo_1 = {{2{maskForGroupWire[93]}}, {2{maskForGroupWire[92]}}};
  wire [3:0]        fillBySeg_hi_lo_hi_hi_hi_hi_1 = {{2{maskForGroupWire[95]}}, {2{maskForGroupWire[94]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_hi_hi_1 = {fillBySeg_hi_lo_hi_hi_hi_hi_1, fillBySeg_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]       fillBySeg_hi_lo_hi_hi_1 = {fillBySeg_hi_lo_hi_hi_hi_1, fillBySeg_hi_lo_hi_hi_lo_1};
  wire [31:0]       fillBySeg_hi_lo_hi_1 = {fillBySeg_hi_lo_hi_hi_1, fillBySeg_hi_lo_hi_lo_1};
  wire [63:0]       fillBySeg_hi_lo_1 = {fillBySeg_hi_lo_hi_1, fillBySeg_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_lo_lo_lo_lo_1 = {{2{maskForGroupWire[97]}}, {2{maskForGroupWire[96]}}};
  wire [3:0]        fillBySeg_hi_hi_lo_lo_lo_hi_1 = {{2{maskForGroupWire[99]}}, {2{maskForGroupWire[98]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_lo_lo_1 = {fillBySeg_hi_hi_lo_lo_lo_hi_1, fillBySeg_hi_hi_lo_lo_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_lo_lo_hi_lo_1 = {{2{maskForGroupWire[101]}}, {2{maskForGroupWire[100]}}};
  wire [3:0]        fillBySeg_hi_hi_lo_lo_hi_hi_1 = {{2{maskForGroupWire[103]}}, {2{maskForGroupWire[102]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_lo_hi_1 = {fillBySeg_hi_hi_lo_lo_hi_hi_1, fillBySeg_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]       fillBySeg_hi_hi_lo_lo_1 = {fillBySeg_hi_hi_lo_lo_hi_1, fillBySeg_hi_hi_lo_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_lo_hi_lo_lo_1 = {{2{maskForGroupWire[105]}}, {2{maskForGroupWire[104]}}};
  wire [3:0]        fillBySeg_hi_hi_lo_hi_lo_hi_1 = {{2{maskForGroupWire[107]}}, {2{maskForGroupWire[106]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_hi_lo_1 = {fillBySeg_hi_hi_lo_hi_lo_hi_1, fillBySeg_hi_hi_lo_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_lo_hi_hi_lo_1 = {{2{maskForGroupWire[109]}}, {2{maskForGroupWire[108]}}};
  wire [3:0]        fillBySeg_hi_hi_lo_hi_hi_hi_1 = {{2{maskForGroupWire[111]}}, {2{maskForGroupWire[110]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_hi_hi_1 = {fillBySeg_hi_hi_lo_hi_hi_hi_1, fillBySeg_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]       fillBySeg_hi_hi_lo_hi_1 = {fillBySeg_hi_hi_lo_hi_hi_1, fillBySeg_hi_hi_lo_hi_lo_1};
  wire [31:0]       fillBySeg_hi_hi_lo_1 = {fillBySeg_hi_hi_lo_hi_1, fillBySeg_hi_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_hi_lo_lo_lo_1 = {{2{maskForGroupWire[113]}}, {2{maskForGroupWire[112]}}};
  wire [3:0]        fillBySeg_hi_hi_hi_lo_lo_hi_1 = {{2{maskForGroupWire[115]}}, {2{maskForGroupWire[114]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_lo_lo_1 = {fillBySeg_hi_hi_hi_lo_lo_hi_1, fillBySeg_hi_hi_hi_lo_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_hi_lo_hi_lo_1 = {{2{maskForGroupWire[117]}}, {2{maskForGroupWire[116]}}};
  wire [3:0]        fillBySeg_hi_hi_hi_lo_hi_hi_1 = {{2{maskForGroupWire[119]}}, {2{maskForGroupWire[118]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_lo_hi_1 = {fillBySeg_hi_hi_hi_lo_hi_hi_1, fillBySeg_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]       fillBySeg_hi_hi_hi_lo_1 = {fillBySeg_hi_hi_hi_lo_hi_1, fillBySeg_hi_hi_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_hi_hi_lo_lo_1 = {{2{maskForGroupWire[121]}}, {2{maskForGroupWire[120]}}};
  wire [3:0]        fillBySeg_hi_hi_hi_hi_lo_hi_1 = {{2{maskForGroupWire[123]}}, {2{maskForGroupWire[122]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_hi_lo_1 = {fillBySeg_hi_hi_hi_hi_lo_hi_1, fillBySeg_hi_hi_hi_hi_lo_lo_1};
  wire [3:0]        fillBySeg_hi_hi_hi_hi_hi_lo_1 = {{2{maskForGroupWire[125]}}, {2{maskForGroupWire[124]}}};
  wire [3:0]        fillBySeg_hi_hi_hi_hi_hi_hi_1 = {{2{maskForGroupWire[127]}}, {2{maskForGroupWire[126]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_hi_hi_1 = {fillBySeg_hi_hi_hi_hi_hi_hi_1, fillBySeg_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]       fillBySeg_hi_hi_hi_hi_1 = {fillBySeg_hi_hi_hi_hi_hi_1, fillBySeg_hi_hi_hi_hi_lo_1};
  wire [31:0]       fillBySeg_hi_hi_hi_1 = {fillBySeg_hi_hi_hi_hi_1, fillBySeg_hi_hi_hi_lo_1};
  wire [63:0]       fillBySeg_hi_hi_1 = {fillBySeg_hi_hi_hi_1, fillBySeg_hi_hi_lo_1};
  wire [127:0]      fillBySeg_hi_1 = {fillBySeg_hi_hi_1, fillBySeg_hi_lo_1};
  wire [5:0]        fillBySeg_lo_lo_lo_lo_lo_lo_2 = {{3{maskForGroupWire[1]}}, {3{maskForGroupWire[0]}}};
  wire [5:0]        fillBySeg_lo_lo_lo_lo_lo_hi_2 = {{3{maskForGroupWire[3]}}, {3{maskForGroupWire[2]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_lo_lo_2 = {fillBySeg_lo_lo_lo_lo_lo_hi_2, fillBySeg_lo_lo_lo_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_lo_lo_lo_hi_lo_2 = {{3{maskForGroupWire[5]}}, {3{maskForGroupWire[4]}}};
  wire [5:0]        fillBySeg_lo_lo_lo_lo_hi_hi_2 = {{3{maskForGroupWire[7]}}, {3{maskForGroupWire[6]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_lo_hi_2 = {fillBySeg_lo_lo_lo_lo_hi_hi_2, fillBySeg_lo_lo_lo_lo_hi_lo_2};
  wire [23:0]       fillBySeg_lo_lo_lo_lo_2 = {fillBySeg_lo_lo_lo_lo_hi_2, fillBySeg_lo_lo_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_lo_lo_hi_lo_lo_2 = {{3{maskForGroupWire[9]}}, {3{maskForGroupWire[8]}}};
  wire [5:0]        fillBySeg_lo_lo_lo_hi_lo_hi_2 = {{3{maskForGroupWire[11]}}, {3{maskForGroupWire[10]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_hi_lo_2 = {fillBySeg_lo_lo_lo_hi_lo_hi_2, fillBySeg_lo_lo_lo_hi_lo_lo_2};
  wire [5:0]        fillBySeg_lo_lo_lo_hi_hi_lo_2 = {{3{maskForGroupWire[13]}}, {3{maskForGroupWire[12]}}};
  wire [5:0]        fillBySeg_lo_lo_lo_hi_hi_hi_2 = {{3{maskForGroupWire[15]}}, {3{maskForGroupWire[14]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_hi_hi_2 = {fillBySeg_lo_lo_lo_hi_hi_hi_2, fillBySeg_lo_lo_lo_hi_hi_lo_2};
  wire [23:0]       fillBySeg_lo_lo_lo_hi_2 = {fillBySeg_lo_lo_lo_hi_hi_2, fillBySeg_lo_lo_lo_hi_lo_2};
  wire [47:0]       fillBySeg_lo_lo_lo_2 = {fillBySeg_lo_lo_lo_hi_2, fillBySeg_lo_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_lo_hi_lo_lo_lo_2 = {{3{maskForGroupWire[17]}}, {3{maskForGroupWire[16]}}};
  wire [5:0]        fillBySeg_lo_lo_hi_lo_lo_hi_2 = {{3{maskForGroupWire[19]}}, {3{maskForGroupWire[18]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_lo_lo_2 = {fillBySeg_lo_lo_hi_lo_lo_hi_2, fillBySeg_lo_lo_hi_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_lo_hi_lo_hi_lo_2 = {{3{maskForGroupWire[21]}}, {3{maskForGroupWire[20]}}};
  wire [5:0]        fillBySeg_lo_lo_hi_lo_hi_hi_2 = {{3{maskForGroupWire[23]}}, {3{maskForGroupWire[22]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_lo_hi_2 = {fillBySeg_lo_lo_hi_lo_hi_hi_2, fillBySeg_lo_lo_hi_lo_hi_lo_2};
  wire [23:0]       fillBySeg_lo_lo_hi_lo_2 = {fillBySeg_lo_lo_hi_lo_hi_2, fillBySeg_lo_lo_hi_lo_lo_2};
  wire [5:0]        fillBySeg_lo_lo_hi_hi_lo_lo_2 = {{3{maskForGroupWire[25]}}, {3{maskForGroupWire[24]}}};
  wire [5:0]        fillBySeg_lo_lo_hi_hi_lo_hi_2 = {{3{maskForGroupWire[27]}}, {3{maskForGroupWire[26]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_hi_lo_2 = {fillBySeg_lo_lo_hi_hi_lo_hi_2, fillBySeg_lo_lo_hi_hi_lo_lo_2};
  wire [5:0]        fillBySeg_lo_lo_hi_hi_hi_lo_2 = {{3{maskForGroupWire[29]}}, {3{maskForGroupWire[28]}}};
  wire [5:0]        fillBySeg_lo_lo_hi_hi_hi_hi_2 = {{3{maskForGroupWire[31]}}, {3{maskForGroupWire[30]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_hi_hi_2 = {fillBySeg_lo_lo_hi_hi_hi_hi_2, fillBySeg_lo_lo_hi_hi_hi_lo_2};
  wire [23:0]       fillBySeg_lo_lo_hi_hi_2 = {fillBySeg_lo_lo_hi_hi_hi_2, fillBySeg_lo_lo_hi_hi_lo_2};
  wire [47:0]       fillBySeg_lo_lo_hi_2 = {fillBySeg_lo_lo_hi_hi_2, fillBySeg_lo_lo_hi_lo_2};
  wire [95:0]       fillBySeg_lo_lo_2 = {fillBySeg_lo_lo_hi_2, fillBySeg_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_lo_lo_lo_lo_2 = {{3{maskForGroupWire[33]}}, {3{maskForGroupWire[32]}}};
  wire [5:0]        fillBySeg_lo_hi_lo_lo_lo_hi_2 = {{3{maskForGroupWire[35]}}, {3{maskForGroupWire[34]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_lo_lo_2 = {fillBySeg_lo_hi_lo_lo_lo_hi_2, fillBySeg_lo_hi_lo_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_lo_lo_hi_lo_2 = {{3{maskForGroupWire[37]}}, {3{maskForGroupWire[36]}}};
  wire [5:0]        fillBySeg_lo_hi_lo_lo_hi_hi_2 = {{3{maskForGroupWire[39]}}, {3{maskForGroupWire[38]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_lo_hi_2 = {fillBySeg_lo_hi_lo_lo_hi_hi_2, fillBySeg_lo_hi_lo_lo_hi_lo_2};
  wire [23:0]       fillBySeg_lo_hi_lo_lo_2 = {fillBySeg_lo_hi_lo_lo_hi_2, fillBySeg_lo_hi_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_lo_hi_lo_lo_2 = {{3{maskForGroupWire[41]}}, {3{maskForGroupWire[40]}}};
  wire [5:0]        fillBySeg_lo_hi_lo_hi_lo_hi_2 = {{3{maskForGroupWire[43]}}, {3{maskForGroupWire[42]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_hi_lo_2 = {fillBySeg_lo_hi_lo_hi_lo_hi_2, fillBySeg_lo_hi_lo_hi_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_lo_hi_hi_lo_2 = {{3{maskForGroupWire[45]}}, {3{maskForGroupWire[44]}}};
  wire [5:0]        fillBySeg_lo_hi_lo_hi_hi_hi_2 = {{3{maskForGroupWire[47]}}, {3{maskForGroupWire[46]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_hi_hi_2 = {fillBySeg_lo_hi_lo_hi_hi_hi_2, fillBySeg_lo_hi_lo_hi_hi_lo_2};
  wire [23:0]       fillBySeg_lo_hi_lo_hi_2 = {fillBySeg_lo_hi_lo_hi_hi_2, fillBySeg_lo_hi_lo_hi_lo_2};
  wire [47:0]       fillBySeg_lo_hi_lo_2 = {fillBySeg_lo_hi_lo_hi_2, fillBySeg_lo_hi_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_hi_lo_lo_lo_2 = {{3{maskForGroupWire[49]}}, {3{maskForGroupWire[48]}}};
  wire [5:0]        fillBySeg_lo_hi_hi_lo_lo_hi_2 = {{3{maskForGroupWire[51]}}, {3{maskForGroupWire[50]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_lo_lo_2 = {fillBySeg_lo_hi_hi_lo_lo_hi_2, fillBySeg_lo_hi_hi_lo_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_hi_lo_hi_lo_2 = {{3{maskForGroupWire[53]}}, {3{maskForGroupWire[52]}}};
  wire [5:0]        fillBySeg_lo_hi_hi_lo_hi_hi_2 = {{3{maskForGroupWire[55]}}, {3{maskForGroupWire[54]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_lo_hi_2 = {fillBySeg_lo_hi_hi_lo_hi_hi_2, fillBySeg_lo_hi_hi_lo_hi_lo_2};
  wire [23:0]       fillBySeg_lo_hi_hi_lo_2 = {fillBySeg_lo_hi_hi_lo_hi_2, fillBySeg_lo_hi_hi_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_hi_hi_lo_lo_2 = {{3{maskForGroupWire[57]}}, {3{maskForGroupWire[56]}}};
  wire [5:0]        fillBySeg_lo_hi_hi_hi_lo_hi_2 = {{3{maskForGroupWire[59]}}, {3{maskForGroupWire[58]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_hi_lo_2 = {fillBySeg_lo_hi_hi_hi_lo_hi_2, fillBySeg_lo_hi_hi_hi_lo_lo_2};
  wire [5:0]        fillBySeg_lo_hi_hi_hi_hi_lo_2 = {{3{maskForGroupWire[61]}}, {3{maskForGroupWire[60]}}};
  wire [5:0]        fillBySeg_lo_hi_hi_hi_hi_hi_2 = {{3{maskForGroupWire[63]}}, {3{maskForGroupWire[62]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_hi_hi_2 = {fillBySeg_lo_hi_hi_hi_hi_hi_2, fillBySeg_lo_hi_hi_hi_hi_lo_2};
  wire [23:0]       fillBySeg_lo_hi_hi_hi_2 = {fillBySeg_lo_hi_hi_hi_hi_2, fillBySeg_lo_hi_hi_hi_lo_2};
  wire [47:0]       fillBySeg_lo_hi_hi_2 = {fillBySeg_lo_hi_hi_hi_2, fillBySeg_lo_hi_hi_lo_2};
  wire [95:0]       fillBySeg_lo_hi_2 = {fillBySeg_lo_hi_hi_2, fillBySeg_lo_hi_lo_2};
  wire [191:0]      fillBySeg_lo_2 = {fillBySeg_lo_hi_2, fillBySeg_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_lo_lo_lo_lo_2 = {{3{maskForGroupWire[65]}}, {3{maskForGroupWire[64]}}};
  wire [5:0]        fillBySeg_hi_lo_lo_lo_lo_hi_2 = {{3{maskForGroupWire[67]}}, {3{maskForGroupWire[66]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_lo_lo_2 = {fillBySeg_hi_lo_lo_lo_lo_hi_2, fillBySeg_hi_lo_lo_lo_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_lo_lo_hi_lo_2 = {{3{maskForGroupWire[69]}}, {3{maskForGroupWire[68]}}};
  wire [5:0]        fillBySeg_hi_lo_lo_lo_hi_hi_2 = {{3{maskForGroupWire[71]}}, {3{maskForGroupWire[70]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_lo_hi_2 = {fillBySeg_hi_lo_lo_lo_hi_hi_2, fillBySeg_hi_lo_lo_lo_hi_lo_2};
  wire [23:0]       fillBySeg_hi_lo_lo_lo_2 = {fillBySeg_hi_lo_lo_lo_hi_2, fillBySeg_hi_lo_lo_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_lo_hi_lo_lo_2 = {{3{maskForGroupWire[73]}}, {3{maskForGroupWire[72]}}};
  wire [5:0]        fillBySeg_hi_lo_lo_hi_lo_hi_2 = {{3{maskForGroupWire[75]}}, {3{maskForGroupWire[74]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_hi_lo_2 = {fillBySeg_hi_lo_lo_hi_lo_hi_2, fillBySeg_hi_lo_lo_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_lo_hi_hi_lo_2 = {{3{maskForGroupWire[77]}}, {3{maskForGroupWire[76]}}};
  wire [5:0]        fillBySeg_hi_lo_lo_hi_hi_hi_2 = {{3{maskForGroupWire[79]}}, {3{maskForGroupWire[78]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_hi_hi_2 = {fillBySeg_hi_lo_lo_hi_hi_hi_2, fillBySeg_hi_lo_lo_hi_hi_lo_2};
  wire [23:0]       fillBySeg_hi_lo_lo_hi_2 = {fillBySeg_hi_lo_lo_hi_hi_2, fillBySeg_hi_lo_lo_hi_lo_2};
  wire [47:0]       fillBySeg_hi_lo_lo_2 = {fillBySeg_hi_lo_lo_hi_2, fillBySeg_hi_lo_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_hi_lo_lo_lo_2 = {{3{maskForGroupWire[81]}}, {3{maskForGroupWire[80]}}};
  wire [5:0]        fillBySeg_hi_lo_hi_lo_lo_hi_2 = {{3{maskForGroupWire[83]}}, {3{maskForGroupWire[82]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_lo_lo_2 = {fillBySeg_hi_lo_hi_lo_lo_hi_2, fillBySeg_hi_lo_hi_lo_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_hi_lo_hi_lo_2 = {{3{maskForGroupWire[85]}}, {3{maskForGroupWire[84]}}};
  wire [5:0]        fillBySeg_hi_lo_hi_lo_hi_hi_2 = {{3{maskForGroupWire[87]}}, {3{maskForGroupWire[86]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_lo_hi_2 = {fillBySeg_hi_lo_hi_lo_hi_hi_2, fillBySeg_hi_lo_hi_lo_hi_lo_2};
  wire [23:0]       fillBySeg_hi_lo_hi_lo_2 = {fillBySeg_hi_lo_hi_lo_hi_2, fillBySeg_hi_lo_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_hi_hi_lo_lo_2 = {{3{maskForGroupWire[89]}}, {3{maskForGroupWire[88]}}};
  wire [5:0]        fillBySeg_hi_lo_hi_hi_lo_hi_2 = {{3{maskForGroupWire[91]}}, {3{maskForGroupWire[90]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_hi_lo_2 = {fillBySeg_hi_lo_hi_hi_lo_hi_2, fillBySeg_hi_lo_hi_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_lo_hi_hi_hi_lo_2 = {{3{maskForGroupWire[93]}}, {3{maskForGroupWire[92]}}};
  wire [5:0]        fillBySeg_hi_lo_hi_hi_hi_hi_2 = {{3{maskForGroupWire[95]}}, {3{maskForGroupWire[94]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_hi_hi_2 = {fillBySeg_hi_lo_hi_hi_hi_hi_2, fillBySeg_hi_lo_hi_hi_hi_lo_2};
  wire [23:0]       fillBySeg_hi_lo_hi_hi_2 = {fillBySeg_hi_lo_hi_hi_hi_2, fillBySeg_hi_lo_hi_hi_lo_2};
  wire [47:0]       fillBySeg_hi_lo_hi_2 = {fillBySeg_hi_lo_hi_hi_2, fillBySeg_hi_lo_hi_lo_2};
  wire [95:0]       fillBySeg_hi_lo_2 = {fillBySeg_hi_lo_hi_2, fillBySeg_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_lo_lo_lo_lo_2 = {{3{maskForGroupWire[97]}}, {3{maskForGroupWire[96]}}};
  wire [5:0]        fillBySeg_hi_hi_lo_lo_lo_hi_2 = {{3{maskForGroupWire[99]}}, {3{maskForGroupWire[98]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_lo_lo_2 = {fillBySeg_hi_hi_lo_lo_lo_hi_2, fillBySeg_hi_hi_lo_lo_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_lo_lo_hi_lo_2 = {{3{maskForGroupWire[101]}}, {3{maskForGroupWire[100]}}};
  wire [5:0]        fillBySeg_hi_hi_lo_lo_hi_hi_2 = {{3{maskForGroupWire[103]}}, {3{maskForGroupWire[102]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_lo_hi_2 = {fillBySeg_hi_hi_lo_lo_hi_hi_2, fillBySeg_hi_hi_lo_lo_hi_lo_2};
  wire [23:0]       fillBySeg_hi_hi_lo_lo_2 = {fillBySeg_hi_hi_lo_lo_hi_2, fillBySeg_hi_hi_lo_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_lo_hi_lo_lo_2 = {{3{maskForGroupWire[105]}}, {3{maskForGroupWire[104]}}};
  wire [5:0]        fillBySeg_hi_hi_lo_hi_lo_hi_2 = {{3{maskForGroupWire[107]}}, {3{maskForGroupWire[106]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_hi_lo_2 = {fillBySeg_hi_hi_lo_hi_lo_hi_2, fillBySeg_hi_hi_lo_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_lo_hi_hi_lo_2 = {{3{maskForGroupWire[109]}}, {3{maskForGroupWire[108]}}};
  wire [5:0]        fillBySeg_hi_hi_lo_hi_hi_hi_2 = {{3{maskForGroupWire[111]}}, {3{maskForGroupWire[110]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_hi_hi_2 = {fillBySeg_hi_hi_lo_hi_hi_hi_2, fillBySeg_hi_hi_lo_hi_hi_lo_2};
  wire [23:0]       fillBySeg_hi_hi_lo_hi_2 = {fillBySeg_hi_hi_lo_hi_hi_2, fillBySeg_hi_hi_lo_hi_lo_2};
  wire [47:0]       fillBySeg_hi_hi_lo_2 = {fillBySeg_hi_hi_lo_hi_2, fillBySeg_hi_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_hi_lo_lo_lo_2 = {{3{maskForGroupWire[113]}}, {3{maskForGroupWire[112]}}};
  wire [5:0]        fillBySeg_hi_hi_hi_lo_lo_hi_2 = {{3{maskForGroupWire[115]}}, {3{maskForGroupWire[114]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_lo_lo_2 = {fillBySeg_hi_hi_hi_lo_lo_hi_2, fillBySeg_hi_hi_hi_lo_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_hi_lo_hi_lo_2 = {{3{maskForGroupWire[117]}}, {3{maskForGroupWire[116]}}};
  wire [5:0]        fillBySeg_hi_hi_hi_lo_hi_hi_2 = {{3{maskForGroupWire[119]}}, {3{maskForGroupWire[118]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_lo_hi_2 = {fillBySeg_hi_hi_hi_lo_hi_hi_2, fillBySeg_hi_hi_hi_lo_hi_lo_2};
  wire [23:0]       fillBySeg_hi_hi_hi_lo_2 = {fillBySeg_hi_hi_hi_lo_hi_2, fillBySeg_hi_hi_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_hi_hi_lo_lo_2 = {{3{maskForGroupWire[121]}}, {3{maskForGroupWire[120]}}};
  wire [5:0]        fillBySeg_hi_hi_hi_hi_lo_hi_2 = {{3{maskForGroupWire[123]}}, {3{maskForGroupWire[122]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_hi_lo_2 = {fillBySeg_hi_hi_hi_hi_lo_hi_2, fillBySeg_hi_hi_hi_hi_lo_lo_2};
  wire [5:0]        fillBySeg_hi_hi_hi_hi_hi_lo_2 = {{3{maskForGroupWire[125]}}, {3{maskForGroupWire[124]}}};
  wire [5:0]        fillBySeg_hi_hi_hi_hi_hi_hi_2 = {{3{maskForGroupWire[127]}}, {3{maskForGroupWire[126]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_hi_hi_2 = {fillBySeg_hi_hi_hi_hi_hi_hi_2, fillBySeg_hi_hi_hi_hi_hi_lo_2};
  wire [23:0]       fillBySeg_hi_hi_hi_hi_2 = {fillBySeg_hi_hi_hi_hi_hi_2, fillBySeg_hi_hi_hi_hi_lo_2};
  wire [47:0]       fillBySeg_hi_hi_hi_2 = {fillBySeg_hi_hi_hi_hi_2, fillBySeg_hi_hi_hi_lo_2};
  wire [95:0]       fillBySeg_hi_hi_2 = {fillBySeg_hi_hi_hi_2, fillBySeg_hi_hi_lo_2};
  wire [191:0]      fillBySeg_hi_2 = {fillBySeg_hi_hi_2, fillBySeg_hi_lo_2};
  wire [7:0]        fillBySeg_lo_lo_lo_lo_lo_lo_3 = {{4{maskForGroupWire[1]}}, {4{maskForGroupWire[0]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_lo_lo_hi_3 = {{4{maskForGroupWire[3]}}, {4{maskForGroupWire[2]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_lo_lo_3 = {fillBySeg_lo_lo_lo_lo_lo_hi_3, fillBySeg_lo_lo_lo_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_lo_lo_lo_hi_lo_3 = {{4{maskForGroupWire[5]}}, {4{maskForGroupWire[4]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_lo_hi_hi_3 = {{4{maskForGroupWire[7]}}, {4{maskForGroupWire[6]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_lo_hi_3 = {fillBySeg_lo_lo_lo_lo_hi_hi_3, fillBySeg_lo_lo_lo_lo_hi_lo_3};
  wire [31:0]       fillBySeg_lo_lo_lo_lo_3 = {fillBySeg_lo_lo_lo_lo_hi_3, fillBySeg_lo_lo_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_lo_lo_hi_lo_lo_3 = {{4{maskForGroupWire[9]}}, {4{maskForGroupWire[8]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_hi_lo_hi_3 = {{4{maskForGroupWire[11]}}, {4{maskForGroupWire[10]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_hi_lo_3 = {fillBySeg_lo_lo_lo_hi_lo_hi_3, fillBySeg_lo_lo_lo_hi_lo_lo_3};
  wire [7:0]        fillBySeg_lo_lo_lo_hi_hi_lo_3 = {{4{maskForGroupWire[13]}}, {4{maskForGroupWire[12]}}};
  wire [7:0]        fillBySeg_lo_lo_lo_hi_hi_hi_3 = {{4{maskForGroupWire[15]}}, {4{maskForGroupWire[14]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_hi_hi_3 = {fillBySeg_lo_lo_lo_hi_hi_hi_3, fillBySeg_lo_lo_lo_hi_hi_lo_3};
  wire [31:0]       fillBySeg_lo_lo_lo_hi_3 = {fillBySeg_lo_lo_lo_hi_hi_3, fillBySeg_lo_lo_lo_hi_lo_3};
  wire [63:0]       fillBySeg_lo_lo_lo_3 = {fillBySeg_lo_lo_lo_hi_3, fillBySeg_lo_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_lo_hi_lo_lo_lo_3 = {{4{maskForGroupWire[17]}}, {4{maskForGroupWire[16]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_lo_lo_hi_3 = {{4{maskForGroupWire[19]}}, {4{maskForGroupWire[18]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_lo_lo_3 = {fillBySeg_lo_lo_hi_lo_lo_hi_3, fillBySeg_lo_lo_hi_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_lo_hi_lo_hi_lo_3 = {{4{maskForGroupWire[21]}}, {4{maskForGroupWire[20]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_lo_hi_hi_3 = {{4{maskForGroupWire[23]}}, {4{maskForGroupWire[22]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_lo_hi_3 = {fillBySeg_lo_lo_hi_lo_hi_hi_3, fillBySeg_lo_lo_hi_lo_hi_lo_3};
  wire [31:0]       fillBySeg_lo_lo_hi_lo_3 = {fillBySeg_lo_lo_hi_lo_hi_3, fillBySeg_lo_lo_hi_lo_lo_3};
  wire [7:0]        fillBySeg_lo_lo_hi_hi_lo_lo_3 = {{4{maskForGroupWire[25]}}, {4{maskForGroupWire[24]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_hi_lo_hi_3 = {{4{maskForGroupWire[27]}}, {4{maskForGroupWire[26]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_hi_lo_3 = {fillBySeg_lo_lo_hi_hi_lo_hi_3, fillBySeg_lo_lo_hi_hi_lo_lo_3};
  wire [7:0]        fillBySeg_lo_lo_hi_hi_hi_lo_3 = {{4{maskForGroupWire[29]}}, {4{maskForGroupWire[28]}}};
  wire [7:0]        fillBySeg_lo_lo_hi_hi_hi_hi_3 = {{4{maskForGroupWire[31]}}, {4{maskForGroupWire[30]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_hi_hi_3 = {fillBySeg_lo_lo_hi_hi_hi_hi_3, fillBySeg_lo_lo_hi_hi_hi_lo_3};
  wire [31:0]       fillBySeg_lo_lo_hi_hi_3 = {fillBySeg_lo_lo_hi_hi_hi_3, fillBySeg_lo_lo_hi_hi_lo_3};
  wire [63:0]       fillBySeg_lo_lo_hi_3 = {fillBySeg_lo_lo_hi_hi_3, fillBySeg_lo_lo_hi_lo_3};
  wire [127:0]      fillBySeg_lo_lo_3 = {fillBySeg_lo_lo_hi_3, fillBySeg_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_lo_lo_lo_lo_3 = {{4{maskForGroupWire[33]}}, {4{maskForGroupWire[32]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_lo_lo_hi_3 = {{4{maskForGroupWire[35]}}, {4{maskForGroupWire[34]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_lo_lo_3 = {fillBySeg_lo_hi_lo_lo_lo_hi_3, fillBySeg_lo_hi_lo_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_lo_lo_hi_lo_3 = {{4{maskForGroupWire[37]}}, {4{maskForGroupWire[36]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_lo_hi_hi_3 = {{4{maskForGroupWire[39]}}, {4{maskForGroupWire[38]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_lo_hi_3 = {fillBySeg_lo_hi_lo_lo_hi_hi_3, fillBySeg_lo_hi_lo_lo_hi_lo_3};
  wire [31:0]       fillBySeg_lo_hi_lo_lo_3 = {fillBySeg_lo_hi_lo_lo_hi_3, fillBySeg_lo_hi_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_lo_hi_lo_lo_3 = {{4{maskForGroupWire[41]}}, {4{maskForGroupWire[40]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_hi_lo_hi_3 = {{4{maskForGroupWire[43]}}, {4{maskForGroupWire[42]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_hi_lo_3 = {fillBySeg_lo_hi_lo_hi_lo_hi_3, fillBySeg_lo_hi_lo_hi_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_lo_hi_hi_lo_3 = {{4{maskForGroupWire[45]}}, {4{maskForGroupWire[44]}}};
  wire [7:0]        fillBySeg_lo_hi_lo_hi_hi_hi_3 = {{4{maskForGroupWire[47]}}, {4{maskForGroupWire[46]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_hi_hi_3 = {fillBySeg_lo_hi_lo_hi_hi_hi_3, fillBySeg_lo_hi_lo_hi_hi_lo_3};
  wire [31:0]       fillBySeg_lo_hi_lo_hi_3 = {fillBySeg_lo_hi_lo_hi_hi_3, fillBySeg_lo_hi_lo_hi_lo_3};
  wire [63:0]       fillBySeg_lo_hi_lo_3 = {fillBySeg_lo_hi_lo_hi_3, fillBySeg_lo_hi_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_hi_lo_lo_lo_3 = {{4{maskForGroupWire[49]}}, {4{maskForGroupWire[48]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_lo_lo_hi_3 = {{4{maskForGroupWire[51]}}, {4{maskForGroupWire[50]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_lo_lo_3 = {fillBySeg_lo_hi_hi_lo_lo_hi_3, fillBySeg_lo_hi_hi_lo_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_hi_lo_hi_lo_3 = {{4{maskForGroupWire[53]}}, {4{maskForGroupWire[52]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_lo_hi_hi_3 = {{4{maskForGroupWire[55]}}, {4{maskForGroupWire[54]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_lo_hi_3 = {fillBySeg_lo_hi_hi_lo_hi_hi_3, fillBySeg_lo_hi_hi_lo_hi_lo_3};
  wire [31:0]       fillBySeg_lo_hi_hi_lo_3 = {fillBySeg_lo_hi_hi_lo_hi_3, fillBySeg_lo_hi_hi_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_hi_hi_lo_lo_3 = {{4{maskForGroupWire[57]}}, {4{maskForGroupWire[56]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_hi_lo_hi_3 = {{4{maskForGroupWire[59]}}, {4{maskForGroupWire[58]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_hi_lo_3 = {fillBySeg_lo_hi_hi_hi_lo_hi_3, fillBySeg_lo_hi_hi_hi_lo_lo_3};
  wire [7:0]        fillBySeg_lo_hi_hi_hi_hi_lo_3 = {{4{maskForGroupWire[61]}}, {4{maskForGroupWire[60]}}};
  wire [7:0]        fillBySeg_lo_hi_hi_hi_hi_hi_3 = {{4{maskForGroupWire[63]}}, {4{maskForGroupWire[62]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_hi_hi_3 = {fillBySeg_lo_hi_hi_hi_hi_hi_3, fillBySeg_lo_hi_hi_hi_hi_lo_3};
  wire [31:0]       fillBySeg_lo_hi_hi_hi_3 = {fillBySeg_lo_hi_hi_hi_hi_3, fillBySeg_lo_hi_hi_hi_lo_3};
  wire [63:0]       fillBySeg_lo_hi_hi_3 = {fillBySeg_lo_hi_hi_hi_3, fillBySeg_lo_hi_hi_lo_3};
  wire [127:0]      fillBySeg_lo_hi_3 = {fillBySeg_lo_hi_hi_3, fillBySeg_lo_hi_lo_3};
  wire [255:0]      fillBySeg_lo_3 = {fillBySeg_lo_hi_3, fillBySeg_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_lo_lo_lo_lo_3 = {{4{maskForGroupWire[65]}}, {4{maskForGroupWire[64]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_lo_lo_hi_3 = {{4{maskForGroupWire[67]}}, {4{maskForGroupWire[66]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_lo_lo_3 = {fillBySeg_hi_lo_lo_lo_lo_hi_3, fillBySeg_hi_lo_lo_lo_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_lo_lo_hi_lo_3 = {{4{maskForGroupWire[69]}}, {4{maskForGroupWire[68]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_lo_hi_hi_3 = {{4{maskForGroupWire[71]}}, {4{maskForGroupWire[70]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_lo_hi_3 = {fillBySeg_hi_lo_lo_lo_hi_hi_3, fillBySeg_hi_lo_lo_lo_hi_lo_3};
  wire [31:0]       fillBySeg_hi_lo_lo_lo_3 = {fillBySeg_hi_lo_lo_lo_hi_3, fillBySeg_hi_lo_lo_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_lo_hi_lo_lo_3 = {{4{maskForGroupWire[73]}}, {4{maskForGroupWire[72]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_hi_lo_hi_3 = {{4{maskForGroupWire[75]}}, {4{maskForGroupWire[74]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_hi_lo_3 = {fillBySeg_hi_lo_lo_hi_lo_hi_3, fillBySeg_hi_lo_lo_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_lo_hi_hi_lo_3 = {{4{maskForGroupWire[77]}}, {4{maskForGroupWire[76]}}};
  wire [7:0]        fillBySeg_hi_lo_lo_hi_hi_hi_3 = {{4{maskForGroupWire[79]}}, {4{maskForGroupWire[78]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_hi_hi_3 = {fillBySeg_hi_lo_lo_hi_hi_hi_3, fillBySeg_hi_lo_lo_hi_hi_lo_3};
  wire [31:0]       fillBySeg_hi_lo_lo_hi_3 = {fillBySeg_hi_lo_lo_hi_hi_3, fillBySeg_hi_lo_lo_hi_lo_3};
  wire [63:0]       fillBySeg_hi_lo_lo_3 = {fillBySeg_hi_lo_lo_hi_3, fillBySeg_hi_lo_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_hi_lo_lo_lo_3 = {{4{maskForGroupWire[81]}}, {4{maskForGroupWire[80]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_lo_lo_hi_3 = {{4{maskForGroupWire[83]}}, {4{maskForGroupWire[82]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_lo_lo_3 = {fillBySeg_hi_lo_hi_lo_lo_hi_3, fillBySeg_hi_lo_hi_lo_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_hi_lo_hi_lo_3 = {{4{maskForGroupWire[85]}}, {4{maskForGroupWire[84]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_lo_hi_hi_3 = {{4{maskForGroupWire[87]}}, {4{maskForGroupWire[86]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_lo_hi_3 = {fillBySeg_hi_lo_hi_lo_hi_hi_3, fillBySeg_hi_lo_hi_lo_hi_lo_3};
  wire [31:0]       fillBySeg_hi_lo_hi_lo_3 = {fillBySeg_hi_lo_hi_lo_hi_3, fillBySeg_hi_lo_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_hi_hi_lo_lo_3 = {{4{maskForGroupWire[89]}}, {4{maskForGroupWire[88]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_hi_lo_hi_3 = {{4{maskForGroupWire[91]}}, {4{maskForGroupWire[90]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_hi_lo_3 = {fillBySeg_hi_lo_hi_hi_lo_hi_3, fillBySeg_hi_lo_hi_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_lo_hi_hi_hi_lo_3 = {{4{maskForGroupWire[93]}}, {4{maskForGroupWire[92]}}};
  wire [7:0]        fillBySeg_hi_lo_hi_hi_hi_hi_3 = {{4{maskForGroupWire[95]}}, {4{maskForGroupWire[94]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_hi_hi_3 = {fillBySeg_hi_lo_hi_hi_hi_hi_3, fillBySeg_hi_lo_hi_hi_hi_lo_3};
  wire [31:0]       fillBySeg_hi_lo_hi_hi_3 = {fillBySeg_hi_lo_hi_hi_hi_3, fillBySeg_hi_lo_hi_hi_lo_3};
  wire [63:0]       fillBySeg_hi_lo_hi_3 = {fillBySeg_hi_lo_hi_hi_3, fillBySeg_hi_lo_hi_lo_3};
  wire [127:0]      fillBySeg_hi_lo_3 = {fillBySeg_hi_lo_hi_3, fillBySeg_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_lo_lo_lo_lo_3 = {{4{maskForGroupWire[97]}}, {4{maskForGroupWire[96]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_lo_lo_hi_3 = {{4{maskForGroupWire[99]}}, {4{maskForGroupWire[98]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_lo_lo_3 = {fillBySeg_hi_hi_lo_lo_lo_hi_3, fillBySeg_hi_hi_lo_lo_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_lo_lo_hi_lo_3 = {{4{maskForGroupWire[101]}}, {4{maskForGroupWire[100]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_lo_hi_hi_3 = {{4{maskForGroupWire[103]}}, {4{maskForGroupWire[102]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_lo_hi_3 = {fillBySeg_hi_hi_lo_lo_hi_hi_3, fillBySeg_hi_hi_lo_lo_hi_lo_3};
  wire [31:0]       fillBySeg_hi_hi_lo_lo_3 = {fillBySeg_hi_hi_lo_lo_hi_3, fillBySeg_hi_hi_lo_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_lo_hi_lo_lo_3 = {{4{maskForGroupWire[105]}}, {4{maskForGroupWire[104]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_hi_lo_hi_3 = {{4{maskForGroupWire[107]}}, {4{maskForGroupWire[106]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_hi_lo_3 = {fillBySeg_hi_hi_lo_hi_lo_hi_3, fillBySeg_hi_hi_lo_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_lo_hi_hi_lo_3 = {{4{maskForGroupWire[109]}}, {4{maskForGroupWire[108]}}};
  wire [7:0]        fillBySeg_hi_hi_lo_hi_hi_hi_3 = {{4{maskForGroupWire[111]}}, {4{maskForGroupWire[110]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_hi_hi_3 = {fillBySeg_hi_hi_lo_hi_hi_hi_3, fillBySeg_hi_hi_lo_hi_hi_lo_3};
  wire [31:0]       fillBySeg_hi_hi_lo_hi_3 = {fillBySeg_hi_hi_lo_hi_hi_3, fillBySeg_hi_hi_lo_hi_lo_3};
  wire [63:0]       fillBySeg_hi_hi_lo_3 = {fillBySeg_hi_hi_lo_hi_3, fillBySeg_hi_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_hi_lo_lo_lo_3 = {{4{maskForGroupWire[113]}}, {4{maskForGroupWire[112]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_lo_lo_hi_3 = {{4{maskForGroupWire[115]}}, {4{maskForGroupWire[114]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_lo_lo_3 = {fillBySeg_hi_hi_hi_lo_lo_hi_3, fillBySeg_hi_hi_hi_lo_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_hi_lo_hi_lo_3 = {{4{maskForGroupWire[117]}}, {4{maskForGroupWire[116]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_lo_hi_hi_3 = {{4{maskForGroupWire[119]}}, {4{maskForGroupWire[118]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_lo_hi_3 = {fillBySeg_hi_hi_hi_lo_hi_hi_3, fillBySeg_hi_hi_hi_lo_hi_lo_3};
  wire [31:0]       fillBySeg_hi_hi_hi_lo_3 = {fillBySeg_hi_hi_hi_lo_hi_3, fillBySeg_hi_hi_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_hi_hi_lo_lo_3 = {{4{maskForGroupWire[121]}}, {4{maskForGroupWire[120]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_hi_lo_hi_3 = {{4{maskForGroupWire[123]}}, {4{maskForGroupWire[122]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_hi_lo_3 = {fillBySeg_hi_hi_hi_hi_lo_hi_3, fillBySeg_hi_hi_hi_hi_lo_lo_3};
  wire [7:0]        fillBySeg_hi_hi_hi_hi_hi_lo_3 = {{4{maskForGroupWire[125]}}, {4{maskForGroupWire[124]}}};
  wire [7:0]        fillBySeg_hi_hi_hi_hi_hi_hi_3 = {{4{maskForGroupWire[127]}}, {4{maskForGroupWire[126]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_hi_hi_3 = {fillBySeg_hi_hi_hi_hi_hi_hi_3, fillBySeg_hi_hi_hi_hi_hi_lo_3};
  wire [31:0]       fillBySeg_hi_hi_hi_hi_3 = {fillBySeg_hi_hi_hi_hi_hi_3, fillBySeg_hi_hi_hi_hi_lo_3};
  wire [63:0]       fillBySeg_hi_hi_hi_3 = {fillBySeg_hi_hi_hi_hi_3, fillBySeg_hi_hi_hi_lo_3};
  wire [127:0]      fillBySeg_hi_hi_3 = {fillBySeg_hi_hi_hi_3, fillBySeg_hi_hi_lo_3};
  wire [255:0]      fillBySeg_hi_3 = {fillBySeg_hi_hi_3, fillBySeg_hi_lo_3};
  wire [9:0]        fillBySeg_lo_lo_lo_lo_lo_lo_4 = {{5{maskForGroupWire[1]}}, {5{maskForGroupWire[0]}}};
  wire [9:0]        fillBySeg_lo_lo_lo_lo_lo_hi_4 = {{5{maskForGroupWire[3]}}, {5{maskForGroupWire[2]}}};
  wire [19:0]       fillBySeg_lo_lo_lo_lo_lo_4 = {fillBySeg_lo_lo_lo_lo_lo_hi_4, fillBySeg_lo_lo_lo_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_lo_lo_lo_hi_lo_4 = {{5{maskForGroupWire[5]}}, {5{maskForGroupWire[4]}}};
  wire [9:0]        fillBySeg_lo_lo_lo_lo_hi_hi_4 = {{5{maskForGroupWire[7]}}, {5{maskForGroupWire[6]}}};
  wire [19:0]       fillBySeg_lo_lo_lo_lo_hi_4 = {fillBySeg_lo_lo_lo_lo_hi_hi_4, fillBySeg_lo_lo_lo_lo_hi_lo_4};
  wire [39:0]       fillBySeg_lo_lo_lo_lo_4 = {fillBySeg_lo_lo_lo_lo_hi_4, fillBySeg_lo_lo_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_lo_lo_hi_lo_lo_4 = {{5{maskForGroupWire[9]}}, {5{maskForGroupWire[8]}}};
  wire [9:0]        fillBySeg_lo_lo_lo_hi_lo_hi_4 = {{5{maskForGroupWire[11]}}, {5{maskForGroupWire[10]}}};
  wire [19:0]       fillBySeg_lo_lo_lo_hi_lo_4 = {fillBySeg_lo_lo_lo_hi_lo_hi_4, fillBySeg_lo_lo_lo_hi_lo_lo_4};
  wire [9:0]        fillBySeg_lo_lo_lo_hi_hi_lo_4 = {{5{maskForGroupWire[13]}}, {5{maskForGroupWire[12]}}};
  wire [9:0]        fillBySeg_lo_lo_lo_hi_hi_hi_4 = {{5{maskForGroupWire[15]}}, {5{maskForGroupWire[14]}}};
  wire [19:0]       fillBySeg_lo_lo_lo_hi_hi_4 = {fillBySeg_lo_lo_lo_hi_hi_hi_4, fillBySeg_lo_lo_lo_hi_hi_lo_4};
  wire [39:0]       fillBySeg_lo_lo_lo_hi_4 = {fillBySeg_lo_lo_lo_hi_hi_4, fillBySeg_lo_lo_lo_hi_lo_4};
  wire [79:0]       fillBySeg_lo_lo_lo_4 = {fillBySeg_lo_lo_lo_hi_4, fillBySeg_lo_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_lo_hi_lo_lo_lo_4 = {{5{maskForGroupWire[17]}}, {5{maskForGroupWire[16]}}};
  wire [9:0]        fillBySeg_lo_lo_hi_lo_lo_hi_4 = {{5{maskForGroupWire[19]}}, {5{maskForGroupWire[18]}}};
  wire [19:0]       fillBySeg_lo_lo_hi_lo_lo_4 = {fillBySeg_lo_lo_hi_lo_lo_hi_4, fillBySeg_lo_lo_hi_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_lo_hi_lo_hi_lo_4 = {{5{maskForGroupWire[21]}}, {5{maskForGroupWire[20]}}};
  wire [9:0]        fillBySeg_lo_lo_hi_lo_hi_hi_4 = {{5{maskForGroupWire[23]}}, {5{maskForGroupWire[22]}}};
  wire [19:0]       fillBySeg_lo_lo_hi_lo_hi_4 = {fillBySeg_lo_lo_hi_lo_hi_hi_4, fillBySeg_lo_lo_hi_lo_hi_lo_4};
  wire [39:0]       fillBySeg_lo_lo_hi_lo_4 = {fillBySeg_lo_lo_hi_lo_hi_4, fillBySeg_lo_lo_hi_lo_lo_4};
  wire [9:0]        fillBySeg_lo_lo_hi_hi_lo_lo_4 = {{5{maskForGroupWire[25]}}, {5{maskForGroupWire[24]}}};
  wire [9:0]        fillBySeg_lo_lo_hi_hi_lo_hi_4 = {{5{maskForGroupWire[27]}}, {5{maskForGroupWire[26]}}};
  wire [19:0]       fillBySeg_lo_lo_hi_hi_lo_4 = {fillBySeg_lo_lo_hi_hi_lo_hi_4, fillBySeg_lo_lo_hi_hi_lo_lo_4};
  wire [9:0]        fillBySeg_lo_lo_hi_hi_hi_lo_4 = {{5{maskForGroupWire[29]}}, {5{maskForGroupWire[28]}}};
  wire [9:0]        fillBySeg_lo_lo_hi_hi_hi_hi_4 = {{5{maskForGroupWire[31]}}, {5{maskForGroupWire[30]}}};
  wire [19:0]       fillBySeg_lo_lo_hi_hi_hi_4 = {fillBySeg_lo_lo_hi_hi_hi_hi_4, fillBySeg_lo_lo_hi_hi_hi_lo_4};
  wire [39:0]       fillBySeg_lo_lo_hi_hi_4 = {fillBySeg_lo_lo_hi_hi_hi_4, fillBySeg_lo_lo_hi_hi_lo_4};
  wire [79:0]       fillBySeg_lo_lo_hi_4 = {fillBySeg_lo_lo_hi_hi_4, fillBySeg_lo_lo_hi_lo_4};
  wire [159:0]      fillBySeg_lo_lo_4 = {fillBySeg_lo_lo_hi_4, fillBySeg_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_lo_lo_lo_lo_4 = {{5{maskForGroupWire[33]}}, {5{maskForGroupWire[32]}}};
  wire [9:0]        fillBySeg_lo_hi_lo_lo_lo_hi_4 = {{5{maskForGroupWire[35]}}, {5{maskForGroupWire[34]}}};
  wire [19:0]       fillBySeg_lo_hi_lo_lo_lo_4 = {fillBySeg_lo_hi_lo_lo_lo_hi_4, fillBySeg_lo_hi_lo_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_lo_lo_hi_lo_4 = {{5{maskForGroupWire[37]}}, {5{maskForGroupWire[36]}}};
  wire [9:0]        fillBySeg_lo_hi_lo_lo_hi_hi_4 = {{5{maskForGroupWire[39]}}, {5{maskForGroupWire[38]}}};
  wire [19:0]       fillBySeg_lo_hi_lo_lo_hi_4 = {fillBySeg_lo_hi_lo_lo_hi_hi_4, fillBySeg_lo_hi_lo_lo_hi_lo_4};
  wire [39:0]       fillBySeg_lo_hi_lo_lo_4 = {fillBySeg_lo_hi_lo_lo_hi_4, fillBySeg_lo_hi_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_lo_hi_lo_lo_4 = {{5{maskForGroupWire[41]}}, {5{maskForGroupWire[40]}}};
  wire [9:0]        fillBySeg_lo_hi_lo_hi_lo_hi_4 = {{5{maskForGroupWire[43]}}, {5{maskForGroupWire[42]}}};
  wire [19:0]       fillBySeg_lo_hi_lo_hi_lo_4 = {fillBySeg_lo_hi_lo_hi_lo_hi_4, fillBySeg_lo_hi_lo_hi_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_lo_hi_hi_lo_4 = {{5{maskForGroupWire[45]}}, {5{maskForGroupWire[44]}}};
  wire [9:0]        fillBySeg_lo_hi_lo_hi_hi_hi_4 = {{5{maskForGroupWire[47]}}, {5{maskForGroupWire[46]}}};
  wire [19:0]       fillBySeg_lo_hi_lo_hi_hi_4 = {fillBySeg_lo_hi_lo_hi_hi_hi_4, fillBySeg_lo_hi_lo_hi_hi_lo_4};
  wire [39:0]       fillBySeg_lo_hi_lo_hi_4 = {fillBySeg_lo_hi_lo_hi_hi_4, fillBySeg_lo_hi_lo_hi_lo_4};
  wire [79:0]       fillBySeg_lo_hi_lo_4 = {fillBySeg_lo_hi_lo_hi_4, fillBySeg_lo_hi_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_hi_lo_lo_lo_4 = {{5{maskForGroupWire[49]}}, {5{maskForGroupWire[48]}}};
  wire [9:0]        fillBySeg_lo_hi_hi_lo_lo_hi_4 = {{5{maskForGroupWire[51]}}, {5{maskForGroupWire[50]}}};
  wire [19:0]       fillBySeg_lo_hi_hi_lo_lo_4 = {fillBySeg_lo_hi_hi_lo_lo_hi_4, fillBySeg_lo_hi_hi_lo_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_hi_lo_hi_lo_4 = {{5{maskForGroupWire[53]}}, {5{maskForGroupWire[52]}}};
  wire [9:0]        fillBySeg_lo_hi_hi_lo_hi_hi_4 = {{5{maskForGroupWire[55]}}, {5{maskForGroupWire[54]}}};
  wire [19:0]       fillBySeg_lo_hi_hi_lo_hi_4 = {fillBySeg_lo_hi_hi_lo_hi_hi_4, fillBySeg_lo_hi_hi_lo_hi_lo_4};
  wire [39:0]       fillBySeg_lo_hi_hi_lo_4 = {fillBySeg_lo_hi_hi_lo_hi_4, fillBySeg_lo_hi_hi_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_hi_hi_lo_lo_4 = {{5{maskForGroupWire[57]}}, {5{maskForGroupWire[56]}}};
  wire [9:0]        fillBySeg_lo_hi_hi_hi_lo_hi_4 = {{5{maskForGroupWire[59]}}, {5{maskForGroupWire[58]}}};
  wire [19:0]       fillBySeg_lo_hi_hi_hi_lo_4 = {fillBySeg_lo_hi_hi_hi_lo_hi_4, fillBySeg_lo_hi_hi_hi_lo_lo_4};
  wire [9:0]        fillBySeg_lo_hi_hi_hi_hi_lo_4 = {{5{maskForGroupWire[61]}}, {5{maskForGroupWire[60]}}};
  wire [9:0]        fillBySeg_lo_hi_hi_hi_hi_hi_4 = {{5{maskForGroupWire[63]}}, {5{maskForGroupWire[62]}}};
  wire [19:0]       fillBySeg_lo_hi_hi_hi_hi_4 = {fillBySeg_lo_hi_hi_hi_hi_hi_4, fillBySeg_lo_hi_hi_hi_hi_lo_4};
  wire [39:0]       fillBySeg_lo_hi_hi_hi_4 = {fillBySeg_lo_hi_hi_hi_hi_4, fillBySeg_lo_hi_hi_hi_lo_4};
  wire [79:0]       fillBySeg_lo_hi_hi_4 = {fillBySeg_lo_hi_hi_hi_4, fillBySeg_lo_hi_hi_lo_4};
  wire [159:0]      fillBySeg_lo_hi_4 = {fillBySeg_lo_hi_hi_4, fillBySeg_lo_hi_lo_4};
  wire [319:0]      fillBySeg_lo_4 = {fillBySeg_lo_hi_4, fillBySeg_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_lo_lo_lo_lo_4 = {{5{maskForGroupWire[65]}}, {5{maskForGroupWire[64]}}};
  wire [9:0]        fillBySeg_hi_lo_lo_lo_lo_hi_4 = {{5{maskForGroupWire[67]}}, {5{maskForGroupWire[66]}}};
  wire [19:0]       fillBySeg_hi_lo_lo_lo_lo_4 = {fillBySeg_hi_lo_lo_lo_lo_hi_4, fillBySeg_hi_lo_lo_lo_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_lo_lo_hi_lo_4 = {{5{maskForGroupWire[69]}}, {5{maskForGroupWire[68]}}};
  wire [9:0]        fillBySeg_hi_lo_lo_lo_hi_hi_4 = {{5{maskForGroupWire[71]}}, {5{maskForGroupWire[70]}}};
  wire [19:0]       fillBySeg_hi_lo_lo_lo_hi_4 = {fillBySeg_hi_lo_lo_lo_hi_hi_4, fillBySeg_hi_lo_lo_lo_hi_lo_4};
  wire [39:0]       fillBySeg_hi_lo_lo_lo_4 = {fillBySeg_hi_lo_lo_lo_hi_4, fillBySeg_hi_lo_lo_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_lo_hi_lo_lo_4 = {{5{maskForGroupWire[73]}}, {5{maskForGroupWire[72]}}};
  wire [9:0]        fillBySeg_hi_lo_lo_hi_lo_hi_4 = {{5{maskForGroupWire[75]}}, {5{maskForGroupWire[74]}}};
  wire [19:0]       fillBySeg_hi_lo_lo_hi_lo_4 = {fillBySeg_hi_lo_lo_hi_lo_hi_4, fillBySeg_hi_lo_lo_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_lo_hi_hi_lo_4 = {{5{maskForGroupWire[77]}}, {5{maskForGroupWire[76]}}};
  wire [9:0]        fillBySeg_hi_lo_lo_hi_hi_hi_4 = {{5{maskForGroupWire[79]}}, {5{maskForGroupWire[78]}}};
  wire [19:0]       fillBySeg_hi_lo_lo_hi_hi_4 = {fillBySeg_hi_lo_lo_hi_hi_hi_4, fillBySeg_hi_lo_lo_hi_hi_lo_4};
  wire [39:0]       fillBySeg_hi_lo_lo_hi_4 = {fillBySeg_hi_lo_lo_hi_hi_4, fillBySeg_hi_lo_lo_hi_lo_4};
  wire [79:0]       fillBySeg_hi_lo_lo_4 = {fillBySeg_hi_lo_lo_hi_4, fillBySeg_hi_lo_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_hi_lo_lo_lo_4 = {{5{maskForGroupWire[81]}}, {5{maskForGroupWire[80]}}};
  wire [9:0]        fillBySeg_hi_lo_hi_lo_lo_hi_4 = {{5{maskForGroupWire[83]}}, {5{maskForGroupWire[82]}}};
  wire [19:0]       fillBySeg_hi_lo_hi_lo_lo_4 = {fillBySeg_hi_lo_hi_lo_lo_hi_4, fillBySeg_hi_lo_hi_lo_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_hi_lo_hi_lo_4 = {{5{maskForGroupWire[85]}}, {5{maskForGroupWire[84]}}};
  wire [9:0]        fillBySeg_hi_lo_hi_lo_hi_hi_4 = {{5{maskForGroupWire[87]}}, {5{maskForGroupWire[86]}}};
  wire [19:0]       fillBySeg_hi_lo_hi_lo_hi_4 = {fillBySeg_hi_lo_hi_lo_hi_hi_4, fillBySeg_hi_lo_hi_lo_hi_lo_4};
  wire [39:0]       fillBySeg_hi_lo_hi_lo_4 = {fillBySeg_hi_lo_hi_lo_hi_4, fillBySeg_hi_lo_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_hi_hi_lo_lo_4 = {{5{maskForGroupWire[89]}}, {5{maskForGroupWire[88]}}};
  wire [9:0]        fillBySeg_hi_lo_hi_hi_lo_hi_4 = {{5{maskForGroupWire[91]}}, {5{maskForGroupWire[90]}}};
  wire [19:0]       fillBySeg_hi_lo_hi_hi_lo_4 = {fillBySeg_hi_lo_hi_hi_lo_hi_4, fillBySeg_hi_lo_hi_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_lo_hi_hi_hi_lo_4 = {{5{maskForGroupWire[93]}}, {5{maskForGroupWire[92]}}};
  wire [9:0]        fillBySeg_hi_lo_hi_hi_hi_hi_4 = {{5{maskForGroupWire[95]}}, {5{maskForGroupWire[94]}}};
  wire [19:0]       fillBySeg_hi_lo_hi_hi_hi_4 = {fillBySeg_hi_lo_hi_hi_hi_hi_4, fillBySeg_hi_lo_hi_hi_hi_lo_4};
  wire [39:0]       fillBySeg_hi_lo_hi_hi_4 = {fillBySeg_hi_lo_hi_hi_hi_4, fillBySeg_hi_lo_hi_hi_lo_4};
  wire [79:0]       fillBySeg_hi_lo_hi_4 = {fillBySeg_hi_lo_hi_hi_4, fillBySeg_hi_lo_hi_lo_4};
  wire [159:0]      fillBySeg_hi_lo_4 = {fillBySeg_hi_lo_hi_4, fillBySeg_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_lo_lo_lo_lo_4 = {{5{maskForGroupWire[97]}}, {5{maskForGroupWire[96]}}};
  wire [9:0]        fillBySeg_hi_hi_lo_lo_lo_hi_4 = {{5{maskForGroupWire[99]}}, {5{maskForGroupWire[98]}}};
  wire [19:0]       fillBySeg_hi_hi_lo_lo_lo_4 = {fillBySeg_hi_hi_lo_lo_lo_hi_4, fillBySeg_hi_hi_lo_lo_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_lo_lo_hi_lo_4 = {{5{maskForGroupWire[101]}}, {5{maskForGroupWire[100]}}};
  wire [9:0]        fillBySeg_hi_hi_lo_lo_hi_hi_4 = {{5{maskForGroupWire[103]}}, {5{maskForGroupWire[102]}}};
  wire [19:0]       fillBySeg_hi_hi_lo_lo_hi_4 = {fillBySeg_hi_hi_lo_lo_hi_hi_4, fillBySeg_hi_hi_lo_lo_hi_lo_4};
  wire [39:0]       fillBySeg_hi_hi_lo_lo_4 = {fillBySeg_hi_hi_lo_lo_hi_4, fillBySeg_hi_hi_lo_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_lo_hi_lo_lo_4 = {{5{maskForGroupWire[105]}}, {5{maskForGroupWire[104]}}};
  wire [9:0]        fillBySeg_hi_hi_lo_hi_lo_hi_4 = {{5{maskForGroupWire[107]}}, {5{maskForGroupWire[106]}}};
  wire [19:0]       fillBySeg_hi_hi_lo_hi_lo_4 = {fillBySeg_hi_hi_lo_hi_lo_hi_4, fillBySeg_hi_hi_lo_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_lo_hi_hi_lo_4 = {{5{maskForGroupWire[109]}}, {5{maskForGroupWire[108]}}};
  wire [9:0]        fillBySeg_hi_hi_lo_hi_hi_hi_4 = {{5{maskForGroupWire[111]}}, {5{maskForGroupWire[110]}}};
  wire [19:0]       fillBySeg_hi_hi_lo_hi_hi_4 = {fillBySeg_hi_hi_lo_hi_hi_hi_4, fillBySeg_hi_hi_lo_hi_hi_lo_4};
  wire [39:0]       fillBySeg_hi_hi_lo_hi_4 = {fillBySeg_hi_hi_lo_hi_hi_4, fillBySeg_hi_hi_lo_hi_lo_4};
  wire [79:0]       fillBySeg_hi_hi_lo_4 = {fillBySeg_hi_hi_lo_hi_4, fillBySeg_hi_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_hi_lo_lo_lo_4 = {{5{maskForGroupWire[113]}}, {5{maskForGroupWire[112]}}};
  wire [9:0]        fillBySeg_hi_hi_hi_lo_lo_hi_4 = {{5{maskForGroupWire[115]}}, {5{maskForGroupWire[114]}}};
  wire [19:0]       fillBySeg_hi_hi_hi_lo_lo_4 = {fillBySeg_hi_hi_hi_lo_lo_hi_4, fillBySeg_hi_hi_hi_lo_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_hi_lo_hi_lo_4 = {{5{maskForGroupWire[117]}}, {5{maskForGroupWire[116]}}};
  wire [9:0]        fillBySeg_hi_hi_hi_lo_hi_hi_4 = {{5{maskForGroupWire[119]}}, {5{maskForGroupWire[118]}}};
  wire [19:0]       fillBySeg_hi_hi_hi_lo_hi_4 = {fillBySeg_hi_hi_hi_lo_hi_hi_4, fillBySeg_hi_hi_hi_lo_hi_lo_4};
  wire [39:0]       fillBySeg_hi_hi_hi_lo_4 = {fillBySeg_hi_hi_hi_lo_hi_4, fillBySeg_hi_hi_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_hi_hi_lo_lo_4 = {{5{maskForGroupWire[121]}}, {5{maskForGroupWire[120]}}};
  wire [9:0]        fillBySeg_hi_hi_hi_hi_lo_hi_4 = {{5{maskForGroupWire[123]}}, {5{maskForGroupWire[122]}}};
  wire [19:0]       fillBySeg_hi_hi_hi_hi_lo_4 = {fillBySeg_hi_hi_hi_hi_lo_hi_4, fillBySeg_hi_hi_hi_hi_lo_lo_4};
  wire [9:0]        fillBySeg_hi_hi_hi_hi_hi_lo_4 = {{5{maskForGroupWire[125]}}, {5{maskForGroupWire[124]}}};
  wire [9:0]        fillBySeg_hi_hi_hi_hi_hi_hi_4 = {{5{maskForGroupWire[127]}}, {5{maskForGroupWire[126]}}};
  wire [19:0]       fillBySeg_hi_hi_hi_hi_hi_4 = {fillBySeg_hi_hi_hi_hi_hi_hi_4, fillBySeg_hi_hi_hi_hi_hi_lo_4};
  wire [39:0]       fillBySeg_hi_hi_hi_hi_4 = {fillBySeg_hi_hi_hi_hi_hi_4, fillBySeg_hi_hi_hi_hi_lo_4};
  wire [79:0]       fillBySeg_hi_hi_hi_4 = {fillBySeg_hi_hi_hi_hi_4, fillBySeg_hi_hi_hi_lo_4};
  wire [159:0]      fillBySeg_hi_hi_4 = {fillBySeg_hi_hi_hi_4, fillBySeg_hi_hi_lo_4};
  wire [319:0]      fillBySeg_hi_4 = {fillBySeg_hi_hi_4, fillBySeg_hi_lo_4};
  wire [11:0]       fillBySeg_lo_lo_lo_lo_lo_lo_5 = {{6{maskForGroupWire[1]}}, {6{maskForGroupWire[0]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_lo_lo_hi_5 = {{6{maskForGroupWire[3]}}, {6{maskForGroupWire[2]}}};
  wire [23:0]       fillBySeg_lo_lo_lo_lo_lo_5 = {fillBySeg_lo_lo_lo_lo_lo_hi_5, fillBySeg_lo_lo_lo_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_lo_lo_lo_hi_lo_5 = {{6{maskForGroupWire[5]}}, {6{maskForGroupWire[4]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_lo_hi_hi_5 = {{6{maskForGroupWire[7]}}, {6{maskForGroupWire[6]}}};
  wire [23:0]       fillBySeg_lo_lo_lo_lo_hi_5 = {fillBySeg_lo_lo_lo_lo_hi_hi_5, fillBySeg_lo_lo_lo_lo_hi_lo_5};
  wire [47:0]       fillBySeg_lo_lo_lo_lo_5 = {fillBySeg_lo_lo_lo_lo_hi_5, fillBySeg_lo_lo_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_lo_lo_hi_lo_lo_5 = {{6{maskForGroupWire[9]}}, {6{maskForGroupWire[8]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_hi_lo_hi_5 = {{6{maskForGroupWire[11]}}, {6{maskForGroupWire[10]}}};
  wire [23:0]       fillBySeg_lo_lo_lo_hi_lo_5 = {fillBySeg_lo_lo_lo_hi_lo_hi_5, fillBySeg_lo_lo_lo_hi_lo_lo_5};
  wire [11:0]       fillBySeg_lo_lo_lo_hi_hi_lo_5 = {{6{maskForGroupWire[13]}}, {6{maskForGroupWire[12]}}};
  wire [11:0]       fillBySeg_lo_lo_lo_hi_hi_hi_5 = {{6{maskForGroupWire[15]}}, {6{maskForGroupWire[14]}}};
  wire [23:0]       fillBySeg_lo_lo_lo_hi_hi_5 = {fillBySeg_lo_lo_lo_hi_hi_hi_5, fillBySeg_lo_lo_lo_hi_hi_lo_5};
  wire [47:0]       fillBySeg_lo_lo_lo_hi_5 = {fillBySeg_lo_lo_lo_hi_hi_5, fillBySeg_lo_lo_lo_hi_lo_5};
  wire [95:0]       fillBySeg_lo_lo_lo_5 = {fillBySeg_lo_lo_lo_hi_5, fillBySeg_lo_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_lo_hi_lo_lo_lo_5 = {{6{maskForGroupWire[17]}}, {6{maskForGroupWire[16]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_lo_lo_hi_5 = {{6{maskForGroupWire[19]}}, {6{maskForGroupWire[18]}}};
  wire [23:0]       fillBySeg_lo_lo_hi_lo_lo_5 = {fillBySeg_lo_lo_hi_lo_lo_hi_5, fillBySeg_lo_lo_hi_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_lo_hi_lo_hi_lo_5 = {{6{maskForGroupWire[21]}}, {6{maskForGroupWire[20]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_lo_hi_hi_5 = {{6{maskForGroupWire[23]}}, {6{maskForGroupWire[22]}}};
  wire [23:0]       fillBySeg_lo_lo_hi_lo_hi_5 = {fillBySeg_lo_lo_hi_lo_hi_hi_5, fillBySeg_lo_lo_hi_lo_hi_lo_5};
  wire [47:0]       fillBySeg_lo_lo_hi_lo_5 = {fillBySeg_lo_lo_hi_lo_hi_5, fillBySeg_lo_lo_hi_lo_lo_5};
  wire [11:0]       fillBySeg_lo_lo_hi_hi_lo_lo_5 = {{6{maskForGroupWire[25]}}, {6{maskForGroupWire[24]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_hi_lo_hi_5 = {{6{maskForGroupWire[27]}}, {6{maskForGroupWire[26]}}};
  wire [23:0]       fillBySeg_lo_lo_hi_hi_lo_5 = {fillBySeg_lo_lo_hi_hi_lo_hi_5, fillBySeg_lo_lo_hi_hi_lo_lo_5};
  wire [11:0]       fillBySeg_lo_lo_hi_hi_hi_lo_5 = {{6{maskForGroupWire[29]}}, {6{maskForGroupWire[28]}}};
  wire [11:0]       fillBySeg_lo_lo_hi_hi_hi_hi_5 = {{6{maskForGroupWire[31]}}, {6{maskForGroupWire[30]}}};
  wire [23:0]       fillBySeg_lo_lo_hi_hi_hi_5 = {fillBySeg_lo_lo_hi_hi_hi_hi_5, fillBySeg_lo_lo_hi_hi_hi_lo_5};
  wire [47:0]       fillBySeg_lo_lo_hi_hi_5 = {fillBySeg_lo_lo_hi_hi_hi_5, fillBySeg_lo_lo_hi_hi_lo_5};
  wire [95:0]       fillBySeg_lo_lo_hi_5 = {fillBySeg_lo_lo_hi_hi_5, fillBySeg_lo_lo_hi_lo_5};
  wire [191:0]      fillBySeg_lo_lo_5 = {fillBySeg_lo_lo_hi_5, fillBySeg_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_lo_lo_lo_lo_5 = {{6{maskForGroupWire[33]}}, {6{maskForGroupWire[32]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_lo_lo_hi_5 = {{6{maskForGroupWire[35]}}, {6{maskForGroupWire[34]}}};
  wire [23:0]       fillBySeg_lo_hi_lo_lo_lo_5 = {fillBySeg_lo_hi_lo_lo_lo_hi_5, fillBySeg_lo_hi_lo_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_lo_lo_hi_lo_5 = {{6{maskForGroupWire[37]}}, {6{maskForGroupWire[36]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_lo_hi_hi_5 = {{6{maskForGroupWire[39]}}, {6{maskForGroupWire[38]}}};
  wire [23:0]       fillBySeg_lo_hi_lo_lo_hi_5 = {fillBySeg_lo_hi_lo_lo_hi_hi_5, fillBySeg_lo_hi_lo_lo_hi_lo_5};
  wire [47:0]       fillBySeg_lo_hi_lo_lo_5 = {fillBySeg_lo_hi_lo_lo_hi_5, fillBySeg_lo_hi_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_lo_hi_lo_lo_5 = {{6{maskForGroupWire[41]}}, {6{maskForGroupWire[40]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_hi_lo_hi_5 = {{6{maskForGroupWire[43]}}, {6{maskForGroupWire[42]}}};
  wire [23:0]       fillBySeg_lo_hi_lo_hi_lo_5 = {fillBySeg_lo_hi_lo_hi_lo_hi_5, fillBySeg_lo_hi_lo_hi_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_lo_hi_hi_lo_5 = {{6{maskForGroupWire[45]}}, {6{maskForGroupWire[44]}}};
  wire [11:0]       fillBySeg_lo_hi_lo_hi_hi_hi_5 = {{6{maskForGroupWire[47]}}, {6{maskForGroupWire[46]}}};
  wire [23:0]       fillBySeg_lo_hi_lo_hi_hi_5 = {fillBySeg_lo_hi_lo_hi_hi_hi_5, fillBySeg_lo_hi_lo_hi_hi_lo_5};
  wire [47:0]       fillBySeg_lo_hi_lo_hi_5 = {fillBySeg_lo_hi_lo_hi_hi_5, fillBySeg_lo_hi_lo_hi_lo_5};
  wire [95:0]       fillBySeg_lo_hi_lo_5 = {fillBySeg_lo_hi_lo_hi_5, fillBySeg_lo_hi_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_hi_lo_lo_lo_5 = {{6{maskForGroupWire[49]}}, {6{maskForGroupWire[48]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_lo_lo_hi_5 = {{6{maskForGroupWire[51]}}, {6{maskForGroupWire[50]}}};
  wire [23:0]       fillBySeg_lo_hi_hi_lo_lo_5 = {fillBySeg_lo_hi_hi_lo_lo_hi_5, fillBySeg_lo_hi_hi_lo_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_hi_lo_hi_lo_5 = {{6{maskForGroupWire[53]}}, {6{maskForGroupWire[52]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_lo_hi_hi_5 = {{6{maskForGroupWire[55]}}, {6{maskForGroupWire[54]}}};
  wire [23:0]       fillBySeg_lo_hi_hi_lo_hi_5 = {fillBySeg_lo_hi_hi_lo_hi_hi_5, fillBySeg_lo_hi_hi_lo_hi_lo_5};
  wire [47:0]       fillBySeg_lo_hi_hi_lo_5 = {fillBySeg_lo_hi_hi_lo_hi_5, fillBySeg_lo_hi_hi_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_hi_hi_lo_lo_5 = {{6{maskForGroupWire[57]}}, {6{maskForGroupWire[56]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_hi_lo_hi_5 = {{6{maskForGroupWire[59]}}, {6{maskForGroupWire[58]}}};
  wire [23:0]       fillBySeg_lo_hi_hi_hi_lo_5 = {fillBySeg_lo_hi_hi_hi_lo_hi_5, fillBySeg_lo_hi_hi_hi_lo_lo_5};
  wire [11:0]       fillBySeg_lo_hi_hi_hi_hi_lo_5 = {{6{maskForGroupWire[61]}}, {6{maskForGroupWire[60]}}};
  wire [11:0]       fillBySeg_lo_hi_hi_hi_hi_hi_5 = {{6{maskForGroupWire[63]}}, {6{maskForGroupWire[62]}}};
  wire [23:0]       fillBySeg_lo_hi_hi_hi_hi_5 = {fillBySeg_lo_hi_hi_hi_hi_hi_5, fillBySeg_lo_hi_hi_hi_hi_lo_5};
  wire [47:0]       fillBySeg_lo_hi_hi_hi_5 = {fillBySeg_lo_hi_hi_hi_hi_5, fillBySeg_lo_hi_hi_hi_lo_5};
  wire [95:0]       fillBySeg_lo_hi_hi_5 = {fillBySeg_lo_hi_hi_hi_5, fillBySeg_lo_hi_hi_lo_5};
  wire [191:0]      fillBySeg_lo_hi_5 = {fillBySeg_lo_hi_hi_5, fillBySeg_lo_hi_lo_5};
  wire [383:0]      fillBySeg_lo_5 = {fillBySeg_lo_hi_5, fillBySeg_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_lo_lo_lo_lo_5 = {{6{maskForGroupWire[65]}}, {6{maskForGroupWire[64]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_lo_lo_hi_5 = {{6{maskForGroupWire[67]}}, {6{maskForGroupWire[66]}}};
  wire [23:0]       fillBySeg_hi_lo_lo_lo_lo_5 = {fillBySeg_hi_lo_lo_lo_lo_hi_5, fillBySeg_hi_lo_lo_lo_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_lo_lo_hi_lo_5 = {{6{maskForGroupWire[69]}}, {6{maskForGroupWire[68]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_lo_hi_hi_5 = {{6{maskForGroupWire[71]}}, {6{maskForGroupWire[70]}}};
  wire [23:0]       fillBySeg_hi_lo_lo_lo_hi_5 = {fillBySeg_hi_lo_lo_lo_hi_hi_5, fillBySeg_hi_lo_lo_lo_hi_lo_5};
  wire [47:0]       fillBySeg_hi_lo_lo_lo_5 = {fillBySeg_hi_lo_lo_lo_hi_5, fillBySeg_hi_lo_lo_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_lo_hi_lo_lo_5 = {{6{maskForGroupWire[73]}}, {6{maskForGroupWire[72]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_hi_lo_hi_5 = {{6{maskForGroupWire[75]}}, {6{maskForGroupWire[74]}}};
  wire [23:0]       fillBySeg_hi_lo_lo_hi_lo_5 = {fillBySeg_hi_lo_lo_hi_lo_hi_5, fillBySeg_hi_lo_lo_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_lo_hi_hi_lo_5 = {{6{maskForGroupWire[77]}}, {6{maskForGroupWire[76]}}};
  wire [11:0]       fillBySeg_hi_lo_lo_hi_hi_hi_5 = {{6{maskForGroupWire[79]}}, {6{maskForGroupWire[78]}}};
  wire [23:0]       fillBySeg_hi_lo_lo_hi_hi_5 = {fillBySeg_hi_lo_lo_hi_hi_hi_5, fillBySeg_hi_lo_lo_hi_hi_lo_5};
  wire [47:0]       fillBySeg_hi_lo_lo_hi_5 = {fillBySeg_hi_lo_lo_hi_hi_5, fillBySeg_hi_lo_lo_hi_lo_5};
  wire [95:0]       fillBySeg_hi_lo_lo_5 = {fillBySeg_hi_lo_lo_hi_5, fillBySeg_hi_lo_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_hi_lo_lo_lo_5 = {{6{maskForGroupWire[81]}}, {6{maskForGroupWire[80]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_lo_lo_hi_5 = {{6{maskForGroupWire[83]}}, {6{maskForGroupWire[82]}}};
  wire [23:0]       fillBySeg_hi_lo_hi_lo_lo_5 = {fillBySeg_hi_lo_hi_lo_lo_hi_5, fillBySeg_hi_lo_hi_lo_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_hi_lo_hi_lo_5 = {{6{maskForGroupWire[85]}}, {6{maskForGroupWire[84]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_lo_hi_hi_5 = {{6{maskForGroupWire[87]}}, {6{maskForGroupWire[86]}}};
  wire [23:0]       fillBySeg_hi_lo_hi_lo_hi_5 = {fillBySeg_hi_lo_hi_lo_hi_hi_5, fillBySeg_hi_lo_hi_lo_hi_lo_5};
  wire [47:0]       fillBySeg_hi_lo_hi_lo_5 = {fillBySeg_hi_lo_hi_lo_hi_5, fillBySeg_hi_lo_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_hi_hi_lo_lo_5 = {{6{maskForGroupWire[89]}}, {6{maskForGroupWire[88]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_hi_lo_hi_5 = {{6{maskForGroupWire[91]}}, {6{maskForGroupWire[90]}}};
  wire [23:0]       fillBySeg_hi_lo_hi_hi_lo_5 = {fillBySeg_hi_lo_hi_hi_lo_hi_5, fillBySeg_hi_lo_hi_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_lo_hi_hi_hi_lo_5 = {{6{maskForGroupWire[93]}}, {6{maskForGroupWire[92]}}};
  wire [11:0]       fillBySeg_hi_lo_hi_hi_hi_hi_5 = {{6{maskForGroupWire[95]}}, {6{maskForGroupWire[94]}}};
  wire [23:0]       fillBySeg_hi_lo_hi_hi_hi_5 = {fillBySeg_hi_lo_hi_hi_hi_hi_5, fillBySeg_hi_lo_hi_hi_hi_lo_5};
  wire [47:0]       fillBySeg_hi_lo_hi_hi_5 = {fillBySeg_hi_lo_hi_hi_hi_5, fillBySeg_hi_lo_hi_hi_lo_5};
  wire [95:0]       fillBySeg_hi_lo_hi_5 = {fillBySeg_hi_lo_hi_hi_5, fillBySeg_hi_lo_hi_lo_5};
  wire [191:0]      fillBySeg_hi_lo_5 = {fillBySeg_hi_lo_hi_5, fillBySeg_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_lo_lo_lo_lo_5 = {{6{maskForGroupWire[97]}}, {6{maskForGroupWire[96]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_lo_lo_hi_5 = {{6{maskForGroupWire[99]}}, {6{maskForGroupWire[98]}}};
  wire [23:0]       fillBySeg_hi_hi_lo_lo_lo_5 = {fillBySeg_hi_hi_lo_lo_lo_hi_5, fillBySeg_hi_hi_lo_lo_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_lo_lo_hi_lo_5 = {{6{maskForGroupWire[101]}}, {6{maskForGroupWire[100]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_lo_hi_hi_5 = {{6{maskForGroupWire[103]}}, {6{maskForGroupWire[102]}}};
  wire [23:0]       fillBySeg_hi_hi_lo_lo_hi_5 = {fillBySeg_hi_hi_lo_lo_hi_hi_5, fillBySeg_hi_hi_lo_lo_hi_lo_5};
  wire [47:0]       fillBySeg_hi_hi_lo_lo_5 = {fillBySeg_hi_hi_lo_lo_hi_5, fillBySeg_hi_hi_lo_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_lo_hi_lo_lo_5 = {{6{maskForGroupWire[105]}}, {6{maskForGroupWire[104]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_hi_lo_hi_5 = {{6{maskForGroupWire[107]}}, {6{maskForGroupWire[106]}}};
  wire [23:0]       fillBySeg_hi_hi_lo_hi_lo_5 = {fillBySeg_hi_hi_lo_hi_lo_hi_5, fillBySeg_hi_hi_lo_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_lo_hi_hi_lo_5 = {{6{maskForGroupWire[109]}}, {6{maskForGroupWire[108]}}};
  wire [11:0]       fillBySeg_hi_hi_lo_hi_hi_hi_5 = {{6{maskForGroupWire[111]}}, {6{maskForGroupWire[110]}}};
  wire [23:0]       fillBySeg_hi_hi_lo_hi_hi_5 = {fillBySeg_hi_hi_lo_hi_hi_hi_5, fillBySeg_hi_hi_lo_hi_hi_lo_5};
  wire [47:0]       fillBySeg_hi_hi_lo_hi_5 = {fillBySeg_hi_hi_lo_hi_hi_5, fillBySeg_hi_hi_lo_hi_lo_5};
  wire [95:0]       fillBySeg_hi_hi_lo_5 = {fillBySeg_hi_hi_lo_hi_5, fillBySeg_hi_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_hi_lo_lo_lo_5 = {{6{maskForGroupWire[113]}}, {6{maskForGroupWire[112]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_lo_lo_hi_5 = {{6{maskForGroupWire[115]}}, {6{maskForGroupWire[114]}}};
  wire [23:0]       fillBySeg_hi_hi_hi_lo_lo_5 = {fillBySeg_hi_hi_hi_lo_lo_hi_5, fillBySeg_hi_hi_hi_lo_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_hi_lo_hi_lo_5 = {{6{maskForGroupWire[117]}}, {6{maskForGroupWire[116]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_lo_hi_hi_5 = {{6{maskForGroupWire[119]}}, {6{maskForGroupWire[118]}}};
  wire [23:0]       fillBySeg_hi_hi_hi_lo_hi_5 = {fillBySeg_hi_hi_hi_lo_hi_hi_5, fillBySeg_hi_hi_hi_lo_hi_lo_5};
  wire [47:0]       fillBySeg_hi_hi_hi_lo_5 = {fillBySeg_hi_hi_hi_lo_hi_5, fillBySeg_hi_hi_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_hi_hi_lo_lo_5 = {{6{maskForGroupWire[121]}}, {6{maskForGroupWire[120]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_hi_lo_hi_5 = {{6{maskForGroupWire[123]}}, {6{maskForGroupWire[122]}}};
  wire [23:0]       fillBySeg_hi_hi_hi_hi_lo_5 = {fillBySeg_hi_hi_hi_hi_lo_hi_5, fillBySeg_hi_hi_hi_hi_lo_lo_5};
  wire [11:0]       fillBySeg_hi_hi_hi_hi_hi_lo_5 = {{6{maskForGroupWire[125]}}, {6{maskForGroupWire[124]}}};
  wire [11:0]       fillBySeg_hi_hi_hi_hi_hi_hi_5 = {{6{maskForGroupWire[127]}}, {6{maskForGroupWire[126]}}};
  wire [23:0]       fillBySeg_hi_hi_hi_hi_hi_5 = {fillBySeg_hi_hi_hi_hi_hi_hi_5, fillBySeg_hi_hi_hi_hi_hi_lo_5};
  wire [47:0]       fillBySeg_hi_hi_hi_hi_5 = {fillBySeg_hi_hi_hi_hi_hi_5, fillBySeg_hi_hi_hi_hi_lo_5};
  wire [95:0]       fillBySeg_hi_hi_hi_5 = {fillBySeg_hi_hi_hi_hi_5, fillBySeg_hi_hi_hi_lo_5};
  wire [191:0]      fillBySeg_hi_hi_5 = {fillBySeg_hi_hi_hi_5, fillBySeg_hi_hi_lo_5};
  wire [383:0]      fillBySeg_hi_5 = {fillBySeg_hi_hi_5, fillBySeg_hi_lo_5};
  wire [13:0]       fillBySeg_lo_lo_lo_lo_lo_lo_6 = {{7{maskForGroupWire[1]}}, {7{maskForGroupWire[0]}}};
  wire [13:0]       fillBySeg_lo_lo_lo_lo_lo_hi_6 = {{7{maskForGroupWire[3]}}, {7{maskForGroupWire[2]}}};
  wire [27:0]       fillBySeg_lo_lo_lo_lo_lo_6 = {fillBySeg_lo_lo_lo_lo_lo_hi_6, fillBySeg_lo_lo_lo_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_lo_lo_lo_hi_lo_6 = {{7{maskForGroupWire[5]}}, {7{maskForGroupWire[4]}}};
  wire [13:0]       fillBySeg_lo_lo_lo_lo_hi_hi_6 = {{7{maskForGroupWire[7]}}, {7{maskForGroupWire[6]}}};
  wire [27:0]       fillBySeg_lo_lo_lo_lo_hi_6 = {fillBySeg_lo_lo_lo_lo_hi_hi_6, fillBySeg_lo_lo_lo_lo_hi_lo_6};
  wire [55:0]       fillBySeg_lo_lo_lo_lo_6 = {fillBySeg_lo_lo_lo_lo_hi_6, fillBySeg_lo_lo_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_lo_lo_hi_lo_lo_6 = {{7{maskForGroupWire[9]}}, {7{maskForGroupWire[8]}}};
  wire [13:0]       fillBySeg_lo_lo_lo_hi_lo_hi_6 = {{7{maskForGroupWire[11]}}, {7{maskForGroupWire[10]}}};
  wire [27:0]       fillBySeg_lo_lo_lo_hi_lo_6 = {fillBySeg_lo_lo_lo_hi_lo_hi_6, fillBySeg_lo_lo_lo_hi_lo_lo_6};
  wire [13:0]       fillBySeg_lo_lo_lo_hi_hi_lo_6 = {{7{maskForGroupWire[13]}}, {7{maskForGroupWire[12]}}};
  wire [13:0]       fillBySeg_lo_lo_lo_hi_hi_hi_6 = {{7{maskForGroupWire[15]}}, {7{maskForGroupWire[14]}}};
  wire [27:0]       fillBySeg_lo_lo_lo_hi_hi_6 = {fillBySeg_lo_lo_lo_hi_hi_hi_6, fillBySeg_lo_lo_lo_hi_hi_lo_6};
  wire [55:0]       fillBySeg_lo_lo_lo_hi_6 = {fillBySeg_lo_lo_lo_hi_hi_6, fillBySeg_lo_lo_lo_hi_lo_6};
  wire [111:0]      fillBySeg_lo_lo_lo_6 = {fillBySeg_lo_lo_lo_hi_6, fillBySeg_lo_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_lo_hi_lo_lo_lo_6 = {{7{maskForGroupWire[17]}}, {7{maskForGroupWire[16]}}};
  wire [13:0]       fillBySeg_lo_lo_hi_lo_lo_hi_6 = {{7{maskForGroupWire[19]}}, {7{maskForGroupWire[18]}}};
  wire [27:0]       fillBySeg_lo_lo_hi_lo_lo_6 = {fillBySeg_lo_lo_hi_lo_lo_hi_6, fillBySeg_lo_lo_hi_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_lo_hi_lo_hi_lo_6 = {{7{maskForGroupWire[21]}}, {7{maskForGroupWire[20]}}};
  wire [13:0]       fillBySeg_lo_lo_hi_lo_hi_hi_6 = {{7{maskForGroupWire[23]}}, {7{maskForGroupWire[22]}}};
  wire [27:0]       fillBySeg_lo_lo_hi_lo_hi_6 = {fillBySeg_lo_lo_hi_lo_hi_hi_6, fillBySeg_lo_lo_hi_lo_hi_lo_6};
  wire [55:0]       fillBySeg_lo_lo_hi_lo_6 = {fillBySeg_lo_lo_hi_lo_hi_6, fillBySeg_lo_lo_hi_lo_lo_6};
  wire [13:0]       fillBySeg_lo_lo_hi_hi_lo_lo_6 = {{7{maskForGroupWire[25]}}, {7{maskForGroupWire[24]}}};
  wire [13:0]       fillBySeg_lo_lo_hi_hi_lo_hi_6 = {{7{maskForGroupWire[27]}}, {7{maskForGroupWire[26]}}};
  wire [27:0]       fillBySeg_lo_lo_hi_hi_lo_6 = {fillBySeg_lo_lo_hi_hi_lo_hi_6, fillBySeg_lo_lo_hi_hi_lo_lo_6};
  wire [13:0]       fillBySeg_lo_lo_hi_hi_hi_lo_6 = {{7{maskForGroupWire[29]}}, {7{maskForGroupWire[28]}}};
  wire [13:0]       fillBySeg_lo_lo_hi_hi_hi_hi_6 = {{7{maskForGroupWire[31]}}, {7{maskForGroupWire[30]}}};
  wire [27:0]       fillBySeg_lo_lo_hi_hi_hi_6 = {fillBySeg_lo_lo_hi_hi_hi_hi_6, fillBySeg_lo_lo_hi_hi_hi_lo_6};
  wire [55:0]       fillBySeg_lo_lo_hi_hi_6 = {fillBySeg_lo_lo_hi_hi_hi_6, fillBySeg_lo_lo_hi_hi_lo_6};
  wire [111:0]      fillBySeg_lo_lo_hi_6 = {fillBySeg_lo_lo_hi_hi_6, fillBySeg_lo_lo_hi_lo_6};
  wire [223:0]      fillBySeg_lo_lo_6 = {fillBySeg_lo_lo_hi_6, fillBySeg_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_lo_lo_lo_lo_6 = {{7{maskForGroupWire[33]}}, {7{maskForGroupWire[32]}}};
  wire [13:0]       fillBySeg_lo_hi_lo_lo_lo_hi_6 = {{7{maskForGroupWire[35]}}, {7{maskForGroupWire[34]}}};
  wire [27:0]       fillBySeg_lo_hi_lo_lo_lo_6 = {fillBySeg_lo_hi_lo_lo_lo_hi_6, fillBySeg_lo_hi_lo_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_lo_lo_hi_lo_6 = {{7{maskForGroupWire[37]}}, {7{maskForGroupWire[36]}}};
  wire [13:0]       fillBySeg_lo_hi_lo_lo_hi_hi_6 = {{7{maskForGroupWire[39]}}, {7{maskForGroupWire[38]}}};
  wire [27:0]       fillBySeg_lo_hi_lo_lo_hi_6 = {fillBySeg_lo_hi_lo_lo_hi_hi_6, fillBySeg_lo_hi_lo_lo_hi_lo_6};
  wire [55:0]       fillBySeg_lo_hi_lo_lo_6 = {fillBySeg_lo_hi_lo_lo_hi_6, fillBySeg_lo_hi_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_lo_hi_lo_lo_6 = {{7{maskForGroupWire[41]}}, {7{maskForGroupWire[40]}}};
  wire [13:0]       fillBySeg_lo_hi_lo_hi_lo_hi_6 = {{7{maskForGroupWire[43]}}, {7{maskForGroupWire[42]}}};
  wire [27:0]       fillBySeg_lo_hi_lo_hi_lo_6 = {fillBySeg_lo_hi_lo_hi_lo_hi_6, fillBySeg_lo_hi_lo_hi_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_lo_hi_hi_lo_6 = {{7{maskForGroupWire[45]}}, {7{maskForGroupWire[44]}}};
  wire [13:0]       fillBySeg_lo_hi_lo_hi_hi_hi_6 = {{7{maskForGroupWire[47]}}, {7{maskForGroupWire[46]}}};
  wire [27:0]       fillBySeg_lo_hi_lo_hi_hi_6 = {fillBySeg_lo_hi_lo_hi_hi_hi_6, fillBySeg_lo_hi_lo_hi_hi_lo_6};
  wire [55:0]       fillBySeg_lo_hi_lo_hi_6 = {fillBySeg_lo_hi_lo_hi_hi_6, fillBySeg_lo_hi_lo_hi_lo_6};
  wire [111:0]      fillBySeg_lo_hi_lo_6 = {fillBySeg_lo_hi_lo_hi_6, fillBySeg_lo_hi_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_hi_lo_lo_lo_6 = {{7{maskForGroupWire[49]}}, {7{maskForGroupWire[48]}}};
  wire [13:0]       fillBySeg_lo_hi_hi_lo_lo_hi_6 = {{7{maskForGroupWire[51]}}, {7{maskForGroupWire[50]}}};
  wire [27:0]       fillBySeg_lo_hi_hi_lo_lo_6 = {fillBySeg_lo_hi_hi_lo_lo_hi_6, fillBySeg_lo_hi_hi_lo_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_hi_lo_hi_lo_6 = {{7{maskForGroupWire[53]}}, {7{maskForGroupWire[52]}}};
  wire [13:0]       fillBySeg_lo_hi_hi_lo_hi_hi_6 = {{7{maskForGroupWire[55]}}, {7{maskForGroupWire[54]}}};
  wire [27:0]       fillBySeg_lo_hi_hi_lo_hi_6 = {fillBySeg_lo_hi_hi_lo_hi_hi_6, fillBySeg_lo_hi_hi_lo_hi_lo_6};
  wire [55:0]       fillBySeg_lo_hi_hi_lo_6 = {fillBySeg_lo_hi_hi_lo_hi_6, fillBySeg_lo_hi_hi_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_hi_hi_lo_lo_6 = {{7{maskForGroupWire[57]}}, {7{maskForGroupWire[56]}}};
  wire [13:0]       fillBySeg_lo_hi_hi_hi_lo_hi_6 = {{7{maskForGroupWire[59]}}, {7{maskForGroupWire[58]}}};
  wire [27:0]       fillBySeg_lo_hi_hi_hi_lo_6 = {fillBySeg_lo_hi_hi_hi_lo_hi_6, fillBySeg_lo_hi_hi_hi_lo_lo_6};
  wire [13:0]       fillBySeg_lo_hi_hi_hi_hi_lo_6 = {{7{maskForGroupWire[61]}}, {7{maskForGroupWire[60]}}};
  wire [13:0]       fillBySeg_lo_hi_hi_hi_hi_hi_6 = {{7{maskForGroupWire[63]}}, {7{maskForGroupWire[62]}}};
  wire [27:0]       fillBySeg_lo_hi_hi_hi_hi_6 = {fillBySeg_lo_hi_hi_hi_hi_hi_6, fillBySeg_lo_hi_hi_hi_hi_lo_6};
  wire [55:0]       fillBySeg_lo_hi_hi_hi_6 = {fillBySeg_lo_hi_hi_hi_hi_6, fillBySeg_lo_hi_hi_hi_lo_6};
  wire [111:0]      fillBySeg_lo_hi_hi_6 = {fillBySeg_lo_hi_hi_hi_6, fillBySeg_lo_hi_hi_lo_6};
  wire [223:0]      fillBySeg_lo_hi_6 = {fillBySeg_lo_hi_hi_6, fillBySeg_lo_hi_lo_6};
  wire [447:0]      fillBySeg_lo_6 = {fillBySeg_lo_hi_6, fillBySeg_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_lo_lo_lo_lo_6 = {{7{maskForGroupWire[65]}}, {7{maskForGroupWire[64]}}};
  wire [13:0]       fillBySeg_hi_lo_lo_lo_lo_hi_6 = {{7{maskForGroupWire[67]}}, {7{maskForGroupWire[66]}}};
  wire [27:0]       fillBySeg_hi_lo_lo_lo_lo_6 = {fillBySeg_hi_lo_lo_lo_lo_hi_6, fillBySeg_hi_lo_lo_lo_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_lo_lo_hi_lo_6 = {{7{maskForGroupWire[69]}}, {7{maskForGroupWire[68]}}};
  wire [13:0]       fillBySeg_hi_lo_lo_lo_hi_hi_6 = {{7{maskForGroupWire[71]}}, {7{maskForGroupWire[70]}}};
  wire [27:0]       fillBySeg_hi_lo_lo_lo_hi_6 = {fillBySeg_hi_lo_lo_lo_hi_hi_6, fillBySeg_hi_lo_lo_lo_hi_lo_6};
  wire [55:0]       fillBySeg_hi_lo_lo_lo_6 = {fillBySeg_hi_lo_lo_lo_hi_6, fillBySeg_hi_lo_lo_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_lo_hi_lo_lo_6 = {{7{maskForGroupWire[73]}}, {7{maskForGroupWire[72]}}};
  wire [13:0]       fillBySeg_hi_lo_lo_hi_lo_hi_6 = {{7{maskForGroupWire[75]}}, {7{maskForGroupWire[74]}}};
  wire [27:0]       fillBySeg_hi_lo_lo_hi_lo_6 = {fillBySeg_hi_lo_lo_hi_lo_hi_6, fillBySeg_hi_lo_lo_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_lo_hi_hi_lo_6 = {{7{maskForGroupWire[77]}}, {7{maskForGroupWire[76]}}};
  wire [13:0]       fillBySeg_hi_lo_lo_hi_hi_hi_6 = {{7{maskForGroupWire[79]}}, {7{maskForGroupWire[78]}}};
  wire [27:0]       fillBySeg_hi_lo_lo_hi_hi_6 = {fillBySeg_hi_lo_lo_hi_hi_hi_6, fillBySeg_hi_lo_lo_hi_hi_lo_6};
  wire [55:0]       fillBySeg_hi_lo_lo_hi_6 = {fillBySeg_hi_lo_lo_hi_hi_6, fillBySeg_hi_lo_lo_hi_lo_6};
  wire [111:0]      fillBySeg_hi_lo_lo_6 = {fillBySeg_hi_lo_lo_hi_6, fillBySeg_hi_lo_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_hi_lo_lo_lo_6 = {{7{maskForGroupWire[81]}}, {7{maskForGroupWire[80]}}};
  wire [13:0]       fillBySeg_hi_lo_hi_lo_lo_hi_6 = {{7{maskForGroupWire[83]}}, {7{maskForGroupWire[82]}}};
  wire [27:0]       fillBySeg_hi_lo_hi_lo_lo_6 = {fillBySeg_hi_lo_hi_lo_lo_hi_6, fillBySeg_hi_lo_hi_lo_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_hi_lo_hi_lo_6 = {{7{maskForGroupWire[85]}}, {7{maskForGroupWire[84]}}};
  wire [13:0]       fillBySeg_hi_lo_hi_lo_hi_hi_6 = {{7{maskForGroupWire[87]}}, {7{maskForGroupWire[86]}}};
  wire [27:0]       fillBySeg_hi_lo_hi_lo_hi_6 = {fillBySeg_hi_lo_hi_lo_hi_hi_6, fillBySeg_hi_lo_hi_lo_hi_lo_6};
  wire [55:0]       fillBySeg_hi_lo_hi_lo_6 = {fillBySeg_hi_lo_hi_lo_hi_6, fillBySeg_hi_lo_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_hi_hi_lo_lo_6 = {{7{maskForGroupWire[89]}}, {7{maskForGroupWire[88]}}};
  wire [13:0]       fillBySeg_hi_lo_hi_hi_lo_hi_6 = {{7{maskForGroupWire[91]}}, {7{maskForGroupWire[90]}}};
  wire [27:0]       fillBySeg_hi_lo_hi_hi_lo_6 = {fillBySeg_hi_lo_hi_hi_lo_hi_6, fillBySeg_hi_lo_hi_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_lo_hi_hi_hi_lo_6 = {{7{maskForGroupWire[93]}}, {7{maskForGroupWire[92]}}};
  wire [13:0]       fillBySeg_hi_lo_hi_hi_hi_hi_6 = {{7{maskForGroupWire[95]}}, {7{maskForGroupWire[94]}}};
  wire [27:0]       fillBySeg_hi_lo_hi_hi_hi_6 = {fillBySeg_hi_lo_hi_hi_hi_hi_6, fillBySeg_hi_lo_hi_hi_hi_lo_6};
  wire [55:0]       fillBySeg_hi_lo_hi_hi_6 = {fillBySeg_hi_lo_hi_hi_hi_6, fillBySeg_hi_lo_hi_hi_lo_6};
  wire [111:0]      fillBySeg_hi_lo_hi_6 = {fillBySeg_hi_lo_hi_hi_6, fillBySeg_hi_lo_hi_lo_6};
  wire [223:0]      fillBySeg_hi_lo_6 = {fillBySeg_hi_lo_hi_6, fillBySeg_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_lo_lo_lo_lo_6 = {{7{maskForGroupWire[97]}}, {7{maskForGroupWire[96]}}};
  wire [13:0]       fillBySeg_hi_hi_lo_lo_lo_hi_6 = {{7{maskForGroupWire[99]}}, {7{maskForGroupWire[98]}}};
  wire [27:0]       fillBySeg_hi_hi_lo_lo_lo_6 = {fillBySeg_hi_hi_lo_lo_lo_hi_6, fillBySeg_hi_hi_lo_lo_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_lo_lo_hi_lo_6 = {{7{maskForGroupWire[101]}}, {7{maskForGroupWire[100]}}};
  wire [13:0]       fillBySeg_hi_hi_lo_lo_hi_hi_6 = {{7{maskForGroupWire[103]}}, {7{maskForGroupWire[102]}}};
  wire [27:0]       fillBySeg_hi_hi_lo_lo_hi_6 = {fillBySeg_hi_hi_lo_lo_hi_hi_6, fillBySeg_hi_hi_lo_lo_hi_lo_6};
  wire [55:0]       fillBySeg_hi_hi_lo_lo_6 = {fillBySeg_hi_hi_lo_lo_hi_6, fillBySeg_hi_hi_lo_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_lo_hi_lo_lo_6 = {{7{maskForGroupWire[105]}}, {7{maskForGroupWire[104]}}};
  wire [13:0]       fillBySeg_hi_hi_lo_hi_lo_hi_6 = {{7{maskForGroupWire[107]}}, {7{maskForGroupWire[106]}}};
  wire [27:0]       fillBySeg_hi_hi_lo_hi_lo_6 = {fillBySeg_hi_hi_lo_hi_lo_hi_6, fillBySeg_hi_hi_lo_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_lo_hi_hi_lo_6 = {{7{maskForGroupWire[109]}}, {7{maskForGroupWire[108]}}};
  wire [13:0]       fillBySeg_hi_hi_lo_hi_hi_hi_6 = {{7{maskForGroupWire[111]}}, {7{maskForGroupWire[110]}}};
  wire [27:0]       fillBySeg_hi_hi_lo_hi_hi_6 = {fillBySeg_hi_hi_lo_hi_hi_hi_6, fillBySeg_hi_hi_lo_hi_hi_lo_6};
  wire [55:0]       fillBySeg_hi_hi_lo_hi_6 = {fillBySeg_hi_hi_lo_hi_hi_6, fillBySeg_hi_hi_lo_hi_lo_6};
  wire [111:0]      fillBySeg_hi_hi_lo_6 = {fillBySeg_hi_hi_lo_hi_6, fillBySeg_hi_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_hi_lo_lo_lo_6 = {{7{maskForGroupWire[113]}}, {7{maskForGroupWire[112]}}};
  wire [13:0]       fillBySeg_hi_hi_hi_lo_lo_hi_6 = {{7{maskForGroupWire[115]}}, {7{maskForGroupWire[114]}}};
  wire [27:0]       fillBySeg_hi_hi_hi_lo_lo_6 = {fillBySeg_hi_hi_hi_lo_lo_hi_6, fillBySeg_hi_hi_hi_lo_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_hi_lo_hi_lo_6 = {{7{maskForGroupWire[117]}}, {7{maskForGroupWire[116]}}};
  wire [13:0]       fillBySeg_hi_hi_hi_lo_hi_hi_6 = {{7{maskForGroupWire[119]}}, {7{maskForGroupWire[118]}}};
  wire [27:0]       fillBySeg_hi_hi_hi_lo_hi_6 = {fillBySeg_hi_hi_hi_lo_hi_hi_6, fillBySeg_hi_hi_hi_lo_hi_lo_6};
  wire [55:0]       fillBySeg_hi_hi_hi_lo_6 = {fillBySeg_hi_hi_hi_lo_hi_6, fillBySeg_hi_hi_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_hi_hi_lo_lo_6 = {{7{maskForGroupWire[121]}}, {7{maskForGroupWire[120]}}};
  wire [13:0]       fillBySeg_hi_hi_hi_hi_lo_hi_6 = {{7{maskForGroupWire[123]}}, {7{maskForGroupWire[122]}}};
  wire [27:0]       fillBySeg_hi_hi_hi_hi_lo_6 = {fillBySeg_hi_hi_hi_hi_lo_hi_6, fillBySeg_hi_hi_hi_hi_lo_lo_6};
  wire [13:0]       fillBySeg_hi_hi_hi_hi_hi_lo_6 = {{7{maskForGroupWire[125]}}, {7{maskForGroupWire[124]}}};
  wire [13:0]       fillBySeg_hi_hi_hi_hi_hi_hi_6 = {{7{maskForGroupWire[127]}}, {7{maskForGroupWire[126]}}};
  wire [27:0]       fillBySeg_hi_hi_hi_hi_hi_6 = {fillBySeg_hi_hi_hi_hi_hi_hi_6, fillBySeg_hi_hi_hi_hi_hi_lo_6};
  wire [55:0]       fillBySeg_hi_hi_hi_hi_6 = {fillBySeg_hi_hi_hi_hi_hi_6, fillBySeg_hi_hi_hi_hi_lo_6};
  wire [111:0]      fillBySeg_hi_hi_hi_6 = {fillBySeg_hi_hi_hi_hi_6, fillBySeg_hi_hi_hi_lo_6};
  wire [223:0]      fillBySeg_hi_hi_6 = {fillBySeg_hi_hi_hi_6, fillBySeg_hi_hi_lo_6};
  wire [447:0]      fillBySeg_hi_6 = {fillBySeg_hi_hi_6, fillBySeg_hi_lo_6};
  wire [15:0]       fillBySeg_lo_lo_lo_lo_lo_lo_7 = {{8{maskForGroupWire[1]}}, {8{maskForGroupWire[0]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_lo_lo_hi_7 = {{8{maskForGroupWire[3]}}, {8{maskForGroupWire[2]}}};
  wire [31:0]       fillBySeg_lo_lo_lo_lo_lo_7 = {fillBySeg_lo_lo_lo_lo_lo_hi_7, fillBySeg_lo_lo_lo_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_lo_lo_lo_hi_lo_7 = {{8{maskForGroupWire[5]}}, {8{maskForGroupWire[4]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_lo_hi_hi_7 = {{8{maskForGroupWire[7]}}, {8{maskForGroupWire[6]}}};
  wire [31:0]       fillBySeg_lo_lo_lo_lo_hi_7 = {fillBySeg_lo_lo_lo_lo_hi_hi_7, fillBySeg_lo_lo_lo_lo_hi_lo_7};
  wire [63:0]       fillBySeg_lo_lo_lo_lo_7 = {fillBySeg_lo_lo_lo_lo_hi_7, fillBySeg_lo_lo_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_lo_lo_hi_lo_lo_7 = {{8{maskForGroupWire[9]}}, {8{maskForGroupWire[8]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_hi_lo_hi_7 = {{8{maskForGroupWire[11]}}, {8{maskForGroupWire[10]}}};
  wire [31:0]       fillBySeg_lo_lo_lo_hi_lo_7 = {fillBySeg_lo_lo_lo_hi_lo_hi_7, fillBySeg_lo_lo_lo_hi_lo_lo_7};
  wire [15:0]       fillBySeg_lo_lo_lo_hi_hi_lo_7 = {{8{maskForGroupWire[13]}}, {8{maskForGroupWire[12]}}};
  wire [15:0]       fillBySeg_lo_lo_lo_hi_hi_hi_7 = {{8{maskForGroupWire[15]}}, {8{maskForGroupWire[14]}}};
  wire [31:0]       fillBySeg_lo_lo_lo_hi_hi_7 = {fillBySeg_lo_lo_lo_hi_hi_hi_7, fillBySeg_lo_lo_lo_hi_hi_lo_7};
  wire [63:0]       fillBySeg_lo_lo_lo_hi_7 = {fillBySeg_lo_lo_lo_hi_hi_7, fillBySeg_lo_lo_lo_hi_lo_7};
  wire [127:0]      fillBySeg_lo_lo_lo_7 = {fillBySeg_lo_lo_lo_hi_7, fillBySeg_lo_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_lo_hi_lo_lo_lo_7 = {{8{maskForGroupWire[17]}}, {8{maskForGroupWire[16]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_lo_lo_hi_7 = {{8{maskForGroupWire[19]}}, {8{maskForGroupWire[18]}}};
  wire [31:0]       fillBySeg_lo_lo_hi_lo_lo_7 = {fillBySeg_lo_lo_hi_lo_lo_hi_7, fillBySeg_lo_lo_hi_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_lo_hi_lo_hi_lo_7 = {{8{maskForGroupWire[21]}}, {8{maskForGroupWire[20]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_lo_hi_hi_7 = {{8{maskForGroupWire[23]}}, {8{maskForGroupWire[22]}}};
  wire [31:0]       fillBySeg_lo_lo_hi_lo_hi_7 = {fillBySeg_lo_lo_hi_lo_hi_hi_7, fillBySeg_lo_lo_hi_lo_hi_lo_7};
  wire [63:0]       fillBySeg_lo_lo_hi_lo_7 = {fillBySeg_lo_lo_hi_lo_hi_7, fillBySeg_lo_lo_hi_lo_lo_7};
  wire [15:0]       fillBySeg_lo_lo_hi_hi_lo_lo_7 = {{8{maskForGroupWire[25]}}, {8{maskForGroupWire[24]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_hi_lo_hi_7 = {{8{maskForGroupWire[27]}}, {8{maskForGroupWire[26]}}};
  wire [31:0]       fillBySeg_lo_lo_hi_hi_lo_7 = {fillBySeg_lo_lo_hi_hi_lo_hi_7, fillBySeg_lo_lo_hi_hi_lo_lo_7};
  wire [15:0]       fillBySeg_lo_lo_hi_hi_hi_lo_7 = {{8{maskForGroupWire[29]}}, {8{maskForGroupWire[28]}}};
  wire [15:0]       fillBySeg_lo_lo_hi_hi_hi_hi_7 = {{8{maskForGroupWire[31]}}, {8{maskForGroupWire[30]}}};
  wire [31:0]       fillBySeg_lo_lo_hi_hi_hi_7 = {fillBySeg_lo_lo_hi_hi_hi_hi_7, fillBySeg_lo_lo_hi_hi_hi_lo_7};
  wire [63:0]       fillBySeg_lo_lo_hi_hi_7 = {fillBySeg_lo_lo_hi_hi_hi_7, fillBySeg_lo_lo_hi_hi_lo_7};
  wire [127:0]      fillBySeg_lo_lo_hi_7 = {fillBySeg_lo_lo_hi_hi_7, fillBySeg_lo_lo_hi_lo_7};
  wire [255:0]      fillBySeg_lo_lo_7 = {fillBySeg_lo_lo_hi_7, fillBySeg_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_lo_lo_lo_lo_7 = {{8{maskForGroupWire[33]}}, {8{maskForGroupWire[32]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_lo_lo_hi_7 = {{8{maskForGroupWire[35]}}, {8{maskForGroupWire[34]}}};
  wire [31:0]       fillBySeg_lo_hi_lo_lo_lo_7 = {fillBySeg_lo_hi_lo_lo_lo_hi_7, fillBySeg_lo_hi_lo_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_lo_lo_hi_lo_7 = {{8{maskForGroupWire[37]}}, {8{maskForGroupWire[36]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_lo_hi_hi_7 = {{8{maskForGroupWire[39]}}, {8{maskForGroupWire[38]}}};
  wire [31:0]       fillBySeg_lo_hi_lo_lo_hi_7 = {fillBySeg_lo_hi_lo_lo_hi_hi_7, fillBySeg_lo_hi_lo_lo_hi_lo_7};
  wire [63:0]       fillBySeg_lo_hi_lo_lo_7 = {fillBySeg_lo_hi_lo_lo_hi_7, fillBySeg_lo_hi_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_lo_hi_lo_lo_7 = {{8{maskForGroupWire[41]}}, {8{maskForGroupWire[40]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_hi_lo_hi_7 = {{8{maskForGroupWire[43]}}, {8{maskForGroupWire[42]}}};
  wire [31:0]       fillBySeg_lo_hi_lo_hi_lo_7 = {fillBySeg_lo_hi_lo_hi_lo_hi_7, fillBySeg_lo_hi_lo_hi_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_lo_hi_hi_lo_7 = {{8{maskForGroupWire[45]}}, {8{maskForGroupWire[44]}}};
  wire [15:0]       fillBySeg_lo_hi_lo_hi_hi_hi_7 = {{8{maskForGroupWire[47]}}, {8{maskForGroupWire[46]}}};
  wire [31:0]       fillBySeg_lo_hi_lo_hi_hi_7 = {fillBySeg_lo_hi_lo_hi_hi_hi_7, fillBySeg_lo_hi_lo_hi_hi_lo_7};
  wire [63:0]       fillBySeg_lo_hi_lo_hi_7 = {fillBySeg_lo_hi_lo_hi_hi_7, fillBySeg_lo_hi_lo_hi_lo_7};
  wire [127:0]      fillBySeg_lo_hi_lo_7 = {fillBySeg_lo_hi_lo_hi_7, fillBySeg_lo_hi_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_hi_lo_lo_lo_7 = {{8{maskForGroupWire[49]}}, {8{maskForGroupWire[48]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_lo_lo_hi_7 = {{8{maskForGroupWire[51]}}, {8{maskForGroupWire[50]}}};
  wire [31:0]       fillBySeg_lo_hi_hi_lo_lo_7 = {fillBySeg_lo_hi_hi_lo_lo_hi_7, fillBySeg_lo_hi_hi_lo_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_hi_lo_hi_lo_7 = {{8{maskForGroupWire[53]}}, {8{maskForGroupWire[52]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_lo_hi_hi_7 = {{8{maskForGroupWire[55]}}, {8{maskForGroupWire[54]}}};
  wire [31:0]       fillBySeg_lo_hi_hi_lo_hi_7 = {fillBySeg_lo_hi_hi_lo_hi_hi_7, fillBySeg_lo_hi_hi_lo_hi_lo_7};
  wire [63:0]       fillBySeg_lo_hi_hi_lo_7 = {fillBySeg_lo_hi_hi_lo_hi_7, fillBySeg_lo_hi_hi_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_hi_hi_lo_lo_7 = {{8{maskForGroupWire[57]}}, {8{maskForGroupWire[56]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_hi_lo_hi_7 = {{8{maskForGroupWire[59]}}, {8{maskForGroupWire[58]}}};
  wire [31:0]       fillBySeg_lo_hi_hi_hi_lo_7 = {fillBySeg_lo_hi_hi_hi_lo_hi_7, fillBySeg_lo_hi_hi_hi_lo_lo_7};
  wire [15:0]       fillBySeg_lo_hi_hi_hi_hi_lo_7 = {{8{maskForGroupWire[61]}}, {8{maskForGroupWire[60]}}};
  wire [15:0]       fillBySeg_lo_hi_hi_hi_hi_hi_7 = {{8{maskForGroupWire[63]}}, {8{maskForGroupWire[62]}}};
  wire [31:0]       fillBySeg_lo_hi_hi_hi_hi_7 = {fillBySeg_lo_hi_hi_hi_hi_hi_7, fillBySeg_lo_hi_hi_hi_hi_lo_7};
  wire [63:0]       fillBySeg_lo_hi_hi_hi_7 = {fillBySeg_lo_hi_hi_hi_hi_7, fillBySeg_lo_hi_hi_hi_lo_7};
  wire [127:0]      fillBySeg_lo_hi_hi_7 = {fillBySeg_lo_hi_hi_hi_7, fillBySeg_lo_hi_hi_lo_7};
  wire [255:0]      fillBySeg_lo_hi_7 = {fillBySeg_lo_hi_hi_7, fillBySeg_lo_hi_lo_7};
  wire [511:0]      fillBySeg_lo_7 = {fillBySeg_lo_hi_7, fillBySeg_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_lo_lo_lo_lo_7 = {{8{maskForGroupWire[65]}}, {8{maskForGroupWire[64]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_lo_lo_hi_7 = {{8{maskForGroupWire[67]}}, {8{maskForGroupWire[66]}}};
  wire [31:0]       fillBySeg_hi_lo_lo_lo_lo_7 = {fillBySeg_hi_lo_lo_lo_lo_hi_7, fillBySeg_hi_lo_lo_lo_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_lo_lo_hi_lo_7 = {{8{maskForGroupWire[69]}}, {8{maskForGroupWire[68]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_lo_hi_hi_7 = {{8{maskForGroupWire[71]}}, {8{maskForGroupWire[70]}}};
  wire [31:0]       fillBySeg_hi_lo_lo_lo_hi_7 = {fillBySeg_hi_lo_lo_lo_hi_hi_7, fillBySeg_hi_lo_lo_lo_hi_lo_7};
  wire [63:0]       fillBySeg_hi_lo_lo_lo_7 = {fillBySeg_hi_lo_lo_lo_hi_7, fillBySeg_hi_lo_lo_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_lo_hi_lo_lo_7 = {{8{maskForGroupWire[73]}}, {8{maskForGroupWire[72]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_hi_lo_hi_7 = {{8{maskForGroupWire[75]}}, {8{maskForGroupWire[74]}}};
  wire [31:0]       fillBySeg_hi_lo_lo_hi_lo_7 = {fillBySeg_hi_lo_lo_hi_lo_hi_7, fillBySeg_hi_lo_lo_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_lo_hi_hi_lo_7 = {{8{maskForGroupWire[77]}}, {8{maskForGroupWire[76]}}};
  wire [15:0]       fillBySeg_hi_lo_lo_hi_hi_hi_7 = {{8{maskForGroupWire[79]}}, {8{maskForGroupWire[78]}}};
  wire [31:0]       fillBySeg_hi_lo_lo_hi_hi_7 = {fillBySeg_hi_lo_lo_hi_hi_hi_7, fillBySeg_hi_lo_lo_hi_hi_lo_7};
  wire [63:0]       fillBySeg_hi_lo_lo_hi_7 = {fillBySeg_hi_lo_lo_hi_hi_7, fillBySeg_hi_lo_lo_hi_lo_7};
  wire [127:0]      fillBySeg_hi_lo_lo_7 = {fillBySeg_hi_lo_lo_hi_7, fillBySeg_hi_lo_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_hi_lo_lo_lo_7 = {{8{maskForGroupWire[81]}}, {8{maskForGroupWire[80]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_lo_lo_hi_7 = {{8{maskForGroupWire[83]}}, {8{maskForGroupWire[82]}}};
  wire [31:0]       fillBySeg_hi_lo_hi_lo_lo_7 = {fillBySeg_hi_lo_hi_lo_lo_hi_7, fillBySeg_hi_lo_hi_lo_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_hi_lo_hi_lo_7 = {{8{maskForGroupWire[85]}}, {8{maskForGroupWire[84]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_lo_hi_hi_7 = {{8{maskForGroupWire[87]}}, {8{maskForGroupWire[86]}}};
  wire [31:0]       fillBySeg_hi_lo_hi_lo_hi_7 = {fillBySeg_hi_lo_hi_lo_hi_hi_7, fillBySeg_hi_lo_hi_lo_hi_lo_7};
  wire [63:0]       fillBySeg_hi_lo_hi_lo_7 = {fillBySeg_hi_lo_hi_lo_hi_7, fillBySeg_hi_lo_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_hi_hi_lo_lo_7 = {{8{maskForGroupWire[89]}}, {8{maskForGroupWire[88]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_hi_lo_hi_7 = {{8{maskForGroupWire[91]}}, {8{maskForGroupWire[90]}}};
  wire [31:0]       fillBySeg_hi_lo_hi_hi_lo_7 = {fillBySeg_hi_lo_hi_hi_lo_hi_7, fillBySeg_hi_lo_hi_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_lo_hi_hi_hi_lo_7 = {{8{maskForGroupWire[93]}}, {8{maskForGroupWire[92]}}};
  wire [15:0]       fillBySeg_hi_lo_hi_hi_hi_hi_7 = {{8{maskForGroupWire[95]}}, {8{maskForGroupWire[94]}}};
  wire [31:0]       fillBySeg_hi_lo_hi_hi_hi_7 = {fillBySeg_hi_lo_hi_hi_hi_hi_7, fillBySeg_hi_lo_hi_hi_hi_lo_7};
  wire [63:0]       fillBySeg_hi_lo_hi_hi_7 = {fillBySeg_hi_lo_hi_hi_hi_7, fillBySeg_hi_lo_hi_hi_lo_7};
  wire [127:0]      fillBySeg_hi_lo_hi_7 = {fillBySeg_hi_lo_hi_hi_7, fillBySeg_hi_lo_hi_lo_7};
  wire [255:0]      fillBySeg_hi_lo_7 = {fillBySeg_hi_lo_hi_7, fillBySeg_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_lo_lo_lo_lo_7 = {{8{maskForGroupWire[97]}}, {8{maskForGroupWire[96]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_lo_lo_hi_7 = {{8{maskForGroupWire[99]}}, {8{maskForGroupWire[98]}}};
  wire [31:0]       fillBySeg_hi_hi_lo_lo_lo_7 = {fillBySeg_hi_hi_lo_lo_lo_hi_7, fillBySeg_hi_hi_lo_lo_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_lo_lo_hi_lo_7 = {{8{maskForGroupWire[101]}}, {8{maskForGroupWire[100]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_lo_hi_hi_7 = {{8{maskForGroupWire[103]}}, {8{maskForGroupWire[102]}}};
  wire [31:0]       fillBySeg_hi_hi_lo_lo_hi_7 = {fillBySeg_hi_hi_lo_lo_hi_hi_7, fillBySeg_hi_hi_lo_lo_hi_lo_7};
  wire [63:0]       fillBySeg_hi_hi_lo_lo_7 = {fillBySeg_hi_hi_lo_lo_hi_7, fillBySeg_hi_hi_lo_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_lo_hi_lo_lo_7 = {{8{maskForGroupWire[105]}}, {8{maskForGroupWire[104]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_hi_lo_hi_7 = {{8{maskForGroupWire[107]}}, {8{maskForGroupWire[106]}}};
  wire [31:0]       fillBySeg_hi_hi_lo_hi_lo_7 = {fillBySeg_hi_hi_lo_hi_lo_hi_7, fillBySeg_hi_hi_lo_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_lo_hi_hi_lo_7 = {{8{maskForGroupWire[109]}}, {8{maskForGroupWire[108]}}};
  wire [15:0]       fillBySeg_hi_hi_lo_hi_hi_hi_7 = {{8{maskForGroupWire[111]}}, {8{maskForGroupWire[110]}}};
  wire [31:0]       fillBySeg_hi_hi_lo_hi_hi_7 = {fillBySeg_hi_hi_lo_hi_hi_hi_7, fillBySeg_hi_hi_lo_hi_hi_lo_7};
  wire [63:0]       fillBySeg_hi_hi_lo_hi_7 = {fillBySeg_hi_hi_lo_hi_hi_7, fillBySeg_hi_hi_lo_hi_lo_7};
  wire [127:0]      fillBySeg_hi_hi_lo_7 = {fillBySeg_hi_hi_lo_hi_7, fillBySeg_hi_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_hi_lo_lo_lo_7 = {{8{maskForGroupWire[113]}}, {8{maskForGroupWire[112]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_lo_lo_hi_7 = {{8{maskForGroupWire[115]}}, {8{maskForGroupWire[114]}}};
  wire [31:0]       fillBySeg_hi_hi_hi_lo_lo_7 = {fillBySeg_hi_hi_hi_lo_lo_hi_7, fillBySeg_hi_hi_hi_lo_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_hi_lo_hi_lo_7 = {{8{maskForGroupWire[117]}}, {8{maskForGroupWire[116]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_lo_hi_hi_7 = {{8{maskForGroupWire[119]}}, {8{maskForGroupWire[118]}}};
  wire [31:0]       fillBySeg_hi_hi_hi_lo_hi_7 = {fillBySeg_hi_hi_hi_lo_hi_hi_7, fillBySeg_hi_hi_hi_lo_hi_lo_7};
  wire [63:0]       fillBySeg_hi_hi_hi_lo_7 = {fillBySeg_hi_hi_hi_lo_hi_7, fillBySeg_hi_hi_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_hi_hi_lo_lo_7 = {{8{maskForGroupWire[121]}}, {8{maskForGroupWire[120]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_hi_lo_hi_7 = {{8{maskForGroupWire[123]}}, {8{maskForGroupWire[122]}}};
  wire [31:0]       fillBySeg_hi_hi_hi_hi_lo_7 = {fillBySeg_hi_hi_hi_hi_lo_hi_7, fillBySeg_hi_hi_hi_hi_lo_lo_7};
  wire [15:0]       fillBySeg_hi_hi_hi_hi_hi_lo_7 = {{8{maskForGroupWire[125]}}, {8{maskForGroupWire[124]}}};
  wire [15:0]       fillBySeg_hi_hi_hi_hi_hi_hi_7 = {{8{maskForGroupWire[127]}}, {8{maskForGroupWire[126]}}};
  wire [31:0]       fillBySeg_hi_hi_hi_hi_hi_7 = {fillBySeg_hi_hi_hi_hi_hi_hi_7, fillBySeg_hi_hi_hi_hi_hi_lo_7};
  wire [63:0]       fillBySeg_hi_hi_hi_hi_7 = {fillBySeg_hi_hi_hi_hi_hi_7, fillBySeg_hi_hi_hi_hi_lo_7};
  wire [127:0]      fillBySeg_hi_hi_hi_7 = {fillBySeg_hi_hi_hi_hi_7, fillBySeg_hi_hi_hi_lo_7};
  wire [255:0]      fillBySeg_hi_hi_7 = {fillBySeg_hi_hi_hi_7, fillBySeg_hi_hi_lo_7};
  wire [511:0]      fillBySeg_hi_7 = {fillBySeg_hi_hi_7, fillBySeg_hi_lo_7};
  wire [1023:0]     fillBySeg =
    {128'h0,
     {128'h0,
      {128'h0,
       {128'h0,
        {128'h0, {128'h0, {128'h0, _fillBySeg_T[0] ? {fillBySeg_hi, fillBySeg_lo} : 128'h0} | (_fillBySeg_T[1] ? {fillBySeg_hi_1, fillBySeg_lo_1} : 256'h0)} | (_fillBySeg_T[2] ? {fillBySeg_hi_2, fillBySeg_lo_2} : 384'h0)}
          | (_fillBySeg_T[3] ? {fillBySeg_hi_3, fillBySeg_lo_3} : 512'h0)} | (_fillBySeg_T[4] ? {fillBySeg_hi_4, fillBySeg_lo_4} : 640'h0)} | (_fillBySeg_T[5] ? {fillBySeg_hi_5, fillBySeg_lo_5} : 768'h0)}
       | (_fillBySeg_T[6] ? {fillBySeg_hi_6, fillBySeg_lo_6} : 896'h0)} | (_fillBySeg_T[7] ? {fillBySeg_hi_7, fillBySeg_lo_7} : 1024'h0);
  wire [7:0]        dataRegroupBySew_0_0 = bufferStageEnqueueData_0[7:0];
  wire [7:0]        dataRegroupBySew_0_1 = bufferStageEnqueueData_0[15:8];
  wire [7:0]        dataRegroupBySew_0_2 = bufferStageEnqueueData_0[23:16];
  wire [7:0]        dataRegroupBySew_0_3 = bufferStageEnqueueData_0[31:24];
  wire [7:0]        dataRegroupBySew_0_4 = bufferStageEnqueueData_0[39:32];
  wire [7:0]        dataRegroupBySew_0_5 = bufferStageEnqueueData_0[47:40];
  wire [7:0]        dataRegroupBySew_0_6 = bufferStageEnqueueData_0[55:48];
  wire [7:0]        dataRegroupBySew_0_7 = bufferStageEnqueueData_0[63:56];
  wire [7:0]        dataRegroupBySew_0_8 = bufferStageEnqueueData_0[71:64];
  wire [7:0]        dataRegroupBySew_0_9 = bufferStageEnqueueData_0[79:72];
  wire [7:0]        dataRegroupBySew_0_10 = bufferStageEnqueueData_0[87:80];
  wire [7:0]        dataRegroupBySew_0_11 = bufferStageEnqueueData_0[95:88];
  wire [7:0]        dataRegroupBySew_0_12 = bufferStageEnqueueData_0[103:96];
  wire [7:0]        dataRegroupBySew_0_13 = bufferStageEnqueueData_0[111:104];
  wire [7:0]        dataRegroupBySew_0_14 = bufferStageEnqueueData_0[119:112];
  wire [7:0]        dataRegroupBySew_0_15 = bufferStageEnqueueData_0[127:120];
  wire [7:0]        dataRegroupBySew_0_16 = bufferStageEnqueueData_0[135:128];
  wire [7:0]        dataRegroupBySew_0_17 = bufferStageEnqueueData_0[143:136];
  wire [7:0]        dataRegroupBySew_0_18 = bufferStageEnqueueData_0[151:144];
  wire [7:0]        dataRegroupBySew_0_19 = bufferStageEnqueueData_0[159:152];
  wire [7:0]        dataRegroupBySew_0_20 = bufferStageEnqueueData_0[167:160];
  wire [7:0]        dataRegroupBySew_0_21 = bufferStageEnqueueData_0[175:168];
  wire [7:0]        dataRegroupBySew_0_22 = bufferStageEnqueueData_0[183:176];
  wire [7:0]        dataRegroupBySew_0_23 = bufferStageEnqueueData_0[191:184];
  wire [7:0]        dataRegroupBySew_0_24 = bufferStageEnqueueData_0[199:192];
  wire [7:0]        dataRegroupBySew_0_25 = bufferStageEnqueueData_0[207:200];
  wire [7:0]        dataRegroupBySew_0_26 = bufferStageEnqueueData_0[215:208];
  wire [7:0]        dataRegroupBySew_0_27 = bufferStageEnqueueData_0[223:216];
  wire [7:0]        dataRegroupBySew_0_28 = bufferStageEnqueueData_0[231:224];
  wire [7:0]        dataRegroupBySew_0_29 = bufferStageEnqueueData_0[239:232];
  wire [7:0]        dataRegroupBySew_0_30 = bufferStageEnqueueData_0[247:240];
  wire [7:0]        dataRegroupBySew_0_31 = bufferStageEnqueueData_0[255:248];
  wire [7:0]        dataRegroupBySew_0_32 = bufferStageEnqueueData_0[263:256];
  wire [7:0]        dataRegroupBySew_0_33 = bufferStageEnqueueData_0[271:264];
  wire [7:0]        dataRegroupBySew_0_34 = bufferStageEnqueueData_0[279:272];
  wire [7:0]        dataRegroupBySew_0_35 = bufferStageEnqueueData_0[287:280];
  wire [7:0]        dataRegroupBySew_0_36 = bufferStageEnqueueData_0[295:288];
  wire [7:0]        dataRegroupBySew_0_37 = bufferStageEnqueueData_0[303:296];
  wire [7:0]        dataRegroupBySew_0_38 = bufferStageEnqueueData_0[311:304];
  wire [7:0]        dataRegroupBySew_0_39 = bufferStageEnqueueData_0[319:312];
  wire [7:0]        dataRegroupBySew_0_40 = bufferStageEnqueueData_0[327:320];
  wire [7:0]        dataRegroupBySew_0_41 = bufferStageEnqueueData_0[335:328];
  wire [7:0]        dataRegroupBySew_0_42 = bufferStageEnqueueData_0[343:336];
  wire [7:0]        dataRegroupBySew_0_43 = bufferStageEnqueueData_0[351:344];
  wire [7:0]        dataRegroupBySew_0_44 = bufferStageEnqueueData_0[359:352];
  wire [7:0]        dataRegroupBySew_0_45 = bufferStageEnqueueData_0[367:360];
  wire [7:0]        dataRegroupBySew_0_46 = bufferStageEnqueueData_0[375:368];
  wire [7:0]        dataRegroupBySew_0_47 = bufferStageEnqueueData_0[383:376];
  wire [7:0]        dataRegroupBySew_0_48 = bufferStageEnqueueData_0[391:384];
  wire [7:0]        dataRegroupBySew_0_49 = bufferStageEnqueueData_0[399:392];
  wire [7:0]        dataRegroupBySew_0_50 = bufferStageEnqueueData_0[407:400];
  wire [7:0]        dataRegroupBySew_0_51 = bufferStageEnqueueData_0[415:408];
  wire [7:0]        dataRegroupBySew_0_52 = bufferStageEnqueueData_0[423:416];
  wire [7:0]        dataRegroupBySew_0_53 = bufferStageEnqueueData_0[431:424];
  wire [7:0]        dataRegroupBySew_0_54 = bufferStageEnqueueData_0[439:432];
  wire [7:0]        dataRegroupBySew_0_55 = bufferStageEnqueueData_0[447:440];
  wire [7:0]        dataRegroupBySew_0_56 = bufferStageEnqueueData_0[455:448];
  wire [7:0]        dataRegroupBySew_0_57 = bufferStageEnqueueData_0[463:456];
  wire [7:0]        dataRegroupBySew_0_58 = bufferStageEnqueueData_0[471:464];
  wire [7:0]        dataRegroupBySew_0_59 = bufferStageEnqueueData_0[479:472];
  wire [7:0]        dataRegroupBySew_0_60 = bufferStageEnqueueData_0[487:480];
  wire [7:0]        dataRegroupBySew_0_61 = bufferStageEnqueueData_0[495:488];
  wire [7:0]        dataRegroupBySew_0_62 = bufferStageEnqueueData_0[503:496];
  wire [7:0]        dataRegroupBySew_0_63 = bufferStageEnqueueData_0[511:504];
  wire [7:0]        dataRegroupBySew_0_64 = bufferStageEnqueueData_0[519:512];
  wire [7:0]        dataRegroupBySew_0_65 = bufferStageEnqueueData_0[527:520];
  wire [7:0]        dataRegroupBySew_0_66 = bufferStageEnqueueData_0[535:528];
  wire [7:0]        dataRegroupBySew_0_67 = bufferStageEnqueueData_0[543:536];
  wire [7:0]        dataRegroupBySew_0_68 = bufferStageEnqueueData_0[551:544];
  wire [7:0]        dataRegroupBySew_0_69 = bufferStageEnqueueData_0[559:552];
  wire [7:0]        dataRegroupBySew_0_70 = bufferStageEnqueueData_0[567:560];
  wire [7:0]        dataRegroupBySew_0_71 = bufferStageEnqueueData_0[575:568];
  wire [7:0]        dataRegroupBySew_0_72 = bufferStageEnqueueData_0[583:576];
  wire [7:0]        dataRegroupBySew_0_73 = bufferStageEnqueueData_0[591:584];
  wire [7:0]        dataRegroupBySew_0_74 = bufferStageEnqueueData_0[599:592];
  wire [7:0]        dataRegroupBySew_0_75 = bufferStageEnqueueData_0[607:600];
  wire [7:0]        dataRegroupBySew_0_76 = bufferStageEnqueueData_0[615:608];
  wire [7:0]        dataRegroupBySew_0_77 = bufferStageEnqueueData_0[623:616];
  wire [7:0]        dataRegroupBySew_0_78 = bufferStageEnqueueData_0[631:624];
  wire [7:0]        dataRegroupBySew_0_79 = bufferStageEnqueueData_0[639:632];
  wire [7:0]        dataRegroupBySew_0_80 = bufferStageEnqueueData_0[647:640];
  wire [7:0]        dataRegroupBySew_0_81 = bufferStageEnqueueData_0[655:648];
  wire [7:0]        dataRegroupBySew_0_82 = bufferStageEnqueueData_0[663:656];
  wire [7:0]        dataRegroupBySew_0_83 = bufferStageEnqueueData_0[671:664];
  wire [7:0]        dataRegroupBySew_0_84 = bufferStageEnqueueData_0[679:672];
  wire [7:0]        dataRegroupBySew_0_85 = bufferStageEnqueueData_0[687:680];
  wire [7:0]        dataRegroupBySew_0_86 = bufferStageEnqueueData_0[695:688];
  wire [7:0]        dataRegroupBySew_0_87 = bufferStageEnqueueData_0[703:696];
  wire [7:0]        dataRegroupBySew_0_88 = bufferStageEnqueueData_0[711:704];
  wire [7:0]        dataRegroupBySew_0_89 = bufferStageEnqueueData_0[719:712];
  wire [7:0]        dataRegroupBySew_0_90 = bufferStageEnqueueData_0[727:720];
  wire [7:0]        dataRegroupBySew_0_91 = bufferStageEnqueueData_0[735:728];
  wire [7:0]        dataRegroupBySew_0_92 = bufferStageEnqueueData_0[743:736];
  wire [7:0]        dataRegroupBySew_0_93 = bufferStageEnqueueData_0[751:744];
  wire [7:0]        dataRegroupBySew_0_94 = bufferStageEnqueueData_0[759:752];
  wire [7:0]        dataRegroupBySew_0_95 = bufferStageEnqueueData_0[767:760];
  wire [7:0]        dataRegroupBySew_0_96 = bufferStageEnqueueData_0[775:768];
  wire [7:0]        dataRegroupBySew_0_97 = bufferStageEnqueueData_0[783:776];
  wire [7:0]        dataRegroupBySew_0_98 = bufferStageEnqueueData_0[791:784];
  wire [7:0]        dataRegroupBySew_0_99 = bufferStageEnqueueData_0[799:792];
  wire [7:0]        dataRegroupBySew_0_100 = bufferStageEnqueueData_0[807:800];
  wire [7:0]        dataRegroupBySew_0_101 = bufferStageEnqueueData_0[815:808];
  wire [7:0]        dataRegroupBySew_0_102 = bufferStageEnqueueData_0[823:816];
  wire [7:0]        dataRegroupBySew_0_103 = bufferStageEnqueueData_0[831:824];
  wire [7:0]        dataRegroupBySew_0_104 = bufferStageEnqueueData_0[839:832];
  wire [7:0]        dataRegroupBySew_0_105 = bufferStageEnqueueData_0[847:840];
  wire [7:0]        dataRegroupBySew_0_106 = bufferStageEnqueueData_0[855:848];
  wire [7:0]        dataRegroupBySew_0_107 = bufferStageEnqueueData_0[863:856];
  wire [7:0]        dataRegroupBySew_0_108 = bufferStageEnqueueData_0[871:864];
  wire [7:0]        dataRegroupBySew_0_109 = bufferStageEnqueueData_0[879:872];
  wire [7:0]        dataRegroupBySew_0_110 = bufferStageEnqueueData_0[887:880];
  wire [7:0]        dataRegroupBySew_0_111 = bufferStageEnqueueData_0[895:888];
  wire [7:0]        dataRegroupBySew_0_112 = bufferStageEnqueueData_0[903:896];
  wire [7:0]        dataRegroupBySew_0_113 = bufferStageEnqueueData_0[911:904];
  wire [7:0]        dataRegroupBySew_0_114 = bufferStageEnqueueData_0[919:912];
  wire [7:0]        dataRegroupBySew_0_115 = bufferStageEnqueueData_0[927:920];
  wire [7:0]        dataRegroupBySew_0_116 = bufferStageEnqueueData_0[935:928];
  wire [7:0]        dataRegroupBySew_0_117 = bufferStageEnqueueData_0[943:936];
  wire [7:0]        dataRegroupBySew_0_118 = bufferStageEnqueueData_0[951:944];
  wire [7:0]        dataRegroupBySew_0_119 = bufferStageEnqueueData_0[959:952];
  wire [7:0]        dataRegroupBySew_0_120 = bufferStageEnqueueData_0[967:960];
  wire [7:0]        dataRegroupBySew_0_121 = bufferStageEnqueueData_0[975:968];
  wire [7:0]        dataRegroupBySew_0_122 = bufferStageEnqueueData_0[983:976];
  wire [7:0]        dataRegroupBySew_0_123 = bufferStageEnqueueData_0[991:984];
  wire [7:0]        dataRegroupBySew_0_124 = bufferStageEnqueueData_0[999:992];
  wire [7:0]        dataRegroupBySew_0_125 = bufferStageEnqueueData_0[1007:1000];
  wire [7:0]        dataRegroupBySew_0_126 = bufferStageEnqueueData_0[1015:1008];
  wire [7:0]        dataRegroupBySew_0_127 = bufferStageEnqueueData_0[1023:1016];
  wire [7:0]        dataRegroupBySew_1_0 = bufferStageEnqueueData_1[7:0];
  wire [7:0]        dataRegroupBySew_1_1 = bufferStageEnqueueData_1[15:8];
  wire [7:0]        dataRegroupBySew_1_2 = bufferStageEnqueueData_1[23:16];
  wire [7:0]        dataRegroupBySew_1_3 = bufferStageEnqueueData_1[31:24];
  wire [7:0]        dataRegroupBySew_1_4 = bufferStageEnqueueData_1[39:32];
  wire [7:0]        dataRegroupBySew_1_5 = bufferStageEnqueueData_1[47:40];
  wire [7:0]        dataRegroupBySew_1_6 = bufferStageEnqueueData_1[55:48];
  wire [7:0]        dataRegroupBySew_1_7 = bufferStageEnqueueData_1[63:56];
  wire [7:0]        dataRegroupBySew_1_8 = bufferStageEnqueueData_1[71:64];
  wire [7:0]        dataRegroupBySew_1_9 = bufferStageEnqueueData_1[79:72];
  wire [7:0]        dataRegroupBySew_1_10 = bufferStageEnqueueData_1[87:80];
  wire [7:0]        dataRegroupBySew_1_11 = bufferStageEnqueueData_1[95:88];
  wire [7:0]        dataRegroupBySew_1_12 = bufferStageEnqueueData_1[103:96];
  wire [7:0]        dataRegroupBySew_1_13 = bufferStageEnqueueData_1[111:104];
  wire [7:0]        dataRegroupBySew_1_14 = bufferStageEnqueueData_1[119:112];
  wire [7:0]        dataRegroupBySew_1_15 = bufferStageEnqueueData_1[127:120];
  wire [7:0]        dataRegroupBySew_1_16 = bufferStageEnqueueData_1[135:128];
  wire [7:0]        dataRegroupBySew_1_17 = bufferStageEnqueueData_1[143:136];
  wire [7:0]        dataRegroupBySew_1_18 = bufferStageEnqueueData_1[151:144];
  wire [7:0]        dataRegroupBySew_1_19 = bufferStageEnqueueData_1[159:152];
  wire [7:0]        dataRegroupBySew_1_20 = bufferStageEnqueueData_1[167:160];
  wire [7:0]        dataRegroupBySew_1_21 = bufferStageEnqueueData_1[175:168];
  wire [7:0]        dataRegroupBySew_1_22 = bufferStageEnqueueData_1[183:176];
  wire [7:0]        dataRegroupBySew_1_23 = bufferStageEnqueueData_1[191:184];
  wire [7:0]        dataRegroupBySew_1_24 = bufferStageEnqueueData_1[199:192];
  wire [7:0]        dataRegroupBySew_1_25 = bufferStageEnqueueData_1[207:200];
  wire [7:0]        dataRegroupBySew_1_26 = bufferStageEnqueueData_1[215:208];
  wire [7:0]        dataRegroupBySew_1_27 = bufferStageEnqueueData_1[223:216];
  wire [7:0]        dataRegroupBySew_1_28 = bufferStageEnqueueData_1[231:224];
  wire [7:0]        dataRegroupBySew_1_29 = bufferStageEnqueueData_1[239:232];
  wire [7:0]        dataRegroupBySew_1_30 = bufferStageEnqueueData_1[247:240];
  wire [7:0]        dataRegroupBySew_1_31 = bufferStageEnqueueData_1[255:248];
  wire [7:0]        dataRegroupBySew_1_32 = bufferStageEnqueueData_1[263:256];
  wire [7:0]        dataRegroupBySew_1_33 = bufferStageEnqueueData_1[271:264];
  wire [7:0]        dataRegroupBySew_1_34 = bufferStageEnqueueData_1[279:272];
  wire [7:0]        dataRegroupBySew_1_35 = bufferStageEnqueueData_1[287:280];
  wire [7:0]        dataRegroupBySew_1_36 = bufferStageEnqueueData_1[295:288];
  wire [7:0]        dataRegroupBySew_1_37 = bufferStageEnqueueData_1[303:296];
  wire [7:0]        dataRegroupBySew_1_38 = bufferStageEnqueueData_1[311:304];
  wire [7:0]        dataRegroupBySew_1_39 = bufferStageEnqueueData_1[319:312];
  wire [7:0]        dataRegroupBySew_1_40 = bufferStageEnqueueData_1[327:320];
  wire [7:0]        dataRegroupBySew_1_41 = bufferStageEnqueueData_1[335:328];
  wire [7:0]        dataRegroupBySew_1_42 = bufferStageEnqueueData_1[343:336];
  wire [7:0]        dataRegroupBySew_1_43 = bufferStageEnqueueData_1[351:344];
  wire [7:0]        dataRegroupBySew_1_44 = bufferStageEnqueueData_1[359:352];
  wire [7:0]        dataRegroupBySew_1_45 = bufferStageEnqueueData_1[367:360];
  wire [7:0]        dataRegroupBySew_1_46 = bufferStageEnqueueData_1[375:368];
  wire [7:0]        dataRegroupBySew_1_47 = bufferStageEnqueueData_1[383:376];
  wire [7:0]        dataRegroupBySew_1_48 = bufferStageEnqueueData_1[391:384];
  wire [7:0]        dataRegroupBySew_1_49 = bufferStageEnqueueData_1[399:392];
  wire [7:0]        dataRegroupBySew_1_50 = bufferStageEnqueueData_1[407:400];
  wire [7:0]        dataRegroupBySew_1_51 = bufferStageEnqueueData_1[415:408];
  wire [7:0]        dataRegroupBySew_1_52 = bufferStageEnqueueData_1[423:416];
  wire [7:0]        dataRegroupBySew_1_53 = bufferStageEnqueueData_1[431:424];
  wire [7:0]        dataRegroupBySew_1_54 = bufferStageEnqueueData_1[439:432];
  wire [7:0]        dataRegroupBySew_1_55 = bufferStageEnqueueData_1[447:440];
  wire [7:0]        dataRegroupBySew_1_56 = bufferStageEnqueueData_1[455:448];
  wire [7:0]        dataRegroupBySew_1_57 = bufferStageEnqueueData_1[463:456];
  wire [7:0]        dataRegroupBySew_1_58 = bufferStageEnqueueData_1[471:464];
  wire [7:0]        dataRegroupBySew_1_59 = bufferStageEnqueueData_1[479:472];
  wire [7:0]        dataRegroupBySew_1_60 = bufferStageEnqueueData_1[487:480];
  wire [7:0]        dataRegroupBySew_1_61 = bufferStageEnqueueData_1[495:488];
  wire [7:0]        dataRegroupBySew_1_62 = bufferStageEnqueueData_1[503:496];
  wire [7:0]        dataRegroupBySew_1_63 = bufferStageEnqueueData_1[511:504];
  wire [7:0]        dataRegroupBySew_1_64 = bufferStageEnqueueData_1[519:512];
  wire [7:0]        dataRegroupBySew_1_65 = bufferStageEnqueueData_1[527:520];
  wire [7:0]        dataRegroupBySew_1_66 = bufferStageEnqueueData_1[535:528];
  wire [7:0]        dataRegroupBySew_1_67 = bufferStageEnqueueData_1[543:536];
  wire [7:0]        dataRegroupBySew_1_68 = bufferStageEnqueueData_1[551:544];
  wire [7:0]        dataRegroupBySew_1_69 = bufferStageEnqueueData_1[559:552];
  wire [7:0]        dataRegroupBySew_1_70 = bufferStageEnqueueData_1[567:560];
  wire [7:0]        dataRegroupBySew_1_71 = bufferStageEnqueueData_1[575:568];
  wire [7:0]        dataRegroupBySew_1_72 = bufferStageEnqueueData_1[583:576];
  wire [7:0]        dataRegroupBySew_1_73 = bufferStageEnqueueData_1[591:584];
  wire [7:0]        dataRegroupBySew_1_74 = bufferStageEnqueueData_1[599:592];
  wire [7:0]        dataRegroupBySew_1_75 = bufferStageEnqueueData_1[607:600];
  wire [7:0]        dataRegroupBySew_1_76 = bufferStageEnqueueData_1[615:608];
  wire [7:0]        dataRegroupBySew_1_77 = bufferStageEnqueueData_1[623:616];
  wire [7:0]        dataRegroupBySew_1_78 = bufferStageEnqueueData_1[631:624];
  wire [7:0]        dataRegroupBySew_1_79 = bufferStageEnqueueData_1[639:632];
  wire [7:0]        dataRegroupBySew_1_80 = bufferStageEnqueueData_1[647:640];
  wire [7:0]        dataRegroupBySew_1_81 = bufferStageEnqueueData_1[655:648];
  wire [7:0]        dataRegroupBySew_1_82 = bufferStageEnqueueData_1[663:656];
  wire [7:0]        dataRegroupBySew_1_83 = bufferStageEnqueueData_1[671:664];
  wire [7:0]        dataRegroupBySew_1_84 = bufferStageEnqueueData_1[679:672];
  wire [7:0]        dataRegroupBySew_1_85 = bufferStageEnqueueData_1[687:680];
  wire [7:0]        dataRegroupBySew_1_86 = bufferStageEnqueueData_1[695:688];
  wire [7:0]        dataRegroupBySew_1_87 = bufferStageEnqueueData_1[703:696];
  wire [7:0]        dataRegroupBySew_1_88 = bufferStageEnqueueData_1[711:704];
  wire [7:0]        dataRegroupBySew_1_89 = bufferStageEnqueueData_1[719:712];
  wire [7:0]        dataRegroupBySew_1_90 = bufferStageEnqueueData_1[727:720];
  wire [7:0]        dataRegroupBySew_1_91 = bufferStageEnqueueData_1[735:728];
  wire [7:0]        dataRegroupBySew_1_92 = bufferStageEnqueueData_1[743:736];
  wire [7:0]        dataRegroupBySew_1_93 = bufferStageEnqueueData_1[751:744];
  wire [7:0]        dataRegroupBySew_1_94 = bufferStageEnqueueData_1[759:752];
  wire [7:0]        dataRegroupBySew_1_95 = bufferStageEnqueueData_1[767:760];
  wire [7:0]        dataRegroupBySew_1_96 = bufferStageEnqueueData_1[775:768];
  wire [7:0]        dataRegroupBySew_1_97 = bufferStageEnqueueData_1[783:776];
  wire [7:0]        dataRegroupBySew_1_98 = bufferStageEnqueueData_1[791:784];
  wire [7:0]        dataRegroupBySew_1_99 = bufferStageEnqueueData_1[799:792];
  wire [7:0]        dataRegroupBySew_1_100 = bufferStageEnqueueData_1[807:800];
  wire [7:0]        dataRegroupBySew_1_101 = bufferStageEnqueueData_1[815:808];
  wire [7:0]        dataRegroupBySew_1_102 = bufferStageEnqueueData_1[823:816];
  wire [7:0]        dataRegroupBySew_1_103 = bufferStageEnqueueData_1[831:824];
  wire [7:0]        dataRegroupBySew_1_104 = bufferStageEnqueueData_1[839:832];
  wire [7:0]        dataRegroupBySew_1_105 = bufferStageEnqueueData_1[847:840];
  wire [7:0]        dataRegroupBySew_1_106 = bufferStageEnqueueData_1[855:848];
  wire [7:0]        dataRegroupBySew_1_107 = bufferStageEnqueueData_1[863:856];
  wire [7:0]        dataRegroupBySew_1_108 = bufferStageEnqueueData_1[871:864];
  wire [7:0]        dataRegroupBySew_1_109 = bufferStageEnqueueData_1[879:872];
  wire [7:0]        dataRegroupBySew_1_110 = bufferStageEnqueueData_1[887:880];
  wire [7:0]        dataRegroupBySew_1_111 = bufferStageEnqueueData_1[895:888];
  wire [7:0]        dataRegroupBySew_1_112 = bufferStageEnqueueData_1[903:896];
  wire [7:0]        dataRegroupBySew_1_113 = bufferStageEnqueueData_1[911:904];
  wire [7:0]        dataRegroupBySew_1_114 = bufferStageEnqueueData_1[919:912];
  wire [7:0]        dataRegroupBySew_1_115 = bufferStageEnqueueData_1[927:920];
  wire [7:0]        dataRegroupBySew_1_116 = bufferStageEnqueueData_1[935:928];
  wire [7:0]        dataRegroupBySew_1_117 = bufferStageEnqueueData_1[943:936];
  wire [7:0]        dataRegroupBySew_1_118 = bufferStageEnqueueData_1[951:944];
  wire [7:0]        dataRegroupBySew_1_119 = bufferStageEnqueueData_1[959:952];
  wire [7:0]        dataRegroupBySew_1_120 = bufferStageEnqueueData_1[967:960];
  wire [7:0]        dataRegroupBySew_1_121 = bufferStageEnqueueData_1[975:968];
  wire [7:0]        dataRegroupBySew_1_122 = bufferStageEnqueueData_1[983:976];
  wire [7:0]        dataRegroupBySew_1_123 = bufferStageEnqueueData_1[991:984];
  wire [7:0]        dataRegroupBySew_1_124 = bufferStageEnqueueData_1[999:992];
  wire [7:0]        dataRegroupBySew_1_125 = bufferStageEnqueueData_1[1007:1000];
  wire [7:0]        dataRegroupBySew_1_126 = bufferStageEnqueueData_1[1015:1008];
  wire [7:0]        dataRegroupBySew_1_127 = bufferStageEnqueueData_1[1023:1016];
  wire [7:0]        dataRegroupBySew_2_0 = bufferStageEnqueueData_2[7:0];
  wire [7:0]        dataRegroupBySew_2_1 = bufferStageEnqueueData_2[15:8];
  wire [7:0]        dataRegroupBySew_2_2 = bufferStageEnqueueData_2[23:16];
  wire [7:0]        dataRegroupBySew_2_3 = bufferStageEnqueueData_2[31:24];
  wire [7:0]        dataRegroupBySew_2_4 = bufferStageEnqueueData_2[39:32];
  wire [7:0]        dataRegroupBySew_2_5 = bufferStageEnqueueData_2[47:40];
  wire [7:0]        dataRegroupBySew_2_6 = bufferStageEnqueueData_2[55:48];
  wire [7:0]        dataRegroupBySew_2_7 = bufferStageEnqueueData_2[63:56];
  wire [7:0]        dataRegroupBySew_2_8 = bufferStageEnqueueData_2[71:64];
  wire [7:0]        dataRegroupBySew_2_9 = bufferStageEnqueueData_2[79:72];
  wire [7:0]        dataRegroupBySew_2_10 = bufferStageEnqueueData_2[87:80];
  wire [7:0]        dataRegroupBySew_2_11 = bufferStageEnqueueData_2[95:88];
  wire [7:0]        dataRegroupBySew_2_12 = bufferStageEnqueueData_2[103:96];
  wire [7:0]        dataRegroupBySew_2_13 = bufferStageEnqueueData_2[111:104];
  wire [7:0]        dataRegroupBySew_2_14 = bufferStageEnqueueData_2[119:112];
  wire [7:0]        dataRegroupBySew_2_15 = bufferStageEnqueueData_2[127:120];
  wire [7:0]        dataRegroupBySew_2_16 = bufferStageEnqueueData_2[135:128];
  wire [7:0]        dataRegroupBySew_2_17 = bufferStageEnqueueData_2[143:136];
  wire [7:0]        dataRegroupBySew_2_18 = bufferStageEnqueueData_2[151:144];
  wire [7:0]        dataRegroupBySew_2_19 = bufferStageEnqueueData_2[159:152];
  wire [7:0]        dataRegroupBySew_2_20 = bufferStageEnqueueData_2[167:160];
  wire [7:0]        dataRegroupBySew_2_21 = bufferStageEnqueueData_2[175:168];
  wire [7:0]        dataRegroupBySew_2_22 = bufferStageEnqueueData_2[183:176];
  wire [7:0]        dataRegroupBySew_2_23 = bufferStageEnqueueData_2[191:184];
  wire [7:0]        dataRegroupBySew_2_24 = bufferStageEnqueueData_2[199:192];
  wire [7:0]        dataRegroupBySew_2_25 = bufferStageEnqueueData_2[207:200];
  wire [7:0]        dataRegroupBySew_2_26 = bufferStageEnqueueData_2[215:208];
  wire [7:0]        dataRegroupBySew_2_27 = bufferStageEnqueueData_2[223:216];
  wire [7:0]        dataRegroupBySew_2_28 = bufferStageEnqueueData_2[231:224];
  wire [7:0]        dataRegroupBySew_2_29 = bufferStageEnqueueData_2[239:232];
  wire [7:0]        dataRegroupBySew_2_30 = bufferStageEnqueueData_2[247:240];
  wire [7:0]        dataRegroupBySew_2_31 = bufferStageEnqueueData_2[255:248];
  wire [7:0]        dataRegroupBySew_2_32 = bufferStageEnqueueData_2[263:256];
  wire [7:0]        dataRegroupBySew_2_33 = bufferStageEnqueueData_2[271:264];
  wire [7:0]        dataRegroupBySew_2_34 = bufferStageEnqueueData_2[279:272];
  wire [7:0]        dataRegroupBySew_2_35 = bufferStageEnqueueData_2[287:280];
  wire [7:0]        dataRegroupBySew_2_36 = bufferStageEnqueueData_2[295:288];
  wire [7:0]        dataRegroupBySew_2_37 = bufferStageEnqueueData_2[303:296];
  wire [7:0]        dataRegroupBySew_2_38 = bufferStageEnqueueData_2[311:304];
  wire [7:0]        dataRegroupBySew_2_39 = bufferStageEnqueueData_2[319:312];
  wire [7:0]        dataRegroupBySew_2_40 = bufferStageEnqueueData_2[327:320];
  wire [7:0]        dataRegroupBySew_2_41 = bufferStageEnqueueData_2[335:328];
  wire [7:0]        dataRegroupBySew_2_42 = bufferStageEnqueueData_2[343:336];
  wire [7:0]        dataRegroupBySew_2_43 = bufferStageEnqueueData_2[351:344];
  wire [7:0]        dataRegroupBySew_2_44 = bufferStageEnqueueData_2[359:352];
  wire [7:0]        dataRegroupBySew_2_45 = bufferStageEnqueueData_2[367:360];
  wire [7:0]        dataRegroupBySew_2_46 = bufferStageEnqueueData_2[375:368];
  wire [7:0]        dataRegroupBySew_2_47 = bufferStageEnqueueData_2[383:376];
  wire [7:0]        dataRegroupBySew_2_48 = bufferStageEnqueueData_2[391:384];
  wire [7:0]        dataRegroupBySew_2_49 = bufferStageEnqueueData_2[399:392];
  wire [7:0]        dataRegroupBySew_2_50 = bufferStageEnqueueData_2[407:400];
  wire [7:0]        dataRegroupBySew_2_51 = bufferStageEnqueueData_2[415:408];
  wire [7:0]        dataRegroupBySew_2_52 = bufferStageEnqueueData_2[423:416];
  wire [7:0]        dataRegroupBySew_2_53 = bufferStageEnqueueData_2[431:424];
  wire [7:0]        dataRegroupBySew_2_54 = bufferStageEnqueueData_2[439:432];
  wire [7:0]        dataRegroupBySew_2_55 = bufferStageEnqueueData_2[447:440];
  wire [7:0]        dataRegroupBySew_2_56 = bufferStageEnqueueData_2[455:448];
  wire [7:0]        dataRegroupBySew_2_57 = bufferStageEnqueueData_2[463:456];
  wire [7:0]        dataRegroupBySew_2_58 = bufferStageEnqueueData_2[471:464];
  wire [7:0]        dataRegroupBySew_2_59 = bufferStageEnqueueData_2[479:472];
  wire [7:0]        dataRegroupBySew_2_60 = bufferStageEnqueueData_2[487:480];
  wire [7:0]        dataRegroupBySew_2_61 = bufferStageEnqueueData_2[495:488];
  wire [7:0]        dataRegroupBySew_2_62 = bufferStageEnqueueData_2[503:496];
  wire [7:0]        dataRegroupBySew_2_63 = bufferStageEnqueueData_2[511:504];
  wire [7:0]        dataRegroupBySew_2_64 = bufferStageEnqueueData_2[519:512];
  wire [7:0]        dataRegroupBySew_2_65 = bufferStageEnqueueData_2[527:520];
  wire [7:0]        dataRegroupBySew_2_66 = bufferStageEnqueueData_2[535:528];
  wire [7:0]        dataRegroupBySew_2_67 = bufferStageEnqueueData_2[543:536];
  wire [7:0]        dataRegroupBySew_2_68 = bufferStageEnqueueData_2[551:544];
  wire [7:0]        dataRegroupBySew_2_69 = bufferStageEnqueueData_2[559:552];
  wire [7:0]        dataRegroupBySew_2_70 = bufferStageEnqueueData_2[567:560];
  wire [7:0]        dataRegroupBySew_2_71 = bufferStageEnqueueData_2[575:568];
  wire [7:0]        dataRegroupBySew_2_72 = bufferStageEnqueueData_2[583:576];
  wire [7:0]        dataRegroupBySew_2_73 = bufferStageEnqueueData_2[591:584];
  wire [7:0]        dataRegroupBySew_2_74 = bufferStageEnqueueData_2[599:592];
  wire [7:0]        dataRegroupBySew_2_75 = bufferStageEnqueueData_2[607:600];
  wire [7:0]        dataRegroupBySew_2_76 = bufferStageEnqueueData_2[615:608];
  wire [7:0]        dataRegroupBySew_2_77 = bufferStageEnqueueData_2[623:616];
  wire [7:0]        dataRegroupBySew_2_78 = bufferStageEnqueueData_2[631:624];
  wire [7:0]        dataRegroupBySew_2_79 = bufferStageEnqueueData_2[639:632];
  wire [7:0]        dataRegroupBySew_2_80 = bufferStageEnqueueData_2[647:640];
  wire [7:0]        dataRegroupBySew_2_81 = bufferStageEnqueueData_2[655:648];
  wire [7:0]        dataRegroupBySew_2_82 = bufferStageEnqueueData_2[663:656];
  wire [7:0]        dataRegroupBySew_2_83 = bufferStageEnqueueData_2[671:664];
  wire [7:0]        dataRegroupBySew_2_84 = bufferStageEnqueueData_2[679:672];
  wire [7:0]        dataRegroupBySew_2_85 = bufferStageEnqueueData_2[687:680];
  wire [7:0]        dataRegroupBySew_2_86 = bufferStageEnqueueData_2[695:688];
  wire [7:0]        dataRegroupBySew_2_87 = bufferStageEnqueueData_2[703:696];
  wire [7:0]        dataRegroupBySew_2_88 = bufferStageEnqueueData_2[711:704];
  wire [7:0]        dataRegroupBySew_2_89 = bufferStageEnqueueData_2[719:712];
  wire [7:0]        dataRegroupBySew_2_90 = bufferStageEnqueueData_2[727:720];
  wire [7:0]        dataRegroupBySew_2_91 = bufferStageEnqueueData_2[735:728];
  wire [7:0]        dataRegroupBySew_2_92 = bufferStageEnqueueData_2[743:736];
  wire [7:0]        dataRegroupBySew_2_93 = bufferStageEnqueueData_2[751:744];
  wire [7:0]        dataRegroupBySew_2_94 = bufferStageEnqueueData_2[759:752];
  wire [7:0]        dataRegroupBySew_2_95 = bufferStageEnqueueData_2[767:760];
  wire [7:0]        dataRegroupBySew_2_96 = bufferStageEnqueueData_2[775:768];
  wire [7:0]        dataRegroupBySew_2_97 = bufferStageEnqueueData_2[783:776];
  wire [7:0]        dataRegroupBySew_2_98 = bufferStageEnqueueData_2[791:784];
  wire [7:0]        dataRegroupBySew_2_99 = bufferStageEnqueueData_2[799:792];
  wire [7:0]        dataRegroupBySew_2_100 = bufferStageEnqueueData_2[807:800];
  wire [7:0]        dataRegroupBySew_2_101 = bufferStageEnqueueData_2[815:808];
  wire [7:0]        dataRegroupBySew_2_102 = bufferStageEnqueueData_2[823:816];
  wire [7:0]        dataRegroupBySew_2_103 = bufferStageEnqueueData_2[831:824];
  wire [7:0]        dataRegroupBySew_2_104 = bufferStageEnqueueData_2[839:832];
  wire [7:0]        dataRegroupBySew_2_105 = bufferStageEnqueueData_2[847:840];
  wire [7:0]        dataRegroupBySew_2_106 = bufferStageEnqueueData_2[855:848];
  wire [7:0]        dataRegroupBySew_2_107 = bufferStageEnqueueData_2[863:856];
  wire [7:0]        dataRegroupBySew_2_108 = bufferStageEnqueueData_2[871:864];
  wire [7:0]        dataRegroupBySew_2_109 = bufferStageEnqueueData_2[879:872];
  wire [7:0]        dataRegroupBySew_2_110 = bufferStageEnqueueData_2[887:880];
  wire [7:0]        dataRegroupBySew_2_111 = bufferStageEnqueueData_2[895:888];
  wire [7:0]        dataRegroupBySew_2_112 = bufferStageEnqueueData_2[903:896];
  wire [7:0]        dataRegroupBySew_2_113 = bufferStageEnqueueData_2[911:904];
  wire [7:0]        dataRegroupBySew_2_114 = bufferStageEnqueueData_2[919:912];
  wire [7:0]        dataRegroupBySew_2_115 = bufferStageEnqueueData_2[927:920];
  wire [7:0]        dataRegroupBySew_2_116 = bufferStageEnqueueData_2[935:928];
  wire [7:0]        dataRegroupBySew_2_117 = bufferStageEnqueueData_2[943:936];
  wire [7:0]        dataRegroupBySew_2_118 = bufferStageEnqueueData_2[951:944];
  wire [7:0]        dataRegroupBySew_2_119 = bufferStageEnqueueData_2[959:952];
  wire [7:0]        dataRegroupBySew_2_120 = bufferStageEnqueueData_2[967:960];
  wire [7:0]        dataRegroupBySew_2_121 = bufferStageEnqueueData_2[975:968];
  wire [7:0]        dataRegroupBySew_2_122 = bufferStageEnqueueData_2[983:976];
  wire [7:0]        dataRegroupBySew_2_123 = bufferStageEnqueueData_2[991:984];
  wire [7:0]        dataRegroupBySew_2_124 = bufferStageEnqueueData_2[999:992];
  wire [7:0]        dataRegroupBySew_2_125 = bufferStageEnqueueData_2[1007:1000];
  wire [7:0]        dataRegroupBySew_2_126 = bufferStageEnqueueData_2[1015:1008];
  wire [7:0]        dataRegroupBySew_2_127 = bufferStageEnqueueData_2[1023:1016];
  wire [7:0]        dataRegroupBySew_3_0 = bufferStageEnqueueData_3[7:0];
  wire [7:0]        dataRegroupBySew_3_1 = bufferStageEnqueueData_3[15:8];
  wire [7:0]        dataRegroupBySew_3_2 = bufferStageEnqueueData_3[23:16];
  wire [7:0]        dataRegroupBySew_3_3 = bufferStageEnqueueData_3[31:24];
  wire [7:0]        dataRegroupBySew_3_4 = bufferStageEnqueueData_3[39:32];
  wire [7:0]        dataRegroupBySew_3_5 = bufferStageEnqueueData_3[47:40];
  wire [7:0]        dataRegroupBySew_3_6 = bufferStageEnqueueData_3[55:48];
  wire [7:0]        dataRegroupBySew_3_7 = bufferStageEnqueueData_3[63:56];
  wire [7:0]        dataRegroupBySew_3_8 = bufferStageEnqueueData_3[71:64];
  wire [7:0]        dataRegroupBySew_3_9 = bufferStageEnqueueData_3[79:72];
  wire [7:0]        dataRegroupBySew_3_10 = bufferStageEnqueueData_3[87:80];
  wire [7:0]        dataRegroupBySew_3_11 = bufferStageEnqueueData_3[95:88];
  wire [7:0]        dataRegroupBySew_3_12 = bufferStageEnqueueData_3[103:96];
  wire [7:0]        dataRegroupBySew_3_13 = bufferStageEnqueueData_3[111:104];
  wire [7:0]        dataRegroupBySew_3_14 = bufferStageEnqueueData_3[119:112];
  wire [7:0]        dataRegroupBySew_3_15 = bufferStageEnqueueData_3[127:120];
  wire [7:0]        dataRegroupBySew_3_16 = bufferStageEnqueueData_3[135:128];
  wire [7:0]        dataRegroupBySew_3_17 = bufferStageEnqueueData_3[143:136];
  wire [7:0]        dataRegroupBySew_3_18 = bufferStageEnqueueData_3[151:144];
  wire [7:0]        dataRegroupBySew_3_19 = bufferStageEnqueueData_3[159:152];
  wire [7:0]        dataRegroupBySew_3_20 = bufferStageEnqueueData_3[167:160];
  wire [7:0]        dataRegroupBySew_3_21 = bufferStageEnqueueData_3[175:168];
  wire [7:0]        dataRegroupBySew_3_22 = bufferStageEnqueueData_3[183:176];
  wire [7:0]        dataRegroupBySew_3_23 = bufferStageEnqueueData_3[191:184];
  wire [7:0]        dataRegroupBySew_3_24 = bufferStageEnqueueData_3[199:192];
  wire [7:0]        dataRegroupBySew_3_25 = bufferStageEnqueueData_3[207:200];
  wire [7:0]        dataRegroupBySew_3_26 = bufferStageEnqueueData_3[215:208];
  wire [7:0]        dataRegroupBySew_3_27 = bufferStageEnqueueData_3[223:216];
  wire [7:0]        dataRegroupBySew_3_28 = bufferStageEnqueueData_3[231:224];
  wire [7:0]        dataRegroupBySew_3_29 = bufferStageEnqueueData_3[239:232];
  wire [7:0]        dataRegroupBySew_3_30 = bufferStageEnqueueData_3[247:240];
  wire [7:0]        dataRegroupBySew_3_31 = bufferStageEnqueueData_3[255:248];
  wire [7:0]        dataRegroupBySew_3_32 = bufferStageEnqueueData_3[263:256];
  wire [7:0]        dataRegroupBySew_3_33 = bufferStageEnqueueData_3[271:264];
  wire [7:0]        dataRegroupBySew_3_34 = bufferStageEnqueueData_3[279:272];
  wire [7:0]        dataRegroupBySew_3_35 = bufferStageEnqueueData_3[287:280];
  wire [7:0]        dataRegroupBySew_3_36 = bufferStageEnqueueData_3[295:288];
  wire [7:0]        dataRegroupBySew_3_37 = bufferStageEnqueueData_3[303:296];
  wire [7:0]        dataRegroupBySew_3_38 = bufferStageEnqueueData_3[311:304];
  wire [7:0]        dataRegroupBySew_3_39 = bufferStageEnqueueData_3[319:312];
  wire [7:0]        dataRegroupBySew_3_40 = bufferStageEnqueueData_3[327:320];
  wire [7:0]        dataRegroupBySew_3_41 = bufferStageEnqueueData_3[335:328];
  wire [7:0]        dataRegroupBySew_3_42 = bufferStageEnqueueData_3[343:336];
  wire [7:0]        dataRegroupBySew_3_43 = bufferStageEnqueueData_3[351:344];
  wire [7:0]        dataRegroupBySew_3_44 = bufferStageEnqueueData_3[359:352];
  wire [7:0]        dataRegroupBySew_3_45 = bufferStageEnqueueData_3[367:360];
  wire [7:0]        dataRegroupBySew_3_46 = bufferStageEnqueueData_3[375:368];
  wire [7:0]        dataRegroupBySew_3_47 = bufferStageEnqueueData_3[383:376];
  wire [7:0]        dataRegroupBySew_3_48 = bufferStageEnqueueData_3[391:384];
  wire [7:0]        dataRegroupBySew_3_49 = bufferStageEnqueueData_3[399:392];
  wire [7:0]        dataRegroupBySew_3_50 = bufferStageEnqueueData_3[407:400];
  wire [7:0]        dataRegroupBySew_3_51 = bufferStageEnqueueData_3[415:408];
  wire [7:0]        dataRegroupBySew_3_52 = bufferStageEnqueueData_3[423:416];
  wire [7:0]        dataRegroupBySew_3_53 = bufferStageEnqueueData_3[431:424];
  wire [7:0]        dataRegroupBySew_3_54 = bufferStageEnqueueData_3[439:432];
  wire [7:0]        dataRegroupBySew_3_55 = bufferStageEnqueueData_3[447:440];
  wire [7:0]        dataRegroupBySew_3_56 = bufferStageEnqueueData_3[455:448];
  wire [7:0]        dataRegroupBySew_3_57 = bufferStageEnqueueData_3[463:456];
  wire [7:0]        dataRegroupBySew_3_58 = bufferStageEnqueueData_3[471:464];
  wire [7:0]        dataRegroupBySew_3_59 = bufferStageEnqueueData_3[479:472];
  wire [7:0]        dataRegroupBySew_3_60 = bufferStageEnqueueData_3[487:480];
  wire [7:0]        dataRegroupBySew_3_61 = bufferStageEnqueueData_3[495:488];
  wire [7:0]        dataRegroupBySew_3_62 = bufferStageEnqueueData_3[503:496];
  wire [7:0]        dataRegroupBySew_3_63 = bufferStageEnqueueData_3[511:504];
  wire [7:0]        dataRegroupBySew_3_64 = bufferStageEnqueueData_3[519:512];
  wire [7:0]        dataRegroupBySew_3_65 = bufferStageEnqueueData_3[527:520];
  wire [7:0]        dataRegroupBySew_3_66 = bufferStageEnqueueData_3[535:528];
  wire [7:0]        dataRegroupBySew_3_67 = bufferStageEnqueueData_3[543:536];
  wire [7:0]        dataRegroupBySew_3_68 = bufferStageEnqueueData_3[551:544];
  wire [7:0]        dataRegroupBySew_3_69 = bufferStageEnqueueData_3[559:552];
  wire [7:0]        dataRegroupBySew_3_70 = bufferStageEnqueueData_3[567:560];
  wire [7:0]        dataRegroupBySew_3_71 = bufferStageEnqueueData_3[575:568];
  wire [7:0]        dataRegroupBySew_3_72 = bufferStageEnqueueData_3[583:576];
  wire [7:0]        dataRegroupBySew_3_73 = bufferStageEnqueueData_3[591:584];
  wire [7:0]        dataRegroupBySew_3_74 = bufferStageEnqueueData_3[599:592];
  wire [7:0]        dataRegroupBySew_3_75 = bufferStageEnqueueData_3[607:600];
  wire [7:0]        dataRegroupBySew_3_76 = bufferStageEnqueueData_3[615:608];
  wire [7:0]        dataRegroupBySew_3_77 = bufferStageEnqueueData_3[623:616];
  wire [7:0]        dataRegroupBySew_3_78 = bufferStageEnqueueData_3[631:624];
  wire [7:0]        dataRegroupBySew_3_79 = bufferStageEnqueueData_3[639:632];
  wire [7:0]        dataRegroupBySew_3_80 = bufferStageEnqueueData_3[647:640];
  wire [7:0]        dataRegroupBySew_3_81 = bufferStageEnqueueData_3[655:648];
  wire [7:0]        dataRegroupBySew_3_82 = bufferStageEnqueueData_3[663:656];
  wire [7:0]        dataRegroupBySew_3_83 = bufferStageEnqueueData_3[671:664];
  wire [7:0]        dataRegroupBySew_3_84 = bufferStageEnqueueData_3[679:672];
  wire [7:0]        dataRegroupBySew_3_85 = bufferStageEnqueueData_3[687:680];
  wire [7:0]        dataRegroupBySew_3_86 = bufferStageEnqueueData_3[695:688];
  wire [7:0]        dataRegroupBySew_3_87 = bufferStageEnqueueData_3[703:696];
  wire [7:0]        dataRegroupBySew_3_88 = bufferStageEnqueueData_3[711:704];
  wire [7:0]        dataRegroupBySew_3_89 = bufferStageEnqueueData_3[719:712];
  wire [7:0]        dataRegroupBySew_3_90 = bufferStageEnqueueData_3[727:720];
  wire [7:0]        dataRegroupBySew_3_91 = bufferStageEnqueueData_3[735:728];
  wire [7:0]        dataRegroupBySew_3_92 = bufferStageEnqueueData_3[743:736];
  wire [7:0]        dataRegroupBySew_3_93 = bufferStageEnqueueData_3[751:744];
  wire [7:0]        dataRegroupBySew_3_94 = bufferStageEnqueueData_3[759:752];
  wire [7:0]        dataRegroupBySew_3_95 = bufferStageEnqueueData_3[767:760];
  wire [7:0]        dataRegroupBySew_3_96 = bufferStageEnqueueData_3[775:768];
  wire [7:0]        dataRegroupBySew_3_97 = bufferStageEnqueueData_3[783:776];
  wire [7:0]        dataRegroupBySew_3_98 = bufferStageEnqueueData_3[791:784];
  wire [7:0]        dataRegroupBySew_3_99 = bufferStageEnqueueData_3[799:792];
  wire [7:0]        dataRegroupBySew_3_100 = bufferStageEnqueueData_3[807:800];
  wire [7:0]        dataRegroupBySew_3_101 = bufferStageEnqueueData_3[815:808];
  wire [7:0]        dataRegroupBySew_3_102 = bufferStageEnqueueData_3[823:816];
  wire [7:0]        dataRegroupBySew_3_103 = bufferStageEnqueueData_3[831:824];
  wire [7:0]        dataRegroupBySew_3_104 = bufferStageEnqueueData_3[839:832];
  wire [7:0]        dataRegroupBySew_3_105 = bufferStageEnqueueData_3[847:840];
  wire [7:0]        dataRegroupBySew_3_106 = bufferStageEnqueueData_3[855:848];
  wire [7:0]        dataRegroupBySew_3_107 = bufferStageEnqueueData_3[863:856];
  wire [7:0]        dataRegroupBySew_3_108 = bufferStageEnqueueData_3[871:864];
  wire [7:0]        dataRegroupBySew_3_109 = bufferStageEnqueueData_3[879:872];
  wire [7:0]        dataRegroupBySew_3_110 = bufferStageEnqueueData_3[887:880];
  wire [7:0]        dataRegroupBySew_3_111 = bufferStageEnqueueData_3[895:888];
  wire [7:0]        dataRegroupBySew_3_112 = bufferStageEnqueueData_3[903:896];
  wire [7:0]        dataRegroupBySew_3_113 = bufferStageEnqueueData_3[911:904];
  wire [7:0]        dataRegroupBySew_3_114 = bufferStageEnqueueData_3[919:912];
  wire [7:0]        dataRegroupBySew_3_115 = bufferStageEnqueueData_3[927:920];
  wire [7:0]        dataRegroupBySew_3_116 = bufferStageEnqueueData_3[935:928];
  wire [7:0]        dataRegroupBySew_3_117 = bufferStageEnqueueData_3[943:936];
  wire [7:0]        dataRegroupBySew_3_118 = bufferStageEnqueueData_3[951:944];
  wire [7:0]        dataRegroupBySew_3_119 = bufferStageEnqueueData_3[959:952];
  wire [7:0]        dataRegroupBySew_3_120 = bufferStageEnqueueData_3[967:960];
  wire [7:0]        dataRegroupBySew_3_121 = bufferStageEnqueueData_3[975:968];
  wire [7:0]        dataRegroupBySew_3_122 = bufferStageEnqueueData_3[983:976];
  wire [7:0]        dataRegroupBySew_3_123 = bufferStageEnqueueData_3[991:984];
  wire [7:0]        dataRegroupBySew_3_124 = bufferStageEnqueueData_3[999:992];
  wire [7:0]        dataRegroupBySew_3_125 = bufferStageEnqueueData_3[1007:1000];
  wire [7:0]        dataRegroupBySew_3_126 = bufferStageEnqueueData_3[1015:1008];
  wire [7:0]        dataRegroupBySew_3_127 = bufferStageEnqueueData_3[1023:1016];
  wire [7:0]        dataRegroupBySew_4_0 = bufferStageEnqueueData_4[7:0];
  wire [7:0]        dataRegroupBySew_4_1 = bufferStageEnqueueData_4[15:8];
  wire [7:0]        dataRegroupBySew_4_2 = bufferStageEnqueueData_4[23:16];
  wire [7:0]        dataRegroupBySew_4_3 = bufferStageEnqueueData_4[31:24];
  wire [7:0]        dataRegroupBySew_4_4 = bufferStageEnqueueData_4[39:32];
  wire [7:0]        dataRegroupBySew_4_5 = bufferStageEnqueueData_4[47:40];
  wire [7:0]        dataRegroupBySew_4_6 = bufferStageEnqueueData_4[55:48];
  wire [7:0]        dataRegroupBySew_4_7 = bufferStageEnqueueData_4[63:56];
  wire [7:0]        dataRegroupBySew_4_8 = bufferStageEnqueueData_4[71:64];
  wire [7:0]        dataRegroupBySew_4_9 = bufferStageEnqueueData_4[79:72];
  wire [7:0]        dataRegroupBySew_4_10 = bufferStageEnqueueData_4[87:80];
  wire [7:0]        dataRegroupBySew_4_11 = bufferStageEnqueueData_4[95:88];
  wire [7:0]        dataRegroupBySew_4_12 = bufferStageEnqueueData_4[103:96];
  wire [7:0]        dataRegroupBySew_4_13 = bufferStageEnqueueData_4[111:104];
  wire [7:0]        dataRegroupBySew_4_14 = bufferStageEnqueueData_4[119:112];
  wire [7:0]        dataRegroupBySew_4_15 = bufferStageEnqueueData_4[127:120];
  wire [7:0]        dataRegroupBySew_4_16 = bufferStageEnqueueData_4[135:128];
  wire [7:0]        dataRegroupBySew_4_17 = bufferStageEnqueueData_4[143:136];
  wire [7:0]        dataRegroupBySew_4_18 = bufferStageEnqueueData_4[151:144];
  wire [7:0]        dataRegroupBySew_4_19 = bufferStageEnqueueData_4[159:152];
  wire [7:0]        dataRegroupBySew_4_20 = bufferStageEnqueueData_4[167:160];
  wire [7:0]        dataRegroupBySew_4_21 = bufferStageEnqueueData_4[175:168];
  wire [7:0]        dataRegroupBySew_4_22 = bufferStageEnqueueData_4[183:176];
  wire [7:0]        dataRegroupBySew_4_23 = bufferStageEnqueueData_4[191:184];
  wire [7:0]        dataRegroupBySew_4_24 = bufferStageEnqueueData_4[199:192];
  wire [7:0]        dataRegroupBySew_4_25 = bufferStageEnqueueData_4[207:200];
  wire [7:0]        dataRegroupBySew_4_26 = bufferStageEnqueueData_4[215:208];
  wire [7:0]        dataRegroupBySew_4_27 = bufferStageEnqueueData_4[223:216];
  wire [7:0]        dataRegroupBySew_4_28 = bufferStageEnqueueData_4[231:224];
  wire [7:0]        dataRegroupBySew_4_29 = bufferStageEnqueueData_4[239:232];
  wire [7:0]        dataRegroupBySew_4_30 = bufferStageEnqueueData_4[247:240];
  wire [7:0]        dataRegroupBySew_4_31 = bufferStageEnqueueData_4[255:248];
  wire [7:0]        dataRegroupBySew_4_32 = bufferStageEnqueueData_4[263:256];
  wire [7:0]        dataRegroupBySew_4_33 = bufferStageEnqueueData_4[271:264];
  wire [7:0]        dataRegroupBySew_4_34 = bufferStageEnqueueData_4[279:272];
  wire [7:0]        dataRegroupBySew_4_35 = bufferStageEnqueueData_4[287:280];
  wire [7:0]        dataRegroupBySew_4_36 = bufferStageEnqueueData_4[295:288];
  wire [7:0]        dataRegroupBySew_4_37 = bufferStageEnqueueData_4[303:296];
  wire [7:0]        dataRegroupBySew_4_38 = bufferStageEnqueueData_4[311:304];
  wire [7:0]        dataRegroupBySew_4_39 = bufferStageEnqueueData_4[319:312];
  wire [7:0]        dataRegroupBySew_4_40 = bufferStageEnqueueData_4[327:320];
  wire [7:0]        dataRegroupBySew_4_41 = bufferStageEnqueueData_4[335:328];
  wire [7:0]        dataRegroupBySew_4_42 = bufferStageEnqueueData_4[343:336];
  wire [7:0]        dataRegroupBySew_4_43 = bufferStageEnqueueData_4[351:344];
  wire [7:0]        dataRegroupBySew_4_44 = bufferStageEnqueueData_4[359:352];
  wire [7:0]        dataRegroupBySew_4_45 = bufferStageEnqueueData_4[367:360];
  wire [7:0]        dataRegroupBySew_4_46 = bufferStageEnqueueData_4[375:368];
  wire [7:0]        dataRegroupBySew_4_47 = bufferStageEnqueueData_4[383:376];
  wire [7:0]        dataRegroupBySew_4_48 = bufferStageEnqueueData_4[391:384];
  wire [7:0]        dataRegroupBySew_4_49 = bufferStageEnqueueData_4[399:392];
  wire [7:0]        dataRegroupBySew_4_50 = bufferStageEnqueueData_4[407:400];
  wire [7:0]        dataRegroupBySew_4_51 = bufferStageEnqueueData_4[415:408];
  wire [7:0]        dataRegroupBySew_4_52 = bufferStageEnqueueData_4[423:416];
  wire [7:0]        dataRegroupBySew_4_53 = bufferStageEnqueueData_4[431:424];
  wire [7:0]        dataRegroupBySew_4_54 = bufferStageEnqueueData_4[439:432];
  wire [7:0]        dataRegroupBySew_4_55 = bufferStageEnqueueData_4[447:440];
  wire [7:0]        dataRegroupBySew_4_56 = bufferStageEnqueueData_4[455:448];
  wire [7:0]        dataRegroupBySew_4_57 = bufferStageEnqueueData_4[463:456];
  wire [7:0]        dataRegroupBySew_4_58 = bufferStageEnqueueData_4[471:464];
  wire [7:0]        dataRegroupBySew_4_59 = bufferStageEnqueueData_4[479:472];
  wire [7:0]        dataRegroupBySew_4_60 = bufferStageEnqueueData_4[487:480];
  wire [7:0]        dataRegroupBySew_4_61 = bufferStageEnqueueData_4[495:488];
  wire [7:0]        dataRegroupBySew_4_62 = bufferStageEnqueueData_4[503:496];
  wire [7:0]        dataRegroupBySew_4_63 = bufferStageEnqueueData_4[511:504];
  wire [7:0]        dataRegroupBySew_4_64 = bufferStageEnqueueData_4[519:512];
  wire [7:0]        dataRegroupBySew_4_65 = bufferStageEnqueueData_4[527:520];
  wire [7:0]        dataRegroupBySew_4_66 = bufferStageEnqueueData_4[535:528];
  wire [7:0]        dataRegroupBySew_4_67 = bufferStageEnqueueData_4[543:536];
  wire [7:0]        dataRegroupBySew_4_68 = bufferStageEnqueueData_4[551:544];
  wire [7:0]        dataRegroupBySew_4_69 = bufferStageEnqueueData_4[559:552];
  wire [7:0]        dataRegroupBySew_4_70 = bufferStageEnqueueData_4[567:560];
  wire [7:0]        dataRegroupBySew_4_71 = bufferStageEnqueueData_4[575:568];
  wire [7:0]        dataRegroupBySew_4_72 = bufferStageEnqueueData_4[583:576];
  wire [7:0]        dataRegroupBySew_4_73 = bufferStageEnqueueData_4[591:584];
  wire [7:0]        dataRegroupBySew_4_74 = bufferStageEnqueueData_4[599:592];
  wire [7:0]        dataRegroupBySew_4_75 = bufferStageEnqueueData_4[607:600];
  wire [7:0]        dataRegroupBySew_4_76 = bufferStageEnqueueData_4[615:608];
  wire [7:0]        dataRegroupBySew_4_77 = bufferStageEnqueueData_4[623:616];
  wire [7:0]        dataRegroupBySew_4_78 = bufferStageEnqueueData_4[631:624];
  wire [7:0]        dataRegroupBySew_4_79 = bufferStageEnqueueData_4[639:632];
  wire [7:0]        dataRegroupBySew_4_80 = bufferStageEnqueueData_4[647:640];
  wire [7:0]        dataRegroupBySew_4_81 = bufferStageEnqueueData_4[655:648];
  wire [7:0]        dataRegroupBySew_4_82 = bufferStageEnqueueData_4[663:656];
  wire [7:0]        dataRegroupBySew_4_83 = bufferStageEnqueueData_4[671:664];
  wire [7:0]        dataRegroupBySew_4_84 = bufferStageEnqueueData_4[679:672];
  wire [7:0]        dataRegroupBySew_4_85 = bufferStageEnqueueData_4[687:680];
  wire [7:0]        dataRegroupBySew_4_86 = bufferStageEnqueueData_4[695:688];
  wire [7:0]        dataRegroupBySew_4_87 = bufferStageEnqueueData_4[703:696];
  wire [7:0]        dataRegroupBySew_4_88 = bufferStageEnqueueData_4[711:704];
  wire [7:0]        dataRegroupBySew_4_89 = bufferStageEnqueueData_4[719:712];
  wire [7:0]        dataRegroupBySew_4_90 = bufferStageEnqueueData_4[727:720];
  wire [7:0]        dataRegroupBySew_4_91 = bufferStageEnqueueData_4[735:728];
  wire [7:0]        dataRegroupBySew_4_92 = bufferStageEnqueueData_4[743:736];
  wire [7:0]        dataRegroupBySew_4_93 = bufferStageEnqueueData_4[751:744];
  wire [7:0]        dataRegroupBySew_4_94 = bufferStageEnqueueData_4[759:752];
  wire [7:0]        dataRegroupBySew_4_95 = bufferStageEnqueueData_4[767:760];
  wire [7:0]        dataRegroupBySew_4_96 = bufferStageEnqueueData_4[775:768];
  wire [7:0]        dataRegroupBySew_4_97 = bufferStageEnqueueData_4[783:776];
  wire [7:0]        dataRegroupBySew_4_98 = bufferStageEnqueueData_4[791:784];
  wire [7:0]        dataRegroupBySew_4_99 = bufferStageEnqueueData_4[799:792];
  wire [7:0]        dataRegroupBySew_4_100 = bufferStageEnqueueData_4[807:800];
  wire [7:0]        dataRegroupBySew_4_101 = bufferStageEnqueueData_4[815:808];
  wire [7:0]        dataRegroupBySew_4_102 = bufferStageEnqueueData_4[823:816];
  wire [7:0]        dataRegroupBySew_4_103 = bufferStageEnqueueData_4[831:824];
  wire [7:0]        dataRegroupBySew_4_104 = bufferStageEnqueueData_4[839:832];
  wire [7:0]        dataRegroupBySew_4_105 = bufferStageEnqueueData_4[847:840];
  wire [7:0]        dataRegroupBySew_4_106 = bufferStageEnqueueData_4[855:848];
  wire [7:0]        dataRegroupBySew_4_107 = bufferStageEnqueueData_4[863:856];
  wire [7:0]        dataRegroupBySew_4_108 = bufferStageEnqueueData_4[871:864];
  wire [7:0]        dataRegroupBySew_4_109 = bufferStageEnqueueData_4[879:872];
  wire [7:0]        dataRegroupBySew_4_110 = bufferStageEnqueueData_4[887:880];
  wire [7:0]        dataRegroupBySew_4_111 = bufferStageEnqueueData_4[895:888];
  wire [7:0]        dataRegroupBySew_4_112 = bufferStageEnqueueData_4[903:896];
  wire [7:0]        dataRegroupBySew_4_113 = bufferStageEnqueueData_4[911:904];
  wire [7:0]        dataRegroupBySew_4_114 = bufferStageEnqueueData_4[919:912];
  wire [7:0]        dataRegroupBySew_4_115 = bufferStageEnqueueData_4[927:920];
  wire [7:0]        dataRegroupBySew_4_116 = bufferStageEnqueueData_4[935:928];
  wire [7:0]        dataRegroupBySew_4_117 = bufferStageEnqueueData_4[943:936];
  wire [7:0]        dataRegroupBySew_4_118 = bufferStageEnqueueData_4[951:944];
  wire [7:0]        dataRegroupBySew_4_119 = bufferStageEnqueueData_4[959:952];
  wire [7:0]        dataRegroupBySew_4_120 = bufferStageEnqueueData_4[967:960];
  wire [7:0]        dataRegroupBySew_4_121 = bufferStageEnqueueData_4[975:968];
  wire [7:0]        dataRegroupBySew_4_122 = bufferStageEnqueueData_4[983:976];
  wire [7:0]        dataRegroupBySew_4_123 = bufferStageEnqueueData_4[991:984];
  wire [7:0]        dataRegroupBySew_4_124 = bufferStageEnqueueData_4[999:992];
  wire [7:0]        dataRegroupBySew_4_125 = bufferStageEnqueueData_4[1007:1000];
  wire [7:0]        dataRegroupBySew_4_126 = bufferStageEnqueueData_4[1015:1008];
  wire [7:0]        dataRegroupBySew_4_127 = bufferStageEnqueueData_4[1023:1016];
  wire [7:0]        dataRegroupBySew_5_0 = bufferStageEnqueueData_5[7:0];
  wire [7:0]        dataRegroupBySew_5_1 = bufferStageEnqueueData_5[15:8];
  wire [7:0]        dataRegroupBySew_5_2 = bufferStageEnqueueData_5[23:16];
  wire [7:0]        dataRegroupBySew_5_3 = bufferStageEnqueueData_5[31:24];
  wire [7:0]        dataRegroupBySew_5_4 = bufferStageEnqueueData_5[39:32];
  wire [7:0]        dataRegroupBySew_5_5 = bufferStageEnqueueData_5[47:40];
  wire [7:0]        dataRegroupBySew_5_6 = bufferStageEnqueueData_5[55:48];
  wire [7:0]        dataRegroupBySew_5_7 = bufferStageEnqueueData_5[63:56];
  wire [7:0]        dataRegroupBySew_5_8 = bufferStageEnqueueData_5[71:64];
  wire [7:0]        dataRegroupBySew_5_9 = bufferStageEnqueueData_5[79:72];
  wire [7:0]        dataRegroupBySew_5_10 = bufferStageEnqueueData_5[87:80];
  wire [7:0]        dataRegroupBySew_5_11 = bufferStageEnqueueData_5[95:88];
  wire [7:0]        dataRegroupBySew_5_12 = bufferStageEnqueueData_5[103:96];
  wire [7:0]        dataRegroupBySew_5_13 = bufferStageEnqueueData_5[111:104];
  wire [7:0]        dataRegroupBySew_5_14 = bufferStageEnqueueData_5[119:112];
  wire [7:0]        dataRegroupBySew_5_15 = bufferStageEnqueueData_5[127:120];
  wire [7:0]        dataRegroupBySew_5_16 = bufferStageEnqueueData_5[135:128];
  wire [7:0]        dataRegroupBySew_5_17 = bufferStageEnqueueData_5[143:136];
  wire [7:0]        dataRegroupBySew_5_18 = bufferStageEnqueueData_5[151:144];
  wire [7:0]        dataRegroupBySew_5_19 = bufferStageEnqueueData_5[159:152];
  wire [7:0]        dataRegroupBySew_5_20 = bufferStageEnqueueData_5[167:160];
  wire [7:0]        dataRegroupBySew_5_21 = bufferStageEnqueueData_5[175:168];
  wire [7:0]        dataRegroupBySew_5_22 = bufferStageEnqueueData_5[183:176];
  wire [7:0]        dataRegroupBySew_5_23 = bufferStageEnqueueData_5[191:184];
  wire [7:0]        dataRegroupBySew_5_24 = bufferStageEnqueueData_5[199:192];
  wire [7:0]        dataRegroupBySew_5_25 = bufferStageEnqueueData_5[207:200];
  wire [7:0]        dataRegroupBySew_5_26 = bufferStageEnqueueData_5[215:208];
  wire [7:0]        dataRegroupBySew_5_27 = bufferStageEnqueueData_5[223:216];
  wire [7:0]        dataRegroupBySew_5_28 = bufferStageEnqueueData_5[231:224];
  wire [7:0]        dataRegroupBySew_5_29 = bufferStageEnqueueData_5[239:232];
  wire [7:0]        dataRegroupBySew_5_30 = bufferStageEnqueueData_5[247:240];
  wire [7:0]        dataRegroupBySew_5_31 = bufferStageEnqueueData_5[255:248];
  wire [7:0]        dataRegroupBySew_5_32 = bufferStageEnqueueData_5[263:256];
  wire [7:0]        dataRegroupBySew_5_33 = bufferStageEnqueueData_5[271:264];
  wire [7:0]        dataRegroupBySew_5_34 = bufferStageEnqueueData_5[279:272];
  wire [7:0]        dataRegroupBySew_5_35 = bufferStageEnqueueData_5[287:280];
  wire [7:0]        dataRegroupBySew_5_36 = bufferStageEnqueueData_5[295:288];
  wire [7:0]        dataRegroupBySew_5_37 = bufferStageEnqueueData_5[303:296];
  wire [7:0]        dataRegroupBySew_5_38 = bufferStageEnqueueData_5[311:304];
  wire [7:0]        dataRegroupBySew_5_39 = bufferStageEnqueueData_5[319:312];
  wire [7:0]        dataRegroupBySew_5_40 = bufferStageEnqueueData_5[327:320];
  wire [7:0]        dataRegroupBySew_5_41 = bufferStageEnqueueData_5[335:328];
  wire [7:0]        dataRegroupBySew_5_42 = bufferStageEnqueueData_5[343:336];
  wire [7:0]        dataRegroupBySew_5_43 = bufferStageEnqueueData_5[351:344];
  wire [7:0]        dataRegroupBySew_5_44 = bufferStageEnqueueData_5[359:352];
  wire [7:0]        dataRegroupBySew_5_45 = bufferStageEnqueueData_5[367:360];
  wire [7:0]        dataRegroupBySew_5_46 = bufferStageEnqueueData_5[375:368];
  wire [7:0]        dataRegroupBySew_5_47 = bufferStageEnqueueData_5[383:376];
  wire [7:0]        dataRegroupBySew_5_48 = bufferStageEnqueueData_5[391:384];
  wire [7:0]        dataRegroupBySew_5_49 = bufferStageEnqueueData_5[399:392];
  wire [7:0]        dataRegroupBySew_5_50 = bufferStageEnqueueData_5[407:400];
  wire [7:0]        dataRegroupBySew_5_51 = bufferStageEnqueueData_5[415:408];
  wire [7:0]        dataRegroupBySew_5_52 = bufferStageEnqueueData_5[423:416];
  wire [7:0]        dataRegroupBySew_5_53 = bufferStageEnqueueData_5[431:424];
  wire [7:0]        dataRegroupBySew_5_54 = bufferStageEnqueueData_5[439:432];
  wire [7:0]        dataRegroupBySew_5_55 = bufferStageEnqueueData_5[447:440];
  wire [7:0]        dataRegroupBySew_5_56 = bufferStageEnqueueData_5[455:448];
  wire [7:0]        dataRegroupBySew_5_57 = bufferStageEnqueueData_5[463:456];
  wire [7:0]        dataRegroupBySew_5_58 = bufferStageEnqueueData_5[471:464];
  wire [7:0]        dataRegroupBySew_5_59 = bufferStageEnqueueData_5[479:472];
  wire [7:0]        dataRegroupBySew_5_60 = bufferStageEnqueueData_5[487:480];
  wire [7:0]        dataRegroupBySew_5_61 = bufferStageEnqueueData_5[495:488];
  wire [7:0]        dataRegroupBySew_5_62 = bufferStageEnqueueData_5[503:496];
  wire [7:0]        dataRegroupBySew_5_63 = bufferStageEnqueueData_5[511:504];
  wire [7:0]        dataRegroupBySew_5_64 = bufferStageEnqueueData_5[519:512];
  wire [7:0]        dataRegroupBySew_5_65 = bufferStageEnqueueData_5[527:520];
  wire [7:0]        dataRegroupBySew_5_66 = bufferStageEnqueueData_5[535:528];
  wire [7:0]        dataRegroupBySew_5_67 = bufferStageEnqueueData_5[543:536];
  wire [7:0]        dataRegroupBySew_5_68 = bufferStageEnqueueData_5[551:544];
  wire [7:0]        dataRegroupBySew_5_69 = bufferStageEnqueueData_5[559:552];
  wire [7:0]        dataRegroupBySew_5_70 = bufferStageEnqueueData_5[567:560];
  wire [7:0]        dataRegroupBySew_5_71 = bufferStageEnqueueData_5[575:568];
  wire [7:0]        dataRegroupBySew_5_72 = bufferStageEnqueueData_5[583:576];
  wire [7:0]        dataRegroupBySew_5_73 = bufferStageEnqueueData_5[591:584];
  wire [7:0]        dataRegroupBySew_5_74 = bufferStageEnqueueData_5[599:592];
  wire [7:0]        dataRegroupBySew_5_75 = bufferStageEnqueueData_5[607:600];
  wire [7:0]        dataRegroupBySew_5_76 = bufferStageEnqueueData_5[615:608];
  wire [7:0]        dataRegroupBySew_5_77 = bufferStageEnqueueData_5[623:616];
  wire [7:0]        dataRegroupBySew_5_78 = bufferStageEnqueueData_5[631:624];
  wire [7:0]        dataRegroupBySew_5_79 = bufferStageEnqueueData_5[639:632];
  wire [7:0]        dataRegroupBySew_5_80 = bufferStageEnqueueData_5[647:640];
  wire [7:0]        dataRegroupBySew_5_81 = bufferStageEnqueueData_5[655:648];
  wire [7:0]        dataRegroupBySew_5_82 = bufferStageEnqueueData_5[663:656];
  wire [7:0]        dataRegroupBySew_5_83 = bufferStageEnqueueData_5[671:664];
  wire [7:0]        dataRegroupBySew_5_84 = bufferStageEnqueueData_5[679:672];
  wire [7:0]        dataRegroupBySew_5_85 = bufferStageEnqueueData_5[687:680];
  wire [7:0]        dataRegroupBySew_5_86 = bufferStageEnqueueData_5[695:688];
  wire [7:0]        dataRegroupBySew_5_87 = bufferStageEnqueueData_5[703:696];
  wire [7:0]        dataRegroupBySew_5_88 = bufferStageEnqueueData_5[711:704];
  wire [7:0]        dataRegroupBySew_5_89 = bufferStageEnqueueData_5[719:712];
  wire [7:0]        dataRegroupBySew_5_90 = bufferStageEnqueueData_5[727:720];
  wire [7:0]        dataRegroupBySew_5_91 = bufferStageEnqueueData_5[735:728];
  wire [7:0]        dataRegroupBySew_5_92 = bufferStageEnqueueData_5[743:736];
  wire [7:0]        dataRegroupBySew_5_93 = bufferStageEnqueueData_5[751:744];
  wire [7:0]        dataRegroupBySew_5_94 = bufferStageEnqueueData_5[759:752];
  wire [7:0]        dataRegroupBySew_5_95 = bufferStageEnqueueData_5[767:760];
  wire [7:0]        dataRegroupBySew_5_96 = bufferStageEnqueueData_5[775:768];
  wire [7:0]        dataRegroupBySew_5_97 = bufferStageEnqueueData_5[783:776];
  wire [7:0]        dataRegroupBySew_5_98 = bufferStageEnqueueData_5[791:784];
  wire [7:0]        dataRegroupBySew_5_99 = bufferStageEnqueueData_5[799:792];
  wire [7:0]        dataRegroupBySew_5_100 = bufferStageEnqueueData_5[807:800];
  wire [7:0]        dataRegroupBySew_5_101 = bufferStageEnqueueData_5[815:808];
  wire [7:0]        dataRegroupBySew_5_102 = bufferStageEnqueueData_5[823:816];
  wire [7:0]        dataRegroupBySew_5_103 = bufferStageEnqueueData_5[831:824];
  wire [7:0]        dataRegroupBySew_5_104 = bufferStageEnqueueData_5[839:832];
  wire [7:0]        dataRegroupBySew_5_105 = bufferStageEnqueueData_5[847:840];
  wire [7:0]        dataRegroupBySew_5_106 = bufferStageEnqueueData_5[855:848];
  wire [7:0]        dataRegroupBySew_5_107 = bufferStageEnqueueData_5[863:856];
  wire [7:0]        dataRegroupBySew_5_108 = bufferStageEnqueueData_5[871:864];
  wire [7:0]        dataRegroupBySew_5_109 = bufferStageEnqueueData_5[879:872];
  wire [7:0]        dataRegroupBySew_5_110 = bufferStageEnqueueData_5[887:880];
  wire [7:0]        dataRegroupBySew_5_111 = bufferStageEnqueueData_5[895:888];
  wire [7:0]        dataRegroupBySew_5_112 = bufferStageEnqueueData_5[903:896];
  wire [7:0]        dataRegroupBySew_5_113 = bufferStageEnqueueData_5[911:904];
  wire [7:0]        dataRegroupBySew_5_114 = bufferStageEnqueueData_5[919:912];
  wire [7:0]        dataRegroupBySew_5_115 = bufferStageEnqueueData_5[927:920];
  wire [7:0]        dataRegroupBySew_5_116 = bufferStageEnqueueData_5[935:928];
  wire [7:0]        dataRegroupBySew_5_117 = bufferStageEnqueueData_5[943:936];
  wire [7:0]        dataRegroupBySew_5_118 = bufferStageEnqueueData_5[951:944];
  wire [7:0]        dataRegroupBySew_5_119 = bufferStageEnqueueData_5[959:952];
  wire [7:0]        dataRegroupBySew_5_120 = bufferStageEnqueueData_5[967:960];
  wire [7:0]        dataRegroupBySew_5_121 = bufferStageEnqueueData_5[975:968];
  wire [7:0]        dataRegroupBySew_5_122 = bufferStageEnqueueData_5[983:976];
  wire [7:0]        dataRegroupBySew_5_123 = bufferStageEnqueueData_5[991:984];
  wire [7:0]        dataRegroupBySew_5_124 = bufferStageEnqueueData_5[999:992];
  wire [7:0]        dataRegroupBySew_5_125 = bufferStageEnqueueData_5[1007:1000];
  wire [7:0]        dataRegroupBySew_5_126 = bufferStageEnqueueData_5[1015:1008];
  wire [7:0]        dataRegroupBySew_5_127 = bufferStageEnqueueData_5[1023:1016];
  wire [7:0]        dataRegroupBySew_6_0 = bufferStageEnqueueData_6[7:0];
  wire [7:0]        dataRegroupBySew_6_1 = bufferStageEnqueueData_6[15:8];
  wire [7:0]        dataRegroupBySew_6_2 = bufferStageEnqueueData_6[23:16];
  wire [7:0]        dataRegroupBySew_6_3 = bufferStageEnqueueData_6[31:24];
  wire [7:0]        dataRegroupBySew_6_4 = bufferStageEnqueueData_6[39:32];
  wire [7:0]        dataRegroupBySew_6_5 = bufferStageEnqueueData_6[47:40];
  wire [7:0]        dataRegroupBySew_6_6 = bufferStageEnqueueData_6[55:48];
  wire [7:0]        dataRegroupBySew_6_7 = bufferStageEnqueueData_6[63:56];
  wire [7:0]        dataRegroupBySew_6_8 = bufferStageEnqueueData_6[71:64];
  wire [7:0]        dataRegroupBySew_6_9 = bufferStageEnqueueData_6[79:72];
  wire [7:0]        dataRegroupBySew_6_10 = bufferStageEnqueueData_6[87:80];
  wire [7:0]        dataRegroupBySew_6_11 = bufferStageEnqueueData_6[95:88];
  wire [7:0]        dataRegroupBySew_6_12 = bufferStageEnqueueData_6[103:96];
  wire [7:0]        dataRegroupBySew_6_13 = bufferStageEnqueueData_6[111:104];
  wire [7:0]        dataRegroupBySew_6_14 = bufferStageEnqueueData_6[119:112];
  wire [7:0]        dataRegroupBySew_6_15 = bufferStageEnqueueData_6[127:120];
  wire [7:0]        dataRegroupBySew_6_16 = bufferStageEnqueueData_6[135:128];
  wire [7:0]        dataRegroupBySew_6_17 = bufferStageEnqueueData_6[143:136];
  wire [7:0]        dataRegroupBySew_6_18 = bufferStageEnqueueData_6[151:144];
  wire [7:0]        dataRegroupBySew_6_19 = bufferStageEnqueueData_6[159:152];
  wire [7:0]        dataRegroupBySew_6_20 = bufferStageEnqueueData_6[167:160];
  wire [7:0]        dataRegroupBySew_6_21 = bufferStageEnqueueData_6[175:168];
  wire [7:0]        dataRegroupBySew_6_22 = bufferStageEnqueueData_6[183:176];
  wire [7:0]        dataRegroupBySew_6_23 = bufferStageEnqueueData_6[191:184];
  wire [7:0]        dataRegroupBySew_6_24 = bufferStageEnqueueData_6[199:192];
  wire [7:0]        dataRegroupBySew_6_25 = bufferStageEnqueueData_6[207:200];
  wire [7:0]        dataRegroupBySew_6_26 = bufferStageEnqueueData_6[215:208];
  wire [7:0]        dataRegroupBySew_6_27 = bufferStageEnqueueData_6[223:216];
  wire [7:0]        dataRegroupBySew_6_28 = bufferStageEnqueueData_6[231:224];
  wire [7:0]        dataRegroupBySew_6_29 = bufferStageEnqueueData_6[239:232];
  wire [7:0]        dataRegroupBySew_6_30 = bufferStageEnqueueData_6[247:240];
  wire [7:0]        dataRegroupBySew_6_31 = bufferStageEnqueueData_6[255:248];
  wire [7:0]        dataRegroupBySew_6_32 = bufferStageEnqueueData_6[263:256];
  wire [7:0]        dataRegroupBySew_6_33 = bufferStageEnqueueData_6[271:264];
  wire [7:0]        dataRegroupBySew_6_34 = bufferStageEnqueueData_6[279:272];
  wire [7:0]        dataRegroupBySew_6_35 = bufferStageEnqueueData_6[287:280];
  wire [7:0]        dataRegroupBySew_6_36 = bufferStageEnqueueData_6[295:288];
  wire [7:0]        dataRegroupBySew_6_37 = bufferStageEnqueueData_6[303:296];
  wire [7:0]        dataRegroupBySew_6_38 = bufferStageEnqueueData_6[311:304];
  wire [7:0]        dataRegroupBySew_6_39 = bufferStageEnqueueData_6[319:312];
  wire [7:0]        dataRegroupBySew_6_40 = bufferStageEnqueueData_6[327:320];
  wire [7:0]        dataRegroupBySew_6_41 = bufferStageEnqueueData_6[335:328];
  wire [7:0]        dataRegroupBySew_6_42 = bufferStageEnqueueData_6[343:336];
  wire [7:0]        dataRegroupBySew_6_43 = bufferStageEnqueueData_6[351:344];
  wire [7:0]        dataRegroupBySew_6_44 = bufferStageEnqueueData_6[359:352];
  wire [7:0]        dataRegroupBySew_6_45 = bufferStageEnqueueData_6[367:360];
  wire [7:0]        dataRegroupBySew_6_46 = bufferStageEnqueueData_6[375:368];
  wire [7:0]        dataRegroupBySew_6_47 = bufferStageEnqueueData_6[383:376];
  wire [7:0]        dataRegroupBySew_6_48 = bufferStageEnqueueData_6[391:384];
  wire [7:0]        dataRegroupBySew_6_49 = bufferStageEnqueueData_6[399:392];
  wire [7:0]        dataRegroupBySew_6_50 = bufferStageEnqueueData_6[407:400];
  wire [7:0]        dataRegroupBySew_6_51 = bufferStageEnqueueData_6[415:408];
  wire [7:0]        dataRegroupBySew_6_52 = bufferStageEnqueueData_6[423:416];
  wire [7:0]        dataRegroupBySew_6_53 = bufferStageEnqueueData_6[431:424];
  wire [7:0]        dataRegroupBySew_6_54 = bufferStageEnqueueData_6[439:432];
  wire [7:0]        dataRegroupBySew_6_55 = bufferStageEnqueueData_6[447:440];
  wire [7:0]        dataRegroupBySew_6_56 = bufferStageEnqueueData_6[455:448];
  wire [7:0]        dataRegroupBySew_6_57 = bufferStageEnqueueData_6[463:456];
  wire [7:0]        dataRegroupBySew_6_58 = bufferStageEnqueueData_6[471:464];
  wire [7:0]        dataRegroupBySew_6_59 = bufferStageEnqueueData_6[479:472];
  wire [7:0]        dataRegroupBySew_6_60 = bufferStageEnqueueData_6[487:480];
  wire [7:0]        dataRegroupBySew_6_61 = bufferStageEnqueueData_6[495:488];
  wire [7:0]        dataRegroupBySew_6_62 = bufferStageEnqueueData_6[503:496];
  wire [7:0]        dataRegroupBySew_6_63 = bufferStageEnqueueData_6[511:504];
  wire [7:0]        dataRegroupBySew_6_64 = bufferStageEnqueueData_6[519:512];
  wire [7:0]        dataRegroupBySew_6_65 = bufferStageEnqueueData_6[527:520];
  wire [7:0]        dataRegroupBySew_6_66 = bufferStageEnqueueData_6[535:528];
  wire [7:0]        dataRegroupBySew_6_67 = bufferStageEnqueueData_6[543:536];
  wire [7:0]        dataRegroupBySew_6_68 = bufferStageEnqueueData_6[551:544];
  wire [7:0]        dataRegroupBySew_6_69 = bufferStageEnqueueData_6[559:552];
  wire [7:0]        dataRegroupBySew_6_70 = bufferStageEnqueueData_6[567:560];
  wire [7:0]        dataRegroupBySew_6_71 = bufferStageEnqueueData_6[575:568];
  wire [7:0]        dataRegroupBySew_6_72 = bufferStageEnqueueData_6[583:576];
  wire [7:0]        dataRegroupBySew_6_73 = bufferStageEnqueueData_6[591:584];
  wire [7:0]        dataRegroupBySew_6_74 = bufferStageEnqueueData_6[599:592];
  wire [7:0]        dataRegroupBySew_6_75 = bufferStageEnqueueData_6[607:600];
  wire [7:0]        dataRegroupBySew_6_76 = bufferStageEnqueueData_6[615:608];
  wire [7:0]        dataRegroupBySew_6_77 = bufferStageEnqueueData_6[623:616];
  wire [7:0]        dataRegroupBySew_6_78 = bufferStageEnqueueData_6[631:624];
  wire [7:0]        dataRegroupBySew_6_79 = bufferStageEnqueueData_6[639:632];
  wire [7:0]        dataRegroupBySew_6_80 = bufferStageEnqueueData_6[647:640];
  wire [7:0]        dataRegroupBySew_6_81 = bufferStageEnqueueData_6[655:648];
  wire [7:0]        dataRegroupBySew_6_82 = bufferStageEnqueueData_6[663:656];
  wire [7:0]        dataRegroupBySew_6_83 = bufferStageEnqueueData_6[671:664];
  wire [7:0]        dataRegroupBySew_6_84 = bufferStageEnqueueData_6[679:672];
  wire [7:0]        dataRegroupBySew_6_85 = bufferStageEnqueueData_6[687:680];
  wire [7:0]        dataRegroupBySew_6_86 = bufferStageEnqueueData_6[695:688];
  wire [7:0]        dataRegroupBySew_6_87 = bufferStageEnqueueData_6[703:696];
  wire [7:0]        dataRegroupBySew_6_88 = bufferStageEnqueueData_6[711:704];
  wire [7:0]        dataRegroupBySew_6_89 = bufferStageEnqueueData_6[719:712];
  wire [7:0]        dataRegroupBySew_6_90 = bufferStageEnqueueData_6[727:720];
  wire [7:0]        dataRegroupBySew_6_91 = bufferStageEnqueueData_6[735:728];
  wire [7:0]        dataRegroupBySew_6_92 = bufferStageEnqueueData_6[743:736];
  wire [7:0]        dataRegroupBySew_6_93 = bufferStageEnqueueData_6[751:744];
  wire [7:0]        dataRegroupBySew_6_94 = bufferStageEnqueueData_6[759:752];
  wire [7:0]        dataRegroupBySew_6_95 = bufferStageEnqueueData_6[767:760];
  wire [7:0]        dataRegroupBySew_6_96 = bufferStageEnqueueData_6[775:768];
  wire [7:0]        dataRegroupBySew_6_97 = bufferStageEnqueueData_6[783:776];
  wire [7:0]        dataRegroupBySew_6_98 = bufferStageEnqueueData_6[791:784];
  wire [7:0]        dataRegroupBySew_6_99 = bufferStageEnqueueData_6[799:792];
  wire [7:0]        dataRegroupBySew_6_100 = bufferStageEnqueueData_6[807:800];
  wire [7:0]        dataRegroupBySew_6_101 = bufferStageEnqueueData_6[815:808];
  wire [7:0]        dataRegroupBySew_6_102 = bufferStageEnqueueData_6[823:816];
  wire [7:0]        dataRegroupBySew_6_103 = bufferStageEnqueueData_6[831:824];
  wire [7:0]        dataRegroupBySew_6_104 = bufferStageEnqueueData_6[839:832];
  wire [7:0]        dataRegroupBySew_6_105 = bufferStageEnqueueData_6[847:840];
  wire [7:0]        dataRegroupBySew_6_106 = bufferStageEnqueueData_6[855:848];
  wire [7:0]        dataRegroupBySew_6_107 = bufferStageEnqueueData_6[863:856];
  wire [7:0]        dataRegroupBySew_6_108 = bufferStageEnqueueData_6[871:864];
  wire [7:0]        dataRegroupBySew_6_109 = bufferStageEnqueueData_6[879:872];
  wire [7:0]        dataRegroupBySew_6_110 = bufferStageEnqueueData_6[887:880];
  wire [7:0]        dataRegroupBySew_6_111 = bufferStageEnqueueData_6[895:888];
  wire [7:0]        dataRegroupBySew_6_112 = bufferStageEnqueueData_6[903:896];
  wire [7:0]        dataRegroupBySew_6_113 = bufferStageEnqueueData_6[911:904];
  wire [7:0]        dataRegroupBySew_6_114 = bufferStageEnqueueData_6[919:912];
  wire [7:0]        dataRegroupBySew_6_115 = bufferStageEnqueueData_6[927:920];
  wire [7:0]        dataRegroupBySew_6_116 = bufferStageEnqueueData_6[935:928];
  wire [7:0]        dataRegroupBySew_6_117 = bufferStageEnqueueData_6[943:936];
  wire [7:0]        dataRegroupBySew_6_118 = bufferStageEnqueueData_6[951:944];
  wire [7:0]        dataRegroupBySew_6_119 = bufferStageEnqueueData_6[959:952];
  wire [7:0]        dataRegroupBySew_6_120 = bufferStageEnqueueData_6[967:960];
  wire [7:0]        dataRegroupBySew_6_121 = bufferStageEnqueueData_6[975:968];
  wire [7:0]        dataRegroupBySew_6_122 = bufferStageEnqueueData_6[983:976];
  wire [7:0]        dataRegroupBySew_6_123 = bufferStageEnqueueData_6[991:984];
  wire [7:0]        dataRegroupBySew_6_124 = bufferStageEnqueueData_6[999:992];
  wire [7:0]        dataRegroupBySew_6_125 = bufferStageEnqueueData_6[1007:1000];
  wire [7:0]        dataRegroupBySew_6_126 = bufferStageEnqueueData_6[1015:1008];
  wire [7:0]        dataRegroupBySew_6_127 = bufferStageEnqueueData_6[1023:1016];
  wire [7:0]        dataRegroupBySew_7_0 = bufferStageEnqueueData_7[7:0];
  wire [7:0]        dataRegroupBySew_7_1 = bufferStageEnqueueData_7[15:8];
  wire [7:0]        dataRegroupBySew_7_2 = bufferStageEnqueueData_7[23:16];
  wire [7:0]        dataRegroupBySew_7_3 = bufferStageEnqueueData_7[31:24];
  wire [7:0]        dataRegroupBySew_7_4 = bufferStageEnqueueData_7[39:32];
  wire [7:0]        dataRegroupBySew_7_5 = bufferStageEnqueueData_7[47:40];
  wire [7:0]        dataRegroupBySew_7_6 = bufferStageEnqueueData_7[55:48];
  wire [7:0]        dataRegroupBySew_7_7 = bufferStageEnqueueData_7[63:56];
  wire [7:0]        dataRegroupBySew_7_8 = bufferStageEnqueueData_7[71:64];
  wire [7:0]        dataRegroupBySew_7_9 = bufferStageEnqueueData_7[79:72];
  wire [7:0]        dataRegroupBySew_7_10 = bufferStageEnqueueData_7[87:80];
  wire [7:0]        dataRegroupBySew_7_11 = bufferStageEnqueueData_7[95:88];
  wire [7:0]        dataRegroupBySew_7_12 = bufferStageEnqueueData_7[103:96];
  wire [7:0]        dataRegroupBySew_7_13 = bufferStageEnqueueData_7[111:104];
  wire [7:0]        dataRegroupBySew_7_14 = bufferStageEnqueueData_7[119:112];
  wire [7:0]        dataRegroupBySew_7_15 = bufferStageEnqueueData_7[127:120];
  wire [7:0]        dataRegroupBySew_7_16 = bufferStageEnqueueData_7[135:128];
  wire [7:0]        dataRegroupBySew_7_17 = bufferStageEnqueueData_7[143:136];
  wire [7:0]        dataRegroupBySew_7_18 = bufferStageEnqueueData_7[151:144];
  wire [7:0]        dataRegroupBySew_7_19 = bufferStageEnqueueData_7[159:152];
  wire [7:0]        dataRegroupBySew_7_20 = bufferStageEnqueueData_7[167:160];
  wire [7:0]        dataRegroupBySew_7_21 = bufferStageEnqueueData_7[175:168];
  wire [7:0]        dataRegroupBySew_7_22 = bufferStageEnqueueData_7[183:176];
  wire [7:0]        dataRegroupBySew_7_23 = bufferStageEnqueueData_7[191:184];
  wire [7:0]        dataRegroupBySew_7_24 = bufferStageEnqueueData_7[199:192];
  wire [7:0]        dataRegroupBySew_7_25 = bufferStageEnqueueData_7[207:200];
  wire [7:0]        dataRegroupBySew_7_26 = bufferStageEnqueueData_7[215:208];
  wire [7:0]        dataRegroupBySew_7_27 = bufferStageEnqueueData_7[223:216];
  wire [7:0]        dataRegroupBySew_7_28 = bufferStageEnqueueData_7[231:224];
  wire [7:0]        dataRegroupBySew_7_29 = bufferStageEnqueueData_7[239:232];
  wire [7:0]        dataRegroupBySew_7_30 = bufferStageEnqueueData_7[247:240];
  wire [7:0]        dataRegroupBySew_7_31 = bufferStageEnqueueData_7[255:248];
  wire [7:0]        dataRegroupBySew_7_32 = bufferStageEnqueueData_7[263:256];
  wire [7:0]        dataRegroupBySew_7_33 = bufferStageEnqueueData_7[271:264];
  wire [7:0]        dataRegroupBySew_7_34 = bufferStageEnqueueData_7[279:272];
  wire [7:0]        dataRegroupBySew_7_35 = bufferStageEnqueueData_7[287:280];
  wire [7:0]        dataRegroupBySew_7_36 = bufferStageEnqueueData_7[295:288];
  wire [7:0]        dataRegroupBySew_7_37 = bufferStageEnqueueData_7[303:296];
  wire [7:0]        dataRegroupBySew_7_38 = bufferStageEnqueueData_7[311:304];
  wire [7:0]        dataRegroupBySew_7_39 = bufferStageEnqueueData_7[319:312];
  wire [7:0]        dataRegroupBySew_7_40 = bufferStageEnqueueData_7[327:320];
  wire [7:0]        dataRegroupBySew_7_41 = bufferStageEnqueueData_7[335:328];
  wire [7:0]        dataRegroupBySew_7_42 = bufferStageEnqueueData_7[343:336];
  wire [7:0]        dataRegroupBySew_7_43 = bufferStageEnqueueData_7[351:344];
  wire [7:0]        dataRegroupBySew_7_44 = bufferStageEnqueueData_7[359:352];
  wire [7:0]        dataRegroupBySew_7_45 = bufferStageEnqueueData_7[367:360];
  wire [7:0]        dataRegroupBySew_7_46 = bufferStageEnqueueData_7[375:368];
  wire [7:0]        dataRegroupBySew_7_47 = bufferStageEnqueueData_7[383:376];
  wire [7:0]        dataRegroupBySew_7_48 = bufferStageEnqueueData_7[391:384];
  wire [7:0]        dataRegroupBySew_7_49 = bufferStageEnqueueData_7[399:392];
  wire [7:0]        dataRegroupBySew_7_50 = bufferStageEnqueueData_7[407:400];
  wire [7:0]        dataRegroupBySew_7_51 = bufferStageEnqueueData_7[415:408];
  wire [7:0]        dataRegroupBySew_7_52 = bufferStageEnqueueData_7[423:416];
  wire [7:0]        dataRegroupBySew_7_53 = bufferStageEnqueueData_7[431:424];
  wire [7:0]        dataRegroupBySew_7_54 = bufferStageEnqueueData_7[439:432];
  wire [7:0]        dataRegroupBySew_7_55 = bufferStageEnqueueData_7[447:440];
  wire [7:0]        dataRegroupBySew_7_56 = bufferStageEnqueueData_7[455:448];
  wire [7:0]        dataRegroupBySew_7_57 = bufferStageEnqueueData_7[463:456];
  wire [7:0]        dataRegroupBySew_7_58 = bufferStageEnqueueData_7[471:464];
  wire [7:0]        dataRegroupBySew_7_59 = bufferStageEnqueueData_7[479:472];
  wire [7:0]        dataRegroupBySew_7_60 = bufferStageEnqueueData_7[487:480];
  wire [7:0]        dataRegroupBySew_7_61 = bufferStageEnqueueData_7[495:488];
  wire [7:0]        dataRegroupBySew_7_62 = bufferStageEnqueueData_7[503:496];
  wire [7:0]        dataRegroupBySew_7_63 = bufferStageEnqueueData_7[511:504];
  wire [7:0]        dataRegroupBySew_7_64 = bufferStageEnqueueData_7[519:512];
  wire [7:0]        dataRegroupBySew_7_65 = bufferStageEnqueueData_7[527:520];
  wire [7:0]        dataRegroupBySew_7_66 = bufferStageEnqueueData_7[535:528];
  wire [7:0]        dataRegroupBySew_7_67 = bufferStageEnqueueData_7[543:536];
  wire [7:0]        dataRegroupBySew_7_68 = bufferStageEnqueueData_7[551:544];
  wire [7:0]        dataRegroupBySew_7_69 = bufferStageEnqueueData_7[559:552];
  wire [7:0]        dataRegroupBySew_7_70 = bufferStageEnqueueData_7[567:560];
  wire [7:0]        dataRegroupBySew_7_71 = bufferStageEnqueueData_7[575:568];
  wire [7:0]        dataRegroupBySew_7_72 = bufferStageEnqueueData_7[583:576];
  wire [7:0]        dataRegroupBySew_7_73 = bufferStageEnqueueData_7[591:584];
  wire [7:0]        dataRegroupBySew_7_74 = bufferStageEnqueueData_7[599:592];
  wire [7:0]        dataRegroupBySew_7_75 = bufferStageEnqueueData_7[607:600];
  wire [7:0]        dataRegroupBySew_7_76 = bufferStageEnqueueData_7[615:608];
  wire [7:0]        dataRegroupBySew_7_77 = bufferStageEnqueueData_7[623:616];
  wire [7:0]        dataRegroupBySew_7_78 = bufferStageEnqueueData_7[631:624];
  wire [7:0]        dataRegroupBySew_7_79 = bufferStageEnqueueData_7[639:632];
  wire [7:0]        dataRegroupBySew_7_80 = bufferStageEnqueueData_7[647:640];
  wire [7:0]        dataRegroupBySew_7_81 = bufferStageEnqueueData_7[655:648];
  wire [7:0]        dataRegroupBySew_7_82 = bufferStageEnqueueData_7[663:656];
  wire [7:0]        dataRegroupBySew_7_83 = bufferStageEnqueueData_7[671:664];
  wire [7:0]        dataRegroupBySew_7_84 = bufferStageEnqueueData_7[679:672];
  wire [7:0]        dataRegroupBySew_7_85 = bufferStageEnqueueData_7[687:680];
  wire [7:0]        dataRegroupBySew_7_86 = bufferStageEnqueueData_7[695:688];
  wire [7:0]        dataRegroupBySew_7_87 = bufferStageEnqueueData_7[703:696];
  wire [7:0]        dataRegroupBySew_7_88 = bufferStageEnqueueData_7[711:704];
  wire [7:0]        dataRegroupBySew_7_89 = bufferStageEnqueueData_7[719:712];
  wire [7:0]        dataRegroupBySew_7_90 = bufferStageEnqueueData_7[727:720];
  wire [7:0]        dataRegroupBySew_7_91 = bufferStageEnqueueData_7[735:728];
  wire [7:0]        dataRegroupBySew_7_92 = bufferStageEnqueueData_7[743:736];
  wire [7:0]        dataRegroupBySew_7_93 = bufferStageEnqueueData_7[751:744];
  wire [7:0]        dataRegroupBySew_7_94 = bufferStageEnqueueData_7[759:752];
  wire [7:0]        dataRegroupBySew_7_95 = bufferStageEnqueueData_7[767:760];
  wire [7:0]        dataRegroupBySew_7_96 = bufferStageEnqueueData_7[775:768];
  wire [7:0]        dataRegroupBySew_7_97 = bufferStageEnqueueData_7[783:776];
  wire [7:0]        dataRegroupBySew_7_98 = bufferStageEnqueueData_7[791:784];
  wire [7:0]        dataRegroupBySew_7_99 = bufferStageEnqueueData_7[799:792];
  wire [7:0]        dataRegroupBySew_7_100 = bufferStageEnqueueData_7[807:800];
  wire [7:0]        dataRegroupBySew_7_101 = bufferStageEnqueueData_7[815:808];
  wire [7:0]        dataRegroupBySew_7_102 = bufferStageEnqueueData_7[823:816];
  wire [7:0]        dataRegroupBySew_7_103 = bufferStageEnqueueData_7[831:824];
  wire [7:0]        dataRegroupBySew_7_104 = bufferStageEnqueueData_7[839:832];
  wire [7:0]        dataRegroupBySew_7_105 = bufferStageEnqueueData_7[847:840];
  wire [7:0]        dataRegroupBySew_7_106 = bufferStageEnqueueData_7[855:848];
  wire [7:0]        dataRegroupBySew_7_107 = bufferStageEnqueueData_7[863:856];
  wire [7:0]        dataRegroupBySew_7_108 = bufferStageEnqueueData_7[871:864];
  wire [7:0]        dataRegroupBySew_7_109 = bufferStageEnqueueData_7[879:872];
  wire [7:0]        dataRegroupBySew_7_110 = bufferStageEnqueueData_7[887:880];
  wire [7:0]        dataRegroupBySew_7_111 = bufferStageEnqueueData_7[895:888];
  wire [7:0]        dataRegroupBySew_7_112 = bufferStageEnqueueData_7[903:896];
  wire [7:0]        dataRegroupBySew_7_113 = bufferStageEnqueueData_7[911:904];
  wire [7:0]        dataRegroupBySew_7_114 = bufferStageEnqueueData_7[919:912];
  wire [7:0]        dataRegroupBySew_7_115 = bufferStageEnqueueData_7[927:920];
  wire [7:0]        dataRegroupBySew_7_116 = bufferStageEnqueueData_7[935:928];
  wire [7:0]        dataRegroupBySew_7_117 = bufferStageEnqueueData_7[943:936];
  wire [7:0]        dataRegroupBySew_7_118 = bufferStageEnqueueData_7[951:944];
  wire [7:0]        dataRegroupBySew_7_119 = bufferStageEnqueueData_7[959:952];
  wire [7:0]        dataRegroupBySew_7_120 = bufferStageEnqueueData_7[967:960];
  wire [7:0]        dataRegroupBySew_7_121 = bufferStageEnqueueData_7[975:968];
  wire [7:0]        dataRegroupBySew_7_122 = bufferStageEnqueueData_7[983:976];
  wire [7:0]        dataRegroupBySew_7_123 = bufferStageEnqueueData_7[991:984];
  wire [7:0]        dataRegroupBySew_7_124 = bufferStageEnqueueData_7[999:992];
  wire [7:0]        dataRegroupBySew_7_125 = bufferStageEnqueueData_7[1007:1000];
  wire [7:0]        dataRegroupBySew_7_126 = bufferStageEnqueueData_7[1015:1008];
  wire [7:0]        dataRegroupBySew_7_127 = bufferStageEnqueueData_7[1023:1016];
  wire [15:0]       dataInMem_lo_lo_lo_lo_lo_lo = {dataRegroupBySew_0_1, dataRegroupBySew_0_0};
  wire [15:0]       dataInMem_lo_lo_lo_lo_lo_hi = {dataRegroupBySew_0_3, dataRegroupBySew_0_2};
  wire [31:0]       dataInMem_lo_lo_lo_lo_lo = {dataInMem_lo_lo_lo_lo_lo_hi, dataInMem_lo_lo_lo_lo_lo_lo};
  wire [15:0]       dataInMem_lo_lo_lo_lo_hi_lo = {dataRegroupBySew_0_5, dataRegroupBySew_0_4};
  wire [15:0]       dataInMem_lo_lo_lo_lo_hi_hi = {dataRegroupBySew_0_7, dataRegroupBySew_0_6};
  wire [31:0]       dataInMem_lo_lo_lo_lo_hi = {dataInMem_lo_lo_lo_lo_hi_hi, dataInMem_lo_lo_lo_lo_hi_lo};
  wire [63:0]       dataInMem_lo_lo_lo_lo = {dataInMem_lo_lo_lo_lo_hi, dataInMem_lo_lo_lo_lo_lo};
  wire [15:0]       dataInMem_lo_lo_lo_hi_lo_lo = {dataRegroupBySew_0_9, dataRegroupBySew_0_8};
  wire [15:0]       dataInMem_lo_lo_lo_hi_lo_hi = {dataRegroupBySew_0_11, dataRegroupBySew_0_10};
  wire [31:0]       dataInMem_lo_lo_lo_hi_lo = {dataInMem_lo_lo_lo_hi_lo_hi, dataInMem_lo_lo_lo_hi_lo_lo};
  wire [15:0]       dataInMem_lo_lo_lo_hi_hi_lo = {dataRegroupBySew_0_13, dataRegroupBySew_0_12};
  wire [15:0]       dataInMem_lo_lo_lo_hi_hi_hi = {dataRegroupBySew_0_15, dataRegroupBySew_0_14};
  wire [31:0]       dataInMem_lo_lo_lo_hi_hi = {dataInMem_lo_lo_lo_hi_hi_hi, dataInMem_lo_lo_lo_hi_hi_lo};
  wire [63:0]       dataInMem_lo_lo_lo_hi = {dataInMem_lo_lo_lo_hi_hi, dataInMem_lo_lo_lo_hi_lo};
  wire [127:0]      dataInMem_lo_lo_lo = {dataInMem_lo_lo_lo_hi, dataInMem_lo_lo_lo_lo};
  wire [15:0]       dataInMem_lo_lo_hi_lo_lo_lo = {dataRegroupBySew_0_17, dataRegroupBySew_0_16};
  wire [15:0]       dataInMem_lo_lo_hi_lo_lo_hi = {dataRegroupBySew_0_19, dataRegroupBySew_0_18};
  wire [31:0]       dataInMem_lo_lo_hi_lo_lo = {dataInMem_lo_lo_hi_lo_lo_hi, dataInMem_lo_lo_hi_lo_lo_lo};
  wire [15:0]       dataInMem_lo_lo_hi_lo_hi_lo = {dataRegroupBySew_0_21, dataRegroupBySew_0_20};
  wire [15:0]       dataInMem_lo_lo_hi_lo_hi_hi = {dataRegroupBySew_0_23, dataRegroupBySew_0_22};
  wire [31:0]       dataInMem_lo_lo_hi_lo_hi = {dataInMem_lo_lo_hi_lo_hi_hi, dataInMem_lo_lo_hi_lo_hi_lo};
  wire [63:0]       dataInMem_lo_lo_hi_lo = {dataInMem_lo_lo_hi_lo_hi, dataInMem_lo_lo_hi_lo_lo};
  wire [15:0]       dataInMem_lo_lo_hi_hi_lo_lo = {dataRegroupBySew_0_25, dataRegroupBySew_0_24};
  wire [15:0]       dataInMem_lo_lo_hi_hi_lo_hi = {dataRegroupBySew_0_27, dataRegroupBySew_0_26};
  wire [31:0]       dataInMem_lo_lo_hi_hi_lo = {dataInMem_lo_lo_hi_hi_lo_hi, dataInMem_lo_lo_hi_hi_lo_lo};
  wire [15:0]       dataInMem_lo_lo_hi_hi_hi_lo = {dataRegroupBySew_0_29, dataRegroupBySew_0_28};
  wire [15:0]       dataInMem_lo_lo_hi_hi_hi_hi = {dataRegroupBySew_0_31, dataRegroupBySew_0_30};
  wire [31:0]       dataInMem_lo_lo_hi_hi_hi = {dataInMem_lo_lo_hi_hi_hi_hi, dataInMem_lo_lo_hi_hi_hi_lo};
  wire [63:0]       dataInMem_lo_lo_hi_hi = {dataInMem_lo_lo_hi_hi_hi, dataInMem_lo_lo_hi_hi_lo};
  wire [127:0]      dataInMem_lo_lo_hi = {dataInMem_lo_lo_hi_hi, dataInMem_lo_lo_hi_lo};
  wire [255:0]      dataInMem_lo_lo = {dataInMem_lo_lo_hi, dataInMem_lo_lo_lo};
  wire [15:0]       dataInMem_lo_hi_lo_lo_lo_lo = {dataRegroupBySew_0_33, dataRegroupBySew_0_32};
  wire [15:0]       dataInMem_lo_hi_lo_lo_lo_hi = {dataRegroupBySew_0_35, dataRegroupBySew_0_34};
  wire [31:0]       dataInMem_lo_hi_lo_lo_lo = {dataInMem_lo_hi_lo_lo_lo_hi, dataInMem_lo_hi_lo_lo_lo_lo};
  wire [15:0]       dataInMem_lo_hi_lo_lo_hi_lo = {dataRegroupBySew_0_37, dataRegroupBySew_0_36};
  wire [15:0]       dataInMem_lo_hi_lo_lo_hi_hi = {dataRegroupBySew_0_39, dataRegroupBySew_0_38};
  wire [31:0]       dataInMem_lo_hi_lo_lo_hi = {dataInMem_lo_hi_lo_lo_hi_hi, dataInMem_lo_hi_lo_lo_hi_lo};
  wire [63:0]       dataInMem_lo_hi_lo_lo = {dataInMem_lo_hi_lo_lo_hi, dataInMem_lo_hi_lo_lo_lo};
  wire [15:0]       dataInMem_lo_hi_lo_hi_lo_lo = {dataRegroupBySew_0_41, dataRegroupBySew_0_40};
  wire [15:0]       dataInMem_lo_hi_lo_hi_lo_hi = {dataRegroupBySew_0_43, dataRegroupBySew_0_42};
  wire [31:0]       dataInMem_lo_hi_lo_hi_lo = {dataInMem_lo_hi_lo_hi_lo_hi, dataInMem_lo_hi_lo_hi_lo_lo};
  wire [15:0]       dataInMem_lo_hi_lo_hi_hi_lo = {dataRegroupBySew_0_45, dataRegroupBySew_0_44};
  wire [15:0]       dataInMem_lo_hi_lo_hi_hi_hi = {dataRegroupBySew_0_47, dataRegroupBySew_0_46};
  wire [31:0]       dataInMem_lo_hi_lo_hi_hi = {dataInMem_lo_hi_lo_hi_hi_hi, dataInMem_lo_hi_lo_hi_hi_lo};
  wire [63:0]       dataInMem_lo_hi_lo_hi = {dataInMem_lo_hi_lo_hi_hi, dataInMem_lo_hi_lo_hi_lo};
  wire [127:0]      dataInMem_lo_hi_lo = {dataInMem_lo_hi_lo_hi, dataInMem_lo_hi_lo_lo};
  wire [15:0]       dataInMem_lo_hi_hi_lo_lo_lo = {dataRegroupBySew_0_49, dataRegroupBySew_0_48};
  wire [15:0]       dataInMem_lo_hi_hi_lo_lo_hi = {dataRegroupBySew_0_51, dataRegroupBySew_0_50};
  wire [31:0]       dataInMem_lo_hi_hi_lo_lo = {dataInMem_lo_hi_hi_lo_lo_hi, dataInMem_lo_hi_hi_lo_lo_lo};
  wire [15:0]       dataInMem_lo_hi_hi_lo_hi_lo = {dataRegroupBySew_0_53, dataRegroupBySew_0_52};
  wire [15:0]       dataInMem_lo_hi_hi_lo_hi_hi = {dataRegroupBySew_0_55, dataRegroupBySew_0_54};
  wire [31:0]       dataInMem_lo_hi_hi_lo_hi = {dataInMem_lo_hi_hi_lo_hi_hi, dataInMem_lo_hi_hi_lo_hi_lo};
  wire [63:0]       dataInMem_lo_hi_hi_lo = {dataInMem_lo_hi_hi_lo_hi, dataInMem_lo_hi_hi_lo_lo};
  wire [15:0]       dataInMem_lo_hi_hi_hi_lo_lo = {dataRegroupBySew_0_57, dataRegroupBySew_0_56};
  wire [15:0]       dataInMem_lo_hi_hi_hi_lo_hi = {dataRegroupBySew_0_59, dataRegroupBySew_0_58};
  wire [31:0]       dataInMem_lo_hi_hi_hi_lo = {dataInMem_lo_hi_hi_hi_lo_hi, dataInMem_lo_hi_hi_hi_lo_lo};
  wire [15:0]       dataInMem_lo_hi_hi_hi_hi_lo = {dataRegroupBySew_0_61, dataRegroupBySew_0_60};
  wire [15:0]       dataInMem_lo_hi_hi_hi_hi_hi = {dataRegroupBySew_0_63, dataRegroupBySew_0_62};
  wire [31:0]       dataInMem_lo_hi_hi_hi_hi = {dataInMem_lo_hi_hi_hi_hi_hi, dataInMem_lo_hi_hi_hi_hi_lo};
  wire [63:0]       dataInMem_lo_hi_hi_hi = {dataInMem_lo_hi_hi_hi_hi, dataInMem_lo_hi_hi_hi_lo};
  wire [127:0]      dataInMem_lo_hi_hi = {dataInMem_lo_hi_hi_hi, dataInMem_lo_hi_hi_lo};
  wire [255:0]      dataInMem_lo_hi = {dataInMem_lo_hi_hi, dataInMem_lo_hi_lo};
  wire [511:0]      dataInMem_lo = {dataInMem_lo_hi, dataInMem_lo_lo};
  wire [15:0]       dataInMem_hi_lo_lo_lo_lo_lo = {dataRegroupBySew_0_65, dataRegroupBySew_0_64};
  wire [15:0]       dataInMem_hi_lo_lo_lo_lo_hi = {dataRegroupBySew_0_67, dataRegroupBySew_0_66};
  wire [31:0]       dataInMem_hi_lo_lo_lo_lo = {dataInMem_hi_lo_lo_lo_lo_hi, dataInMem_hi_lo_lo_lo_lo_lo};
  wire [15:0]       dataInMem_hi_lo_lo_lo_hi_lo = {dataRegroupBySew_0_69, dataRegroupBySew_0_68};
  wire [15:0]       dataInMem_hi_lo_lo_lo_hi_hi = {dataRegroupBySew_0_71, dataRegroupBySew_0_70};
  wire [31:0]       dataInMem_hi_lo_lo_lo_hi = {dataInMem_hi_lo_lo_lo_hi_hi, dataInMem_hi_lo_lo_lo_hi_lo};
  wire [63:0]       dataInMem_hi_lo_lo_lo = {dataInMem_hi_lo_lo_lo_hi, dataInMem_hi_lo_lo_lo_lo};
  wire [15:0]       dataInMem_hi_lo_lo_hi_lo_lo = {dataRegroupBySew_0_73, dataRegroupBySew_0_72};
  wire [15:0]       dataInMem_hi_lo_lo_hi_lo_hi = {dataRegroupBySew_0_75, dataRegroupBySew_0_74};
  wire [31:0]       dataInMem_hi_lo_lo_hi_lo = {dataInMem_hi_lo_lo_hi_lo_hi, dataInMem_hi_lo_lo_hi_lo_lo};
  wire [15:0]       dataInMem_hi_lo_lo_hi_hi_lo = {dataRegroupBySew_0_77, dataRegroupBySew_0_76};
  wire [15:0]       dataInMem_hi_lo_lo_hi_hi_hi = {dataRegroupBySew_0_79, dataRegroupBySew_0_78};
  wire [31:0]       dataInMem_hi_lo_lo_hi_hi = {dataInMem_hi_lo_lo_hi_hi_hi, dataInMem_hi_lo_lo_hi_hi_lo};
  wire [63:0]       dataInMem_hi_lo_lo_hi = {dataInMem_hi_lo_lo_hi_hi, dataInMem_hi_lo_lo_hi_lo};
  wire [127:0]      dataInMem_hi_lo_lo = {dataInMem_hi_lo_lo_hi, dataInMem_hi_lo_lo_lo};
  wire [15:0]       dataInMem_hi_lo_hi_lo_lo_lo = {dataRegroupBySew_0_81, dataRegroupBySew_0_80};
  wire [15:0]       dataInMem_hi_lo_hi_lo_lo_hi = {dataRegroupBySew_0_83, dataRegroupBySew_0_82};
  wire [31:0]       dataInMem_hi_lo_hi_lo_lo = {dataInMem_hi_lo_hi_lo_lo_hi, dataInMem_hi_lo_hi_lo_lo_lo};
  wire [15:0]       dataInMem_hi_lo_hi_lo_hi_lo = {dataRegroupBySew_0_85, dataRegroupBySew_0_84};
  wire [15:0]       dataInMem_hi_lo_hi_lo_hi_hi = {dataRegroupBySew_0_87, dataRegroupBySew_0_86};
  wire [31:0]       dataInMem_hi_lo_hi_lo_hi = {dataInMem_hi_lo_hi_lo_hi_hi, dataInMem_hi_lo_hi_lo_hi_lo};
  wire [63:0]       dataInMem_hi_lo_hi_lo = {dataInMem_hi_lo_hi_lo_hi, dataInMem_hi_lo_hi_lo_lo};
  wire [15:0]       dataInMem_hi_lo_hi_hi_lo_lo = {dataRegroupBySew_0_89, dataRegroupBySew_0_88};
  wire [15:0]       dataInMem_hi_lo_hi_hi_lo_hi = {dataRegroupBySew_0_91, dataRegroupBySew_0_90};
  wire [31:0]       dataInMem_hi_lo_hi_hi_lo = {dataInMem_hi_lo_hi_hi_lo_hi, dataInMem_hi_lo_hi_hi_lo_lo};
  wire [15:0]       dataInMem_hi_lo_hi_hi_hi_lo = {dataRegroupBySew_0_93, dataRegroupBySew_0_92};
  wire [15:0]       dataInMem_hi_lo_hi_hi_hi_hi = {dataRegroupBySew_0_95, dataRegroupBySew_0_94};
  wire [31:0]       dataInMem_hi_lo_hi_hi_hi = {dataInMem_hi_lo_hi_hi_hi_hi, dataInMem_hi_lo_hi_hi_hi_lo};
  wire [63:0]       dataInMem_hi_lo_hi_hi = {dataInMem_hi_lo_hi_hi_hi, dataInMem_hi_lo_hi_hi_lo};
  wire [127:0]      dataInMem_hi_lo_hi = {dataInMem_hi_lo_hi_hi, dataInMem_hi_lo_hi_lo};
  wire [255:0]      dataInMem_hi_lo = {dataInMem_hi_lo_hi, dataInMem_hi_lo_lo};
  wire [15:0]       dataInMem_hi_hi_lo_lo_lo_lo = {dataRegroupBySew_0_97, dataRegroupBySew_0_96};
  wire [15:0]       dataInMem_hi_hi_lo_lo_lo_hi = {dataRegroupBySew_0_99, dataRegroupBySew_0_98};
  wire [31:0]       dataInMem_hi_hi_lo_lo_lo = {dataInMem_hi_hi_lo_lo_lo_hi, dataInMem_hi_hi_lo_lo_lo_lo};
  wire [15:0]       dataInMem_hi_hi_lo_lo_hi_lo = {dataRegroupBySew_0_101, dataRegroupBySew_0_100};
  wire [15:0]       dataInMem_hi_hi_lo_lo_hi_hi = {dataRegroupBySew_0_103, dataRegroupBySew_0_102};
  wire [31:0]       dataInMem_hi_hi_lo_lo_hi = {dataInMem_hi_hi_lo_lo_hi_hi, dataInMem_hi_hi_lo_lo_hi_lo};
  wire [63:0]       dataInMem_hi_hi_lo_lo = {dataInMem_hi_hi_lo_lo_hi, dataInMem_hi_hi_lo_lo_lo};
  wire [15:0]       dataInMem_hi_hi_lo_hi_lo_lo = {dataRegroupBySew_0_105, dataRegroupBySew_0_104};
  wire [15:0]       dataInMem_hi_hi_lo_hi_lo_hi = {dataRegroupBySew_0_107, dataRegroupBySew_0_106};
  wire [31:0]       dataInMem_hi_hi_lo_hi_lo = {dataInMem_hi_hi_lo_hi_lo_hi, dataInMem_hi_hi_lo_hi_lo_lo};
  wire [15:0]       dataInMem_hi_hi_lo_hi_hi_lo = {dataRegroupBySew_0_109, dataRegroupBySew_0_108};
  wire [15:0]       dataInMem_hi_hi_lo_hi_hi_hi = {dataRegroupBySew_0_111, dataRegroupBySew_0_110};
  wire [31:0]       dataInMem_hi_hi_lo_hi_hi = {dataInMem_hi_hi_lo_hi_hi_hi, dataInMem_hi_hi_lo_hi_hi_lo};
  wire [63:0]       dataInMem_hi_hi_lo_hi = {dataInMem_hi_hi_lo_hi_hi, dataInMem_hi_hi_lo_hi_lo};
  wire [127:0]      dataInMem_hi_hi_lo = {dataInMem_hi_hi_lo_hi, dataInMem_hi_hi_lo_lo};
  wire [15:0]       dataInMem_hi_hi_hi_lo_lo_lo = {dataRegroupBySew_0_113, dataRegroupBySew_0_112};
  wire [15:0]       dataInMem_hi_hi_hi_lo_lo_hi = {dataRegroupBySew_0_115, dataRegroupBySew_0_114};
  wire [31:0]       dataInMem_hi_hi_hi_lo_lo = {dataInMem_hi_hi_hi_lo_lo_hi, dataInMem_hi_hi_hi_lo_lo_lo};
  wire [15:0]       dataInMem_hi_hi_hi_lo_hi_lo = {dataRegroupBySew_0_117, dataRegroupBySew_0_116};
  wire [15:0]       dataInMem_hi_hi_hi_lo_hi_hi = {dataRegroupBySew_0_119, dataRegroupBySew_0_118};
  wire [31:0]       dataInMem_hi_hi_hi_lo_hi = {dataInMem_hi_hi_hi_lo_hi_hi, dataInMem_hi_hi_hi_lo_hi_lo};
  wire [63:0]       dataInMem_hi_hi_hi_lo = {dataInMem_hi_hi_hi_lo_hi, dataInMem_hi_hi_hi_lo_lo};
  wire [15:0]       dataInMem_hi_hi_hi_hi_lo_lo = {dataRegroupBySew_0_121, dataRegroupBySew_0_120};
  wire [15:0]       dataInMem_hi_hi_hi_hi_lo_hi = {dataRegroupBySew_0_123, dataRegroupBySew_0_122};
  wire [31:0]       dataInMem_hi_hi_hi_hi_lo = {dataInMem_hi_hi_hi_hi_lo_hi, dataInMem_hi_hi_hi_hi_lo_lo};
  wire [15:0]       dataInMem_hi_hi_hi_hi_hi_lo = {dataRegroupBySew_0_125, dataRegroupBySew_0_124};
  wire [15:0]       dataInMem_hi_hi_hi_hi_hi_hi = {dataRegroupBySew_0_127, dataRegroupBySew_0_126};
  wire [31:0]       dataInMem_hi_hi_hi_hi_hi = {dataInMem_hi_hi_hi_hi_hi_hi, dataInMem_hi_hi_hi_hi_hi_lo};
  wire [63:0]       dataInMem_hi_hi_hi_hi = {dataInMem_hi_hi_hi_hi_hi, dataInMem_hi_hi_hi_hi_lo};
  wire [127:0]      dataInMem_hi_hi_hi = {dataInMem_hi_hi_hi_hi, dataInMem_hi_hi_hi_lo};
  wire [255:0]      dataInMem_hi_hi = {dataInMem_hi_hi_hi, dataInMem_hi_hi_lo};
  wire [511:0]      dataInMem_hi = {dataInMem_hi_hi, dataInMem_hi_lo};
  wire [1023:0]     dataInMem = {dataInMem_hi, dataInMem_lo};
  wire [1023:0]     regroupCacheLine_0 = dataInMem;
  wire [1023:0]     res = regroupCacheLine_0;
  wire [2047:0]     lo_lo = {1024'h0, res};
  wire [4095:0]     lo = {2048'h0, lo_lo};
  wire [8191:0]     regroupLoadData_0_0 = {4096'h0, lo};
  wire [31:0]       dataInMem_lo_lo_lo_lo_lo_lo_1 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1, dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [31:0]       dataInMem_lo_lo_lo_lo_lo_hi_1 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3, dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [63:0]       dataInMem_lo_lo_lo_lo_lo_1 = {dataInMem_lo_lo_lo_lo_lo_hi_1, dataInMem_lo_lo_lo_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_lo_lo_lo_hi_lo_1 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5, dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [31:0]       dataInMem_lo_lo_lo_lo_hi_hi_1 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7, dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [63:0]       dataInMem_lo_lo_lo_lo_hi_1 = {dataInMem_lo_lo_lo_lo_hi_hi_1, dataInMem_lo_lo_lo_lo_hi_lo_1};
  wire [127:0]      dataInMem_lo_lo_lo_lo_1 = {dataInMem_lo_lo_lo_lo_hi_1, dataInMem_lo_lo_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_lo_lo_hi_lo_lo_1 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9, dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [31:0]       dataInMem_lo_lo_lo_hi_lo_hi_1 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11, dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [63:0]       dataInMem_lo_lo_lo_hi_lo_1 = {dataInMem_lo_lo_lo_hi_lo_hi_1, dataInMem_lo_lo_lo_hi_lo_lo_1};
  wire [31:0]       dataInMem_lo_lo_lo_hi_hi_lo_1 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13, dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [31:0]       dataInMem_lo_lo_lo_hi_hi_hi_1 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15, dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [63:0]       dataInMem_lo_lo_lo_hi_hi_1 = {dataInMem_lo_lo_lo_hi_hi_hi_1, dataInMem_lo_lo_lo_hi_hi_lo_1};
  wire [127:0]      dataInMem_lo_lo_lo_hi_1 = {dataInMem_lo_lo_lo_hi_hi_1, dataInMem_lo_lo_lo_hi_lo_1};
  wire [255:0]      dataInMem_lo_lo_lo_1 = {dataInMem_lo_lo_lo_hi_1, dataInMem_lo_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_lo_hi_lo_lo_lo_1 = {dataRegroupBySew_1_17, dataRegroupBySew_0_17, dataRegroupBySew_1_16, dataRegroupBySew_0_16};
  wire [31:0]       dataInMem_lo_lo_hi_lo_lo_hi_1 = {dataRegroupBySew_1_19, dataRegroupBySew_0_19, dataRegroupBySew_1_18, dataRegroupBySew_0_18};
  wire [63:0]       dataInMem_lo_lo_hi_lo_lo_1 = {dataInMem_lo_lo_hi_lo_lo_hi_1, dataInMem_lo_lo_hi_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_lo_hi_lo_hi_lo_1 = {dataRegroupBySew_1_21, dataRegroupBySew_0_21, dataRegroupBySew_1_20, dataRegroupBySew_0_20};
  wire [31:0]       dataInMem_lo_lo_hi_lo_hi_hi_1 = {dataRegroupBySew_1_23, dataRegroupBySew_0_23, dataRegroupBySew_1_22, dataRegroupBySew_0_22};
  wire [63:0]       dataInMem_lo_lo_hi_lo_hi_1 = {dataInMem_lo_lo_hi_lo_hi_hi_1, dataInMem_lo_lo_hi_lo_hi_lo_1};
  wire [127:0]      dataInMem_lo_lo_hi_lo_1 = {dataInMem_lo_lo_hi_lo_hi_1, dataInMem_lo_lo_hi_lo_lo_1};
  wire [31:0]       dataInMem_lo_lo_hi_hi_lo_lo_1 = {dataRegroupBySew_1_25, dataRegroupBySew_0_25, dataRegroupBySew_1_24, dataRegroupBySew_0_24};
  wire [31:0]       dataInMem_lo_lo_hi_hi_lo_hi_1 = {dataRegroupBySew_1_27, dataRegroupBySew_0_27, dataRegroupBySew_1_26, dataRegroupBySew_0_26};
  wire [63:0]       dataInMem_lo_lo_hi_hi_lo_1 = {dataInMem_lo_lo_hi_hi_lo_hi_1, dataInMem_lo_lo_hi_hi_lo_lo_1};
  wire [31:0]       dataInMem_lo_lo_hi_hi_hi_lo_1 = {dataRegroupBySew_1_29, dataRegroupBySew_0_29, dataRegroupBySew_1_28, dataRegroupBySew_0_28};
  wire [31:0]       dataInMem_lo_lo_hi_hi_hi_hi_1 = {dataRegroupBySew_1_31, dataRegroupBySew_0_31, dataRegroupBySew_1_30, dataRegroupBySew_0_30};
  wire [63:0]       dataInMem_lo_lo_hi_hi_hi_1 = {dataInMem_lo_lo_hi_hi_hi_hi_1, dataInMem_lo_lo_hi_hi_hi_lo_1};
  wire [127:0]      dataInMem_lo_lo_hi_hi_1 = {dataInMem_lo_lo_hi_hi_hi_1, dataInMem_lo_lo_hi_hi_lo_1};
  wire [255:0]      dataInMem_lo_lo_hi_1 = {dataInMem_lo_lo_hi_hi_1, dataInMem_lo_lo_hi_lo_1};
  wire [511:0]      dataInMem_lo_lo_1 = {dataInMem_lo_lo_hi_1, dataInMem_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_lo_lo_lo_lo_1 = {dataRegroupBySew_1_33, dataRegroupBySew_0_33, dataRegroupBySew_1_32, dataRegroupBySew_0_32};
  wire [31:0]       dataInMem_lo_hi_lo_lo_lo_hi_1 = {dataRegroupBySew_1_35, dataRegroupBySew_0_35, dataRegroupBySew_1_34, dataRegroupBySew_0_34};
  wire [63:0]       dataInMem_lo_hi_lo_lo_lo_1 = {dataInMem_lo_hi_lo_lo_lo_hi_1, dataInMem_lo_hi_lo_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_lo_lo_hi_lo_1 = {dataRegroupBySew_1_37, dataRegroupBySew_0_37, dataRegroupBySew_1_36, dataRegroupBySew_0_36};
  wire [31:0]       dataInMem_lo_hi_lo_lo_hi_hi_1 = {dataRegroupBySew_1_39, dataRegroupBySew_0_39, dataRegroupBySew_1_38, dataRegroupBySew_0_38};
  wire [63:0]       dataInMem_lo_hi_lo_lo_hi_1 = {dataInMem_lo_hi_lo_lo_hi_hi_1, dataInMem_lo_hi_lo_lo_hi_lo_1};
  wire [127:0]      dataInMem_lo_hi_lo_lo_1 = {dataInMem_lo_hi_lo_lo_hi_1, dataInMem_lo_hi_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_lo_hi_lo_lo_1 = {dataRegroupBySew_1_41, dataRegroupBySew_0_41, dataRegroupBySew_1_40, dataRegroupBySew_0_40};
  wire [31:0]       dataInMem_lo_hi_lo_hi_lo_hi_1 = {dataRegroupBySew_1_43, dataRegroupBySew_0_43, dataRegroupBySew_1_42, dataRegroupBySew_0_42};
  wire [63:0]       dataInMem_lo_hi_lo_hi_lo_1 = {dataInMem_lo_hi_lo_hi_lo_hi_1, dataInMem_lo_hi_lo_hi_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_lo_hi_hi_lo_1 = {dataRegroupBySew_1_45, dataRegroupBySew_0_45, dataRegroupBySew_1_44, dataRegroupBySew_0_44};
  wire [31:0]       dataInMem_lo_hi_lo_hi_hi_hi_1 = {dataRegroupBySew_1_47, dataRegroupBySew_0_47, dataRegroupBySew_1_46, dataRegroupBySew_0_46};
  wire [63:0]       dataInMem_lo_hi_lo_hi_hi_1 = {dataInMem_lo_hi_lo_hi_hi_hi_1, dataInMem_lo_hi_lo_hi_hi_lo_1};
  wire [127:0]      dataInMem_lo_hi_lo_hi_1 = {dataInMem_lo_hi_lo_hi_hi_1, dataInMem_lo_hi_lo_hi_lo_1};
  wire [255:0]      dataInMem_lo_hi_lo_1 = {dataInMem_lo_hi_lo_hi_1, dataInMem_lo_hi_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_hi_lo_lo_lo_1 = {dataRegroupBySew_1_49, dataRegroupBySew_0_49, dataRegroupBySew_1_48, dataRegroupBySew_0_48};
  wire [31:0]       dataInMem_lo_hi_hi_lo_lo_hi_1 = {dataRegroupBySew_1_51, dataRegroupBySew_0_51, dataRegroupBySew_1_50, dataRegroupBySew_0_50};
  wire [63:0]       dataInMem_lo_hi_hi_lo_lo_1 = {dataInMem_lo_hi_hi_lo_lo_hi_1, dataInMem_lo_hi_hi_lo_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_hi_lo_hi_lo_1 = {dataRegroupBySew_1_53, dataRegroupBySew_0_53, dataRegroupBySew_1_52, dataRegroupBySew_0_52};
  wire [31:0]       dataInMem_lo_hi_hi_lo_hi_hi_1 = {dataRegroupBySew_1_55, dataRegroupBySew_0_55, dataRegroupBySew_1_54, dataRegroupBySew_0_54};
  wire [63:0]       dataInMem_lo_hi_hi_lo_hi_1 = {dataInMem_lo_hi_hi_lo_hi_hi_1, dataInMem_lo_hi_hi_lo_hi_lo_1};
  wire [127:0]      dataInMem_lo_hi_hi_lo_1 = {dataInMem_lo_hi_hi_lo_hi_1, dataInMem_lo_hi_hi_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_hi_hi_lo_lo_1 = {dataRegroupBySew_1_57, dataRegroupBySew_0_57, dataRegroupBySew_1_56, dataRegroupBySew_0_56};
  wire [31:0]       dataInMem_lo_hi_hi_hi_lo_hi_1 = {dataRegroupBySew_1_59, dataRegroupBySew_0_59, dataRegroupBySew_1_58, dataRegroupBySew_0_58};
  wire [63:0]       dataInMem_lo_hi_hi_hi_lo_1 = {dataInMem_lo_hi_hi_hi_lo_hi_1, dataInMem_lo_hi_hi_hi_lo_lo_1};
  wire [31:0]       dataInMem_lo_hi_hi_hi_hi_lo_1 = {dataRegroupBySew_1_61, dataRegroupBySew_0_61, dataRegroupBySew_1_60, dataRegroupBySew_0_60};
  wire [31:0]       dataInMem_lo_hi_hi_hi_hi_hi_1 = {dataRegroupBySew_1_63, dataRegroupBySew_0_63, dataRegroupBySew_1_62, dataRegroupBySew_0_62};
  wire [63:0]       dataInMem_lo_hi_hi_hi_hi_1 = {dataInMem_lo_hi_hi_hi_hi_hi_1, dataInMem_lo_hi_hi_hi_hi_lo_1};
  wire [127:0]      dataInMem_lo_hi_hi_hi_1 = {dataInMem_lo_hi_hi_hi_hi_1, dataInMem_lo_hi_hi_hi_lo_1};
  wire [255:0]      dataInMem_lo_hi_hi_1 = {dataInMem_lo_hi_hi_hi_1, dataInMem_lo_hi_hi_lo_1};
  wire [511:0]      dataInMem_lo_hi_1 = {dataInMem_lo_hi_hi_1, dataInMem_lo_hi_lo_1};
  wire [1023:0]     dataInMem_lo_1 = {dataInMem_lo_hi_1, dataInMem_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_lo_lo_lo_lo_1 = {dataRegroupBySew_1_65, dataRegroupBySew_0_65, dataRegroupBySew_1_64, dataRegroupBySew_0_64};
  wire [31:0]       dataInMem_hi_lo_lo_lo_lo_hi_1 = {dataRegroupBySew_1_67, dataRegroupBySew_0_67, dataRegroupBySew_1_66, dataRegroupBySew_0_66};
  wire [63:0]       dataInMem_hi_lo_lo_lo_lo_1 = {dataInMem_hi_lo_lo_lo_lo_hi_1, dataInMem_hi_lo_lo_lo_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_lo_lo_hi_lo_1 = {dataRegroupBySew_1_69, dataRegroupBySew_0_69, dataRegroupBySew_1_68, dataRegroupBySew_0_68};
  wire [31:0]       dataInMem_hi_lo_lo_lo_hi_hi_1 = {dataRegroupBySew_1_71, dataRegroupBySew_0_71, dataRegroupBySew_1_70, dataRegroupBySew_0_70};
  wire [63:0]       dataInMem_hi_lo_lo_lo_hi_1 = {dataInMem_hi_lo_lo_lo_hi_hi_1, dataInMem_hi_lo_lo_lo_hi_lo_1};
  wire [127:0]      dataInMem_hi_lo_lo_lo_1 = {dataInMem_hi_lo_lo_lo_hi_1, dataInMem_hi_lo_lo_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_lo_hi_lo_lo_1 = {dataRegroupBySew_1_73, dataRegroupBySew_0_73, dataRegroupBySew_1_72, dataRegroupBySew_0_72};
  wire [31:0]       dataInMem_hi_lo_lo_hi_lo_hi_1 = {dataRegroupBySew_1_75, dataRegroupBySew_0_75, dataRegroupBySew_1_74, dataRegroupBySew_0_74};
  wire [63:0]       dataInMem_hi_lo_lo_hi_lo_1 = {dataInMem_hi_lo_lo_hi_lo_hi_1, dataInMem_hi_lo_lo_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_lo_hi_hi_lo_1 = {dataRegroupBySew_1_77, dataRegroupBySew_0_77, dataRegroupBySew_1_76, dataRegroupBySew_0_76};
  wire [31:0]       dataInMem_hi_lo_lo_hi_hi_hi_1 = {dataRegroupBySew_1_79, dataRegroupBySew_0_79, dataRegroupBySew_1_78, dataRegroupBySew_0_78};
  wire [63:0]       dataInMem_hi_lo_lo_hi_hi_1 = {dataInMem_hi_lo_lo_hi_hi_hi_1, dataInMem_hi_lo_lo_hi_hi_lo_1};
  wire [127:0]      dataInMem_hi_lo_lo_hi_1 = {dataInMem_hi_lo_lo_hi_hi_1, dataInMem_hi_lo_lo_hi_lo_1};
  wire [255:0]      dataInMem_hi_lo_lo_1 = {dataInMem_hi_lo_lo_hi_1, dataInMem_hi_lo_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_hi_lo_lo_lo_1 = {dataRegroupBySew_1_81, dataRegroupBySew_0_81, dataRegroupBySew_1_80, dataRegroupBySew_0_80};
  wire [31:0]       dataInMem_hi_lo_hi_lo_lo_hi_1 = {dataRegroupBySew_1_83, dataRegroupBySew_0_83, dataRegroupBySew_1_82, dataRegroupBySew_0_82};
  wire [63:0]       dataInMem_hi_lo_hi_lo_lo_1 = {dataInMem_hi_lo_hi_lo_lo_hi_1, dataInMem_hi_lo_hi_lo_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_hi_lo_hi_lo_1 = {dataRegroupBySew_1_85, dataRegroupBySew_0_85, dataRegroupBySew_1_84, dataRegroupBySew_0_84};
  wire [31:0]       dataInMem_hi_lo_hi_lo_hi_hi_1 = {dataRegroupBySew_1_87, dataRegroupBySew_0_87, dataRegroupBySew_1_86, dataRegroupBySew_0_86};
  wire [63:0]       dataInMem_hi_lo_hi_lo_hi_1 = {dataInMem_hi_lo_hi_lo_hi_hi_1, dataInMem_hi_lo_hi_lo_hi_lo_1};
  wire [127:0]      dataInMem_hi_lo_hi_lo_1 = {dataInMem_hi_lo_hi_lo_hi_1, dataInMem_hi_lo_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_hi_hi_lo_lo_1 = {dataRegroupBySew_1_89, dataRegroupBySew_0_89, dataRegroupBySew_1_88, dataRegroupBySew_0_88};
  wire [31:0]       dataInMem_hi_lo_hi_hi_lo_hi_1 = {dataRegroupBySew_1_91, dataRegroupBySew_0_91, dataRegroupBySew_1_90, dataRegroupBySew_0_90};
  wire [63:0]       dataInMem_hi_lo_hi_hi_lo_1 = {dataInMem_hi_lo_hi_hi_lo_hi_1, dataInMem_hi_lo_hi_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_lo_hi_hi_hi_lo_1 = {dataRegroupBySew_1_93, dataRegroupBySew_0_93, dataRegroupBySew_1_92, dataRegroupBySew_0_92};
  wire [31:0]       dataInMem_hi_lo_hi_hi_hi_hi_1 = {dataRegroupBySew_1_95, dataRegroupBySew_0_95, dataRegroupBySew_1_94, dataRegroupBySew_0_94};
  wire [63:0]       dataInMem_hi_lo_hi_hi_hi_1 = {dataInMem_hi_lo_hi_hi_hi_hi_1, dataInMem_hi_lo_hi_hi_hi_lo_1};
  wire [127:0]      dataInMem_hi_lo_hi_hi_1 = {dataInMem_hi_lo_hi_hi_hi_1, dataInMem_hi_lo_hi_hi_lo_1};
  wire [255:0]      dataInMem_hi_lo_hi_1 = {dataInMem_hi_lo_hi_hi_1, dataInMem_hi_lo_hi_lo_1};
  wire [511:0]      dataInMem_hi_lo_1 = {dataInMem_hi_lo_hi_1, dataInMem_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_lo_lo_lo_lo_1 = {dataRegroupBySew_1_97, dataRegroupBySew_0_97, dataRegroupBySew_1_96, dataRegroupBySew_0_96};
  wire [31:0]       dataInMem_hi_hi_lo_lo_lo_hi_1 = {dataRegroupBySew_1_99, dataRegroupBySew_0_99, dataRegroupBySew_1_98, dataRegroupBySew_0_98};
  wire [63:0]       dataInMem_hi_hi_lo_lo_lo_1 = {dataInMem_hi_hi_lo_lo_lo_hi_1, dataInMem_hi_hi_lo_lo_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_lo_lo_hi_lo_1 = {dataRegroupBySew_1_101, dataRegroupBySew_0_101, dataRegroupBySew_1_100, dataRegroupBySew_0_100};
  wire [31:0]       dataInMem_hi_hi_lo_lo_hi_hi_1 = {dataRegroupBySew_1_103, dataRegroupBySew_0_103, dataRegroupBySew_1_102, dataRegroupBySew_0_102};
  wire [63:0]       dataInMem_hi_hi_lo_lo_hi_1 = {dataInMem_hi_hi_lo_lo_hi_hi_1, dataInMem_hi_hi_lo_lo_hi_lo_1};
  wire [127:0]      dataInMem_hi_hi_lo_lo_1 = {dataInMem_hi_hi_lo_lo_hi_1, dataInMem_hi_hi_lo_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_lo_hi_lo_lo_1 = {dataRegroupBySew_1_105, dataRegroupBySew_0_105, dataRegroupBySew_1_104, dataRegroupBySew_0_104};
  wire [31:0]       dataInMem_hi_hi_lo_hi_lo_hi_1 = {dataRegroupBySew_1_107, dataRegroupBySew_0_107, dataRegroupBySew_1_106, dataRegroupBySew_0_106};
  wire [63:0]       dataInMem_hi_hi_lo_hi_lo_1 = {dataInMem_hi_hi_lo_hi_lo_hi_1, dataInMem_hi_hi_lo_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_lo_hi_hi_lo_1 = {dataRegroupBySew_1_109, dataRegroupBySew_0_109, dataRegroupBySew_1_108, dataRegroupBySew_0_108};
  wire [31:0]       dataInMem_hi_hi_lo_hi_hi_hi_1 = {dataRegroupBySew_1_111, dataRegroupBySew_0_111, dataRegroupBySew_1_110, dataRegroupBySew_0_110};
  wire [63:0]       dataInMem_hi_hi_lo_hi_hi_1 = {dataInMem_hi_hi_lo_hi_hi_hi_1, dataInMem_hi_hi_lo_hi_hi_lo_1};
  wire [127:0]      dataInMem_hi_hi_lo_hi_1 = {dataInMem_hi_hi_lo_hi_hi_1, dataInMem_hi_hi_lo_hi_lo_1};
  wire [255:0]      dataInMem_hi_hi_lo_1 = {dataInMem_hi_hi_lo_hi_1, dataInMem_hi_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_hi_lo_lo_lo_1 = {dataRegroupBySew_1_113, dataRegroupBySew_0_113, dataRegroupBySew_1_112, dataRegroupBySew_0_112};
  wire [31:0]       dataInMem_hi_hi_hi_lo_lo_hi_1 = {dataRegroupBySew_1_115, dataRegroupBySew_0_115, dataRegroupBySew_1_114, dataRegroupBySew_0_114};
  wire [63:0]       dataInMem_hi_hi_hi_lo_lo_1 = {dataInMem_hi_hi_hi_lo_lo_hi_1, dataInMem_hi_hi_hi_lo_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_hi_lo_hi_lo_1 = {dataRegroupBySew_1_117, dataRegroupBySew_0_117, dataRegroupBySew_1_116, dataRegroupBySew_0_116};
  wire [31:0]       dataInMem_hi_hi_hi_lo_hi_hi_1 = {dataRegroupBySew_1_119, dataRegroupBySew_0_119, dataRegroupBySew_1_118, dataRegroupBySew_0_118};
  wire [63:0]       dataInMem_hi_hi_hi_lo_hi_1 = {dataInMem_hi_hi_hi_lo_hi_hi_1, dataInMem_hi_hi_hi_lo_hi_lo_1};
  wire [127:0]      dataInMem_hi_hi_hi_lo_1 = {dataInMem_hi_hi_hi_lo_hi_1, dataInMem_hi_hi_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_hi_hi_lo_lo_1 = {dataRegroupBySew_1_121, dataRegroupBySew_0_121, dataRegroupBySew_1_120, dataRegroupBySew_0_120};
  wire [31:0]       dataInMem_hi_hi_hi_hi_lo_hi_1 = {dataRegroupBySew_1_123, dataRegroupBySew_0_123, dataRegroupBySew_1_122, dataRegroupBySew_0_122};
  wire [63:0]       dataInMem_hi_hi_hi_hi_lo_1 = {dataInMem_hi_hi_hi_hi_lo_hi_1, dataInMem_hi_hi_hi_hi_lo_lo_1};
  wire [31:0]       dataInMem_hi_hi_hi_hi_hi_lo_1 = {dataRegroupBySew_1_125, dataRegroupBySew_0_125, dataRegroupBySew_1_124, dataRegroupBySew_0_124};
  wire [31:0]       dataInMem_hi_hi_hi_hi_hi_hi_1 = {dataRegroupBySew_1_127, dataRegroupBySew_0_127, dataRegroupBySew_1_126, dataRegroupBySew_0_126};
  wire [63:0]       dataInMem_hi_hi_hi_hi_hi_1 = {dataInMem_hi_hi_hi_hi_hi_hi_1, dataInMem_hi_hi_hi_hi_hi_lo_1};
  wire [127:0]      dataInMem_hi_hi_hi_hi_1 = {dataInMem_hi_hi_hi_hi_hi_1, dataInMem_hi_hi_hi_hi_lo_1};
  wire [255:0]      dataInMem_hi_hi_hi_1 = {dataInMem_hi_hi_hi_hi_1, dataInMem_hi_hi_hi_lo_1};
  wire [511:0]      dataInMem_hi_hi_1 = {dataInMem_hi_hi_hi_1, dataInMem_hi_hi_lo_1};
  wire [1023:0]     dataInMem_hi_1 = {dataInMem_hi_hi_1, dataInMem_hi_lo_1};
  wire [2047:0]     dataInMem_1 = {dataInMem_hi_1, dataInMem_lo_1};
  wire [1023:0]     regroupCacheLine_1_0 = dataInMem_1[1023:0];
  wire [1023:0]     regroupCacheLine_1_1 = dataInMem_1[2047:1024];
  wire [1023:0]     res_8 = regroupCacheLine_1_0;
  wire [1023:0]     res_9 = regroupCacheLine_1_1;
  wire [2047:0]     lo_lo_1 = {res_9, res_8};
  wire [4095:0]     lo_1 = {2048'h0, lo_lo_1};
  wire [8191:0]     regroupLoadData_0_1 = {4096'h0, lo_1};
  wire [15:0]       _GEN_6 = {dataRegroupBySew_2_0, dataRegroupBySew_1_0};
  wire [15:0]       dataInMem_hi_2;
  assign dataInMem_hi_2 = _GEN_6;
  wire [15:0]       dataInMem_lo_hi_5;
  assign dataInMem_lo_hi_5 = _GEN_6;
  wire [15:0]       dataInMem_lo_hi_134;
  assign dataInMem_lo_hi_134 = _GEN_6;
  wire [15:0]       _GEN_7 = {dataRegroupBySew_2_1, dataRegroupBySew_1_1};
  wire [15:0]       dataInMem_hi_3;
  assign dataInMem_hi_3 = _GEN_7;
  wire [15:0]       dataInMem_lo_hi_6;
  assign dataInMem_lo_hi_6 = _GEN_7;
  wire [15:0]       dataInMem_lo_hi_135;
  assign dataInMem_lo_hi_135 = _GEN_7;
  wire [15:0]       _GEN_8 = {dataRegroupBySew_2_2, dataRegroupBySew_1_2};
  wire [15:0]       dataInMem_hi_4;
  assign dataInMem_hi_4 = _GEN_8;
  wire [15:0]       dataInMem_lo_hi_7;
  assign dataInMem_lo_hi_7 = _GEN_8;
  wire [15:0]       dataInMem_lo_hi_136;
  assign dataInMem_lo_hi_136 = _GEN_8;
  wire [15:0]       _GEN_9 = {dataRegroupBySew_2_3, dataRegroupBySew_1_3};
  wire [15:0]       dataInMem_hi_5;
  assign dataInMem_hi_5 = _GEN_9;
  wire [15:0]       dataInMem_lo_hi_8;
  assign dataInMem_lo_hi_8 = _GEN_9;
  wire [15:0]       dataInMem_lo_hi_137;
  assign dataInMem_lo_hi_137 = _GEN_9;
  wire [15:0]       _GEN_10 = {dataRegroupBySew_2_4, dataRegroupBySew_1_4};
  wire [15:0]       dataInMem_hi_6;
  assign dataInMem_hi_6 = _GEN_10;
  wire [15:0]       dataInMem_lo_hi_9;
  assign dataInMem_lo_hi_9 = _GEN_10;
  wire [15:0]       dataInMem_lo_hi_138;
  assign dataInMem_lo_hi_138 = _GEN_10;
  wire [15:0]       _GEN_11 = {dataRegroupBySew_2_5, dataRegroupBySew_1_5};
  wire [15:0]       dataInMem_hi_7;
  assign dataInMem_hi_7 = _GEN_11;
  wire [15:0]       dataInMem_lo_hi_10;
  assign dataInMem_lo_hi_10 = _GEN_11;
  wire [15:0]       dataInMem_lo_hi_139;
  assign dataInMem_lo_hi_139 = _GEN_11;
  wire [15:0]       _GEN_12 = {dataRegroupBySew_2_6, dataRegroupBySew_1_6};
  wire [15:0]       dataInMem_hi_8;
  assign dataInMem_hi_8 = _GEN_12;
  wire [15:0]       dataInMem_lo_hi_11;
  assign dataInMem_lo_hi_11 = _GEN_12;
  wire [15:0]       dataInMem_lo_hi_140;
  assign dataInMem_lo_hi_140 = _GEN_12;
  wire [15:0]       _GEN_13 = {dataRegroupBySew_2_7, dataRegroupBySew_1_7};
  wire [15:0]       dataInMem_hi_9;
  assign dataInMem_hi_9 = _GEN_13;
  wire [15:0]       dataInMem_lo_hi_12;
  assign dataInMem_lo_hi_12 = _GEN_13;
  wire [15:0]       dataInMem_lo_hi_141;
  assign dataInMem_lo_hi_141 = _GEN_13;
  wire [15:0]       _GEN_14 = {dataRegroupBySew_2_8, dataRegroupBySew_1_8};
  wire [15:0]       dataInMem_hi_10;
  assign dataInMem_hi_10 = _GEN_14;
  wire [15:0]       dataInMem_lo_hi_13;
  assign dataInMem_lo_hi_13 = _GEN_14;
  wire [15:0]       dataInMem_lo_hi_142;
  assign dataInMem_lo_hi_142 = _GEN_14;
  wire [15:0]       _GEN_15 = {dataRegroupBySew_2_9, dataRegroupBySew_1_9};
  wire [15:0]       dataInMem_hi_11;
  assign dataInMem_hi_11 = _GEN_15;
  wire [15:0]       dataInMem_lo_hi_14;
  assign dataInMem_lo_hi_14 = _GEN_15;
  wire [15:0]       dataInMem_lo_hi_143;
  assign dataInMem_lo_hi_143 = _GEN_15;
  wire [15:0]       _GEN_16 = {dataRegroupBySew_2_10, dataRegroupBySew_1_10};
  wire [15:0]       dataInMem_hi_12;
  assign dataInMem_hi_12 = _GEN_16;
  wire [15:0]       dataInMem_lo_hi_15;
  assign dataInMem_lo_hi_15 = _GEN_16;
  wire [15:0]       dataInMem_lo_hi_144;
  assign dataInMem_lo_hi_144 = _GEN_16;
  wire [15:0]       _GEN_17 = {dataRegroupBySew_2_11, dataRegroupBySew_1_11};
  wire [15:0]       dataInMem_hi_13;
  assign dataInMem_hi_13 = _GEN_17;
  wire [15:0]       dataInMem_lo_hi_16;
  assign dataInMem_lo_hi_16 = _GEN_17;
  wire [15:0]       dataInMem_lo_hi_145;
  assign dataInMem_lo_hi_145 = _GEN_17;
  wire [15:0]       _GEN_18 = {dataRegroupBySew_2_12, dataRegroupBySew_1_12};
  wire [15:0]       dataInMem_hi_14;
  assign dataInMem_hi_14 = _GEN_18;
  wire [15:0]       dataInMem_lo_hi_17;
  assign dataInMem_lo_hi_17 = _GEN_18;
  wire [15:0]       dataInMem_lo_hi_146;
  assign dataInMem_lo_hi_146 = _GEN_18;
  wire [15:0]       _GEN_19 = {dataRegroupBySew_2_13, dataRegroupBySew_1_13};
  wire [15:0]       dataInMem_hi_15;
  assign dataInMem_hi_15 = _GEN_19;
  wire [15:0]       dataInMem_lo_hi_18;
  assign dataInMem_lo_hi_18 = _GEN_19;
  wire [15:0]       dataInMem_lo_hi_147;
  assign dataInMem_lo_hi_147 = _GEN_19;
  wire [15:0]       _GEN_20 = {dataRegroupBySew_2_14, dataRegroupBySew_1_14};
  wire [15:0]       dataInMem_hi_16;
  assign dataInMem_hi_16 = _GEN_20;
  wire [15:0]       dataInMem_lo_hi_19;
  assign dataInMem_lo_hi_19 = _GEN_20;
  wire [15:0]       dataInMem_lo_hi_148;
  assign dataInMem_lo_hi_148 = _GEN_20;
  wire [15:0]       _GEN_21 = {dataRegroupBySew_2_15, dataRegroupBySew_1_15};
  wire [15:0]       dataInMem_hi_17;
  assign dataInMem_hi_17 = _GEN_21;
  wire [15:0]       dataInMem_lo_hi_20;
  assign dataInMem_lo_hi_20 = _GEN_21;
  wire [15:0]       dataInMem_lo_hi_149;
  assign dataInMem_lo_hi_149 = _GEN_21;
  wire [15:0]       _GEN_22 = {dataRegroupBySew_2_16, dataRegroupBySew_1_16};
  wire [15:0]       dataInMem_hi_18;
  assign dataInMem_hi_18 = _GEN_22;
  wire [15:0]       dataInMem_lo_hi_21;
  assign dataInMem_lo_hi_21 = _GEN_22;
  wire [15:0]       dataInMem_lo_hi_150;
  assign dataInMem_lo_hi_150 = _GEN_22;
  wire [15:0]       _GEN_23 = {dataRegroupBySew_2_17, dataRegroupBySew_1_17};
  wire [15:0]       dataInMem_hi_19;
  assign dataInMem_hi_19 = _GEN_23;
  wire [15:0]       dataInMem_lo_hi_22;
  assign dataInMem_lo_hi_22 = _GEN_23;
  wire [15:0]       dataInMem_lo_hi_151;
  assign dataInMem_lo_hi_151 = _GEN_23;
  wire [15:0]       _GEN_24 = {dataRegroupBySew_2_18, dataRegroupBySew_1_18};
  wire [15:0]       dataInMem_hi_20;
  assign dataInMem_hi_20 = _GEN_24;
  wire [15:0]       dataInMem_lo_hi_23;
  assign dataInMem_lo_hi_23 = _GEN_24;
  wire [15:0]       dataInMem_lo_hi_152;
  assign dataInMem_lo_hi_152 = _GEN_24;
  wire [15:0]       _GEN_25 = {dataRegroupBySew_2_19, dataRegroupBySew_1_19};
  wire [15:0]       dataInMem_hi_21;
  assign dataInMem_hi_21 = _GEN_25;
  wire [15:0]       dataInMem_lo_hi_24;
  assign dataInMem_lo_hi_24 = _GEN_25;
  wire [15:0]       dataInMem_lo_hi_153;
  assign dataInMem_lo_hi_153 = _GEN_25;
  wire [15:0]       _GEN_26 = {dataRegroupBySew_2_20, dataRegroupBySew_1_20};
  wire [15:0]       dataInMem_hi_22;
  assign dataInMem_hi_22 = _GEN_26;
  wire [15:0]       dataInMem_lo_hi_25;
  assign dataInMem_lo_hi_25 = _GEN_26;
  wire [15:0]       dataInMem_lo_hi_154;
  assign dataInMem_lo_hi_154 = _GEN_26;
  wire [15:0]       _GEN_27 = {dataRegroupBySew_2_21, dataRegroupBySew_1_21};
  wire [15:0]       dataInMem_hi_23;
  assign dataInMem_hi_23 = _GEN_27;
  wire [15:0]       dataInMem_lo_hi_26;
  assign dataInMem_lo_hi_26 = _GEN_27;
  wire [15:0]       dataInMem_lo_hi_155;
  assign dataInMem_lo_hi_155 = _GEN_27;
  wire [15:0]       _GEN_28 = {dataRegroupBySew_2_22, dataRegroupBySew_1_22};
  wire [15:0]       dataInMem_hi_24;
  assign dataInMem_hi_24 = _GEN_28;
  wire [15:0]       dataInMem_lo_hi_27;
  assign dataInMem_lo_hi_27 = _GEN_28;
  wire [15:0]       dataInMem_lo_hi_156;
  assign dataInMem_lo_hi_156 = _GEN_28;
  wire [15:0]       _GEN_29 = {dataRegroupBySew_2_23, dataRegroupBySew_1_23};
  wire [15:0]       dataInMem_hi_25;
  assign dataInMem_hi_25 = _GEN_29;
  wire [15:0]       dataInMem_lo_hi_28;
  assign dataInMem_lo_hi_28 = _GEN_29;
  wire [15:0]       dataInMem_lo_hi_157;
  assign dataInMem_lo_hi_157 = _GEN_29;
  wire [15:0]       _GEN_30 = {dataRegroupBySew_2_24, dataRegroupBySew_1_24};
  wire [15:0]       dataInMem_hi_26;
  assign dataInMem_hi_26 = _GEN_30;
  wire [15:0]       dataInMem_lo_hi_29;
  assign dataInMem_lo_hi_29 = _GEN_30;
  wire [15:0]       dataInMem_lo_hi_158;
  assign dataInMem_lo_hi_158 = _GEN_30;
  wire [15:0]       _GEN_31 = {dataRegroupBySew_2_25, dataRegroupBySew_1_25};
  wire [15:0]       dataInMem_hi_27;
  assign dataInMem_hi_27 = _GEN_31;
  wire [15:0]       dataInMem_lo_hi_30;
  assign dataInMem_lo_hi_30 = _GEN_31;
  wire [15:0]       dataInMem_lo_hi_159;
  assign dataInMem_lo_hi_159 = _GEN_31;
  wire [15:0]       _GEN_32 = {dataRegroupBySew_2_26, dataRegroupBySew_1_26};
  wire [15:0]       dataInMem_hi_28;
  assign dataInMem_hi_28 = _GEN_32;
  wire [15:0]       dataInMem_lo_hi_31;
  assign dataInMem_lo_hi_31 = _GEN_32;
  wire [15:0]       dataInMem_lo_hi_160;
  assign dataInMem_lo_hi_160 = _GEN_32;
  wire [15:0]       _GEN_33 = {dataRegroupBySew_2_27, dataRegroupBySew_1_27};
  wire [15:0]       dataInMem_hi_29;
  assign dataInMem_hi_29 = _GEN_33;
  wire [15:0]       dataInMem_lo_hi_32;
  assign dataInMem_lo_hi_32 = _GEN_33;
  wire [15:0]       dataInMem_lo_hi_161;
  assign dataInMem_lo_hi_161 = _GEN_33;
  wire [15:0]       _GEN_34 = {dataRegroupBySew_2_28, dataRegroupBySew_1_28};
  wire [15:0]       dataInMem_hi_30;
  assign dataInMem_hi_30 = _GEN_34;
  wire [15:0]       dataInMem_lo_hi_33;
  assign dataInMem_lo_hi_33 = _GEN_34;
  wire [15:0]       dataInMem_lo_hi_162;
  assign dataInMem_lo_hi_162 = _GEN_34;
  wire [15:0]       _GEN_35 = {dataRegroupBySew_2_29, dataRegroupBySew_1_29};
  wire [15:0]       dataInMem_hi_31;
  assign dataInMem_hi_31 = _GEN_35;
  wire [15:0]       dataInMem_lo_hi_34;
  assign dataInMem_lo_hi_34 = _GEN_35;
  wire [15:0]       dataInMem_lo_hi_163;
  assign dataInMem_lo_hi_163 = _GEN_35;
  wire [15:0]       _GEN_36 = {dataRegroupBySew_2_30, dataRegroupBySew_1_30};
  wire [15:0]       dataInMem_hi_32;
  assign dataInMem_hi_32 = _GEN_36;
  wire [15:0]       dataInMem_lo_hi_35;
  assign dataInMem_lo_hi_35 = _GEN_36;
  wire [15:0]       dataInMem_lo_hi_164;
  assign dataInMem_lo_hi_164 = _GEN_36;
  wire [15:0]       _GEN_37 = {dataRegroupBySew_2_31, dataRegroupBySew_1_31};
  wire [15:0]       dataInMem_hi_33;
  assign dataInMem_hi_33 = _GEN_37;
  wire [15:0]       dataInMem_lo_hi_36;
  assign dataInMem_lo_hi_36 = _GEN_37;
  wire [15:0]       dataInMem_lo_hi_165;
  assign dataInMem_lo_hi_165 = _GEN_37;
  wire [15:0]       _GEN_38 = {dataRegroupBySew_2_32, dataRegroupBySew_1_32};
  wire [15:0]       dataInMem_hi_34;
  assign dataInMem_hi_34 = _GEN_38;
  wire [15:0]       dataInMem_lo_hi_37;
  assign dataInMem_lo_hi_37 = _GEN_38;
  wire [15:0]       dataInMem_lo_hi_166;
  assign dataInMem_lo_hi_166 = _GEN_38;
  wire [15:0]       _GEN_39 = {dataRegroupBySew_2_33, dataRegroupBySew_1_33};
  wire [15:0]       dataInMem_hi_35;
  assign dataInMem_hi_35 = _GEN_39;
  wire [15:0]       dataInMem_lo_hi_38;
  assign dataInMem_lo_hi_38 = _GEN_39;
  wire [15:0]       dataInMem_lo_hi_167;
  assign dataInMem_lo_hi_167 = _GEN_39;
  wire [15:0]       _GEN_40 = {dataRegroupBySew_2_34, dataRegroupBySew_1_34};
  wire [15:0]       dataInMem_hi_36;
  assign dataInMem_hi_36 = _GEN_40;
  wire [15:0]       dataInMem_lo_hi_39;
  assign dataInMem_lo_hi_39 = _GEN_40;
  wire [15:0]       dataInMem_lo_hi_168;
  assign dataInMem_lo_hi_168 = _GEN_40;
  wire [15:0]       _GEN_41 = {dataRegroupBySew_2_35, dataRegroupBySew_1_35};
  wire [15:0]       dataInMem_hi_37;
  assign dataInMem_hi_37 = _GEN_41;
  wire [15:0]       dataInMem_lo_hi_40;
  assign dataInMem_lo_hi_40 = _GEN_41;
  wire [15:0]       dataInMem_lo_hi_169;
  assign dataInMem_lo_hi_169 = _GEN_41;
  wire [15:0]       _GEN_42 = {dataRegroupBySew_2_36, dataRegroupBySew_1_36};
  wire [15:0]       dataInMem_hi_38;
  assign dataInMem_hi_38 = _GEN_42;
  wire [15:0]       dataInMem_lo_hi_41;
  assign dataInMem_lo_hi_41 = _GEN_42;
  wire [15:0]       dataInMem_lo_hi_170;
  assign dataInMem_lo_hi_170 = _GEN_42;
  wire [15:0]       _GEN_43 = {dataRegroupBySew_2_37, dataRegroupBySew_1_37};
  wire [15:0]       dataInMem_hi_39;
  assign dataInMem_hi_39 = _GEN_43;
  wire [15:0]       dataInMem_lo_hi_42;
  assign dataInMem_lo_hi_42 = _GEN_43;
  wire [15:0]       dataInMem_lo_hi_171;
  assign dataInMem_lo_hi_171 = _GEN_43;
  wire [15:0]       _GEN_44 = {dataRegroupBySew_2_38, dataRegroupBySew_1_38};
  wire [15:0]       dataInMem_hi_40;
  assign dataInMem_hi_40 = _GEN_44;
  wire [15:0]       dataInMem_lo_hi_43;
  assign dataInMem_lo_hi_43 = _GEN_44;
  wire [15:0]       dataInMem_lo_hi_172;
  assign dataInMem_lo_hi_172 = _GEN_44;
  wire [15:0]       _GEN_45 = {dataRegroupBySew_2_39, dataRegroupBySew_1_39};
  wire [15:0]       dataInMem_hi_41;
  assign dataInMem_hi_41 = _GEN_45;
  wire [15:0]       dataInMem_lo_hi_44;
  assign dataInMem_lo_hi_44 = _GEN_45;
  wire [15:0]       dataInMem_lo_hi_173;
  assign dataInMem_lo_hi_173 = _GEN_45;
  wire [15:0]       _GEN_46 = {dataRegroupBySew_2_40, dataRegroupBySew_1_40};
  wire [15:0]       dataInMem_hi_42;
  assign dataInMem_hi_42 = _GEN_46;
  wire [15:0]       dataInMem_lo_hi_45;
  assign dataInMem_lo_hi_45 = _GEN_46;
  wire [15:0]       dataInMem_lo_hi_174;
  assign dataInMem_lo_hi_174 = _GEN_46;
  wire [15:0]       _GEN_47 = {dataRegroupBySew_2_41, dataRegroupBySew_1_41};
  wire [15:0]       dataInMem_hi_43;
  assign dataInMem_hi_43 = _GEN_47;
  wire [15:0]       dataInMem_lo_hi_46;
  assign dataInMem_lo_hi_46 = _GEN_47;
  wire [15:0]       dataInMem_lo_hi_175;
  assign dataInMem_lo_hi_175 = _GEN_47;
  wire [15:0]       _GEN_48 = {dataRegroupBySew_2_42, dataRegroupBySew_1_42};
  wire [15:0]       dataInMem_hi_44;
  assign dataInMem_hi_44 = _GEN_48;
  wire [15:0]       dataInMem_lo_hi_47;
  assign dataInMem_lo_hi_47 = _GEN_48;
  wire [15:0]       dataInMem_lo_hi_176;
  assign dataInMem_lo_hi_176 = _GEN_48;
  wire [15:0]       _GEN_49 = {dataRegroupBySew_2_43, dataRegroupBySew_1_43};
  wire [15:0]       dataInMem_hi_45;
  assign dataInMem_hi_45 = _GEN_49;
  wire [15:0]       dataInMem_lo_hi_48;
  assign dataInMem_lo_hi_48 = _GEN_49;
  wire [15:0]       dataInMem_lo_hi_177;
  assign dataInMem_lo_hi_177 = _GEN_49;
  wire [15:0]       _GEN_50 = {dataRegroupBySew_2_44, dataRegroupBySew_1_44};
  wire [15:0]       dataInMem_hi_46;
  assign dataInMem_hi_46 = _GEN_50;
  wire [15:0]       dataInMem_lo_hi_49;
  assign dataInMem_lo_hi_49 = _GEN_50;
  wire [15:0]       dataInMem_lo_hi_178;
  assign dataInMem_lo_hi_178 = _GEN_50;
  wire [15:0]       _GEN_51 = {dataRegroupBySew_2_45, dataRegroupBySew_1_45};
  wire [15:0]       dataInMem_hi_47;
  assign dataInMem_hi_47 = _GEN_51;
  wire [15:0]       dataInMem_lo_hi_50;
  assign dataInMem_lo_hi_50 = _GEN_51;
  wire [15:0]       dataInMem_lo_hi_179;
  assign dataInMem_lo_hi_179 = _GEN_51;
  wire [15:0]       _GEN_52 = {dataRegroupBySew_2_46, dataRegroupBySew_1_46};
  wire [15:0]       dataInMem_hi_48;
  assign dataInMem_hi_48 = _GEN_52;
  wire [15:0]       dataInMem_lo_hi_51;
  assign dataInMem_lo_hi_51 = _GEN_52;
  wire [15:0]       dataInMem_lo_hi_180;
  assign dataInMem_lo_hi_180 = _GEN_52;
  wire [15:0]       _GEN_53 = {dataRegroupBySew_2_47, dataRegroupBySew_1_47};
  wire [15:0]       dataInMem_hi_49;
  assign dataInMem_hi_49 = _GEN_53;
  wire [15:0]       dataInMem_lo_hi_52;
  assign dataInMem_lo_hi_52 = _GEN_53;
  wire [15:0]       dataInMem_lo_hi_181;
  assign dataInMem_lo_hi_181 = _GEN_53;
  wire [15:0]       _GEN_54 = {dataRegroupBySew_2_48, dataRegroupBySew_1_48};
  wire [15:0]       dataInMem_hi_50;
  assign dataInMem_hi_50 = _GEN_54;
  wire [15:0]       dataInMem_lo_hi_53;
  assign dataInMem_lo_hi_53 = _GEN_54;
  wire [15:0]       dataInMem_lo_hi_182;
  assign dataInMem_lo_hi_182 = _GEN_54;
  wire [15:0]       _GEN_55 = {dataRegroupBySew_2_49, dataRegroupBySew_1_49};
  wire [15:0]       dataInMem_hi_51;
  assign dataInMem_hi_51 = _GEN_55;
  wire [15:0]       dataInMem_lo_hi_54;
  assign dataInMem_lo_hi_54 = _GEN_55;
  wire [15:0]       dataInMem_lo_hi_183;
  assign dataInMem_lo_hi_183 = _GEN_55;
  wire [15:0]       _GEN_56 = {dataRegroupBySew_2_50, dataRegroupBySew_1_50};
  wire [15:0]       dataInMem_hi_52;
  assign dataInMem_hi_52 = _GEN_56;
  wire [15:0]       dataInMem_lo_hi_55;
  assign dataInMem_lo_hi_55 = _GEN_56;
  wire [15:0]       dataInMem_lo_hi_184;
  assign dataInMem_lo_hi_184 = _GEN_56;
  wire [15:0]       _GEN_57 = {dataRegroupBySew_2_51, dataRegroupBySew_1_51};
  wire [15:0]       dataInMem_hi_53;
  assign dataInMem_hi_53 = _GEN_57;
  wire [15:0]       dataInMem_lo_hi_56;
  assign dataInMem_lo_hi_56 = _GEN_57;
  wire [15:0]       dataInMem_lo_hi_185;
  assign dataInMem_lo_hi_185 = _GEN_57;
  wire [15:0]       _GEN_58 = {dataRegroupBySew_2_52, dataRegroupBySew_1_52};
  wire [15:0]       dataInMem_hi_54;
  assign dataInMem_hi_54 = _GEN_58;
  wire [15:0]       dataInMem_lo_hi_57;
  assign dataInMem_lo_hi_57 = _GEN_58;
  wire [15:0]       dataInMem_lo_hi_186;
  assign dataInMem_lo_hi_186 = _GEN_58;
  wire [15:0]       _GEN_59 = {dataRegroupBySew_2_53, dataRegroupBySew_1_53};
  wire [15:0]       dataInMem_hi_55;
  assign dataInMem_hi_55 = _GEN_59;
  wire [15:0]       dataInMem_lo_hi_58;
  assign dataInMem_lo_hi_58 = _GEN_59;
  wire [15:0]       dataInMem_lo_hi_187;
  assign dataInMem_lo_hi_187 = _GEN_59;
  wire [15:0]       _GEN_60 = {dataRegroupBySew_2_54, dataRegroupBySew_1_54};
  wire [15:0]       dataInMem_hi_56;
  assign dataInMem_hi_56 = _GEN_60;
  wire [15:0]       dataInMem_lo_hi_59;
  assign dataInMem_lo_hi_59 = _GEN_60;
  wire [15:0]       dataInMem_lo_hi_188;
  assign dataInMem_lo_hi_188 = _GEN_60;
  wire [15:0]       _GEN_61 = {dataRegroupBySew_2_55, dataRegroupBySew_1_55};
  wire [15:0]       dataInMem_hi_57;
  assign dataInMem_hi_57 = _GEN_61;
  wire [15:0]       dataInMem_lo_hi_60;
  assign dataInMem_lo_hi_60 = _GEN_61;
  wire [15:0]       dataInMem_lo_hi_189;
  assign dataInMem_lo_hi_189 = _GEN_61;
  wire [15:0]       _GEN_62 = {dataRegroupBySew_2_56, dataRegroupBySew_1_56};
  wire [15:0]       dataInMem_hi_58;
  assign dataInMem_hi_58 = _GEN_62;
  wire [15:0]       dataInMem_lo_hi_61;
  assign dataInMem_lo_hi_61 = _GEN_62;
  wire [15:0]       dataInMem_lo_hi_190;
  assign dataInMem_lo_hi_190 = _GEN_62;
  wire [15:0]       _GEN_63 = {dataRegroupBySew_2_57, dataRegroupBySew_1_57};
  wire [15:0]       dataInMem_hi_59;
  assign dataInMem_hi_59 = _GEN_63;
  wire [15:0]       dataInMem_lo_hi_62;
  assign dataInMem_lo_hi_62 = _GEN_63;
  wire [15:0]       dataInMem_lo_hi_191;
  assign dataInMem_lo_hi_191 = _GEN_63;
  wire [15:0]       _GEN_64 = {dataRegroupBySew_2_58, dataRegroupBySew_1_58};
  wire [15:0]       dataInMem_hi_60;
  assign dataInMem_hi_60 = _GEN_64;
  wire [15:0]       dataInMem_lo_hi_63;
  assign dataInMem_lo_hi_63 = _GEN_64;
  wire [15:0]       dataInMem_lo_hi_192;
  assign dataInMem_lo_hi_192 = _GEN_64;
  wire [15:0]       _GEN_65 = {dataRegroupBySew_2_59, dataRegroupBySew_1_59};
  wire [15:0]       dataInMem_hi_61;
  assign dataInMem_hi_61 = _GEN_65;
  wire [15:0]       dataInMem_lo_hi_64;
  assign dataInMem_lo_hi_64 = _GEN_65;
  wire [15:0]       dataInMem_lo_hi_193;
  assign dataInMem_lo_hi_193 = _GEN_65;
  wire [15:0]       _GEN_66 = {dataRegroupBySew_2_60, dataRegroupBySew_1_60};
  wire [15:0]       dataInMem_hi_62;
  assign dataInMem_hi_62 = _GEN_66;
  wire [15:0]       dataInMem_lo_hi_65;
  assign dataInMem_lo_hi_65 = _GEN_66;
  wire [15:0]       dataInMem_lo_hi_194;
  assign dataInMem_lo_hi_194 = _GEN_66;
  wire [15:0]       _GEN_67 = {dataRegroupBySew_2_61, dataRegroupBySew_1_61};
  wire [15:0]       dataInMem_hi_63;
  assign dataInMem_hi_63 = _GEN_67;
  wire [15:0]       dataInMem_lo_hi_66;
  assign dataInMem_lo_hi_66 = _GEN_67;
  wire [15:0]       dataInMem_lo_hi_195;
  assign dataInMem_lo_hi_195 = _GEN_67;
  wire [15:0]       _GEN_68 = {dataRegroupBySew_2_62, dataRegroupBySew_1_62};
  wire [15:0]       dataInMem_hi_64;
  assign dataInMem_hi_64 = _GEN_68;
  wire [15:0]       dataInMem_lo_hi_67;
  assign dataInMem_lo_hi_67 = _GEN_68;
  wire [15:0]       dataInMem_lo_hi_196;
  assign dataInMem_lo_hi_196 = _GEN_68;
  wire [15:0]       _GEN_69 = {dataRegroupBySew_2_63, dataRegroupBySew_1_63};
  wire [15:0]       dataInMem_hi_65;
  assign dataInMem_hi_65 = _GEN_69;
  wire [15:0]       dataInMem_lo_hi_68;
  assign dataInMem_lo_hi_68 = _GEN_69;
  wire [15:0]       dataInMem_lo_hi_197;
  assign dataInMem_lo_hi_197 = _GEN_69;
  wire [15:0]       _GEN_70 = {dataRegroupBySew_2_64, dataRegroupBySew_1_64};
  wire [15:0]       dataInMem_hi_66;
  assign dataInMem_hi_66 = _GEN_70;
  wire [15:0]       dataInMem_lo_hi_69;
  assign dataInMem_lo_hi_69 = _GEN_70;
  wire [15:0]       dataInMem_lo_hi_198;
  assign dataInMem_lo_hi_198 = _GEN_70;
  wire [15:0]       _GEN_71 = {dataRegroupBySew_2_65, dataRegroupBySew_1_65};
  wire [15:0]       dataInMem_hi_67;
  assign dataInMem_hi_67 = _GEN_71;
  wire [15:0]       dataInMem_lo_hi_70;
  assign dataInMem_lo_hi_70 = _GEN_71;
  wire [15:0]       dataInMem_lo_hi_199;
  assign dataInMem_lo_hi_199 = _GEN_71;
  wire [15:0]       _GEN_72 = {dataRegroupBySew_2_66, dataRegroupBySew_1_66};
  wire [15:0]       dataInMem_hi_68;
  assign dataInMem_hi_68 = _GEN_72;
  wire [15:0]       dataInMem_lo_hi_71;
  assign dataInMem_lo_hi_71 = _GEN_72;
  wire [15:0]       dataInMem_lo_hi_200;
  assign dataInMem_lo_hi_200 = _GEN_72;
  wire [15:0]       _GEN_73 = {dataRegroupBySew_2_67, dataRegroupBySew_1_67};
  wire [15:0]       dataInMem_hi_69;
  assign dataInMem_hi_69 = _GEN_73;
  wire [15:0]       dataInMem_lo_hi_72;
  assign dataInMem_lo_hi_72 = _GEN_73;
  wire [15:0]       dataInMem_lo_hi_201;
  assign dataInMem_lo_hi_201 = _GEN_73;
  wire [15:0]       _GEN_74 = {dataRegroupBySew_2_68, dataRegroupBySew_1_68};
  wire [15:0]       dataInMem_hi_70;
  assign dataInMem_hi_70 = _GEN_74;
  wire [15:0]       dataInMem_lo_hi_73;
  assign dataInMem_lo_hi_73 = _GEN_74;
  wire [15:0]       dataInMem_lo_hi_202;
  assign dataInMem_lo_hi_202 = _GEN_74;
  wire [15:0]       _GEN_75 = {dataRegroupBySew_2_69, dataRegroupBySew_1_69};
  wire [15:0]       dataInMem_hi_71;
  assign dataInMem_hi_71 = _GEN_75;
  wire [15:0]       dataInMem_lo_hi_74;
  assign dataInMem_lo_hi_74 = _GEN_75;
  wire [15:0]       dataInMem_lo_hi_203;
  assign dataInMem_lo_hi_203 = _GEN_75;
  wire [15:0]       _GEN_76 = {dataRegroupBySew_2_70, dataRegroupBySew_1_70};
  wire [15:0]       dataInMem_hi_72;
  assign dataInMem_hi_72 = _GEN_76;
  wire [15:0]       dataInMem_lo_hi_75;
  assign dataInMem_lo_hi_75 = _GEN_76;
  wire [15:0]       dataInMem_lo_hi_204;
  assign dataInMem_lo_hi_204 = _GEN_76;
  wire [15:0]       _GEN_77 = {dataRegroupBySew_2_71, dataRegroupBySew_1_71};
  wire [15:0]       dataInMem_hi_73;
  assign dataInMem_hi_73 = _GEN_77;
  wire [15:0]       dataInMem_lo_hi_76;
  assign dataInMem_lo_hi_76 = _GEN_77;
  wire [15:0]       dataInMem_lo_hi_205;
  assign dataInMem_lo_hi_205 = _GEN_77;
  wire [15:0]       _GEN_78 = {dataRegroupBySew_2_72, dataRegroupBySew_1_72};
  wire [15:0]       dataInMem_hi_74;
  assign dataInMem_hi_74 = _GEN_78;
  wire [15:0]       dataInMem_lo_hi_77;
  assign dataInMem_lo_hi_77 = _GEN_78;
  wire [15:0]       dataInMem_lo_hi_206;
  assign dataInMem_lo_hi_206 = _GEN_78;
  wire [15:0]       _GEN_79 = {dataRegroupBySew_2_73, dataRegroupBySew_1_73};
  wire [15:0]       dataInMem_hi_75;
  assign dataInMem_hi_75 = _GEN_79;
  wire [15:0]       dataInMem_lo_hi_78;
  assign dataInMem_lo_hi_78 = _GEN_79;
  wire [15:0]       dataInMem_lo_hi_207;
  assign dataInMem_lo_hi_207 = _GEN_79;
  wire [15:0]       _GEN_80 = {dataRegroupBySew_2_74, dataRegroupBySew_1_74};
  wire [15:0]       dataInMem_hi_76;
  assign dataInMem_hi_76 = _GEN_80;
  wire [15:0]       dataInMem_lo_hi_79;
  assign dataInMem_lo_hi_79 = _GEN_80;
  wire [15:0]       dataInMem_lo_hi_208;
  assign dataInMem_lo_hi_208 = _GEN_80;
  wire [15:0]       _GEN_81 = {dataRegroupBySew_2_75, dataRegroupBySew_1_75};
  wire [15:0]       dataInMem_hi_77;
  assign dataInMem_hi_77 = _GEN_81;
  wire [15:0]       dataInMem_lo_hi_80;
  assign dataInMem_lo_hi_80 = _GEN_81;
  wire [15:0]       dataInMem_lo_hi_209;
  assign dataInMem_lo_hi_209 = _GEN_81;
  wire [15:0]       _GEN_82 = {dataRegroupBySew_2_76, dataRegroupBySew_1_76};
  wire [15:0]       dataInMem_hi_78;
  assign dataInMem_hi_78 = _GEN_82;
  wire [15:0]       dataInMem_lo_hi_81;
  assign dataInMem_lo_hi_81 = _GEN_82;
  wire [15:0]       dataInMem_lo_hi_210;
  assign dataInMem_lo_hi_210 = _GEN_82;
  wire [15:0]       _GEN_83 = {dataRegroupBySew_2_77, dataRegroupBySew_1_77};
  wire [15:0]       dataInMem_hi_79;
  assign dataInMem_hi_79 = _GEN_83;
  wire [15:0]       dataInMem_lo_hi_82;
  assign dataInMem_lo_hi_82 = _GEN_83;
  wire [15:0]       dataInMem_lo_hi_211;
  assign dataInMem_lo_hi_211 = _GEN_83;
  wire [15:0]       _GEN_84 = {dataRegroupBySew_2_78, dataRegroupBySew_1_78};
  wire [15:0]       dataInMem_hi_80;
  assign dataInMem_hi_80 = _GEN_84;
  wire [15:0]       dataInMem_lo_hi_83;
  assign dataInMem_lo_hi_83 = _GEN_84;
  wire [15:0]       dataInMem_lo_hi_212;
  assign dataInMem_lo_hi_212 = _GEN_84;
  wire [15:0]       _GEN_85 = {dataRegroupBySew_2_79, dataRegroupBySew_1_79};
  wire [15:0]       dataInMem_hi_81;
  assign dataInMem_hi_81 = _GEN_85;
  wire [15:0]       dataInMem_lo_hi_84;
  assign dataInMem_lo_hi_84 = _GEN_85;
  wire [15:0]       dataInMem_lo_hi_213;
  assign dataInMem_lo_hi_213 = _GEN_85;
  wire [15:0]       _GEN_86 = {dataRegroupBySew_2_80, dataRegroupBySew_1_80};
  wire [15:0]       dataInMem_hi_82;
  assign dataInMem_hi_82 = _GEN_86;
  wire [15:0]       dataInMem_lo_hi_85;
  assign dataInMem_lo_hi_85 = _GEN_86;
  wire [15:0]       dataInMem_lo_hi_214;
  assign dataInMem_lo_hi_214 = _GEN_86;
  wire [15:0]       _GEN_87 = {dataRegroupBySew_2_81, dataRegroupBySew_1_81};
  wire [15:0]       dataInMem_hi_83;
  assign dataInMem_hi_83 = _GEN_87;
  wire [15:0]       dataInMem_lo_hi_86;
  assign dataInMem_lo_hi_86 = _GEN_87;
  wire [15:0]       dataInMem_lo_hi_215;
  assign dataInMem_lo_hi_215 = _GEN_87;
  wire [15:0]       _GEN_88 = {dataRegroupBySew_2_82, dataRegroupBySew_1_82};
  wire [15:0]       dataInMem_hi_84;
  assign dataInMem_hi_84 = _GEN_88;
  wire [15:0]       dataInMem_lo_hi_87;
  assign dataInMem_lo_hi_87 = _GEN_88;
  wire [15:0]       dataInMem_lo_hi_216;
  assign dataInMem_lo_hi_216 = _GEN_88;
  wire [15:0]       _GEN_89 = {dataRegroupBySew_2_83, dataRegroupBySew_1_83};
  wire [15:0]       dataInMem_hi_85;
  assign dataInMem_hi_85 = _GEN_89;
  wire [15:0]       dataInMem_lo_hi_88;
  assign dataInMem_lo_hi_88 = _GEN_89;
  wire [15:0]       dataInMem_lo_hi_217;
  assign dataInMem_lo_hi_217 = _GEN_89;
  wire [15:0]       _GEN_90 = {dataRegroupBySew_2_84, dataRegroupBySew_1_84};
  wire [15:0]       dataInMem_hi_86;
  assign dataInMem_hi_86 = _GEN_90;
  wire [15:0]       dataInMem_lo_hi_89;
  assign dataInMem_lo_hi_89 = _GEN_90;
  wire [15:0]       dataInMem_lo_hi_218;
  assign dataInMem_lo_hi_218 = _GEN_90;
  wire [15:0]       _GEN_91 = {dataRegroupBySew_2_85, dataRegroupBySew_1_85};
  wire [15:0]       dataInMem_hi_87;
  assign dataInMem_hi_87 = _GEN_91;
  wire [15:0]       dataInMem_lo_hi_90;
  assign dataInMem_lo_hi_90 = _GEN_91;
  wire [15:0]       dataInMem_lo_hi_219;
  assign dataInMem_lo_hi_219 = _GEN_91;
  wire [15:0]       _GEN_92 = {dataRegroupBySew_2_86, dataRegroupBySew_1_86};
  wire [15:0]       dataInMem_hi_88;
  assign dataInMem_hi_88 = _GEN_92;
  wire [15:0]       dataInMem_lo_hi_91;
  assign dataInMem_lo_hi_91 = _GEN_92;
  wire [15:0]       dataInMem_lo_hi_220;
  assign dataInMem_lo_hi_220 = _GEN_92;
  wire [15:0]       _GEN_93 = {dataRegroupBySew_2_87, dataRegroupBySew_1_87};
  wire [15:0]       dataInMem_hi_89;
  assign dataInMem_hi_89 = _GEN_93;
  wire [15:0]       dataInMem_lo_hi_92;
  assign dataInMem_lo_hi_92 = _GEN_93;
  wire [15:0]       dataInMem_lo_hi_221;
  assign dataInMem_lo_hi_221 = _GEN_93;
  wire [15:0]       _GEN_94 = {dataRegroupBySew_2_88, dataRegroupBySew_1_88};
  wire [15:0]       dataInMem_hi_90;
  assign dataInMem_hi_90 = _GEN_94;
  wire [15:0]       dataInMem_lo_hi_93;
  assign dataInMem_lo_hi_93 = _GEN_94;
  wire [15:0]       dataInMem_lo_hi_222;
  assign dataInMem_lo_hi_222 = _GEN_94;
  wire [15:0]       _GEN_95 = {dataRegroupBySew_2_89, dataRegroupBySew_1_89};
  wire [15:0]       dataInMem_hi_91;
  assign dataInMem_hi_91 = _GEN_95;
  wire [15:0]       dataInMem_lo_hi_94;
  assign dataInMem_lo_hi_94 = _GEN_95;
  wire [15:0]       dataInMem_lo_hi_223;
  assign dataInMem_lo_hi_223 = _GEN_95;
  wire [15:0]       _GEN_96 = {dataRegroupBySew_2_90, dataRegroupBySew_1_90};
  wire [15:0]       dataInMem_hi_92;
  assign dataInMem_hi_92 = _GEN_96;
  wire [15:0]       dataInMem_lo_hi_95;
  assign dataInMem_lo_hi_95 = _GEN_96;
  wire [15:0]       dataInMem_lo_hi_224;
  assign dataInMem_lo_hi_224 = _GEN_96;
  wire [15:0]       _GEN_97 = {dataRegroupBySew_2_91, dataRegroupBySew_1_91};
  wire [15:0]       dataInMem_hi_93;
  assign dataInMem_hi_93 = _GEN_97;
  wire [15:0]       dataInMem_lo_hi_96;
  assign dataInMem_lo_hi_96 = _GEN_97;
  wire [15:0]       dataInMem_lo_hi_225;
  assign dataInMem_lo_hi_225 = _GEN_97;
  wire [15:0]       _GEN_98 = {dataRegroupBySew_2_92, dataRegroupBySew_1_92};
  wire [15:0]       dataInMem_hi_94;
  assign dataInMem_hi_94 = _GEN_98;
  wire [15:0]       dataInMem_lo_hi_97;
  assign dataInMem_lo_hi_97 = _GEN_98;
  wire [15:0]       dataInMem_lo_hi_226;
  assign dataInMem_lo_hi_226 = _GEN_98;
  wire [15:0]       _GEN_99 = {dataRegroupBySew_2_93, dataRegroupBySew_1_93};
  wire [15:0]       dataInMem_hi_95;
  assign dataInMem_hi_95 = _GEN_99;
  wire [15:0]       dataInMem_lo_hi_98;
  assign dataInMem_lo_hi_98 = _GEN_99;
  wire [15:0]       dataInMem_lo_hi_227;
  assign dataInMem_lo_hi_227 = _GEN_99;
  wire [15:0]       _GEN_100 = {dataRegroupBySew_2_94, dataRegroupBySew_1_94};
  wire [15:0]       dataInMem_hi_96;
  assign dataInMem_hi_96 = _GEN_100;
  wire [15:0]       dataInMem_lo_hi_99;
  assign dataInMem_lo_hi_99 = _GEN_100;
  wire [15:0]       dataInMem_lo_hi_228;
  assign dataInMem_lo_hi_228 = _GEN_100;
  wire [15:0]       _GEN_101 = {dataRegroupBySew_2_95, dataRegroupBySew_1_95};
  wire [15:0]       dataInMem_hi_97;
  assign dataInMem_hi_97 = _GEN_101;
  wire [15:0]       dataInMem_lo_hi_100;
  assign dataInMem_lo_hi_100 = _GEN_101;
  wire [15:0]       dataInMem_lo_hi_229;
  assign dataInMem_lo_hi_229 = _GEN_101;
  wire [15:0]       _GEN_102 = {dataRegroupBySew_2_96, dataRegroupBySew_1_96};
  wire [15:0]       dataInMem_hi_98;
  assign dataInMem_hi_98 = _GEN_102;
  wire [15:0]       dataInMem_lo_hi_101;
  assign dataInMem_lo_hi_101 = _GEN_102;
  wire [15:0]       dataInMem_lo_hi_230;
  assign dataInMem_lo_hi_230 = _GEN_102;
  wire [15:0]       _GEN_103 = {dataRegroupBySew_2_97, dataRegroupBySew_1_97};
  wire [15:0]       dataInMem_hi_99;
  assign dataInMem_hi_99 = _GEN_103;
  wire [15:0]       dataInMem_lo_hi_102;
  assign dataInMem_lo_hi_102 = _GEN_103;
  wire [15:0]       dataInMem_lo_hi_231;
  assign dataInMem_lo_hi_231 = _GEN_103;
  wire [15:0]       _GEN_104 = {dataRegroupBySew_2_98, dataRegroupBySew_1_98};
  wire [15:0]       dataInMem_hi_100;
  assign dataInMem_hi_100 = _GEN_104;
  wire [15:0]       dataInMem_lo_hi_103;
  assign dataInMem_lo_hi_103 = _GEN_104;
  wire [15:0]       dataInMem_lo_hi_232;
  assign dataInMem_lo_hi_232 = _GEN_104;
  wire [15:0]       _GEN_105 = {dataRegroupBySew_2_99, dataRegroupBySew_1_99};
  wire [15:0]       dataInMem_hi_101;
  assign dataInMem_hi_101 = _GEN_105;
  wire [15:0]       dataInMem_lo_hi_104;
  assign dataInMem_lo_hi_104 = _GEN_105;
  wire [15:0]       dataInMem_lo_hi_233;
  assign dataInMem_lo_hi_233 = _GEN_105;
  wire [15:0]       _GEN_106 = {dataRegroupBySew_2_100, dataRegroupBySew_1_100};
  wire [15:0]       dataInMem_hi_102;
  assign dataInMem_hi_102 = _GEN_106;
  wire [15:0]       dataInMem_lo_hi_105;
  assign dataInMem_lo_hi_105 = _GEN_106;
  wire [15:0]       dataInMem_lo_hi_234;
  assign dataInMem_lo_hi_234 = _GEN_106;
  wire [15:0]       _GEN_107 = {dataRegroupBySew_2_101, dataRegroupBySew_1_101};
  wire [15:0]       dataInMem_hi_103;
  assign dataInMem_hi_103 = _GEN_107;
  wire [15:0]       dataInMem_lo_hi_106;
  assign dataInMem_lo_hi_106 = _GEN_107;
  wire [15:0]       dataInMem_lo_hi_235;
  assign dataInMem_lo_hi_235 = _GEN_107;
  wire [15:0]       _GEN_108 = {dataRegroupBySew_2_102, dataRegroupBySew_1_102};
  wire [15:0]       dataInMem_hi_104;
  assign dataInMem_hi_104 = _GEN_108;
  wire [15:0]       dataInMem_lo_hi_107;
  assign dataInMem_lo_hi_107 = _GEN_108;
  wire [15:0]       dataInMem_lo_hi_236;
  assign dataInMem_lo_hi_236 = _GEN_108;
  wire [15:0]       _GEN_109 = {dataRegroupBySew_2_103, dataRegroupBySew_1_103};
  wire [15:0]       dataInMem_hi_105;
  assign dataInMem_hi_105 = _GEN_109;
  wire [15:0]       dataInMem_lo_hi_108;
  assign dataInMem_lo_hi_108 = _GEN_109;
  wire [15:0]       dataInMem_lo_hi_237;
  assign dataInMem_lo_hi_237 = _GEN_109;
  wire [15:0]       _GEN_110 = {dataRegroupBySew_2_104, dataRegroupBySew_1_104};
  wire [15:0]       dataInMem_hi_106;
  assign dataInMem_hi_106 = _GEN_110;
  wire [15:0]       dataInMem_lo_hi_109;
  assign dataInMem_lo_hi_109 = _GEN_110;
  wire [15:0]       dataInMem_lo_hi_238;
  assign dataInMem_lo_hi_238 = _GEN_110;
  wire [15:0]       _GEN_111 = {dataRegroupBySew_2_105, dataRegroupBySew_1_105};
  wire [15:0]       dataInMem_hi_107;
  assign dataInMem_hi_107 = _GEN_111;
  wire [15:0]       dataInMem_lo_hi_110;
  assign dataInMem_lo_hi_110 = _GEN_111;
  wire [15:0]       dataInMem_lo_hi_239;
  assign dataInMem_lo_hi_239 = _GEN_111;
  wire [15:0]       _GEN_112 = {dataRegroupBySew_2_106, dataRegroupBySew_1_106};
  wire [15:0]       dataInMem_hi_108;
  assign dataInMem_hi_108 = _GEN_112;
  wire [15:0]       dataInMem_lo_hi_111;
  assign dataInMem_lo_hi_111 = _GEN_112;
  wire [15:0]       dataInMem_lo_hi_240;
  assign dataInMem_lo_hi_240 = _GEN_112;
  wire [15:0]       _GEN_113 = {dataRegroupBySew_2_107, dataRegroupBySew_1_107};
  wire [15:0]       dataInMem_hi_109;
  assign dataInMem_hi_109 = _GEN_113;
  wire [15:0]       dataInMem_lo_hi_112;
  assign dataInMem_lo_hi_112 = _GEN_113;
  wire [15:0]       dataInMem_lo_hi_241;
  assign dataInMem_lo_hi_241 = _GEN_113;
  wire [15:0]       _GEN_114 = {dataRegroupBySew_2_108, dataRegroupBySew_1_108};
  wire [15:0]       dataInMem_hi_110;
  assign dataInMem_hi_110 = _GEN_114;
  wire [15:0]       dataInMem_lo_hi_113;
  assign dataInMem_lo_hi_113 = _GEN_114;
  wire [15:0]       dataInMem_lo_hi_242;
  assign dataInMem_lo_hi_242 = _GEN_114;
  wire [15:0]       _GEN_115 = {dataRegroupBySew_2_109, dataRegroupBySew_1_109};
  wire [15:0]       dataInMem_hi_111;
  assign dataInMem_hi_111 = _GEN_115;
  wire [15:0]       dataInMem_lo_hi_114;
  assign dataInMem_lo_hi_114 = _GEN_115;
  wire [15:0]       dataInMem_lo_hi_243;
  assign dataInMem_lo_hi_243 = _GEN_115;
  wire [15:0]       _GEN_116 = {dataRegroupBySew_2_110, dataRegroupBySew_1_110};
  wire [15:0]       dataInMem_hi_112;
  assign dataInMem_hi_112 = _GEN_116;
  wire [15:0]       dataInMem_lo_hi_115;
  assign dataInMem_lo_hi_115 = _GEN_116;
  wire [15:0]       dataInMem_lo_hi_244;
  assign dataInMem_lo_hi_244 = _GEN_116;
  wire [15:0]       _GEN_117 = {dataRegroupBySew_2_111, dataRegroupBySew_1_111};
  wire [15:0]       dataInMem_hi_113;
  assign dataInMem_hi_113 = _GEN_117;
  wire [15:0]       dataInMem_lo_hi_116;
  assign dataInMem_lo_hi_116 = _GEN_117;
  wire [15:0]       dataInMem_lo_hi_245;
  assign dataInMem_lo_hi_245 = _GEN_117;
  wire [15:0]       _GEN_118 = {dataRegroupBySew_2_112, dataRegroupBySew_1_112};
  wire [15:0]       dataInMem_hi_114;
  assign dataInMem_hi_114 = _GEN_118;
  wire [15:0]       dataInMem_lo_hi_117;
  assign dataInMem_lo_hi_117 = _GEN_118;
  wire [15:0]       dataInMem_lo_hi_246;
  assign dataInMem_lo_hi_246 = _GEN_118;
  wire [15:0]       _GEN_119 = {dataRegroupBySew_2_113, dataRegroupBySew_1_113};
  wire [15:0]       dataInMem_hi_115;
  assign dataInMem_hi_115 = _GEN_119;
  wire [15:0]       dataInMem_lo_hi_118;
  assign dataInMem_lo_hi_118 = _GEN_119;
  wire [15:0]       dataInMem_lo_hi_247;
  assign dataInMem_lo_hi_247 = _GEN_119;
  wire [15:0]       _GEN_120 = {dataRegroupBySew_2_114, dataRegroupBySew_1_114};
  wire [15:0]       dataInMem_hi_116;
  assign dataInMem_hi_116 = _GEN_120;
  wire [15:0]       dataInMem_lo_hi_119;
  assign dataInMem_lo_hi_119 = _GEN_120;
  wire [15:0]       dataInMem_lo_hi_248;
  assign dataInMem_lo_hi_248 = _GEN_120;
  wire [15:0]       _GEN_121 = {dataRegroupBySew_2_115, dataRegroupBySew_1_115};
  wire [15:0]       dataInMem_hi_117;
  assign dataInMem_hi_117 = _GEN_121;
  wire [15:0]       dataInMem_lo_hi_120;
  assign dataInMem_lo_hi_120 = _GEN_121;
  wire [15:0]       dataInMem_lo_hi_249;
  assign dataInMem_lo_hi_249 = _GEN_121;
  wire [15:0]       _GEN_122 = {dataRegroupBySew_2_116, dataRegroupBySew_1_116};
  wire [15:0]       dataInMem_hi_118;
  assign dataInMem_hi_118 = _GEN_122;
  wire [15:0]       dataInMem_lo_hi_121;
  assign dataInMem_lo_hi_121 = _GEN_122;
  wire [15:0]       dataInMem_lo_hi_250;
  assign dataInMem_lo_hi_250 = _GEN_122;
  wire [15:0]       _GEN_123 = {dataRegroupBySew_2_117, dataRegroupBySew_1_117};
  wire [15:0]       dataInMem_hi_119;
  assign dataInMem_hi_119 = _GEN_123;
  wire [15:0]       dataInMem_lo_hi_122;
  assign dataInMem_lo_hi_122 = _GEN_123;
  wire [15:0]       dataInMem_lo_hi_251;
  assign dataInMem_lo_hi_251 = _GEN_123;
  wire [15:0]       _GEN_124 = {dataRegroupBySew_2_118, dataRegroupBySew_1_118};
  wire [15:0]       dataInMem_hi_120;
  assign dataInMem_hi_120 = _GEN_124;
  wire [15:0]       dataInMem_lo_hi_123;
  assign dataInMem_lo_hi_123 = _GEN_124;
  wire [15:0]       dataInMem_lo_hi_252;
  assign dataInMem_lo_hi_252 = _GEN_124;
  wire [15:0]       _GEN_125 = {dataRegroupBySew_2_119, dataRegroupBySew_1_119};
  wire [15:0]       dataInMem_hi_121;
  assign dataInMem_hi_121 = _GEN_125;
  wire [15:0]       dataInMem_lo_hi_124;
  assign dataInMem_lo_hi_124 = _GEN_125;
  wire [15:0]       dataInMem_lo_hi_253;
  assign dataInMem_lo_hi_253 = _GEN_125;
  wire [15:0]       _GEN_126 = {dataRegroupBySew_2_120, dataRegroupBySew_1_120};
  wire [15:0]       dataInMem_hi_122;
  assign dataInMem_hi_122 = _GEN_126;
  wire [15:0]       dataInMem_lo_hi_125;
  assign dataInMem_lo_hi_125 = _GEN_126;
  wire [15:0]       dataInMem_lo_hi_254;
  assign dataInMem_lo_hi_254 = _GEN_126;
  wire [15:0]       _GEN_127 = {dataRegroupBySew_2_121, dataRegroupBySew_1_121};
  wire [15:0]       dataInMem_hi_123;
  assign dataInMem_hi_123 = _GEN_127;
  wire [15:0]       dataInMem_lo_hi_126;
  assign dataInMem_lo_hi_126 = _GEN_127;
  wire [15:0]       dataInMem_lo_hi_255;
  assign dataInMem_lo_hi_255 = _GEN_127;
  wire [15:0]       _GEN_128 = {dataRegroupBySew_2_122, dataRegroupBySew_1_122};
  wire [15:0]       dataInMem_hi_124;
  assign dataInMem_hi_124 = _GEN_128;
  wire [15:0]       dataInMem_lo_hi_127;
  assign dataInMem_lo_hi_127 = _GEN_128;
  wire [15:0]       dataInMem_lo_hi_256;
  assign dataInMem_lo_hi_256 = _GEN_128;
  wire [15:0]       _GEN_129 = {dataRegroupBySew_2_123, dataRegroupBySew_1_123};
  wire [15:0]       dataInMem_hi_125;
  assign dataInMem_hi_125 = _GEN_129;
  wire [15:0]       dataInMem_lo_hi_128;
  assign dataInMem_lo_hi_128 = _GEN_129;
  wire [15:0]       dataInMem_lo_hi_257;
  assign dataInMem_lo_hi_257 = _GEN_129;
  wire [15:0]       _GEN_130 = {dataRegroupBySew_2_124, dataRegroupBySew_1_124};
  wire [15:0]       dataInMem_hi_126;
  assign dataInMem_hi_126 = _GEN_130;
  wire [15:0]       dataInMem_lo_hi_129;
  assign dataInMem_lo_hi_129 = _GEN_130;
  wire [15:0]       dataInMem_lo_hi_258;
  assign dataInMem_lo_hi_258 = _GEN_130;
  wire [15:0]       _GEN_131 = {dataRegroupBySew_2_125, dataRegroupBySew_1_125};
  wire [15:0]       dataInMem_hi_127;
  assign dataInMem_hi_127 = _GEN_131;
  wire [15:0]       dataInMem_lo_hi_130;
  assign dataInMem_lo_hi_130 = _GEN_131;
  wire [15:0]       dataInMem_lo_hi_259;
  assign dataInMem_lo_hi_259 = _GEN_131;
  wire [15:0]       _GEN_132 = {dataRegroupBySew_2_126, dataRegroupBySew_1_126};
  wire [15:0]       dataInMem_hi_128;
  assign dataInMem_hi_128 = _GEN_132;
  wire [15:0]       dataInMem_lo_hi_131;
  assign dataInMem_lo_hi_131 = _GEN_132;
  wire [15:0]       dataInMem_lo_hi_260;
  assign dataInMem_lo_hi_260 = _GEN_132;
  wire [15:0]       _GEN_133 = {dataRegroupBySew_2_127, dataRegroupBySew_1_127};
  wire [15:0]       dataInMem_hi_129;
  assign dataInMem_hi_129 = _GEN_133;
  wire [15:0]       dataInMem_lo_hi_132;
  assign dataInMem_lo_hi_132 = _GEN_133;
  wire [15:0]       dataInMem_lo_hi_261;
  assign dataInMem_lo_hi_261 = _GEN_133;
  wire [47:0]       dataInMem_lo_lo_lo_lo_lo_lo_2 = {dataInMem_hi_3, dataRegroupBySew_0_1, dataInMem_hi_2, dataRegroupBySew_0_0};
  wire [47:0]       dataInMem_lo_lo_lo_lo_lo_hi_2 = {dataInMem_hi_5, dataRegroupBySew_0_3, dataInMem_hi_4, dataRegroupBySew_0_2};
  wire [95:0]       dataInMem_lo_lo_lo_lo_lo_2 = {dataInMem_lo_lo_lo_lo_lo_hi_2, dataInMem_lo_lo_lo_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_lo_lo_lo_hi_lo_2 = {dataInMem_hi_7, dataRegroupBySew_0_5, dataInMem_hi_6, dataRegroupBySew_0_4};
  wire [47:0]       dataInMem_lo_lo_lo_lo_hi_hi_2 = {dataInMem_hi_9, dataRegroupBySew_0_7, dataInMem_hi_8, dataRegroupBySew_0_6};
  wire [95:0]       dataInMem_lo_lo_lo_lo_hi_2 = {dataInMem_lo_lo_lo_lo_hi_hi_2, dataInMem_lo_lo_lo_lo_hi_lo_2};
  wire [191:0]      dataInMem_lo_lo_lo_lo_2 = {dataInMem_lo_lo_lo_lo_hi_2, dataInMem_lo_lo_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_lo_lo_hi_lo_lo_2 = {dataInMem_hi_11, dataRegroupBySew_0_9, dataInMem_hi_10, dataRegroupBySew_0_8};
  wire [47:0]       dataInMem_lo_lo_lo_hi_lo_hi_2 = {dataInMem_hi_13, dataRegroupBySew_0_11, dataInMem_hi_12, dataRegroupBySew_0_10};
  wire [95:0]       dataInMem_lo_lo_lo_hi_lo_2 = {dataInMem_lo_lo_lo_hi_lo_hi_2, dataInMem_lo_lo_lo_hi_lo_lo_2};
  wire [47:0]       dataInMem_lo_lo_lo_hi_hi_lo_2 = {dataInMem_hi_15, dataRegroupBySew_0_13, dataInMem_hi_14, dataRegroupBySew_0_12};
  wire [47:0]       dataInMem_lo_lo_lo_hi_hi_hi_2 = {dataInMem_hi_17, dataRegroupBySew_0_15, dataInMem_hi_16, dataRegroupBySew_0_14};
  wire [95:0]       dataInMem_lo_lo_lo_hi_hi_2 = {dataInMem_lo_lo_lo_hi_hi_hi_2, dataInMem_lo_lo_lo_hi_hi_lo_2};
  wire [191:0]      dataInMem_lo_lo_lo_hi_2 = {dataInMem_lo_lo_lo_hi_hi_2, dataInMem_lo_lo_lo_hi_lo_2};
  wire [383:0]      dataInMem_lo_lo_lo_2 = {dataInMem_lo_lo_lo_hi_2, dataInMem_lo_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_lo_hi_lo_lo_lo_2 = {dataInMem_hi_19, dataRegroupBySew_0_17, dataInMem_hi_18, dataRegroupBySew_0_16};
  wire [47:0]       dataInMem_lo_lo_hi_lo_lo_hi_2 = {dataInMem_hi_21, dataRegroupBySew_0_19, dataInMem_hi_20, dataRegroupBySew_0_18};
  wire [95:0]       dataInMem_lo_lo_hi_lo_lo_2 = {dataInMem_lo_lo_hi_lo_lo_hi_2, dataInMem_lo_lo_hi_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_lo_hi_lo_hi_lo_2 = {dataInMem_hi_23, dataRegroupBySew_0_21, dataInMem_hi_22, dataRegroupBySew_0_20};
  wire [47:0]       dataInMem_lo_lo_hi_lo_hi_hi_2 = {dataInMem_hi_25, dataRegroupBySew_0_23, dataInMem_hi_24, dataRegroupBySew_0_22};
  wire [95:0]       dataInMem_lo_lo_hi_lo_hi_2 = {dataInMem_lo_lo_hi_lo_hi_hi_2, dataInMem_lo_lo_hi_lo_hi_lo_2};
  wire [191:0]      dataInMem_lo_lo_hi_lo_2 = {dataInMem_lo_lo_hi_lo_hi_2, dataInMem_lo_lo_hi_lo_lo_2};
  wire [47:0]       dataInMem_lo_lo_hi_hi_lo_lo_2 = {dataInMem_hi_27, dataRegroupBySew_0_25, dataInMem_hi_26, dataRegroupBySew_0_24};
  wire [47:0]       dataInMem_lo_lo_hi_hi_lo_hi_2 = {dataInMem_hi_29, dataRegroupBySew_0_27, dataInMem_hi_28, dataRegroupBySew_0_26};
  wire [95:0]       dataInMem_lo_lo_hi_hi_lo_2 = {dataInMem_lo_lo_hi_hi_lo_hi_2, dataInMem_lo_lo_hi_hi_lo_lo_2};
  wire [47:0]       dataInMem_lo_lo_hi_hi_hi_lo_2 = {dataInMem_hi_31, dataRegroupBySew_0_29, dataInMem_hi_30, dataRegroupBySew_0_28};
  wire [47:0]       dataInMem_lo_lo_hi_hi_hi_hi_2 = {dataInMem_hi_33, dataRegroupBySew_0_31, dataInMem_hi_32, dataRegroupBySew_0_30};
  wire [95:0]       dataInMem_lo_lo_hi_hi_hi_2 = {dataInMem_lo_lo_hi_hi_hi_hi_2, dataInMem_lo_lo_hi_hi_hi_lo_2};
  wire [191:0]      dataInMem_lo_lo_hi_hi_2 = {dataInMem_lo_lo_hi_hi_hi_2, dataInMem_lo_lo_hi_hi_lo_2};
  wire [383:0]      dataInMem_lo_lo_hi_2 = {dataInMem_lo_lo_hi_hi_2, dataInMem_lo_lo_hi_lo_2};
  wire [767:0]      dataInMem_lo_lo_2 = {dataInMem_lo_lo_hi_2, dataInMem_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_lo_lo_lo_lo_2 = {dataInMem_hi_35, dataRegroupBySew_0_33, dataInMem_hi_34, dataRegroupBySew_0_32};
  wire [47:0]       dataInMem_lo_hi_lo_lo_lo_hi_2 = {dataInMem_hi_37, dataRegroupBySew_0_35, dataInMem_hi_36, dataRegroupBySew_0_34};
  wire [95:0]       dataInMem_lo_hi_lo_lo_lo_2 = {dataInMem_lo_hi_lo_lo_lo_hi_2, dataInMem_lo_hi_lo_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_lo_lo_hi_lo_2 = {dataInMem_hi_39, dataRegroupBySew_0_37, dataInMem_hi_38, dataRegroupBySew_0_36};
  wire [47:0]       dataInMem_lo_hi_lo_lo_hi_hi_2 = {dataInMem_hi_41, dataRegroupBySew_0_39, dataInMem_hi_40, dataRegroupBySew_0_38};
  wire [95:0]       dataInMem_lo_hi_lo_lo_hi_2 = {dataInMem_lo_hi_lo_lo_hi_hi_2, dataInMem_lo_hi_lo_lo_hi_lo_2};
  wire [191:0]      dataInMem_lo_hi_lo_lo_2 = {dataInMem_lo_hi_lo_lo_hi_2, dataInMem_lo_hi_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_lo_hi_lo_lo_2 = {dataInMem_hi_43, dataRegroupBySew_0_41, dataInMem_hi_42, dataRegroupBySew_0_40};
  wire [47:0]       dataInMem_lo_hi_lo_hi_lo_hi_2 = {dataInMem_hi_45, dataRegroupBySew_0_43, dataInMem_hi_44, dataRegroupBySew_0_42};
  wire [95:0]       dataInMem_lo_hi_lo_hi_lo_2 = {dataInMem_lo_hi_lo_hi_lo_hi_2, dataInMem_lo_hi_lo_hi_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_lo_hi_hi_lo_2 = {dataInMem_hi_47, dataRegroupBySew_0_45, dataInMem_hi_46, dataRegroupBySew_0_44};
  wire [47:0]       dataInMem_lo_hi_lo_hi_hi_hi_2 = {dataInMem_hi_49, dataRegroupBySew_0_47, dataInMem_hi_48, dataRegroupBySew_0_46};
  wire [95:0]       dataInMem_lo_hi_lo_hi_hi_2 = {dataInMem_lo_hi_lo_hi_hi_hi_2, dataInMem_lo_hi_lo_hi_hi_lo_2};
  wire [191:0]      dataInMem_lo_hi_lo_hi_2 = {dataInMem_lo_hi_lo_hi_hi_2, dataInMem_lo_hi_lo_hi_lo_2};
  wire [383:0]      dataInMem_lo_hi_lo_2 = {dataInMem_lo_hi_lo_hi_2, dataInMem_lo_hi_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_hi_lo_lo_lo_2 = {dataInMem_hi_51, dataRegroupBySew_0_49, dataInMem_hi_50, dataRegroupBySew_0_48};
  wire [47:0]       dataInMem_lo_hi_hi_lo_lo_hi_2 = {dataInMem_hi_53, dataRegroupBySew_0_51, dataInMem_hi_52, dataRegroupBySew_0_50};
  wire [95:0]       dataInMem_lo_hi_hi_lo_lo_2 = {dataInMem_lo_hi_hi_lo_lo_hi_2, dataInMem_lo_hi_hi_lo_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_hi_lo_hi_lo_2 = {dataInMem_hi_55, dataRegroupBySew_0_53, dataInMem_hi_54, dataRegroupBySew_0_52};
  wire [47:0]       dataInMem_lo_hi_hi_lo_hi_hi_2 = {dataInMem_hi_57, dataRegroupBySew_0_55, dataInMem_hi_56, dataRegroupBySew_0_54};
  wire [95:0]       dataInMem_lo_hi_hi_lo_hi_2 = {dataInMem_lo_hi_hi_lo_hi_hi_2, dataInMem_lo_hi_hi_lo_hi_lo_2};
  wire [191:0]      dataInMem_lo_hi_hi_lo_2 = {dataInMem_lo_hi_hi_lo_hi_2, dataInMem_lo_hi_hi_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_hi_hi_lo_lo_2 = {dataInMem_hi_59, dataRegroupBySew_0_57, dataInMem_hi_58, dataRegroupBySew_0_56};
  wire [47:0]       dataInMem_lo_hi_hi_hi_lo_hi_2 = {dataInMem_hi_61, dataRegroupBySew_0_59, dataInMem_hi_60, dataRegroupBySew_0_58};
  wire [95:0]       dataInMem_lo_hi_hi_hi_lo_2 = {dataInMem_lo_hi_hi_hi_lo_hi_2, dataInMem_lo_hi_hi_hi_lo_lo_2};
  wire [47:0]       dataInMem_lo_hi_hi_hi_hi_lo_2 = {dataInMem_hi_63, dataRegroupBySew_0_61, dataInMem_hi_62, dataRegroupBySew_0_60};
  wire [47:0]       dataInMem_lo_hi_hi_hi_hi_hi_2 = {dataInMem_hi_65, dataRegroupBySew_0_63, dataInMem_hi_64, dataRegroupBySew_0_62};
  wire [95:0]       dataInMem_lo_hi_hi_hi_hi_2 = {dataInMem_lo_hi_hi_hi_hi_hi_2, dataInMem_lo_hi_hi_hi_hi_lo_2};
  wire [191:0]      dataInMem_lo_hi_hi_hi_2 = {dataInMem_lo_hi_hi_hi_hi_2, dataInMem_lo_hi_hi_hi_lo_2};
  wire [383:0]      dataInMem_lo_hi_hi_2 = {dataInMem_lo_hi_hi_hi_2, dataInMem_lo_hi_hi_lo_2};
  wire [767:0]      dataInMem_lo_hi_2 = {dataInMem_lo_hi_hi_2, dataInMem_lo_hi_lo_2};
  wire [1535:0]     dataInMem_lo_2 = {dataInMem_lo_hi_2, dataInMem_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_lo_lo_lo_lo_2 = {dataInMem_hi_67, dataRegroupBySew_0_65, dataInMem_hi_66, dataRegroupBySew_0_64};
  wire [47:0]       dataInMem_hi_lo_lo_lo_lo_hi_2 = {dataInMem_hi_69, dataRegroupBySew_0_67, dataInMem_hi_68, dataRegroupBySew_0_66};
  wire [95:0]       dataInMem_hi_lo_lo_lo_lo_2 = {dataInMem_hi_lo_lo_lo_lo_hi_2, dataInMem_hi_lo_lo_lo_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_lo_lo_hi_lo_2 = {dataInMem_hi_71, dataRegroupBySew_0_69, dataInMem_hi_70, dataRegroupBySew_0_68};
  wire [47:0]       dataInMem_hi_lo_lo_lo_hi_hi_2 = {dataInMem_hi_73, dataRegroupBySew_0_71, dataInMem_hi_72, dataRegroupBySew_0_70};
  wire [95:0]       dataInMem_hi_lo_lo_lo_hi_2 = {dataInMem_hi_lo_lo_lo_hi_hi_2, dataInMem_hi_lo_lo_lo_hi_lo_2};
  wire [191:0]      dataInMem_hi_lo_lo_lo_2 = {dataInMem_hi_lo_lo_lo_hi_2, dataInMem_hi_lo_lo_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_lo_hi_lo_lo_2 = {dataInMem_hi_75, dataRegroupBySew_0_73, dataInMem_hi_74, dataRegroupBySew_0_72};
  wire [47:0]       dataInMem_hi_lo_lo_hi_lo_hi_2 = {dataInMem_hi_77, dataRegroupBySew_0_75, dataInMem_hi_76, dataRegroupBySew_0_74};
  wire [95:0]       dataInMem_hi_lo_lo_hi_lo_2 = {dataInMem_hi_lo_lo_hi_lo_hi_2, dataInMem_hi_lo_lo_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_lo_hi_hi_lo_2 = {dataInMem_hi_79, dataRegroupBySew_0_77, dataInMem_hi_78, dataRegroupBySew_0_76};
  wire [47:0]       dataInMem_hi_lo_lo_hi_hi_hi_2 = {dataInMem_hi_81, dataRegroupBySew_0_79, dataInMem_hi_80, dataRegroupBySew_0_78};
  wire [95:0]       dataInMem_hi_lo_lo_hi_hi_2 = {dataInMem_hi_lo_lo_hi_hi_hi_2, dataInMem_hi_lo_lo_hi_hi_lo_2};
  wire [191:0]      dataInMem_hi_lo_lo_hi_2 = {dataInMem_hi_lo_lo_hi_hi_2, dataInMem_hi_lo_lo_hi_lo_2};
  wire [383:0]      dataInMem_hi_lo_lo_2 = {dataInMem_hi_lo_lo_hi_2, dataInMem_hi_lo_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_hi_lo_lo_lo_2 = {dataInMem_hi_83, dataRegroupBySew_0_81, dataInMem_hi_82, dataRegroupBySew_0_80};
  wire [47:0]       dataInMem_hi_lo_hi_lo_lo_hi_2 = {dataInMem_hi_85, dataRegroupBySew_0_83, dataInMem_hi_84, dataRegroupBySew_0_82};
  wire [95:0]       dataInMem_hi_lo_hi_lo_lo_2 = {dataInMem_hi_lo_hi_lo_lo_hi_2, dataInMem_hi_lo_hi_lo_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_hi_lo_hi_lo_2 = {dataInMem_hi_87, dataRegroupBySew_0_85, dataInMem_hi_86, dataRegroupBySew_0_84};
  wire [47:0]       dataInMem_hi_lo_hi_lo_hi_hi_2 = {dataInMem_hi_89, dataRegroupBySew_0_87, dataInMem_hi_88, dataRegroupBySew_0_86};
  wire [95:0]       dataInMem_hi_lo_hi_lo_hi_2 = {dataInMem_hi_lo_hi_lo_hi_hi_2, dataInMem_hi_lo_hi_lo_hi_lo_2};
  wire [191:0]      dataInMem_hi_lo_hi_lo_2 = {dataInMem_hi_lo_hi_lo_hi_2, dataInMem_hi_lo_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_hi_hi_lo_lo_2 = {dataInMem_hi_91, dataRegroupBySew_0_89, dataInMem_hi_90, dataRegroupBySew_0_88};
  wire [47:0]       dataInMem_hi_lo_hi_hi_lo_hi_2 = {dataInMem_hi_93, dataRegroupBySew_0_91, dataInMem_hi_92, dataRegroupBySew_0_90};
  wire [95:0]       dataInMem_hi_lo_hi_hi_lo_2 = {dataInMem_hi_lo_hi_hi_lo_hi_2, dataInMem_hi_lo_hi_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_lo_hi_hi_hi_lo_2 = {dataInMem_hi_95, dataRegroupBySew_0_93, dataInMem_hi_94, dataRegroupBySew_0_92};
  wire [47:0]       dataInMem_hi_lo_hi_hi_hi_hi_2 = {dataInMem_hi_97, dataRegroupBySew_0_95, dataInMem_hi_96, dataRegroupBySew_0_94};
  wire [95:0]       dataInMem_hi_lo_hi_hi_hi_2 = {dataInMem_hi_lo_hi_hi_hi_hi_2, dataInMem_hi_lo_hi_hi_hi_lo_2};
  wire [191:0]      dataInMem_hi_lo_hi_hi_2 = {dataInMem_hi_lo_hi_hi_hi_2, dataInMem_hi_lo_hi_hi_lo_2};
  wire [383:0]      dataInMem_hi_lo_hi_2 = {dataInMem_hi_lo_hi_hi_2, dataInMem_hi_lo_hi_lo_2};
  wire [767:0]      dataInMem_hi_lo_2 = {dataInMem_hi_lo_hi_2, dataInMem_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_lo_lo_lo_lo_2 = {dataInMem_hi_99, dataRegroupBySew_0_97, dataInMem_hi_98, dataRegroupBySew_0_96};
  wire [47:0]       dataInMem_hi_hi_lo_lo_lo_hi_2 = {dataInMem_hi_101, dataRegroupBySew_0_99, dataInMem_hi_100, dataRegroupBySew_0_98};
  wire [95:0]       dataInMem_hi_hi_lo_lo_lo_2 = {dataInMem_hi_hi_lo_lo_lo_hi_2, dataInMem_hi_hi_lo_lo_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_lo_lo_hi_lo_2 = {dataInMem_hi_103, dataRegroupBySew_0_101, dataInMem_hi_102, dataRegroupBySew_0_100};
  wire [47:0]       dataInMem_hi_hi_lo_lo_hi_hi_2 = {dataInMem_hi_105, dataRegroupBySew_0_103, dataInMem_hi_104, dataRegroupBySew_0_102};
  wire [95:0]       dataInMem_hi_hi_lo_lo_hi_2 = {dataInMem_hi_hi_lo_lo_hi_hi_2, dataInMem_hi_hi_lo_lo_hi_lo_2};
  wire [191:0]      dataInMem_hi_hi_lo_lo_2 = {dataInMem_hi_hi_lo_lo_hi_2, dataInMem_hi_hi_lo_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_lo_hi_lo_lo_2 = {dataInMem_hi_107, dataRegroupBySew_0_105, dataInMem_hi_106, dataRegroupBySew_0_104};
  wire [47:0]       dataInMem_hi_hi_lo_hi_lo_hi_2 = {dataInMem_hi_109, dataRegroupBySew_0_107, dataInMem_hi_108, dataRegroupBySew_0_106};
  wire [95:0]       dataInMem_hi_hi_lo_hi_lo_2 = {dataInMem_hi_hi_lo_hi_lo_hi_2, dataInMem_hi_hi_lo_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_lo_hi_hi_lo_2 = {dataInMem_hi_111, dataRegroupBySew_0_109, dataInMem_hi_110, dataRegroupBySew_0_108};
  wire [47:0]       dataInMem_hi_hi_lo_hi_hi_hi_2 = {dataInMem_hi_113, dataRegroupBySew_0_111, dataInMem_hi_112, dataRegroupBySew_0_110};
  wire [95:0]       dataInMem_hi_hi_lo_hi_hi_2 = {dataInMem_hi_hi_lo_hi_hi_hi_2, dataInMem_hi_hi_lo_hi_hi_lo_2};
  wire [191:0]      dataInMem_hi_hi_lo_hi_2 = {dataInMem_hi_hi_lo_hi_hi_2, dataInMem_hi_hi_lo_hi_lo_2};
  wire [383:0]      dataInMem_hi_hi_lo_2 = {dataInMem_hi_hi_lo_hi_2, dataInMem_hi_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_hi_lo_lo_lo_2 = {dataInMem_hi_115, dataRegroupBySew_0_113, dataInMem_hi_114, dataRegroupBySew_0_112};
  wire [47:0]       dataInMem_hi_hi_hi_lo_lo_hi_2 = {dataInMem_hi_117, dataRegroupBySew_0_115, dataInMem_hi_116, dataRegroupBySew_0_114};
  wire [95:0]       dataInMem_hi_hi_hi_lo_lo_2 = {dataInMem_hi_hi_hi_lo_lo_hi_2, dataInMem_hi_hi_hi_lo_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_hi_lo_hi_lo_2 = {dataInMem_hi_119, dataRegroupBySew_0_117, dataInMem_hi_118, dataRegroupBySew_0_116};
  wire [47:0]       dataInMem_hi_hi_hi_lo_hi_hi_2 = {dataInMem_hi_121, dataRegroupBySew_0_119, dataInMem_hi_120, dataRegroupBySew_0_118};
  wire [95:0]       dataInMem_hi_hi_hi_lo_hi_2 = {dataInMem_hi_hi_hi_lo_hi_hi_2, dataInMem_hi_hi_hi_lo_hi_lo_2};
  wire [191:0]      dataInMem_hi_hi_hi_lo_2 = {dataInMem_hi_hi_hi_lo_hi_2, dataInMem_hi_hi_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_hi_hi_lo_lo_2 = {dataInMem_hi_123, dataRegroupBySew_0_121, dataInMem_hi_122, dataRegroupBySew_0_120};
  wire [47:0]       dataInMem_hi_hi_hi_hi_lo_hi_2 = {dataInMem_hi_125, dataRegroupBySew_0_123, dataInMem_hi_124, dataRegroupBySew_0_122};
  wire [95:0]       dataInMem_hi_hi_hi_hi_lo_2 = {dataInMem_hi_hi_hi_hi_lo_hi_2, dataInMem_hi_hi_hi_hi_lo_lo_2};
  wire [47:0]       dataInMem_hi_hi_hi_hi_hi_lo_2 = {dataInMem_hi_127, dataRegroupBySew_0_125, dataInMem_hi_126, dataRegroupBySew_0_124};
  wire [47:0]       dataInMem_hi_hi_hi_hi_hi_hi_2 = {dataInMem_hi_129, dataRegroupBySew_0_127, dataInMem_hi_128, dataRegroupBySew_0_126};
  wire [95:0]       dataInMem_hi_hi_hi_hi_hi_2 = {dataInMem_hi_hi_hi_hi_hi_hi_2, dataInMem_hi_hi_hi_hi_hi_lo_2};
  wire [191:0]      dataInMem_hi_hi_hi_hi_2 = {dataInMem_hi_hi_hi_hi_hi_2, dataInMem_hi_hi_hi_hi_lo_2};
  wire [383:0]      dataInMem_hi_hi_hi_2 = {dataInMem_hi_hi_hi_hi_2, dataInMem_hi_hi_hi_lo_2};
  wire [767:0]      dataInMem_hi_hi_2 = {dataInMem_hi_hi_hi_2, dataInMem_hi_hi_lo_2};
  wire [1535:0]     dataInMem_hi_130 = {dataInMem_hi_hi_2, dataInMem_hi_lo_2};
  wire [3071:0]     dataInMem_2 = {dataInMem_hi_130, dataInMem_lo_2};
  wire [1023:0]     regroupCacheLine_2_0 = dataInMem_2[1023:0];
  wire [1023:0]     regroupCacheLine_2_1 = dataInMem_2[2047:1024];
  wire [1023:0]     regroupCacheLine_2_2 = dataInMem_2[3071:2048];
  wire [1023:0]     res_16 = regroupCacheLine_2_0;
  wire [1023:0]     res_17 = regroupCacheLine_2_1;
  wire [1023:0]     res_18 = regroupCacheLine_2_2;
  wire [2047:0]     lo_lo_2 = {res_17, res_16};
  wire [2047:0]     lo_hi_2 = {1024'h0, res_18};
  wire [4095:0]     lo_2 = {lo_hi_2, lo_lo_2};
  wire [8191:0]     regroupLoadData_0_2 = {4096'h0, lo_2};
  wire [15:0]       _GEN_134 = {dataRegroupBySew_1_0, dataRegroupBySew_0_0};
  wire [15:0]       dataInMem_lo_3;
  assign dataInMem_lo_3 = _GEN_134;
  wire [15:0]       dataInMem_lo_132;
  assign dataInMem_lo_132 = _GEN_134;
  wire [15:0]       dataInMem_lo_lo_7;
  assign dataInMem_lo_lo_7 = _GEN_134;
  wire [15:0]       _GEN_135 = {dataRegroupBySew_3_0, dataRegroupBySew_2_0};
  wire [15:0]       dataInMem_hi_131;
  assign dataInMem_hi_131 = _GEN_135;
  wire [15:0]       dataInMem_lo_hi_263;
  assign dataInMem_lo_hi_263 = _GEN_135;
  wire [15:0]       _GEN_136 = {dataRegroupBySew_1_1, dataRegroupBySew_0_1};
  wire [15:0]       dataInMem_lo_4;
  assign dataInMem_lo_4 = _GEN_136;
  wire [15:0]       dataInMem_lo_133;
  assign dataInMem_lo_133 = _GEN_136;
  wire [15:0]       dataInMem_lo_lo_8;
  assign dataInMem_lo_lo_8 = _GEN_136;
  wire [15:0]       _GEN_137 = {dataRegroupBySew_3_1, dataRegroupBySew_2_1};
  wire [15:0]       dataInMem_hi_132;
  assign dataInMem_hi_132 = _GEN_137;
  wire [15:0]       dataInMem_lo_hi_264;
  assign dataInMem_lo_hi_264 = _GEN_137;
  wire [15:0]       _GEN_138 = {dataRegroupBySew_1_2, dataRegroupBySew_0_2};
  wire [15:0]       dataInMem_lo_5;
  assign dataInMem_lo_5 = _GEN_138;
  wire [15:0]       dataInMem_lo_134;
  assign dataInMem_lo_134 = _GEN_138;
  wire [15:0]       dataInMem_lo_lo_9;
  assign dataInMem_lo_lo_9 = _GEN_138;
  wire [15:0]       _GEN_139 = {dataRegroupBySew_3_2, dataRegroupBySew_2_2};
  wire [15:0]       dataInMem_hi_133;
  assign dataInMem_hi_133 = _GEN_139;
  wire [15:0]       dataInMem_lo_hi_265;
  assign dataInMem_lo_hi_265 = _GEN_139;
  wire [15:0]       _GEN_140 = {dataRegroupBySew_1_3, dataRegroupBySew_0_3};
  wire [15:0]       dataInMem_lo_6;
  assign dataInMem_lo_6 = _GEN_140;
  wire [15:0]       dataInMem_lo_135;
  assign dataInMem_lo_135 = _GEN_140;
  wire [15:0]       dataInMem_lo_lo_10;
  assign dataInMem_lo_lo_10 = _GEN_140;
  wire [15:0]       _GEN_141 = {dataRegroupBySew_3_3, dataRegroupBySew_2_3};
  wire [15:0]       dataInMem_hi_134;
  assign dataInMem_hi_134 = _GEN_141;
  wire [15:0]       dataInMem_lo_hi_266;
  assign dataInMem_lo_hi_266 = _GEN_141;
  wire [15:0]       _GEN_142 = {dataRegroupBySew_1_4, dataRegroupBySew_0_4};
  wire [15:0]       dataInMem_lo_7;
  assign dataInMem_lo_7 = _GEN_142;
  wire [15:0]       dataInMem_lo_136;
  assign dataInMem_lo_136 = _GEN_142;
  wire [15:0]       dataInMem_lo_lo_11;
  assign dataInMem_lo_lo_11 = _GEN_142;
  wire [15:0]       _GEN_143 = {dataRegroupBySew_3_4, dataRegroupBySew_2_4};
  wire [15:0]       dataInMem_hi_135;
  assign dataInMem_hi_135 = _GEN_143;
  wire [15:0]       dataInMem_lo_hi_267;
  assign dataInMem_lo_hi_267 = _GEN_143;
  wire [15:0]       _GEN_144 = {dataRegroupBySew_1_5, dataRegroupBySew_0_5};
  wire [15:0]       dataInMem_lo_8;
  assign dataInMem_lo_8 = _GEN_144;
  wire [15:0]       dataInMem_lo_137;
  assign dataInMem_lo_137 = _GEN_144;
  wire [15:0]       dataInMem_lo_lo_12;
  assign dataInMem_lo_lo_12 = _GEN_144;
  wire [15:0]       _GEN_145 = {dataRegroupBySew_3_5, dataRegroupBySew_2_5};
  wire [15:0]       dataInMem_hi_136;
  assign dataInMem_hi_136 = _GEN_145;
  wire [15:0]       dataInMem_lo_hi_268;
  assign dataInMem_lo_hi_268 = _GEN_145;
  wire [15:0]       _GEN_146 = {dataRegroupBySew_1_6, dataRegroupBySew_0_6};
  wire [15:0]       dataInMem_lo_9;
  assign dataInMem_lo_9 = _GEN_146;
  wire [15:0]       dataInMem_lo_138;
  assign dataInMem_lo_138 = _GEN_146;
  wire [15:0]       dataInMem_lo_lo_13;
  assign dataInMem_lo_lo_13 = _GEN_146;
  wire [15:0]       _GEN_147 = {dataRegroupBySew_3_6, dataRegroupBySew_2_6};
  wire [15:0]       dataInMem_hi_137;
  assign dataInMem_hi_137 = _GEN_147;
  wire [15:0]       dataInMem_lo_hi_269;
  assign dataInMem_lo_hi_269 = _GEN_147;
  wire [15:0]       _GEN_148 = {dataRegroupBySew_1_7, dataRegroupBySew_0_7};
  wire [15:0]       dataInMem_lo_10;
  assign dataInMem_lo_10 = _GEN_148;
  wire [15:0]       dataInMem_lo_139;
  assign dataInMem_lo_139 = _GEN_148;
  wire [15:0]       dataInMem_lo_lo_14;
  assign dataInMem_lo_lo_14 = _GEN_148;
  wire [15:0]       _GEN_149 = {dataRegroupBySew_3_7, dataRegroupBySew_2_7};
  wire [15:0]       dataInMem_hi_138;
  assign dataInMem_hi_138 = _GEN_149;
  wire [15:0]       dataInMem_lo_hi_270;
  assign dataInMem_lo_hi_270 = _GEN_149;
  wire [15:0]       _GEN_150 = {dataRegroupBySew_1_8, dataRegroupBySew_0_8};
  wire [15:0]       dataInMem_lo_11;
  assign dataInMem_lo_11 = _GEN_150;
  wire [15:0]       dataInMem_lo_140;
  assign dataInMem_lo_140 = _GEN_150;
  wire [15:0]       dataInMem_lo_lo_15;
  assign dataInMem_lo_lo_15 = _GEN_150;
  wire [15:0]       _GEN_151 = {dataRegroupBySew_3_8, dataRegroupBySew_2_8};
  wire [15:0]       dataInMem_hi_139;
  assign dataInMem_hi_139 = _GEN_151;
  wire [15:0]       dataInMem_lo_hi_271;
  assign dataInMem_lo_hi_271 = _GEN_151;
  wire [15:0]       _GEN_152 = {dataRegroupBySew_1_9, dataRegroupBySew_0_9};
  wire [15:0]       dataInMem_lo_12;
  assign dataInMem_lo_12 = _GEN_152;
  wire [15:0]       dataInMem_lo_141;
  assign dataInMem_lo_141 = _GEN_152;
  wire [15:0]       dataInMem_lo_lo_16;
  assign dataInMem_lo_lo_16 = _GEN_152;
  wire [15:0]       _GEN_153 = {dataRegroupBySew_3_9, dataRegroupBySew_2_9};
  wire [15:0]       dataInMem_hi_140;
  assign dataInMem_hi_140 = _GEN_153;
  wire [15:0]       dataInMem_lo_hi_272;
  assign dataInMem_lo_hi_272 = _GEN_153;
  wire [15:0]       _GEN_154 = {dataRegroupBySew_1_10, dataRegroupBySew_0_10};
  wire [15:0]       dataInMem_lo_13;
  assign dataInMem_lo_13 = _GEN_154;
  wire [15:0]       dataInMem_lo_142;
  assign dataInMem_lo_142 = _GEN_154;
  wire [15:0]       dataInMem_lo_lo_17;
  assign dataInMem_lo_lo_17 = _GEN_154;
  wire [15:0]       _GEN_155 = {dataRegroupBySew_3_10, dataRegroupBySew_2_10};
  wire [15:0]       dataInMem_hi_141;
  assign dataInMem_hi_141 = _GEN_155;
  wire [15:0]       dataInMem_lo_hi_273;
  assign dataInMem_lo_hi_273 = _GEN_155;
  wire [15:0]       _GEN_156 = {dataRegroupBySew_1_11, dataRegroupBySew_0_11};
  wire [15:0]       dataInMem_lo_14;
  assign dataInMem_lo_14 = _GEN_156;
  wire [15:0]       dataInMem_lo_143;
  assign dataInMem_lo_143 = _GEN_156;
  wire [15:0]       dataInMem_lo_lo_18;
  assign dataInMem_lo_lo_18 = _GEN_156;
  wire [15:0]       _GEN_157 = {dataRegroupBySew_3_11, dataRegroupBySew_2_11};
  wire [15:0]       dataInMem_hi_142;
  assign dataInMem_hi_142 = _GEN_157;
  wire [15:0]       dataInMem_lo_hi_274;
  assign dataInMem_lo_hi_274 = _GEN_157;
  wire [15:0]       _GEN_158 = {dataRegroupBySew_1_12, dataRegroupBySew_0_12};
  wire [15:0]       dataInMem_lo_15;
  assign dataInMem_lo_15 = _GEN_158;
  wire [15:0]       dataInMem_lo_144;
  assign dataInMem_lo_144 = _GEN_158;
  wire [15:0]       dataInMem_lo_lo_19;
  assign dataInMem_lo_lo_19 = _GEN_158;
  wire [15:0]       _GEN_159 = {dataRegroupBySew_3_12, dataRegroupBySew_2_12};
  wire [15:0]       dataInMem_hi_143;
  assign dataInMem_hi_143 = _GEN_159;
  wire [15:0]       dataInMem_lo_hi_275;
  assign dataInMem_lo_hi_275 = _GEN_159;
  wire [15:0]       _GEN_160 = {dataRegroupBySew_1_13, dataRegroupBySew_0_13};
  wire [15:0]       dataInMem_lo_16;
  assign dataInMem_lo_16 = _GEN_160;
  wire [15:0]       dataInMem_lo_145;
  assign dataInMem_lo_145 = _GEN_160;
  wire [15:0]       dataInMem_lo_lo_20;
  assign dataInMem_lo_lo_20 = _GEN_160;
  wire [15:0]       _GEN_161 = {dataRegroupBySew_3_13, dataRegroupBySew_2_13};
  wire [15:0]       dataInMem_hi_144;
  assign dataInMem_hi_144 = _GEN_161;
  wire [15:0]       dataInMem_lo_hi_276;
  assign dataInMem_lo_hi_276 = _GEN_161;
  wire [15:0]       _GEN_162 = {dataRegroupBySew_1_14, dataRegroupBySew_0_14};
  wire [15:0]       dataInMem_lo_17;
  assign dataInMem_lo_17 = _GEN_162;
  wire [15:0]       dataInMem_lo_146;
  assign dataInMem_lo_146 = _GEN_162;
  wire [15:0]       dataInMem_lo_lo_21;
  assign dataInMem_lo_lo_21 = _GEN_162;
  wire [15:0]       _GEN_163 = {dataRegroupBySew_3_14, dataRegroupBySew_2_14};
  wire [15:0]       dataInMem_hi_145;
  assign dataInMem_hi_145 = _GEN_163;
  wire [15:0]       dataInMem_lo_hi_277;
  assign dataInMem_lo_hi_277 = _GEN_163;
  wire [15:0]       _GEN_164 = {dataRegroupBySew_1_15, dataRegroupBySew_0_15};
  wire [15:0]       dataInMem_lo_18;
  assign dataInMem_lo_18 = _GEN_164;
  wire [15:0]       dataInMem_lo_147;
  assign dataInMem_lo_147 = _GEN_164;
  wire [15:0]       dataInMem_lo_lo_22;
  assign dataInMem_lo_lo_22 = _GEN_164;
  wire [15:0]       _GEN_165 = {dataRegroupBySew_3_15, dataRegroupBySew_2_15};
  wire [15:0]       dataInMem_hi_146;
  assign dataInMem_hi_146 = _GEN_165;
  wire [15:0]       dataInMem_lo_hi_278;
  assign dataInMem_lo_hi_278 = _GEN_165;
  wire [15:0]       _GEN_166 = {dataRegroupBySew_1_16, dataRegroupBySew_0_16};
  wire [15:0]       dataInMem_lo_19;
  assign dataInMem_lo_19 = _GEN_166;
  wire [15:0]       dataInMem_lo_148;
  assign dataInMem_lo_148 = _GEN_166;
  wire [15:0]       dataInMem_lo_lo_23;
  assign dataInMem_lo_lo_23 = _GEN_166;
  wire [15:0]       _GEN_167 = {dataRegroupBySew_3_16, dataRegroupBySew_2_16};
  wire [15:0]       dataInMem_hi_147;
  assign dataInMem_hi_147 = _GEN_167;
  wire [15:0]       dataInMem_lo_hi_279;
  assign dataInMem_lo_hi_279 = _GEN_167;
  wire [15:0]       _GEN_168 = {dataRegroupBySew_1_17, dataRegroupBySew_0_17};
  wire [15:0]       dataInMem_lo_20;
  assign dataInMem_lo_20 = _GEN_168;
  wire [15:0]       dataInMem_lo_149;
  assign dataInMem_lo_149 = _GEN_168;
  wire [15:0]       dataInMem_lo_lo_24;
  assign dataInMem_lo_lo_24 = _GEN_168;
  wire [15:0]       _GEN_169 = {dataRegroupBySew_3_17, dataRegroupBySew_2_17};
  wire [15:0]       dataInMem_hi_148;
  assign dataInMem_hi_148 = _GEN_169;
  wire [15:0]       dataInMem_lo_hi_280;
  assign dataInMem_lo_hi_280 = _GEN_169;
  wire [15:0]       _GEN_170 = {dataRegroupBySew_1_18, dataRegroupBySew_0_18};
  wire [15:0]       dataInMem_lo_21;
  assign dataInMem_lo_21 = _GEN_170;
  wire [15:0]       dataInMem_lo_150;
  assign dataInMem_lo_150 = _GEN_170;
  wire [15:0]       dataInMem_lo_lo_25;
  assign dataInMem_lo_lo_25 = _GEN_170;
  wire [15:0]       _GEN_171 = {dataRegroupBySew_3_18, dataRegroupBySew_2_18};
  wire [15:0]       dataInMem_hi_149;
  assign dataInMem_hi_149 = _GEN_171;
  wire [15:0]       dataInMem_lo_hi_281;
  assign dataInMem_lo_hi_281 = _GEN_171;
  wire [15:0]       _GEN_172 = {dataRegroupBySew_1_19, dataRegroupBySew_0_19};
  wire [15:0]       dataInMem_lo_22;
  assign dataInMem_lo_22 = _GEN_172;
  wire [15:0]       dataInMem_lo_151;
  assign dataInMem_lo_151 = _GEN_172;
  wire [15:0]       dataInMem_lo_lo_26;
  assign dataInMem_lo_lo_26 = _GEN_172;
  wire [15:0]       _GEN_173 = {dataRegroupBySew_3_19, dataRegroupBySew_2_19};
  wire [15:0]       dataInMem_hi_150;
  assign dataInMem_hi_150 = _GEN_173;
  wire [15:0]       dataInMem_lo_hi_282;
  assign dataInMem_lo_hi_282 = _GEN_173;
  wire [15:0]       _GEN_174 = {dataRegroupBySew_1_20, dataRegroupBySew_0_20};
  wire [15:0]       dataInMem_lo_23;
  assign dataInMem_lo_23 = _GEN_174;
  wire [15:0]       dataInMem_lo_152;
  assign dataInMem_lo_152 = _GEN_174;
  wire [15:0]       dataInMem_lo_lo_27;
  assign dataInMem_lo_lo_27 = _GEN_174;
  wire [15:0]       _GEN_175 = {dataRegroupBySew_3_20, dataRegroupBySew_2_20};
  wire [15:0]       dataInMem_hi_151;
  assign dataInMem_hi_151 = _GEN_175;
  wire [15:0]       dataInMem_lo_hi_283;
  assign dataInMem_lo_hi_283 = _GEN_175;
  wire [15:0]       _GEN_176 = {dataRegroupBySew_1_21, dataRegroupBySew_0_21};
  wire [15:0]       dataInMem_lo_24;
  assign dataInMem_lo_24 = _GEN_176;
  wire [15:0]       dataInMem_lo_153;
  assign dataInMem_lo_153 = _GEN_176;
  wire [15:0]       dataInMem_lo_lo_28;
  assign dataInMem_lo_lo_28 = _GEN_176;
  wire [15:0]       _GEN_177 = {dataRegroupBySew_3_21, dataRegroupBySew_2_21};
  wire [15:0]       dataInMem_hi_152;
  assign dataInMem_hi_152 = _GEN_177;
  wire [15:0]       dataInMem_lo_hi_284;
  assign dataInMem_lo_hi_284 = _GEN_177;
  wire [15:0]       _GEN_178 = {dataRegroupBySew_1_22, dataRegroupBySew_0_22};
  wire [15:0]       dataInMem_lo_25;
  assign dataInMem_lo_25 = _GEN_178;
  wire [15:0]       dataInMem_lo_154;
  assign dataInMem_lo_154 = _GEN_178;
  wire [15:0]       dataInMem_lo_lo_29;
  assign dataInMem_lo_lo_29 = _GEN_178;
  wire [15:0]       _GEN_179 = {dataRegroupBySew_3_22, dataRegroupBySew_2_22};
  wire [15:0]       dataInMem_hi_153;
  assign dataInMem_hi_153 = _GEN_179;
  wire [15:0]       dataInMem_lo_hi_285;
  assign dataInMem_lo_hi_285 = _GEN_179;
  wire [15:0]       _GEN_180 = {dataRegroupBySew_1_23, dataRegroupBySew_0_23};
  wire [15:0]       dataInMem_lo_26;
  assign dataInMem_lo_26 = _GEN_180;
  wire [15:0]       dataInMem_lo_155;
  assign dataInMem_lo_155 = _GEN_180;
  wire [15:0]       dataInMem_lo_lo_30;
  assign dataInMem_lo_lo_30 = _GEN_180;
  wire [15:0]       _GEN_181 = {dataRegroupBySew_3_23, dataRegroupBySew_2_23};
  wire [15:0]       dataInMem_hi_154;
  assign dataInMem_hi_154 = _GEN_181;
  wire [15:0]       dataInMem_lo_hi_286;
  assign dataInMem_lo_hi_286 = _GEN_181;
  wire [15:0]       _GEN_182 = {dataRegroupBySew_1_24, dataRegroupBySew_0_24};
  wire [15:0]       dataInMem_lo_27;
  assign dataInMem_lo_27 = _GEN_182;
  wire [15:0]       dataInMem_lo_156;
  assign dataInMem_lo_156 = _GEN_182;
  wire [15:0]       dataInMem_lo_lo_31;
  assign dataInMem_lo_lo_31 = _GEN_182;
  wire [15:0]       _GEN_183 = {dataRegroupBySew_3_24, dataRegroupBySew_2_24};
  wire [15:0]       dataInMem_hi_155;
  assign dataInMem_hi_155 = _GEN_183;
  wire [15:0]       dataInMem_lo_hi_287;
  assign dataInMem_lo_hi_287 = _GEN_183;
  wire [15:0]       _GEN_184 = {dataRegroupBySew_1_25, dataRegroupBySew_0_25};
  wire [15:0]       dataInMem_lo_28;
  assign dataInMem_lo_28 = _GEN_184;
  wire [15:0]       dataInMem_lo_157;
  assign dataInMem_lo_157 = _GEN_184;
  wire [15:0]       dataInMem_lo_lo_32;
  assign dataInMem_lo_lo_32 = _GEN_184;
  wire [15:0]       _GEN_185 = {dataRegroupBySew_3_25, dataRegroupBySew_2_25};
  wire [15:0]       dataInMem_hi_156;
  assign dataInMem_hi_156 = _GEN_185;
  wire [15:0]       dataInMem_lo_hi_288;
  assign dataInMem_lo_hi_288 = _GEN_185;
  wire [15:0]       _GEN_186 = {dataRegroupBySew_1_26, dataRegroupBySew_0_26};
  wire [15:0]       dataInMem_lo_29;
  assign dataInMem_lo_29 = _GEN_186;
  wire [15:0]       dataInMem_lo_158;
  assign dataInMem_lo_158 = _GEN_186;
  wire [15:0]       dataInMem_lo_lo_33;
  assign dataInMem_lo_lo_33 = _GEN_186;
  wire [15:0]       _GEN_187 = {dataRegroupBySew_3_26, dataRegroupBySew_2_26};
  wire [15:0]       dataInMem_hi_157;
  assign dataInMem_hi_157 = _GEN_187;
  wire [15:0]       dataInMem_lo_hi_289;
  assign dataInMem_lo_hi_289 = _GEN_187;
  wire [15:0]       _GEN_188 = {dataRegroupBySew_1_27, dataRegroupBySew_0_27};
  wire [15:0]       dataInMem_lo_30;
  assign dataInMem_lo_30 = _GEN_188;
  wire [15:0]       dataInMem_lo_159;
  assign dataInMem_lo_159 = _GEN_188;
  wire [15:0]       dataInMem_lo_lo_34;
  assign dataInMem_lo_lo_34 = _GEN_188;
  wire [15:0]       _GEN_189 = {dataRegroupBySew_3_27, dataRegroupBySew_2_27};
  wire [15:0]       dataInMem_hi_158;
  assign dataInMem_hi_158 = _GEN_189;
  wire [15:0]       dataInMem_lo_hi_290;
  assign dataInMem_lo_hi_290 = _GEN_189;
  wire [15:0]       _GEN_190 = {dataRegroupBySew_1_28, dataRegroupBySew_0_28};
  wire [15:0]       dataInMem_lo_31;
  assign dataInMem_lo_31 = _GEN_190;
  wire [15:0]       dataInMem_lo_160;
  assign dataInMem_lo_160 = _GEN_190;
  wire [15:0]       dataInMem_lo_lo_35;
  assign dataInMem_lo_lo_35 = _GEN_190;
  wire [15:0]       _GEN_191 = {dataRegroupBySew_3_28, dataRegroupBySew_2_28};
  wire [15:0]       dataInMem_hi_159;
  assign dataInMem_hi_159 = _GEN_191;
  wire [15:0]       dataInMem_lo_hi_291;
  assign dataInMem_lo_hi_291 = _GEN_191;
  wire [15:0]       _GEN_192 = {dataRegroupBySew_1_29, dataRegroupBySew_0_29};
  wire [15:0]       dataInMem_lo_32;
  assign dataInMem_lo_32 = _GEN_192;
  wire [15:0]       dataInMem_lo_161;
  assign dataInMem_lo_161 = _GEN_192;
  wire [15:0]       dataInMem_lo_lo_36;
  assign dataInMem_lo_lo_36 = _GEN_192;
  wire [15:0]       _GEN_193 = {dataRegroupBySew_3_29, dataRegroupBySew_2_29};
  wire [15:0]       dataInMem_hi_160;
  assign dataInMem_hi_160 = _GEN_193;
  wire [15:0]       dataInMem_lo_hi_292;
  assign dataInMem_lo_hi_292 = _GEN_193;
  wire [15:0]       _GEN_194 = {dataRegroupBySew_1_30, dataRegroupBySew_0_30};
  wire [15:0]       dataInMem_lo_33;
  assign dataInMem_lo_33 = _GEN_194;
  wire [15:0]       dataInMem_lo_162;
  assign dataInMem_lo_162 = _GEN_194;
  wire [15:0]       dataInMem_lo_lo_37;
  assign dataInMem_lo_lo_37 = _GEN_194;
  wire [15:0]       _GEN_195 = {dataRegroupBySew_3_30, dataRegroupBySew_2_30};
  wire [15:0]       dataInMem_hi_161;
  assign dataInMem_hi_161 = _GEN_195;
  wire [15:0]       dataInMem_lo_hi_293;
  assign dataInMem_lo_hi_293 = _GEN_195;
  wire [15:0]       _GEN_196 = {dataRegroupBySew_1_31, dataRegroupBySew_0_31};
  wire [15:0]       dataInMem_lo_34;
  assign dataInMem_lo_34 = _GEN_196;
  wire [15:0]       dataInMem_lo_163;
  assign dataInMem_lo_163 = _GEN_196;
  wire [15:0]       dataInMem_lo_lo_38;
  assign dataInMem_lo_lo_38 = _GEN_196;
  wire [15:0]       _GEN_197 = {dataRegroupBySew_3_31, dataRegroupBySew_2_31};
  wire [15:0]       dataInMem_hi_162;
  assign dataInMem_hi_162 = _GEN_197;
  wire [15:0]       dataInMem_lo_hi_294;
  assign dataInMem_lo_hi_294 = _GEN_197;
  wire [15:0]       _GEN_198 = {dataRegroupBySew_1_32, dataRegroupBySew_0_32};
  wire [15:0]       dataInMem_lo_35;
  assign dataInMem_lo_35 = _GEN_198;
  wire [15:0]       dataInMem_lo_164;
  assign dataInMem_lo_164 = _GEN_198;
  wire [15:0]       dataInMem_lo_lo_39;
  assign dataInMem_lo_lo_39 = _GEN_198;
  wire [15:0]       _GEN_199 = {dataRegroupBySew_3_32, dataRegroupBySew_2_32};
  wire [15:0]       dataInMem_hi_163;
  assign dataInMem_hi_163 = _GEN_199;
  wire [15:0]       dataInMem_lo_hi_295;
  assign dataInMem_lo_hi_295 = _GEN_199;
  wire [15:0]       _GEN_200 = {dataRegroupBySew_1_33, dataRegroupBySew_0_33};
  wire [15:0]       dataInMem_lo_36;
  assign dataInMem_lo_36 = _GEN_200;
  wire [15:0]       dataInMem_lo_165;
  assign dataInMem_lo_165 = _GEN_200;
  wire [15:0]       dataInMem_lo_lo_40;
  assign dataInMem_lo_lo_40 = _GEN_200;
  wire [15:0]       _GEN_201 = {dataRegroupBySew_3_33, dataRegroupBySew_2_33};
  wire [15:0]       dataInMem_hi_164;
  assign dataInMem_hi_164 = _GEN_201;
  wire [15:0]       dataInMem_lo_hi_296;
  assign dataInMem_lo_hi_296 = _GEN_201;
  wire [15:0]       _GEN_202 = {dataRegroupBySew_1_34, dataRegroupBySew_0_34};
  wire [15:0]       dataInMem_lo_37;
  assign dataInMem_lo_37 = _GEN_202;
  wire [15:0]       dataInMem_lo_166;
  assign dataInMem_lo_166 = _GEN_202;
  wire [15:0]       dataInMem_lo_lo_41;
  assign dataInMem_lo_lo_41 = _GEN_202;
  wire [15:0]       _GEN_203 = {dataRegroupBySew_3_34, dataRegroupBySew_2_34};
  wire [15:0]       dataInMem_hi_165;
  assign dataInMem_hi_165 = _GEN_203;
  wire [15:0]       dataInMem_lo_hi_297;
  assign dataInMem_lo_hi_297 = _GEN_203;
  wire [15:0]       _GEN_204 = {dataRegroupBySew_1_35, dataRegroupBySew_0_35};
  wire [15:0]       dataInMem_lo_38;
  assign dataInMem_lo_38 = _GEN_204;
  wire [15:0]       dataInMem_lo_167;
  assign dataInMem_lo_167 = _GEN_204;
  wire [15:0]       dataInMem_lo_lo_42;
  assign dataInMem_lo_lo_42 = _GEN_204;
  wire [15:0]       _GEN_205 = {dataRegroupBySew_3_35, dataRegroupBySew_2_35};
  wire [15:0]       dataInMem_hi_166;
  assign dataInMem_hi_166 = _GEN_205;
  wire [15:0]       dataInMem_lo_hi_298;
  assign dataInMem_lo_hi_298 = _GEN_205;
  wire [15:0]       _GEN_206 = {dataRegroupBySew_1_36, dataRegroupBySew_0_36};
  wire [15:0]       dataInMem_lo_39;
  assign dataInMem_lo_39 = _GEN_206;
  wire [15:0]       dataInMem_lo_168;
  assign dataInMem_lo_168 = _GEN_206;
  wire [15:0]       dataInMem_lo_lo_43;
  assign dataInMem_lo_lo_43 = _GEN_206;
  wire [15:0]       _GEN_207 = {dataRegroupBySew_3_36, dataRegroupBySew_2_36};
  wire [15:0]       dataInMem_hi_167;
  assign dataInMem_hi_167 = _GEN_207;
  wire [15:0]       dataInMem_lo_hi_299;
  assign dataInMem_lo_hi_299 = _GEN_207;
  wire [15:0]       _GEN_208 = {dataRegroupBySew_1_37, dataRegroupBySew_0_37};
  wire [15:0]       dataInMem_lo_40;
  assign dataInMem_lo_40 = _GEN_208;
  wire [15:0]       dataInMem_lo_169;
  assign dataInMem_lo_169 = _GEN_208;
  wire [15:0]       dataInMem_lo_lo_44;
  assign dataInMem_lo_lo_44 = _GEN_208;
  wire [15:0]       _GEN_209 = {dataRegroupBySew_3_37, dataRegroupBySew_2_37};
  wire [15:0]       dataInMem_hi_168;
  assign dataInMem_hi_168 = _GEN_209;
  wire [15:0]       dataInMem_lo_hi_300;
  assign dataInMem_lo_hi_300 = _GEN_209;
  wire [15:0]       _GEN_210 = {dataRegroupBySew_1_38, dataRegroupBySew_0_38};
  wire [15:0]       dataInMem_lo_41;
  assign dataInMem_lo_41 = _GEN_210;
  wire [15:0]       dataInMem_lo_170;
  assign dataInMem_lo_170 = _GEN_210;
  wire [15:0]       dataInMem_lo_lo_45;
  assign dataInMem_lo_lo_45 = _GEN_210;
  wire [15:0]       _GEN_211 = {dataRegroupBySew_3_38, dataRegroupBySew_2_38};
  wire [15:0]       dataInMem_hi_169;
  assign dataInMem_hi_169 = _GEN_211;
  wire [15:0]       dataInMem_lo_hi_301;
  assign dataInMem_lo_hi_301 = _GEN_211;
  wire [15:0]       _GEN_212 = {dataRegroupBySew_1_39, dataRegroupBySew_0_39};
  wire [15:0]       dataInMem_lo_42;
  assign dataInMem_lo_42 = _GEN_212;
  wire [15:0]       dataInMem_lo_171;
  assign dataInMem_lo_171 = _GEN_212;
  wire [15:0]       dataInMem_lo_lo_46;
  assign dataInMem_lo_lo_46 = _GEN_212;
  wire [15:0]       _GEN_213 = {dataRegroupBySew_3_39, dataRegroupBySew_2_39};
  wire [15:0]       dataInMem_hi_170;
  assign dataInMem_hi_170 = _GEN_213;
  wire [15:0]       dataInMem_lo_hi_302;
  assign dataInMem_lo_hi_302 = _GEN_213;
  wire [15:0]       _GEN_214 = {dataRegroupBySew_1_40, dataRegroupBySew_0_40};
  wire [15:0]       dataInMem_lo_43;
  assign dataInMem_lo_43 = _GEN_214;
  wire [15:0]       dataInMem_lo_172;
  assign dataInMem_lo_172 = _GEN_214;
  wire [15:0]       dataInMem_lo_lo_47;
  assign dataInMem_lo_lo_47 = _GEN_214;
  wire [15:0]       _GEN_215 = {dataRegroupBySew_3_40, dataRegroupBySew_2_40};
  wire [15:0]       dataInMem_hi_171;
  assign dataInMem_hi_171 = _GEN_215;
  wire [15:0]       dataInMem_lo_hi_303;
  assign dataInMem_lo_hi_303 = _GEN_215;
  wire [15:0]       _GEN_216 = {dataRegroupBySew_1_41, dataRegroupBySew_0_41};
  wire [15:0]       dataInMem_lo_44;
  assign dataInMem_lo_44 = _GEN_216;
  wire [15:0]       dataInMem_lo_173;
  assign dataInMem_lo_173 = _GEN_216;
  wire [15:0]       dataInMem_lo_lo_48;
  assign dataInMem_lo_lo_48 = _GEN_216;
  wire [15:0]       _GEN_217 = {dataRegroupBySew_3_41, dataRegroupBySew_2_41};
  wire [15:0]       dataInMem_hi_172;
  assign dataInMem_hi_172 = _GEN_217;
  wire [15:0]       dataInMem_lo_hi_304;
  assign dataInMem_lo_hi_304 = _GEN_217;
  wire [15:0]       _GEN_218 = {dataRegroupBySew_1_42, dataRegroupBySew_0_42};
  wire [15:0]       dataInMem_lo_45;
  assign dataInMem_lo_45 = _GEN_218;
  wire [15:0]       dataInMem_lo_174;
  assign dataInMem_lo_174 = _GEN_218;
  wire [15:0]       dataInMem_lo_lo_49;
  assign dataInMem_lo_lo_49 = _GEN_218;
  wire [15:0]       _GEN_219 = {dataRegroupBySew_3_42, dataRegroupBySew_2_42};
  wire [15:0]       dataInMem_hi_173;
  assign dataInMem_hi_173 = _GEN_219;
  wire [15:0]       dataInMem_lo_hi_305;
  assign dataInMem_lo_hi_305 = _GEN_219;
  wire [15:0]       _GEN_220 = {dataRegroupBySew_1_43, dataRegroupBySew_0_43};
  wire [15:0]       dataInMem_lo_46;
  assign dataInMem_lo_46 = _GEN_220;
  wire [15:0]       dataInMem_lo_175;
  assign dataInMem_lo_175 = _GEN_220;
  wire [15:0]       dataInMem_lo_lo_50;
  assign dataInMem_lo_lo_50 = _GEN_220;
  wire [15:0]       _GEN_221 = {dataRegroupBySew_3_43, dataRegroupBySew_2_43};
  wire [15:0]       dataInMem_hi_174;
  assign dataInMem_hi_174 = _GEN_221;
  wire [15:0]       dataInMem_lo_hi_306;
  assign dataInMem_lo_hi_306 = _GEN_221;
  wire [15:0]       _GEN_222 = {dataRegroupBySew_1_44, dataRegroupBySew_0_44};
  wire [15:0]       dataInMem_lo_47;
  assign dataInMem_lo_47 = _GEN_222;
  wire [15:0]       dataInMem_lo_176;
  assign dataInMem_lo_176 = _GEN_222;
  wire [15:0]       dataInMem_lo_lo_51;
  assign dataInMem_lo_lo_51 = _GEN_222;
  wire [15:0]       _GEN_223 = {dataRegroupBySew_3_44, dataRegroupBySew_2_44};
  wire [15:0]       dataInMem_hi_175;
  assign dataInMem_hi_175 = _GEN_223;
  wire [15:0]       dataInMem_lo_hi_307;
  assign dataInMem_lo_hi_307 = _GEN_223;
  wire [15:0]       _GEN_224 = {dataRegroupBySew_1_45, dataRegroupBySew_0_45};
  wire [15:0]       dataInMem_lo_48;
  assign dataInMem_lo_48 = _GEN_224;
  wire [15:0]       dataInMem_lo_177;
  assign dataInMem_lo_177 = _GEN_224;
  wire [15:0]       dataInMem_lo_lo_52;
  assign dataInMem_lo_lo_52 = _GEN_224;
  wire [15:0]       _GEN_225 = {dataRegroupBySew_3_45, dataRegroupBySew_2_45};
  wire [15:0]       dataInMem_hi_176;
  assign dataInMem_hi_176 = _GEN_225;
  wire [15:0]       dataInMem_lo_hi_308;
  assign dataInMem_lo_hi_308 = _GEN_225;
  wire [15:0]       _GEN_226 = {dataRegroupBySew_1_46, dataRegroupBySew_0_46};
  wire [15:0]       dataInMem_lo_49;
  assign dataInMem_lo_49 = _GEN_226;
  wire [15:0]       dataInMem_lo_178;
  assign dataInMem_lo_178 = _GEN_226;
  wire [15:0]       dataInMem_lo_lo_53;
  assign dataInMem_lo_lo_53 = _GEN_226;
  wire [15:0]       _GEN_227 = {dataRegroupBySew_3_46, dataRegroupBySew_2_46};
  wire [15:0]       dataInMem_hi_177;
  assign dataInMem_hi_177 = _GEN_227;
  wire [15:0]       dataInMem_lo_hi_309;
  assign dataInMem_lo_hi_309 = _GEN_227;
  wire [15:0]       _GEN_228 = {dataRegroupBySew_1_47, dataRegroupBySew_0_47};
  wire [15:0]       dataInMem_lo_50;
  assign dataInMem_lo_50 = _GEN_228;
  wire [15:0]       dataInMem_lo_179;
  assign dataInMem_lo_179 = _GEN_228;
  wire [15:0]       dataInMem_lo_lo_54;
  assign dataInMem_lo_lo_54 = _GEN_228;
  wire [15:0]       _GEN_229 = {dataRegroupBySew_3_47, dataRegroupBySew_2_47};
  wire [15:0]       dataInMem_hi_178;
  assign dataInMem_hi_178 = _GEN_229;
  wire [15:0]       dataInMem_lo_hi_310;
  assign dataInMem_lo_hi_310 = _GEN_229;
  wire [15:0]       _GEN_230 = {dataRegroupBySew_1_48, dataRegroupBySew_0_48};
  wire [15:0]       dataInMem_lo_51;
  assign dataInMem_lo_51 = _GEN_230;
  wire [15:0]       dataInMem_lo_180;
  assign dataInMem_lo_180 = _GEN_230;
  wire [15:0]       dataInMem_lo_lo_55;
  assign dataInMem_lo_lo_55 = _GEN_230;
  wire [15:0]       _GEN_231 = {dataRegroupBySew_3_48, dataRegroupBySew_2_48};
  wire [15:0]       dataInMem_hi_179;
  assign dataInMem_hi_179 = _GEN_231;
  wire [15:0]       dataInMem_lo_hi_311;
  assign dataInMem_lo_hi_311 = _GEN_231;
  wire [15:0]       _GEN_232 = {dataRegroupBySew_1_49, dataRegroupBySew_0_49};
  wire [15:0]       dataInMem_lo_52;
  assign dataInMem_lo_52 = _GEN_232;
  wire [15:0]       dataInMem_lo_181;
  assign dataInMem_lo_181 = _GEN_232;
  wire [15:0]       dataInMem_lo_lo_56;
  assign dataInMem_lo_lo_56 = _GEN_232;
  wire [15:0]       _GEN_233 = {dataRegroupBySew_3_49, dataRegroupBySew_2_49};
  wire [15:0]       dataInMem_hi_180;
  assign dataInMem_hi_180 = _GEN_233;
  wire [15:0]       dataInMem_lo_hi_312;
  assign dataInMem_lo_hi_312 = _GEN_233;
  wire [15:0]       _GEN_234 = {dataRegroupBySew_1_50, dataRegroupBySew_0_50};
  wire [15:0]       dataInMem_lo_53;
  assign dataInMem_lo_53 = _GEN_234;
  wire [15:0]       dataInMem_lo_182;
  assign dataInMem_lo_182 = _GEN_234;
  wire [15:0]       dataInMem_lo_lo_57;
  assign dataInMem_lo_lo_57 = _GEN_234;
  wire [15:0]       _GEN_235 = {dataRegroupBySew_3_50, dataRegroupBySew_2_50};
  wire [15:0]       dataInMem_hi_181;
  assign dataInMem_hi_181 = _GEN_235;
  wire [15:0]       dataInMem_lo_hi_313;
  assign dataInMem_lo_hi_313 = _GEN_235;
  wire [15:0]       _GEN_236 = {dataRegroupBySew_1_51, dataRegroupBySew_0_51};
  wire [15:0]       dataInMem_lo_54;
  assign dataInMem_lo_54 = _GEN_236;
  wire [15:0]       dataInMem_lo_183;
  assign dataInMem_lo_183 = _GEN_236;
  wire [15:0]       dataInMem_lo_lo_58;
  assign dataInMem_lo_lo_58 = _GEN_236;
  wire [15:0]       _GEN_237 = {dataRegroupBySew_3_51, dataRegroupBySew_2_51};
  wire [15:0]       dataInMem_hi_182;
  assign dataInMem_hi_182 = _GEN_237;
  wire [15:0]       dataInMem_lo_hi_314;
  assign dataInMem_lo_hi_314 = _GEN_237;
  wire [15:0]       _GEN_238 = {dataRegroupBySew_1_52, dataRegroupBySew_0_52};
  wire [15:0]       dataInMem_lo_55;
  assign dataInMem_lo_55 = _GEN_238;
  wire [15:0]       dataInMem_lo_184;
  assign dataInMem_lo_184 = _GEN_238;
  wire [15:0]       dataInMem_lo_lo_59;
  assign dataInMem_lo_lo_59 = _GEN_238;
  wire [15:0]       _GEN_239 = {dataRegroupBySew_3_52, dataRegroupBySew_2_52};
  wire [15:0]       dataInMem_hi_183;
  assign dataInMem_hi_183 = _GEN_239;
  wire [15:0]       dataInMem_lo_hi_315;
  assign dataInMem_lo_hi_315 = _GEN_239;
  wire [15:0]       _GEN_240 = {dataRegroupBySew_1_53, dataRegroupBySew_0_53};
  wire [15:0]       dataInMem_lo_56;
  assign dataInMem_lo_56 = _GEN_240;
  wire [15:0]       dataInMem_lo_185;
  assign dataInMem_lo_185 = _GEN_240;
  wire [15:0]       dataInMem_lo_lo_60;
  assign dataInMem_lo_lo_60 = _GEN_240;
  wire [15:0]       _GEN_241 = {dataRegroupBySew_3_53, dataRegroupBySew_2_53};
  wire [15:0]       dataInMem_hi_184;
  assign dataInMem_hi_184 = _GEN_241;
  wire [15:0]       dataInMem_lo_hi_316;
  assign dataInMem_lo_hi_316 = _GEN_241;
  wire [15:0]       _GEN_242 = {dataRegroupBySew_1_54, dataRegroupBySew_0_54};
  wire [15:0]       dataInMem_lo_57;
  assign dataInMem_lo_57 = _GEN_242;
  wire [15:0]       dataInMem_lo_186;
  assign dataInMem_lo_186 = _GEN_242;
  wire [15:0]       dataInMem_lo_lo_61;
  assign dataInMem_lo_lo_61 = _GEN_242;
  wire [15:0]       _GEN_243 = {dataRegroupBySew_3_54, dataRegroupBySew_2_54};
  wire [15:0]       dataInMem_hi_185;
  assign dataInMem_hi_185 = _GEN_243;
  wire [15:0]       dataInMem_lo_hi_317;
  assign dataInMem_lo_hi_317 = _GEN_243;
  wire [15:0]       _GEN_244 = {dataRegroupBySew_1_55, dataRegroupBySew_0_55};
  wire [15:0]       dataInMem_lo_58;
  assign dataInMem_lo_58 = _GEN_244;
  wire [15:0]       dataInMem_lo_187;
  assign dataInMem_lo_187 = _GEN_244;
  wire [15:0]       dataInMem_lo_lo_62;
  assign dataInMem_lo_lo_62 = _GEN_244;
  wire [15:0]       _GEN_245 = {dataRegroupBySew_3_55, dataRegroupBySew_2_55};
  wire [15:0]       dataInMem_hi_186;
  assign dataInMem_hi_186 = _GEN_245;
  wire [15:0]       dataInMem_lo_hi_318;
  assign dataInMem_lo_hi_318 = _GEN_245;
  wire [15:0]       _GEN_246 = {dataRegroupBySew_1_56, dataRegroupBySew_0_56};
  wire [15:0]       dataInMem_lo_59;
  assign dataInMem_lo_59 = _GEN_246;
  wire [15:0]       dataInMem_lo_188;
  assign dataInMem_lo_188 = _GEN_246;
  wire [15:0]       dataInMem_lo_lo_63;
  assign dataInMem_lo_lo_63 = _GEN_246;
  wire [15:0]       _GEN_247 = {dataRegroupBySew_3_56, dataRegroupBySew_2_56};
  wire [15:0]       dataInMem_hi_187;
  assign dataInMem_hi_187 = _GEN_247;
  wire [15:0]       dataInMem_lo_hi_319;
  assign dataInMem_lo_hi_319 = _GEN_247;
  wire [15:0]       _GEN_248 = {dataRegroupBySew_1_57, dataRegroupBySew_0_57};
  wire [15:0]       dataInMem_lo_60;
  assign dataInMem_lo_60 = _GEN_248;
  wire [15:0]       dataInMem_lo_189;
  assign dataInMem_lo_189 = _GEN_248;
  wire [15:0]       dataInMem_lo_lo_64;
  assign dataInMem_lo_lo_64 = _GEN_248;
  wire [15:0]       _GEN_249 = {dataRegroupBySew_3_57, dataRegroupBySew_2_57};
  wire [15:0]       dataInMem_hi_188;
  assign dataInMem_hi_188 = _GEN_249;
  wire [15:0]       dataInMem_lo_hi_320;
  assign dataInMem_lo_hi_320 = _GEN_249;
  wire [15:0]       _GEN_250 = {dataRegroupBySew_1_58, dataRegroupBySew_0_58};
  wire [15:0]       dataInMem_lo_61;
  assign dataInMem_lo_61 = _GEN_250;
  wire [15:0]       dataInMem_lo_190;
  assign dataInMem_lo_190 = _GEN_250;
  wire [15:0]       dataInMem_lo_lo_65;
  assign dataInMem_lo_lo_65 = _GEN_250;
  wire [15:0]       _GEN_251 = {dataRegroupBySew_3_58, dataRegroupBySew_2_58};
  wire [15:0]       dataInMem_hi_189;
  assign dataInMem_hi_189 = _GEN_251;
  wire [15:0]       dataInMem_lo_hi_321;
  assign dataInMem_lo_hi_321 = _GEN_251;
  wire [15:0]       _GEN_252 = {dataRegroupBySew_1_59, dataRegroupBySew_0_59};
  wire [15:0]       dataInMem_lo_62;
  assign dataInMem_lo_62 = _GEN_252;
  wire [15:0]       dataInMem_lo_191;
  assign dataInMem_lo_191 = _GEN_252;
  wire [15:0]       dataInMem_lo_lo_66;
  assign dataInMem_lo_lo_66 = _GEN_252;
  wire [15:0]       _GEN_253 = {dataRegroupBySew_3_59, dataRegroupBySew_2_59};
  wire [15:0]       dataInMem_hi_190;
  assign dataInMem_hi_190 = _GEN_253;
  wire [15:0]       dataInMem_lo_hi_322;
  assign dataInMem_lo_hi_322 = _GEN_253;
  wire [15:0]       _GEN_254 = {dataRegroupBySew_1_60, dataRegroupBySew_0_60};
  wire [15:0]       dataInMem_lo_63;
  assign dataInMem_lo_63 = _GEN_254;
  wire [15:0]       dataInMem_lo_192;
  assign dataInMem_lo_192 = _GEN_254;
  wire [15:0]       dataInMem_lo_lo_67;
  assign dataInMem_lo_lo_67 = _GEN_254;
  wire [15:0]       _GEN_255 = {dataRegroupBySew_3_60, dataRegroupBySew_2_60};
  wire [15:0]       dataInMem_hi_191;
  assign dataInMem_hi_191 = _GEN_255;
  wire [15:0]       dataInMem_lo_hi_323;
  assign dataInMem_lo_hi_323 = _GEN_255;
  wire [15:0]       _GEN_256 = {dataRegroupBySew_1_61, dataRegroupBySew_0_61};
  wire [15:0]       dataInMem_lo_64;
  assign dataInMem_lo_64 = _GEN_256;
  wire [15:0]       dataInMem_lo_193;
  assign dataInMem_lo_193 = _GEN_256;
  wire [15:0]       dataInMem_lo_lo_68;
  assign dataInMem_lo_lo_68 = _GEN_256;
  wire [15:0]       _GEN_257 = {dataRegroupBySew_3_61, dataRegroupBySew_2_61};
  wire [15:0]       dataInMem_hi_192;
  assign dataInMem_hi_192 = _GEN_257;
  wire [15:0]       dataInMem_lo_hi_324;
  assign dataInMem_lo_hi_324 = _GEN_257;
  wire [15:0]       _GEN_258 = {dataRegroupBySew_1_62, dataRegroupBySew_0_62};
  wire [15:0]       dataInMem_lo_65;
  assign dataInMem_lo_65 = _GEN_258;
  wire [15:0]       dataInMem_lo_194;
  assign dataInMem_lo_194 = _GEN_258;
  wire [15:0]       dataInMem_lo_lo_69;
  assign dataInMem_lo_lo_69 = _GEN_258;
  wire [15:0]       _GEN_259 = {dataRegroupBySew_3_62, dataRegroupBySew_2_62};
  wire [15:0]       dataInMem_hi_193;
  assign dataInMem_hi_193 = _GEN_259;
  wire [15:0]       dataInMem_lo_hi_325;
  assign dataInMem_lo_hi_325 = _GEN_259;
  wire [15:0]       _GEN_260 = {dataRegroupBySew_1_63, dataRegroupBySew_0_63};
  wire [15:0]       dataInMem_lo_66;
  assign dataInMem_lo_66 = _GEN_260;
  wire [15:0]       dataInMem_lo_195;
  assign dataInMem_lo_195 = _GEN_260;
  wire [15:0]       dataInMem_lo_lo_70;
  assign dataInMem_lo_lo_70 = _GEN_260;
  wire [15:0]       _GEN_261 = {dataRegroupBySew_3_63, dataRegroupBySew_2_63};
  wire [15:0]       dataInMem_hi_194;
  assign dataInMem_hi_194 = _GEN_261;
  wire [15:0]       dataInMem_lo_hi_326;
  assign dataInMem_lo_hi_326 = _GEN_261;
  wire [15:0]       _GEN_262 = {dataRegroupBySew_1_64, dataRegroupBySew_0_64};
  wire [15:0]       dataInMem_lo_67;
  assign dataInMem_lo_67 = _GEN_262;
  wire [15:0]       dataInMem_lo_196;
  assign dataInMem_lo_196 = _GEN_262;
  wire [15:0]       dataInMem_lo_lo_71;
  assign dataInMem_lo_lo_71 = _GEN_262;
  wire [15:0]       _GEN_263 = {dataRegroupBySew_3_64, dataRegroupBySew_2_64};
  wire [15:0]       dataInMem_hi_195;
  assign dataInMem_hi_195 = _GEN_263;
  wire [15:0]       dataInMem_lo_hi_327;
  assign dataInMem_lo_hi_327 = _GEN_263;
  wire [15:0]       _GEN_264 = {dataRegroupBySew_1_65, dataRegroupBySew_0_65};
  wire [15:0]       dataInMem_lo_68;
  assign dataInMem_lo_68 = _GEN_264;
  wire [15:0]       dataInMem_lo_197;
  assign dataInMem_lo_197 = _GEN_264;
  wire [15:0]       dataInMem_lo_lo_72;
  assign dataInMem_lo_lo_72 = _GEN_264;
  wire [15:0]       _GEN_265 = {dataRegroupBySew_3_65, dataRegroupBySew_2_65};
  wire [15:0]       dataInMem_hi_196;
  assign dataInMem_hi_196 = _GEN_265;
  wire [15:0]       dataInMem_lo_hi_328;
  assign dataInMem_lo_hi_328 = _GEN_265;
  wire [15:0]       _GEN_266 = {dataRegroupBySew_1_66, dataRegroupBySew_0_66};
  wire [15:0]       dataInMem_lo_69;
  assign dataInMem_lo_69 = _GEN_266;
  wire [15:0]       dataInMem_lo_198;
  assign dataInMem_lo_198 = _GEN_266;
  wire [15:0]       dataInMem_lo_lo_73;
  assign dataInMem_lo_lo_73 = _GEN_266;
  wire [15:0]       _GEN_267 = {dataRegroupBySew_3_66, dataRegroupBySew_2_66};
  wire [15:0]       dataInMem_hi_197;
  assign dataInMem_hi_197 = _GEN_267;
  wire [15:0]       dataInMem_lo_hi_329;
  assign dataInMem_lo_hi_329 = _GEN_267;
  wire [15:0]       _GEN_268 = {dataRegroupBySew_1_67, dataRegroupBySew_0_67};
  wire [15:0]       dataInMem_lo_70;
  assign dataInMem_lo_70 = _GEN_268;
  wire [15:0]       dataInMem_lo_199;
  assign dataInMem_lo_199 = _GEN_268;
  wire [15:0]       dataInMem_lo_lo_74;
  assign dataInMem_lo_lo_74 = _GEN_268;
  wire [15:0]       _GEN_269 = {dataRegroupBySew_3_67, dataRegroupBySew_2_67};
  wire [15:0]       dataInMem_hi_198;
  assign dataInMem_hi_198 = _GEN_269;
  wire [15:0]       dataInMem_lo_hi_330;
  assign dataInMem_lo_hi_330 = _GEN_269;
  wire [15:0]       _GEN_270 = {dataRegroupBySew_1_68, dataRegroupBySew_0_68};
  wire [15:0]       dataInMem_lo_71;
  assign dataInMem_lo_71 = _GEN_270;
  wire [15:0]       dataInMem_lo_200;
  assign dataInMem_lo_200 = _GEN_270;
  wire [15:0]       dataInMem_lo_lo_75;
  assign dataInMem_lo_lo_75 = _GEN_270;
  wire [15:0]       _GEN_271 = {dataRegroupBySew_3_68, dataRegroupBySew_2_68};
  wire [15:0]       dataInMem_hi_199;
  assign dataInMem_hi_199 = _GEN_271;
  wire [15:0]       dataInMem_lo_hi_331;
  assign dataInMem_lo_hi_331 = _GEN_271;
  wire [15:0]       _GEN_272 = {dataRegroupBySew_1_69, dataRegroupBySew_0_69};
  wire [15:0]       dataInMem_lo_72;
  assign dataInMem_lo_72 = _GEN_272;
  wire [15:0]       dataInMem_lo_201;
  assign dataInMem_lo_201 = _GEN_272;
  wire [15:0]       dataInMem_lo_lo_76;
  assign dataInMem_lo_lo_76 = _GEN_272;
  wire [15:0]       _GEN_273 = {dataRegroupBySew_3_69, dataRegroupBySew_2_69};
  wire [15:0]       dataInMem_hi_200;
  assign dataInMem_hi_200 = _GEN_273;
  wire [15:0]       dataInMem_lo_hi_332;
  assign dataInMem_lo_hi_332 = _GEN_273;
  wire [15:0]       _GEN_274 = {dataRegroupBySew_1_70, dataRegroupBySew_0_70};
  wire [15:0]       dataInMem_lo_73;
  assign dataInMem_lo_73 = _GEN_274;
  wire [15:0]       dataInMem_lo_202;
  assign dataInMem_lo_202 = _GEN_274;
  wire [15:0]       dataInMem_lo_lo_77;
  assign dataInMem_lo_lo_77 = _GEN_274;
  wire [15:0]       _GEN_275 = {dataRegroupBySew_3_70, dataRegroupBySew_2_70};
  wire [15:0]       dataInMem_hi_201;
  assign dataInMem_hi_201 = _GEN_275;
  wire [15:0]       dataInMem_lo_hi_333;
  assign dataInMem_lo_hi_333 = _GEN_275;
  wire [15:0]       _GEN_276 = {dataRegroupBySew_1_71, dataRegroupBySew_0_71};
  wire [15:0]       dataInMem_lo_74;
  assign dataInMem_lo_74 = _GEN_276;
  wire [15:0]       dataInMem_lo_203;
  assign dataInMem_lo_203 = _GEN_276;
  wire [15:0]       dataInMem_lo_lo_78;
  assign dataInMem_lo_lo_78 = _GEN_276;
  wire [15:0]       _GEN_277 = {dataRegroupBySew_3_71, dataRegroupBySew_2_71};
  wire [15:0]       dataInMem_hi_202;
  assign dataInMem_hi_202 = _GEN_277;
  wire [15:0]       dataInMem_lo_hi_334;
  assign dataInMem_lo_hi_334 = _GEN_277;
  wire [15:0]       _GEN_278 = {dataRegroupBySew_1_72, dataRegroupBySew_0_72};
  wire [15:0]       dataInMem_lo_75;
  assign dataInMem_lo_75 = _GEN_278;
  wire [15:0]       dataInMem_lo_204;
  assign dataInMem_lo_204 = _GEN_278;
  wire [15:0]       dataInMem_lo_lo_79;
  assign dataInMem_lo_lo_79 = _GEN_278;
  wire [15:0]       _GEN_279 = {dataRegroupBySew_3_72, dataRegroupBySew_2_72};
  wire [15:0]       dataInMem_hi_203;
  assign dataInMem_hi_203 = _GEN_279;
  wire [15:0]       dataInMem_lo_hi_335;
  assign dataInMem_lo_hi_335 = _GEN_279;
  wire [15:0]       _GEN_280 = {dataRegroupBySew_1_73, dataRegroupBySew_0_73};
  wire [15:0]       dataInMem_lo_76;
  assign dataInMem_lo_76 = _GEN_280;
  wire [15:0]       dataInMem_lo_205;
  assign dataInMem_lo_205 = _GEN_280;
  wire [15:0]       dataInMem_lo_lo_80;
  assign dataInMem_lo_lo_80 = _GEN_280;
  wire [15:0]       _GEN_281 = {dataRegroupBySew_3_73, dataRegroupBySew_2_73};
  wire [15:0]       dataInMem_hi_204;
  assign dataInMem_hi_204 = _GEN_281;
  wire [15:0]       dataInMem_lo_hi_336;
  assign dataInMem_lo_hi_336 = _GEN_281;
  wire [15:0]       _GEN_282 = {dataRegroupBySew_1_74, dataRegroupBySew_0_74};
  wire [15:0]       dataInMem_lo_77;
  assign dataInMem_lo_77 = _GEN_282;
  wire [15:0]       dataInMem_lo_206;
  assign dataInMem_lo_206 = _GEN_282;
  wire [15:0]       dataInMem_lo_lo_81;
  assign dataInMem_lo_lo_81 = _GEN_282;
  wire [15:0]       _GEN_283 = {dataRegroupBySew_3_74, dataRegroupBySew_2_74};
  wire [15:0]       dataInMem_hi_205;
  assign dataInMem_hi_205 = _GEN_283;
  wire [15:0]       dataInMem_lo_hi_337;
  assign dataInMem_lo_hi_337 = _GEN_283;
  wire [15:0]       _GEN_284 = {dataRegroupBySew_1_75, dataRegroupBySew_0_75};
  wire [15:0]       dataInMem_lo_78;
  assign dataInMem_lo_78 = _GEN_284;
  wire [15:0]       dataInMem_lo_207;
  assign dataInMem_lo_207 = _GEN_284;
  wire [15:0]       dataInMem_lo_lo_82;
  assign dataInMem_lo_lo_82 = _GEN_284;
  wire [15:0]       _GEN_285 = {dataRegroupBySew_3_75, dataRegroupBySew_2_75};
  wire [15:0]       dataInMem_hi_206;
  assign dataInMem_hi_206 = _GEN_285;
  wire [15:0]       dataInMem_lo_hi_338;
  assign dataInMem_lo_hi_338 = _GEN_285;
  wire [15:0]       _GEN_286 = {dataRegroupBySew_1_76, dataRegroupBySew_0_76};
  wire [15:0]       dataInMem_lo_79;
  assign dataInMem_lo_79 = _GEN_286;
  wire [15:0]       dataInMem_lo_208;
  assign dataInMem_lo_208 = _GEN_286;
  wire [15:0]       dataInMem_lo_lo_83;
  assign dataInMem_lo_lo_83 = _GEN_286;
  wire [15:0]       _GEN_287 = {dataRegroupBySew_3_76, dataRegroupBySew_2_76};
  wire [15:0]       dataInMem_hi_207;
  assign dataInMem_hi_207 = _GEN_287;
  wire [15:0]       dataInMem_lo_hi_339;
  assign dataInMem_lo_hi_339 = _GEN_287;
  wire [15:0]       _GEN_288 = {dataRegroupBySew_1_77, dataRegroupBySew_0_77};
  wire [15:0]       dataInMem_lo_80;
  assign dataInMem_lo_80 = _GEN_288;
  wire [15:0]       dataInMem_lo_209;
  assign dataInMem_lo_209 = _GEN_288;
  wire [15:0]       dataInMem_lo_lo_84;
  assign dataInMem_lo_lo_84 = _GEN_288;
  wire [15:0]       _GEN_289 = {dataRegroupBySew_3_77, dataRegroupBySew_2_77};
  wire [15:0]       dataInMem_hi_208;
  assign dataInMem_hi_208 = _GEN_289;
  wire [15:0]       dataInMem_lo_hi_340;
  assign dataInMem_lo_hi_340 = _GEN_289;
  wire [15:0]       _GEN_290 = {dataRegroupBySew_1_78, dataRegroupBySew_0_78};
  wire [15:0]       dataInMem_lo_81;
  assign dataInMem_lo_81 = _GEN_290;
  wire [15:0]       dataInMem_lo_210;
  assign dataInMem_lo_210 = _GEN_290;
  wire [15:0]       dataInMem_lo_lo_85;
  assign dataInMem_lo_lo_85 = _GEN_290;
  wire [15:0]       _GEN_291 = {dataRegroupBySew_3_78, dataRegroupBySew_2_78};
  wire [15:0]       dataInMem_hi_209;
  assign dataInMem_hi_209 = _GEN_291;
  wire [15:0]       dataInMem_lo_hi_341;
  assign dataInMem_lo_hi_341 = _GEN_291;
  wire [15:0]       _GEN_292 = {dataRegroupBySew_1_79, dataRegroupBySew_0_79};
  wire [15:0]       dataInMem_lo_82;
  assign dataInMem_lo_82 = _GEN_292;
  wire [15:0]       dataInMem_lo_211;
  assign dataInMem_lo_211 = _GEN_292;
  wire [15:0]       dataInMem_lo_lo_86;
  assign dataInMem_lo_lo_86 = _GEN_292;
  wire [15:0]       _GEN_293 = {dataRegroupBySew_3_79, dataRegroupBySew_2_79};
  wire [15:0]       dataInMem_hi_210;
  assign dataInMem_hi_210 = _GEN_293;
  wire [15:0]       dataInMem_lo_hi_342;
  assign dataInMem_lo_hi_342 = _GEN_293;
  wire [15:0]       _GEN_294 = {dataRegroupBySew_1_80, dataRegroupBySew_0_80};
  wire [15:0]       dataInMem_lo_83;
  assign dataInMem_lo_83 = _GEN_294;
  wire [15:0]       dataInMem_lo_212;
  assign dataInMem_lo_212 = _GEN_294;
  wire [15:0]       dataInMem_lo_lo_87;
  assign dataInMem_lo_lo_87 = _GEN_294;
  wire [15:0]       _GEN_295 = {dataRegroupBySew_3_80, dataRegroupBySew_2_80};
  wire [15:0]       dataInMem_hi_211;
  assign dataInMem_hi_211 = _GEN_295;
  wire [15:0]       dataInMem_lo_hi_343;
  assign dataInMem_lo_hi_343 = _GEN_295;
  wire [15:0]       _GEN_296 = {dataRegroupBySew_1_81, dataRegroupBySew_0_81};
  wire [15:0]       dataInMem_lo_84;
  assign dataInMem_lo_84 = _GEN_296;
  wire [15:0]       dataInMem_lo_213;
  assign dataInMem_lo_213 = _GEN_296;
  wire [15:0]       dataInMem_lo_lo_88;
  assign dataInMem_lo_lo_88 = _GEN_296;
  wire [15:0]       _GEN_297 = {dataRegroupBySew_3_81, dataRegroupBySew_2_81};
  wire [15:0]       dataInMem_hi_212;
  assign dataInMem_hi_212 = _GEN_297;
  wire [15:0]       dataInMem_lo_hi_344;
  assign dataInMem_lo_hi_344 = _GEN_297;
  wire [15:0]       _GEN_298 = {dataRegroupBySew_1_82, dataRegroupBySew_0_82};
  wire [15:0]       dataInMem_lo_85;
  assign dataInMem_lo_85 = _GEN_298;
  wire [15:0]       dataInMem_lo_214;
  assign dataInMem_lo_214 = _GEN_298;
  wire [15:0]       dataInMem_lo_lo_89;
  assign dataInMem_lo_lo_89 = _GEN_298;
  wire [15:0]       _GEN_299 = {dataRegroupBySew_3_82, dataRegroupBySew_2_82};
  wire [15:0]       dataInMem_hi_213;
  assign dataInMem_hi_213 = _GEN_299;
  wire [15:0]       dataInMem_lo_hi_345;
  assign dataInMem_lo_hi_345 = _GEN_299;
  wire [15:0]       _GEN_300 = {dataRegroupBySew_1_83, dataRegroupBySew_0_83};
  wire [15:0]       dataInMem_lo_86;
  assign dataInMem_lo_86 = _GEN_300;
  wire [15:0]       dataInMem_lo_215;
  assign dataInMem_lo_215 = _GEN_300;
  wire [15:0]       dataInMem_lo_lo_90;
  assign dataInMem_lo_lo_90 = _GEN_300;
  wire [15:0]       _GEN_301 = {dataRegroupBySew_3_83, dataRegroupBySew_2_83};
  wire [15:0]       dataInMem_hi_214;
  assign dataInMem_hi_214 = _GEN_301;
  wire [15:0]       dataInMem_lo_hi_346;
  assign dataInMem_lo_hi_346 = _GEN_301;
  wire [15:0]       _GEN_302 = {dataRegroupBySew_1_84, dataRegroupBySew_0_84};
  wire [15:0]       dataInMem_lo_87;
  assign dataInMem_lo_87 = _GEN_302;
  wire [15:0]       dataInMem_lo_216;
  assign dataInMem_lo_216 = _GEN_302;
  wire [15:0]       dataInMem_lo_lo_91;
  assign dataInMem_lo_lo_91 = _GEN_302;
  wire [15:0]       _GEN_303 = {dataRegroupBySew_3_84, dataRegroupBySew_2_84};
  wire [15:0]       dataInMem_hi_215;
  assign dataInMem_hi_215 = _GEN_303;
  wire [15:0]       dataInMem_lo_hi_347;
  assign dataInMem_lo_hi_347 = _GEN_303;
  wire [15:0]       _GEN_304 = {dataRegroupBySew_1_85, dataRegroupBySew_0_85};
  wire [15:0]       dataInMem_lo_88;
  assign dataInMem_lo_88 = _GEN_304;
  wire [15:0]       dataInMem_lo_217;
  assign dataInMem_lo_217 = _GEN_304;
  wire [15:0]       dataInMem_lo_lo_92;
  assign dataInMem_lo_lo_92 = _GEN_304;
  wire [15:0]       _GEN_305 = {dataRegroupBySew_3_85, dataRegroupBySew_2_85};
  wire [15:0]       dataInMem_hi_216;
  assign dataInMem_hi_216 = _GEN_305;
  wire [15:0]       dataInMem_lo_hi_348;
  assign dataInMem_lo_hi_348 = _GEN_305;
  wire [15:0]       _GEN_306 = {dataRegroupBySew_1_86, dataRegroupBySew_0_86};
  wire [15:0]       dataInMem_lo_89;
  assign dataInMem_lo_89 = _GEN_306;
  wire [15:0]       dataInMem_lo_218;
  assign dataInMem_lo_218 = _GEN_306;
  wire [15:0]       dataInMem_lo_lo_93;
  assign dataInMem_lo_lo_93 = _GEN_306;
  wire [15:0]       _GEN_307 = {dataRegroupBySew_3_86, dataRegroupBySew_2_86};
  wire [15:0]       dataInMem_hi_217;
  assign dataInMem_hi_217 = _GEN_307;
  wire [15:0]       dataInMem_lo_hi_349;
  assign dataInMem_lo_hi_349 = _GEN_307;
  wire [15:0]       _GEN_308 = {dataRegroupBySew_1_87, dataRegroupBySew_0_87};
  wire [15:0]       dataInMem_lo_90;
  assign dataInMem_lo_90 = _GEN_308;
  wire [15:0]       dataInMem_lo_219;
  assign dataInMem_lo_219 = _GEN_308;
  wire [15:0]       dataInMem_lo_lo_94;
  assign dataInMem_lo_lo_94 = _GEN_308;
  wire [15:0]       _GEN_309 = {dataRegroupBySew_3_87, dataRegroupBySew_2_87};
  wire [15:0]       dataInMem_hi_218;
  assign dataInMem_hi_218 = _GEN_309;
  wire [15:0]       dataInMem_lo_hi_350;
  assign dataInMem_lo_hi_350 = _GEN_309;
  wire [15:0]       _GEN_310 = {dataRegroupBySew_1_88, dataRegroupBySew_0_88};
  wire [15:0]       dataInMem_lo_91;
  assign dataInMem_lo_91 = _GEN_310;
  wire [15:0]       dataInMem_lo_220;
  assign dataInMem_lo_220 = _GEN_310;
  wire [15:0]       dataInMem_lo_lo_95;
  assign dataInMem_lo_lo_95 = _GEN_310;
  wire [15:0]       _GEN_311 = {dataRegroupBySew_3_88, dataRegroupBySew_2_88};
  wire [15:0]       dataInMem_hi_219;
  assign dataInMem_hi_219 = _GEN_311;
  wire [15:0]       dataInMem_lo_hi_351;
  assign dataInMem_lo_hi_351 = _GEN_311;
  wire [15:0]       _GEN_312 = {dataRegroupBySew_1_89, dataRegroupBySew_0_89};
  wire [15:0]       dataInMem_lo_92;
  assign dataInMem_lo_92 = _GEN_312;
  wire [15:0]       dataInMem_lo_221;
  assign dataInMem_lo_221 = _GEN_312;
  wire [15:0]       dataInMem_lo_lo_96;
  assign dataInMem_lo_lo_96 = _GEN_312;
  wire [15:0]       _GEN_313 = {dataRegroupBySew_3_89, dataRegroupBySew_2_89};
  wire [15:0]       dataInMem_hi_220;
  assign dataInMem_hi_220 = _GEN_313;
  wire [15:0]       dataInMem_lo_hi_352;
  assign dataInMem_lo_hi_352 = _GEN_313;
  wire [15:0]       _GEN_314 = {dataRegroupBySew_1_90, dataRegroupBySew_0_90};
  wire [15:0]       dataInMem_lo_93;
  assign dataInMem_lo_93 = _GEN_314;
  wire [15:0]       dataInMem_lo_222;
  assign dataInMem_lo_222 = _GEN_314;
  wire [15:0]       dataInMem_lo_lo_97;
  assign dataInMem_lo_lo_97 = _GEN_314;
  wire [15:0]       _GEN_315 = {dataRegroupBySew_3_90, dataRegroupBySew_2_90};
  wire [15:0]       dataInMem_hi_221;
  assign dataInMem_hi_221 = _GEN_315;
  wire [15:0]       dataInMem_lo_hi_353;
  assign dataInMem_lo_hi_353 = _GEN_315;
  wire [15:0]       _GEN_316 = {dataRegroupBySew_1_91, dataRegroupBySew_0_91};
  wire [15:0]       dataInMem_lo_94;
  assign dataInMem_lo_94 = _GEN_316;
  wire [15:0]       dataInMem_lo_223;
  assign dataInMem_lo_223 = _GEN_316;
  wire [15:0]       dataInMem_lo_lo_98;
  assign dataInMem_lo_lo_98 = _GEN_316;
  wire [15:0]       _GEN_317 = {dataRegroupBySew_3_91, dataRegroupBySew_2_91};
  wire [15:0]       dataInMem_hi_222;
  assign dataInMem_hi_222 = _GEN_317;
  wire [15:0]       dataInMem_lo_hi_354;
  assign dataInMem_lo_hi_354 = _GEN_317;
  wire [15:0]       _GEN_318 = {dataRegroupBySew_1_92, dataRegroupBySew_0_92};
  wire [15:0]       dataInMem_lo_95;
  assign dataInMem_lo_95 = _GEN_318;
  wire [15:0]       dataInMem_lo_224;
  assign dataInMem_lo_224 = _GEN_318;
  wire [15:0]       dataInMem_lo_lo_99;
  assign dataInMem_lo_lo_99 = _GEN_318;
  wire [15:0]       _GEN_319 = {dataRegroupBySew_3_92, dataRegroupBySew_2_92};
  wire [15:0]       dataInMem_hi_223;
  assign dataInMem_hi_223 = _GEN_319;
  wire [15:0]       dataInMem_lo_hi_355;
  assign dataInMem_lo_hi_355 = _GEN_319;
  wire [15:0]       _GEN_320 = {dataRegroupBySew_1_93, dataRegroupBySew_0_93};
  wire [15:0]       dataInMem_lo_96;
  assign dataInMem_lo_96 = _GEN_320;
  wire [15:0]       dataInMem_lo_225;
  assign dataInMem_lo_225 = _GEN_320;
  wire [15:0]       dataInMem_lo_lo_100;
  assign dataInMem_lo_lo_100 = _GEN_320;
  wire [15:0]       _GEN_321 = {dataRegroupBySew_3_93, dataRegroupBySew_2_93};
  wire [15:0]       dataInMem_hi_224;
  assign dataInMem_hi_224 = _GEN_321;
  wire [15:0]       dataInMem_lo_hi_356;
  assign dataInMem_lo_hi_356 = _GEN_321;
  wire [15:0]       _GEN_322 = {dataRegroupBySew_1_94, dataRegroupBySew_0_94};
  wire [15:0]       dataInMem_lo_97;
  assign dataInMem_lo_97 = _GEN_322;
  wire [15:0]       dataInMem_lo_226;
  assign dataInMem_lo_226 = _GEN_322;
  wire [15:0]       dataInMem_lo_lo_101;
  assign dataInMem_lo_lo_101 = _GEN_322;
  wire [15:0]       _GEN_323 = {dataRegroupBySew_3_94, dataRegroupBySew_2_94};
  wire [15:0]       dataInMem_hi_225;
  assign dataInMem_hi_225 = _GEN_323;
  wire [15:0]       dataInMem_lo_hi_357;
  assign dataInMem_lo_hi_357 = _GEN_323;
  wire [15:0]       _GEN_324 = {dataRegroupBySew_1_95, dataRegroupBySew_0_95};
  wire [15:0]       dataInMem_lo_98;
  assign dataInMem_lo_98 = _GEN_324;
  wire [15:0]       dataInMem_lo_227;
  assign dataInMem_lo_227 = _GEN_324;
  wire [15:0]       dataInMem_lo_lo_102;
  assign dataInMem_lo_lo_102 = _GEN_324;
  wire [15:0]       _GEN_325 = {dataRegroupBySew_3_95, dataRegroupBySew_2_95};
  wire [15:0]       dataInMem_hi_226;
  assign dataInMem_hi_226 = _GEN_325;
  wire [15:0]       dataInMem_lo_hi_358;
  assign dataInMem_lo_hi_358 = _GEN_325;
  wire [15:0]       _GEN_326 = {dataRegroupBySew_1_96, dataRegroupBySew_0_96};
  wire [15:0]       dataInMem_lo_99;
  assign dataInMem_lo_99 = _GEN_326;
  wire [15:0]       dataInMem_lo_228;
  assign dataInMem_lo_228 = _GEN_326;
  wire [15:0]       dataInMem_lo_lo_103;
  assign dataInMem_lo_lo_103 = _GEN_326;
  wire [15:0]       _GEN_327 = {dataRegroupBySew_3_96, dataRegroupBySew_2_96};
  wire [15:0]       dataInMem_hi_227;
  assign dataInMem_hi_227 = _GEN_327;
  wire [15:0]       dataInMem_lo_hi_359;
  assign dataInMem_lo_hi_359 = _GEN_327;
  wire [15:0]       _GEN_328 = {dataRegroupBySew_1_97, dataRegroupBySew_0_97};
  wire [15:0]       dataInMem_lo_100;
  assign dataInMem_lo_100 = _GEN_328;
  wire [15:0]       dataInMem_lo_229;
  assign dataInMem_lo_229 = _GEN_328;
  wire [15:0]       dataInMem_lo_lo_104;
  assign dataInMem_lo_lo_104 = _GEN_328;
  wire [15:0]       _GEN_329 = {dataRegroupBySew_3_97, dataRegroupBySew_2_97};
  wire [15:0]       dataInMem_hi_228;
  assign dataInMem_hi_228 = _GEN_329;
  wire [15:0]       dataInMem_lo_hi_360;
  assign dataInMem_lo_hi_360 = _GEN_329;
  wire [15:0]       _GEN_330 = {dataRegroupBySew_1_98, dataRegroupBySew_0_98};
  wire [15:0]       dataInMem_lo_101;
  assign dataInMem_lo_101 = _GEN_330;
  wire [15:0]       dataInMem_lo_230;
  assign dataInMem_lo_230 = _GEN_330;
  wire [15:0]       dataInMem_lo_lo_105;
  assign dataInMem_lo_lo_105 = _GEN_330;
  wire [15:0]       _GEN_331 = {dataRegroupBySew_3_98, dataRegroupBySew_2_98};
  wire [15:0]       dataInMem_hi_229;
  assign dataInMem_hi_229 = _GEN_331;
  wire [15:0]       dataInMem_lo_hi_361;
  assign dataInMem_lo_hi_361 = _GEN_331;
  wire [15:0]       _GEN_332 = {dataRegroupBySew_1_99, dataRegroupBySew_0_99};
  wire [15:0]       dataInMem_lo_102;
  assign dataInMem_lo_102 = _GEN_332;
  wire [15:0]       dataInMem_lo_231;
  assign dataInMem_lo_231 = _GEN_332;
  wire [15:0]       dataInMem_lo_lo_106;
  assign dataInMem_lo_lo_106 = _GEN_332;
  wire [15:0]       _GEN_333 = {dataRegroupBySew_3_99, dataRegroupBySew_2_99};
  wire [15:0]       dataInMem_hi_230;
  assign dataInMem_hi_230 = _GEN_333;
  wire [15:0]       dataInMem_lo_hi_362;
  assign dataInMem_lo_hi_362 = _GEN_333;
  wire [15:0]       _GEN_334 = {dataRegroupBySew_1_100, dataRegroupBySew_0_100};
  wire [15:0]       dataInMem_lo_103;
  assign dataInMem_lo_103 = _GEN_334;
  wire [15:0]       dataInMem_lo_232;
  assign dataInMem_lo_232 = _GEN_334;
  wire [15:0]       dataInMem_lo_lo_107;
  assign dataInMem_lo_lo_107 = _GEN_334;
  wire [15:0]       _GEN_335 = {dataRegroupBySew_3_100, dataRegroupBySew_2_100};
  wire [15:0]       dataInMem_hi_231;
  assign dataInMem_hi_231 = _GEN_335;
  wire [15:0]       dataInMem_lo_hi_363;
  assign dataInMem_lo_hi_363 = _GEN_335;
  wire [15:0]       _GEN_336 = {dataRegroupBySew_1_101, dataRegroupBySew_0_101};
  wire [15:0]       dataInMem_lo_104;
  assign dataInMem_lo_104 = _GEN_336;
  wire [15:0]       dataInMem_lo_233;
  assign dataInMem_lo_233 = _GEN_336;
  wire [15:0]       dataInMem_lo_lo_108;
  assign dataInMem_lo_lo_108 = _GEN_336;
  wire [15:0]       _GEN_337 = {dataRegroupBySew_3_101, dataRegroupBySew_2_101};
  wire [15:0]       dataInMem_hi_232;
  assign dataInMem_hi_232 = _GEN_337;
  wire [15:0]       dataInMem_lo_hi_364;
  assign dataInMem_lo_hi_364 = _GEN_337;
  wire [15:0]       _GEN_338 = {dataRegroupBySew_1_102, dataRegroupBySew_0_102};
  wire [15:0]       dataInMem_lo_105;
  assign dataInMem_lo_105 = _GEN_338;
  wire [15:0]       dataInMem_lo_234;
  assign dataInMem_lo_234 = _GEN_338;
  wire [15:0]       dataInMem_lo_lo_109;
  assign dataInMem_lo_lo_109 = _GEN_338;
  wire [15:0]       _GEN_339 = {dataRegroupBySew_3_102, dataRegroupBySew_2_102};
  wire [15:0]       dataInMem_hi_233;
  assign dataInMem_hi_233 = _GEN_339;
  wire [15:0]       dataInMem_lo_hi_365;
  assign dataInMem_lo_hi_365 = _GEN_339;
  wire [15:0]       _GEN_340 = {dataRegroupBySew_1_103, dataRegroupBySew_0_103};
  wire [15:0]       dataInMem_lo_106;
  assign dataInMem_lo_106 = _GEN_340;
  wire [15:0]       dataInMem_lo_235;
  assign dataInMem_lo_235 = _GEN_340;
  wire [15:0]       dataInMem_lo_lo_110;
  assign dataInMem_lo_lo_110 = _GEN_340;
  wire [15:0]       _GEN_341 = {dataRegroupBySew_3_103, dataRegroupBySew_2_103};
  wire [15:0]       dataInMem_hi_234;
  assign dataInMem_hi_234 = _GEN_341;
  wire [15:0]       dataInMem_lo_hi_366;
  assign dataInMem_lo_hi_366 = _GEN_341;
  wire [15:0]       _GEN_342 = {dataRegroupBySew_1_104, dataRegroupBySew_0_104};
  wire [15:0]       dataInMem_lo_107;
  assign dataInMem_lo_107 = _GEN_342;
  wire [15:0]       dataInMem_lo_236;
  assign dataInMem_lo_236 = _GEN_342;
  wire [15:0]       dataInMem_lo_lo_111;
  assign dataInMem_lo_lo_111 = _GEN_342;
  wire [15:0]       _GEN_343 = {dataRegroupBySew_3_104, dataRegroupBySew_2_104};
  wire [15:0]       dataInMem_hi_235;
  assign dataInMem_hi_235 = _GEN_343;
  wire [15:0]       dataInMem_lo_hi_367;
  assign dataInMem_lo_hi_367 = _GEN_343;
  wire [15:0]       _GEN_344 = {dataRegroupBySew_1_105, dataRegroupBySew_0_105};
  wire [15:0]       dataInMem_lo_108;
  assign dataInMem_lo_108 = _GEN_344;
  wire [15:0]       dataInMem_lo_237;
  assign dataInMem_lo_237 = _GEN_344;
  wire [15:0]       dataInMem_lo_lo_112;
  assign dataInMem_lo_lo_112 = _GEN_344;
  wire [15:0]       _GEN_345 = {dataRegroupBySew_3_105, dataRegroupBySew_2_105};
  wire [15:0]       dataInMem_hi_236;
  assign dataInMem_hi_236 = _GEN_345;
  wire [15:0]       dataInMem_lo_hi_368;
  assign dataInMem_lo_hi_368 = _GEN_345;
  wire [15:0]       _GEN_346 = {dataRegroupBySew_1_106, dataRegroupBySew_0_106};
  wire [15:0]       dataInMem_lo_109;
  assign dataInMem_lo_109 = _GEN_346;
  wire [15:0]       dataInMem_lo_238;
  assign dataInMem_lo_238 = _GEN_346;
  wire [15:0]       dataInMem_lo_lo_113;
  assign dataInMem_lo_lo_113 = _GEN_346;
  wire [15:0]       _GEN_347 = {dataRegroupBySew_3_106, dataRegroupBySew_2_106};
  wire [15:0]       dataInMem_hi_237;
  assign dataInMem_hi_237 = _GEN_347;
  wire [15:0]       dataInMem_lo_hi_369;
  assign dataInMem_lo_hi_369 = _GEN_347;
  wire [15:0]       _GEN_348 = {dataRegroupBySew_1_107, dataRegroupBySew_0_107};
  wire [15:0]       dataInMem_lo_110;
  assign dataInMem_lo_110 = _GEN_348;
  wire [15:0]       dataInMem_lo_239;
  assign dataInMem_lo_239 = _GEN_348;
  wire [15:0]       dataInMem_lo_lo_114;
  assign dataInMem_lo_lo_114 = _GEN_348;
  wire [15:0]       _GEN_349 = {dataRegroupBySew_3_107, dataRegroupBySew_2_107};
  wire [15:0]       dataInMem_hi_238;
  assign dataInMem_hi_238 = _GEN_349;
  wire [15:0]       dataInMem_lo_hi_370;
  assign dataInMem_lo_hi_370 = _GEN_349;
  wire [15:0]       _GEN_350 = {dataRegroupBySew_1_108, dataRegroupBySew_0_108};
  wire [15:0]       dataInMem_lo_111;
  assign dataInMem_lo_111 = _GEN_350;
  wire [15:0]       dataInMem_lo_240;
  assign dataInMem_lo_240 = _GEN_350;
  wire [15:0]       dataInMem_lo_lo_115;
  assign dataInMem_lo_lo_115 = _GEN_350;
  wire [15:0]       _GEN_351 = {dataRegroupBySew_3_108, dataRegroupBySew_2_108};
  wire [15:0]       dataInMem_hi_239;
  assign dataInMem_hi_239 = _GEN_351;
  wire [15:0]       dataInMem_lo_hi_371;
  assign dataInMem_lo_hi_371 = _GEN_351;
  wire [15:0]       _GEN_352 = {dataRegroupBySew_1_109, dataRegroupBySew_0_109};
  wire [15:0]       dataInMem_lo_112;
  assign dataInMem_lo_112 = _GEN_352;
  wire [15:0]       dataInMem_lo_241;
  assign dataInMem_lo_241 = _GEN_352;
  wire [15:0]       dataInMem_lo_lo_116;
  assign dataInMem_lo_lo_116 = _GEN_352;
  wire [15:0]       _GEN_353 = {dataRegroupBySew_3_109, dataRegroupBySew_2_109};
  wire [15:0]       dataInMem_hi_240;
  assign dataInMem_hi_240 = _GEN_353;
  wire [15:0]       dataInMem_lo_hi_372;
  assign dataInMem_lo_hi_372 = _GEN_353;
  wire [15:0]       _GEN_354 = {dataRegroupBySew_1_110, dataRegroupBySew_0_110};
  wire [15:0]       dataInMem_lo_113;
  assign dataInMem_lo_113 = _GEN_354;
  wire [15:0]       dataInMem_lo_242;
  assign dataInMem_lo_242 = _GEN_354;
  wire [15:0]       dataInMem_lo_lo_117;
  assign dataInMem_lo_lo_117 = _GEN_354;
  wire [15:0]       _GEN_355 = {dataRegroupBySew_3_110, dataRegroupBySew_2_110};
  wire [15:0]       dataInMem_hi_241;
  assign dataInMem_hi_241 = _GEN_355;
  wire [15:0]       dataInMem_lo_hi_373;
  assign dataInMem_lo_hi_373 = _GEN_355;
  wire [15:0]       _GEN_356 = {dataRegroupBySew_1_111, dataRegroupBySew_0_111};
  wire [15:0]       dataInMem_lo_114;
  assign dataInMem_lo_114 = _GEN_356;
  wire [15:0]       dataInMem_lo_243;
  assign dataInMem_lo_243 = _GEN_356;
  wire [15:0]       dataInMem_lo_lo_118;
  assign dataInMem_lo_lo_118 = _GEN_356;
  wire [15:0]       _GEN_357 = {dataRegroupBySew_3_111, dataRegroupBySew_2_111};
  wire [15:0]       dataInMem_hi_242;
  assign dataInMem_hi_242 = _GEN_357;
  wire [15:0]       dataInMem_lo_hi_374;
  assign dataInMem_lo_hi_374 = _GEN_357;
  wire [15:0]       _GEN_358 = {dataRegroupBySew_1_112, dataRegroupBySew_0_112};
  wire [15:0]       dataInMem_lo_115;
  assign dataInMem_lo_115 = _GEN_358;
  wire [15:0]       dataInMem_lo_244;
  assign dataInMem_lo_244 = _GEN_358;
  wire [15:0]       dataInMem_lo_lo_119;
  assign dataInMem_lo_lo_119 = _GEN_358;
  wire [15:0]       _GEN_359 = {dataRegroupBySew_3_112, dataRegroupBySew_2_112};
  wire [15:0]       dataInMem_hi_243;
  assign dataInMem_hi_243 = _GEN_359;
  wire [15:0]       dataInMem_lo_hi_375;
  assign dataInMem_lo_hi_375 = _GEN_359;
  wire [15:0]       _GEN_360 = {dataRegroupBySew_1_113, dataRegroupBySew_0_113};
  wire [15:0]       dataInMem_lo_116;
  assign dataInMem_lo_116 = _GEN_360;
  wire [15:0]       dataInMem_lo_245;
  assign dataInMem_lo_245 = _GEN_360;
  wire [15:0]       dataInMem_lo_lo_120;
  assign dataInMem_lo_lo_120 = _GEN_360;
  wire [15:0]       _GEN_361 = {dataRegroupBySew_3_113, dataRegroupBySew_2_113};
  wire [15:0]       dataInMem_hi_244;
  assign dataInMem_hi_244 = _GEN_361;
  wire [15:0]       dataInMem_lo_hi_376;
  assign dataInMem_lo_hi_376 = _GEN_361;
  wire [15:0]       _GEN_362 = {dataRegroupBySew_1_114, dataRegroupBySew_0_114};
  wire [15:0]       dataInMem_lo_117;
  assign dataInMem_lo_117 = _GEN_362;
  wire [15:0]       dataInMem_lo_246;
  assign dataInMem_lo_246 = _GEN_362;
  wire [15:0]       dataInMem_lo_lo_121;
  assign dataInMem_lo_lo_121 = _GEN_362;
  wire [15:0]       _GEN_363 = {dataRegroupBySew_3_114, dataRegroupBySew_2_114};
  wire [15:0]       dataInMem_hi_245;
  assign dataInMem_hi_245 = _GEN_363;
  wire [15:0]       dataInMem_lo_hi_377;
  assign dataInMem_lo_hi_377 = _GEN_363;
  wire [15:0]       _GEN_364 = {dataRegroupBySew_1_115, dataRegroupBySew_0_115};
  wire [15:0]       dataInMem_lo_118;
  assign dataInMem_lo_118 = _GEN_364;
  wire [15:0]       dataInMem_lo_247;
  assign dataInMem_lo_247 = _GEN_364;
  wire [15:0]       dataInMem_lo_lo_122;
  assign dataInMem_lo_lo_122 = _GEN_364;
  wire [15:0]       _GEN_365 = {dataRegroupBySew_3_115, dataRegroupBySew_2_115};
  wire [15:0]       dataInMem_hi_246;
  assign dataInMem_hi_246 = _GEN_365;
  wire [15:0]       dataInMem_lo_hi_378;
  assign dataInMem_lo_hi_378 = _GEN_365;
  wire [15:0]       _GEN_366 = {dataRegroupBySew_1_116, dataRegroupBySew_0_116};
  wire [15:0]       dataInMem_lo_119;
  assign dataInMem_lo_119 = _GEN_366;
  wire [15:0]       dataInMem_lo_248;
  assign dataInMem_lo_248 = _GEN_366;
  wire [15:0]       dataInMem_lo_lo_123;
  assign dataInMem_lo_lo_123 = _GEN_366;
  wire [15:0]       _GEN_367 = {dataRegroupBySew_3_116, dataRegroupBySew_2_116};
  wire [15:0]       dataInMem_hi_247;
  assign dataInMem_hi_247 = _GEN_367;
  wire [15:0]       dataInMem_lo_hi_379;
  assign dataInMem_lo_hi_379 = _GEN_367;
  wire [15:0]       _GEN_368 = {dataRegroupBySew_1_117, dataRegroupBySew_0_117};
  wire [15:0]       dataInMem_lo_120;
  assign dataInMem_lo_120 = _GEN_368;
  wire [15:0]       dataInMem_lo_249;
  assign dataInMem_lo_249 = _GEN_368;
  wire [15:0]       dataInMem_lo_lo_124;
  assign dataInMem_lo_lo_124 = _GEN_368;
  wire [15:0]       _GEN_369 = {dataRegroupBySew_3_117, dataRegroupBySew_2_117};
  wire [15:0]       dataInMem_hi_248;
  assign dataInMem_hi_248 = _GEN_369;
  wire [15:0]       dataInMem_lo_hi_380;
  assign dataInMem_lo_hi_380 = _GEN_369;
  wire [15:0]       _GEN_370 = {dataRegroupBySew_1_118, dataRegroupBySew_0_118};
  wire [15:0]       dataInMem_lo_121;
  assign dataInMem_lo_121 = _GEN_370;
  wire [15:0]       dataInMem_lo_250;
  assign dataInMem_lo_250 = _GEN_370;
  wire [15:0]       dataInMem_lo_lo_125;
  assign dataInMem_lo_lo_125 = _GEN_370;
  wire [15:0]       _GEN_371 = {dataRegroupBySew_3_118, dataRegroupBySew_2_118};
  wire [15:0]       dataInMem_hi_249;
  assign dataInMem_hi_249 = _GEN_371;
  wire [15:0]       dataInMem_lo_hi_381;
  assign dataInMem_lo_hi_381 = _GEN_371;
  wire [15:0]       _GEN_372 = {dataRegroupBySew_1_119, dataRegroupBySew_0_119};
  wire [15:0]       dataInMem_lo_122;
  assign dataInMem_lo_122 = _GEN_372;
  wire [15:0]       dataInMem_lo_251;
  assign dataInMem_lo_251 = _GEN_372;
  wire [15:0]       dataInMem_lo_lo_126;
  assign dataInMem_lo_lo_126 = _GEN_372;
  wire [15:0]       _GEN_373 = {dataRegroupBySew_3_119, dataRegroupBySew_2_119};
  wire [15:0]       dataInMem_hi_250;
  assign dataInMem_hi_250 = _GEN_373;
  wire [15:0]       dataInMem_lo_hi_382;
  assign dataInMem_lo_hi_382 = _GEN_373;
  wire [15:0]       _GEN_374 = {dataRegroupBySew_1_120, dataRegroupBySew_0_120};
  wire [15:0]       dataInMem_lo_123;
  assign dataInMem_lo_123 = _GEN_374;
  wire [15:0]       dataInMem_lo_252;
  assign dataInMem_lo_252 = _GEN_374;
  wire [15:0]       dataInMem_lo_lo_127;
  assign dataInMem_lo_lo_127 = _GEN_374;
  wire [15:0]       _GEN_375 = {dataRegroupBySew_3_120, dataRegroupBySew_2_120};
  wire [15:0]       dataInMem_hi_251;
  assign dataInMem_hi_251 = _GEN_375;
  wire [15:0]       dataInMem_lo_hi_383;
  assign dataInMem_lo_hi_383 = _GEN_375;
  wire [15:0]       _GEN_376 = {dataRegroupBySew_1_121, dataRegroupBySew_0_121};
  wire [15:0]       dataInMem_lo_124;
  assign dataInMem_lo_124 = _GEN_376;
  wire [15:0]       dataInMem_lo_253;
  assign dataInMem_lo_253 = _GEN_376;
  wire [15:0]       dataInMem_lo_lo_128;
  assign dataInMem_lo_lo_128 = _GEN_376;
  wire [15:0]       _GEN_377 = {dataRegroupBySew_3_121, dataRegroupBySew_2_121};
  wire [15:0]       dataInMem_hi_252;
  assign dataInMem_hi_252 = _GEN_377;
  wire [15:0]       dataInMem_lo_hi_384;
  assign dataInMem_lo_hi_384 = _GEN_377;
  wire [15:0]       _GEN_378 = {dataRegroupBySew_1_122, dataRegroupBySew_0_122};
  wire [15:0]       dataInMem_lo_125;
  assign dataInMem_lo_125 = _GEN_378;
  wire [15:0]       dataInMem_lo_254;
  assign dataInMem_lo_254 = _GEN_378;
  wire [15:0]       dataInMem_lo_lo_129;
  assign dataInMem_lo_lo_129 = _GEN_378;
  wire [15:0]       _GEN_379 = {dataRegroupBySew_3_122, dataRegroupBySew_2_122};
  wire [15:0]       dataInMem_hi_253;
  assign dataInMem_hi_253 = _GEN_379;
  wire [15:0]       dataInMem_lo_hi_385;
  assign dataInMem_lo_hi_385 = _GEN_379;
  wire [15:0]       _GEN_380 = {dataRegroupBySew_1_123, dataRegroupBySew_0_123};
  wire [15:0]       dataInMem_lo_126;
  assign dataInMem_lo_126 = _GEN_380;
  wire [15:0]       dataInMem_lo_255;
  assign dataInMem_lo_255 = _GEN_380;
  wire [15:0]       dataInMem_lo_lo_130;
  assign dataInMem_lo_lo_130 = _GEN_380;
  wire [15:0]       _GEN_381 = {dataRegroupBySew_3_123, dataRegroupBySew_2_123};
  wire [15:0]       dataInMem_hi_254;
  assign dataInMem_hi_254 = _GEN_381;
  wire [15:0]       dataInMem_lo_hi_386;
  assign dataInMem_lo_hi_386 = _GEN_381;
  wire [15:0]       _GEN_382 = {dataRegroupBySew_1_124, dataRegroupBySew_0_124};
  wire [15:0]       dataInMem_lo_127;
  assign dataInMem_lo_127 = _GEN_382;
  wire [15:0]       dataInMem_lo_256;
  assign dataInMem_lo_256 = _GEN_382;
  wire [15:0]       dataInMem_lo_lo_131;
  assign dataInMem_lo_lo_131 = _GEN_382;
  wire [15:0]       _GEN_383 = {dataRegroupBySew_3_124, dataRegroupBySew_2_124};
  wire [15:0]       dataInMem_hi_255;
  assign dataInMem_hi_255 = _GEN_383;
  wire [15:0]       dataInMem_lo_hi_387;
  assign dataInMem_lo_hi_387 = _GEN_383;
  wire [15:0]       _GEN_384 = {dataRegroupBySew_1_125, dataRegroupBySew_0_125};
  wire [15:0]       dataInMem_lo_128;
  assign dataInMem_lo_128 = _GEN_384;
  wire [15:0]       dataInMem_lo_257;
  assign dataInMem_lo_257 = _GEN_384;
  wire [15:0]       dataInMem_lo_lo_132;
  assign dataInMem_lo_lo_132 = _GEN_384;
  wire [15:0]       _GEN_385 = {dataRegroupBySew_3_125, dataRegroupBySew_2_125};
  wire [15:0]       dataInMem_hi_256;
  assign dataInMem_hi_256 = _GEN_385;
  wire [15:0]       dataInMem_lo_hi_388;
  assign dataInMem_lo_hi_388 = _GEN_385;
  wire [15:0]       _GEN_386 = {dataRegroupBySew_1_126, dataRegroupBySew_0_126};
  wire [15:0]       dataInMem_lo_129;
  assign dataInMem_lo_129 = _GEN_386;
  wire [15:0]       dataInMem_lo_258;
  assign dataInMem_lo_258 = _GEN_386;
  wire [15:0]       dataInMem_lo_lo_133;
  assign dataInMem_lo_lo_133 = _GEN_386;
  wire [15:0]       _GEN_387 = {dataRegroupBySew_3_126, dataRegroupBySew_2_126};
  wire [15:0]       dataInMem_hi_257;
  assign dataInMem_hi_257 = _GEN_387;
  wire [15:0]       dataInMem_lo_hi_389;
  assign dataInMem_lo_hi_389 = _GEN_387;
  wire [15:0]       _GEN_388 = {dataRegroupBySew_1_127, dataRegroupBySew_0_127};
  wire [15:0]       dataInMem_lo_130;
  assign dataInMem_lo_130 = _GEN_388;
  wire [15:0]       dataInMem_lo_259;
  assign dataInMem_lo_259 = _GEN_388;
  wire [15:0]       dataInMem_lo_lo_134;
  assign dataInMem_lo_lo_134 = _GEN_388;
  wire [15:0]       _GEN_389 = {dataRegroupBySew_3_127, dataRegroupBySew_2_127};
  wire [15:0]       dataInMem_hi_258;
  assign dataInMem_hi_258 = _GEN_389;
  wire [15:0]       dataInMem_lo_hi_390;
  assign dataInMem_lo_hi_390 = _GEN_389;
  wire [63:0]       dataInMem_lo_lo_lo_lo_lo_lo_3 = {dataInMem_hi_132, dataInMem_lo_4, dataInMem_hi_131, dataInMem_lo_3};
  wire [63:0]       dataInMem_lo_lo_lo_lo_lo_hi_3 = {dataInMem_hi_134, dataInMem_lo_6, dataInMem_hi_133, dataInMem_lo_5};
  wire [127:0]      dataInMem_lo_lo_lo_lo_lo_3 = {dataInMem_lo_lo_lo_lo_lo_hi_3, dataInMem_lo_lo_lo_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_lo_lo_lo_hi_lo_3 = {dataInMem_hi_136, dataInMem_lo_8, dataInMem_hi_135, dataInMem_lo_7};
  wire [63:0]       dataInMem_lo_lo_lo_lo_hi_hi_3 = {dataInMem_hi_138, dataInMem_lo_10, dataInMem_hi_137, dataInMem_lo_9};
  wire [127:0]      dataInMem_lo_lo_lo_lo_hi_3 = {dataInMem_lo_lo_lo_lo_hi_hi_3, dataInMem_lo_lo_lo_lo_hi_lo_3};
  wire [255:0]      dataInMem_lo_lo_lo_lo_3 = {dataInMem_lo_lo_lo_lo_hi_3, dataInMem_lo_lo_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_lo_lo_hi_lo_lo_3 = {dataInMem_hi_140, dataInMem_lo_12, dataInMem_hi_139, dataInMem_lo_11};
  wire [63:0]       dataInMem_lo_lo_lo_hi_lo_hi_3 = {dataInMem_hi_142, dataInMem_lo_14, dataInMem_hi_141, dataInMem_lo_13};
  wire [127:0]      dataInMem_lo_lo_lo_hi_lo_3 = {dataInMem_lo_lo_lo_hi_lo_hi_3, dataInMem_lo_lo_lo_hi_lo_lo_3};
  wire [63:0]       dataInMem_lo_lo_lo_hi_hi_lo_3 = {dataInMem_hi_144, dataInMem_lo_16, dataInMem_hi_143, dataInMem_lo_15};
  wire [63:0]       dataInMem_lo_lo_lo_hi_hi_hi_3 = {dataInMem_hi_146, dataInMem_lo_18, dataInMem_hi_145, dataInMem_lo_17};
  wire [127:0]      dataInMem_lo_lo_lo_hi_hi_3 = {dataInMem_lo_lo_lo_hi_hi_hi_3, dataInMem_lo_lo_lo_hi_hi_lo_3};
  wire [255:0]      dataInMem_lo_lo_lo_hi_3 = {dataInMem_lo_lo_lo_hi_hi_3, dataInMem_lo_lo_lo_hi_lo_3};
  wire [511:0]      dataInMem_lo_lo_lo_3 = {dataInMem_lo_lo_lo_hi_3, dataInMem_lo_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_lo_hi_lo_lo_lo_3 = {dataInMem_hi_148, dataInMem_lo_20, dataInMem_hi_147, dataInMem_lo_19};
  wire [63:0]       dataInMem_lo_lo_hi_lo_lo_hi_3 = {dataInMem_hi_150, dataInMem_lo_22, dataInMem_hi_149, dataInMem_lo_21};
  wire [127:0]      dataInMem_lo_lo_hi_lo_lo_3 = {dataInMem_lo_lo_hi_lo_lo_hi_3, dataInMem_lo_lo_hi_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_lo_hi_lo_hi_lo_3 = {dataInMem_hi_152, dataInMem_lo_24, dataInMem_hi_151, dataInMem_lo_23};
  wire [63:0]       dataInMem_lo_lo_hi_lo_hi_hi_3 = {dataInMem_hi_154, dataInMem_lo_26, dataInMem_hi_153, dataInMem_lo_25};
  wire [127:0]      dataInMem_lo_lo_hi_lo_hi_3 = {dataInMem_lo_lo_hi_lo_hi_hi_3, dataInMem_lo_lo_hi_lo_hi_lo_3};
  wire [255:0]      dataInMem_lo_lo_hi_lo_3 = {dataInMem_lo_lo_hi_lo_hi_3, dataInMem_lo_lo_hi_lo_lo_3};
  wire [63:0]       dataInMem_lo_lo_hi_hi_lo_lo_3 = {dataInMem_hi_156, dataInMem_lo_28, dataInMem_hi_155, dataInMem_lo_27};
  wire [63:0]       dataInMem_lo_lo_hi_hi_lo_hi_3 = {dataInMem_hi_158, dataInMem_lo_30, dataInMem_hi_157, dataInMem_lo_29};
  wire [127:0]      dataInMem_lo_lo_hi_hi_lo_3 = {dataInMem_lo_lo_hi_hi_lo_hi_3, dataInMem_lo_lo_hi_hi_lo_lo_3};
  wire [63:0]       dataInMem_lo_lo_hi_hi_hi_lo_3 = {dataInMem_hi_160, dataInMem_lo_32, dataInMem_hi_159, dataInMem_lo_31};
  wire [63:0]       dataInMem_lo_lo_hi_hi_hi_hi_3 = {dataInMem_hi_162, dataInMem_lo_34, dataInMem_hi_161, dataInMem_lo_33};
  wire [127:0]      dataInMem_lo_lo_hi_hi_hi_3 = {dataInMem_lo_lo_hi_hi_hi_hi_3, dataInMem_lo_lo_hi_hi_hi_lo_3};
  wire [255:0]      dataInMem_lo_lo_hi_hi_3 = {dataInMem_lo_lo_hi_hi_hi_3, dataInMem_lo_lo_hi_hi_lo_3};
  wire [511:0]      dataInMem_lo_lo_hi_3 = {dataInMem_lo_lo_hi_hi_3, dataInMem_lo_lo_hi_lo_3};
  wire [1023:0]     dataInMem_lo_lo_3 = {dataInMem_lo_lo_hi_3, dataInMem_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_lo_lo_lo_lo_3 = {dataInMem_hi_164, dataInMem_lo_36, dataInMem_hi_163, dataInMem_lo_35};
  wire [63:0]       dataInMem_lo_hi_lo_lo_lo_hi_3 = {dataInMem_hi_166, dataInMem_lo_38, dataInMem_hi_165, dataInMem_lo_37};
  wire [127:0]      dataInMem_lo_hi_lo_lo_lo_3 = {dataInMem_lo_hi_lo_lo_lo_hi_3, dataInMem_lo_hi_lo_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_lo_lo_hi_lo_3 = {dataInMem_hi_168, dataInMem_lo_40, dataInMem_hi_167, dataInMem_lo_39};
  wire [63:0]       dataInMem_lo_hi_lo_lo_hi_hi_3 = {dataInMem_hi_170, dataInMem_lo_42, dataInMem_hi_169, dataInMem_lo_41};
  wire [127:0]      dataInMem_lo_hi_lo_lo_hi_3 = {dataInMem_lo_hi_lo_lo_hi_hi_3, dataInMem_lo_hi_lo_lo_hi_lo_3};
  wire [255:0]      dataInMem_lo_hi_lo_lo_3 = {dataInMem_lo_hi_lo_lo_hi_3, dataInMem_lo_hi_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_lo_hi_lo_lo_3 = {dataInMem_hi_172, dataInMem_lo_44, dataInMem_hi_171, dataInMem_lo_43};
  wire [63:0]       dataInMem_lo_hi_lo_hi_lo_hi_3 = {dataInMem_hi_174, dataInMem_lo_46, dataInMem_hi_173, dataInMem_lo_45};
  wire [127:0]      dataInMem_lo_hi_lo_hi_lo_3 = {dataInMem_lo_hi_lo_hi_lo_hi_3, dataInMem_lo_hi_lo_hi_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_lo_hi_hi_lo_3 = {dataInMem_hi_176, dataInMem_lo_48, dataInMem_hi_175, dataInMem_lo_47};
  wire [63:0]       dataInMem_lo_hi_lo_hi_hi_hi_3 = {dataInMem_hi_178, dataInMem_lo_50, dataInMem_hi_177, dataInMem_lo_49};
  wire [127:0]      dataInMem_lo_hi_lo_hi_hi_3 = {dataInMem_lo_hi_lo_hi_hi_hi_3, dataInMem_lo_hi_lo_hi_hi_lo_3};
  wire [255:0]      dataInMem_lo_hi_lo_hi_3 = {dataInMem_lo_hi_lo_hi_hi_3, dataInMem_lo_hi_lo_hi_lo_3};
  wire [511:0]      dataInMem_lo_hi_lo_3 = {dataInMem_lo_hi_lo_hi_3, dataInMem_lo_hi_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_hi_lo_lo_lo_3 = {dataInMem_hi_180, dataInMem_lo_52, dataInMem_hi_179, dataInMem_lo_51};
  wire [63:0]       dataInMem_lo_hi_hi_lo_lo_hi_3 = {dataInMem_hi_182, dataInMem_lo_54, dataInMem_hi_181, dataInMem_lo_53};
  wire [127:0]      dataInMem_lo_hi_hi_lo_lo_3 = {dataInMem_lo_hi_hi_lo_lo_hi_3, dataInMem_lo_hi_hi_lo_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_hi_lo_hi_lo_3 = {dataInMem_hi_184, dataInMem_lo_56, dataInMem_hi_183, dataInMem_lo_55};
  wire [63:0]       dataInMem_lo_hi_hi_lo_hi_hi_3 = {dataInMem_hi_186, dataInMem_lo_58, dataInMem_hi_185, dataInMem_lo_57};
  wire [127:0]      dataInMem_lo_hi_hi_lo_hi_3 = {dataInMem_lo_hi_hi_lo_hi_hi_3, dataInMem_lo_hi_hi_lo_hi_lo_3};
  wire [255:0]      dataInMem_lo_hi_hi_lo_3 = {dataInMem_lo_hi_hi_lo_hi_3, dataInMem_lo_hi_hi_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_hi_hi_lo_lo_3 = {dataInMem_hi_188, dataInMem_lo_60, dataInMem_hi_187, dataInMem_lo_59};
  wire [63:0]       dataInMem_lo_hi_hi_hi_lo_hi_3 = {dataInMem_hi_190, dataInMem_lo_62, dataInMem_hi_189, dataInMem_lo_61};
  wire [127:0]      dataInMem_lo_hi_hi_hi_lo_3 = {dataInMem_lo_hi_hi_hi_lo_hi_3, dataInMem_lo_hi_hi_hi_lo_lo_3};
  wire [63:0]       dataInMem_lo_hi_hi_hi_hi_lo_3 = {dataInMem_hi_192, dataInMem_lo_64, dataInMem_hi_191, dataInMem_lo_63};
  wire [63:0]       dataInMem_lo_hi_hi_hi_hi_hi_3 = {dataInMem_hi_194, dataInMem_lo_66, dataInMem_hi_193, dataInMem_lo_65};
  wire [127:0]      dataInMem_lo_hi_hi_hi_hi_3 = {dataInMem_lo_hi_hi_hi_hi_hi_3, dataInMem_lo_hi_hi_hi_hi_lo_3};
  wire [255:0]      dataInMem_lo_hi_hi_hi_3 = {dataInMem_lo_hi_hi_hi_hi_3, dataInMem_lo_hi_hi_hi_lo_3};
  wire [511:0]      dataInMem_lo_hi_hi_3 = {dataInMem_lo_hi_hi_hi_3, dataInMem_lo_hi_hi_lo_3};
  wire [1023:0]     dataInMem_lo_hi_3 = {dataInMem_lo_hi_hi_3, dataInMem_lo_hi_lo_3};
  wire [2047:0]     dataInMem_lo_131 = {dataInMem_lo_hi_3, dataInMem_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_lo_lo_lo_lo_3 = {dataInMem_hi_196, dataInMem_lo_68, dataInMem_hi_195, dataInMem_lo_67};
  wire [63:0]       dataInMem_hi_lo_lo_lo_lo_hi_3 = {dataInMem_hi_198, dataInMem_lo_70, dataInMem_hi_197, dataInMem_lo_69};
  wire [127:0]      dataInMem_hi_lo_lo_lo_lo_3 = {dataInMem_hi_lo_lo_lo_lo_hi_3, dataInMem_hi_lo_lo_lo_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_lo_lo_hi_lo_3 = {dataInMem_hi_200, dataInMem_lo_72, dataInMem_hi_199, dataInMem_lo_71};
  wire [63:0]       dataInMem_hi_lo_lo_lo_hi_hi_3 = {dataInMem_hi_202, dataInMem_lo_74, dataInMem_hi_201, dataInMem_lo_73};
  wire [127:0]      dataInMem_hi_lo_lo_lo_hi_3 = {dataInMem_hi_lo_lo_lo_hi_hi_3, dataInMem_hi_lo_lo_lo_hi_lo_3};
  wire [255:0]      dataInMem_hi_lo_lo_lo_3 = {dataInMem_hi_lo_lo_lo_hi_3, dataInMem_hi_lo_lo_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_lo_hi_lo_lo_3 = {dataInMem_hi_204, dataInMem_lo_76, dataInMem_hi_203, dataInMem_lo_75};
  wire [63:0]       dataInMem_hi_lo_lo_hi_lo_hi_3 = {dataInMem_hi_206, dataInMem_lo_78, dataInMem_hi_205, dataInMem_lo_77};
  wire [127:0]      dataInMem_hi_lo_lo_hi_lo_3 = {dataInMem_hi_lo_lo_hi_lo_hi_3, dataInMem_hi_lo_lo_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_lo_hi_hi_lo_3 = {dataInMem_hi_208, dataInMem_lo_80, dataInMem_hi_207, dataInMem_lo_79};
  wire [63:0]       dataInMem_hi_lo_lo_hi_hi_hi_3 = {dataInMem_hi_210, dataInMem_lo_82, dataInMem_hi_209, dataInMem_lo_81};
  wire [127:0]      dataInMem_hi_lo_lo_hi_hi_3 = {dataInMem_hi_lo_lo_hi_hi_hi_3, dataInMem_hi_lo_lo_hi_hi_lo_3};
  wire [255:0]      dataInMem_hi_lo_lo_hi_3 = {dataInMem_hi_lo_lo_hi_hi_3, dataInMem_hi_lo_lo_hi_lo_3};
  wire [511:0]      dataInMem_hi_lo_lo_3 = {dataInMem_hi_lo_lo_hi_3, dataInMem_hi_lo_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_hi_lo_lo_lo_3 = {dataInMem_hi_212, dataInMem_lo_84, dataInMem_hi_211, dataInMem_lo_83};
  wire [63:0]       dataInMem_hi_lo_hi_lo_lo_hi_3 = {dataInMem_hi_214, dataInMem_lo_86, dataInMem_hi_213, dataInMem_lo_85};
  wire [127:0]      dataInMem_hi_lo_hi_lo_lo_3 = {dataInMem_hi_lo_hi_lo_lo_hi_3, dataInMem_hi_lo_hi_lo_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_hi_lo_hi_lo_3 = {dataInMem_hi_216, dataInMem_lo_88, dataInMem_hi_215, dataInMem_lo_87};
  wire [63:0]       dataInMem_hi_lo_hi_lo_hi_hi_3 = {dataInMem_hi_218, dataInMem_lo_90, dataInMem_hi_217, dataInMem_lo_89};
  wire [127:0]      dataInMem_hi_lo_hi_lo_hi_3 = {dataInMem_hi_lo_hi_lo_hi_hi_3, dataInMem_hi_lo_hi_lo_hi_lo_3};
  wire [255:0]      dataInMem_hi_lo_hi_lo_3 = {dataInMem_hi_lo_hi_lo_hi_3, dataInMem_hi_lo_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_hi_hi_lo_lo_3 = {dataInMem_hi_220, dataInMem_lo_92, dataInMem_hi_219, dataInMem_lo_91};
  wire [63:0]       dataInMem_hi_lo_hi_hi_lo_hi_3 = {dataInMem_hi_222, dataInMem_lo_94, dataInMem_hi_221, dataInMem_lo_93};
  wire [127:0]      dataInMem_hi_lo_hi_hi_lo_3 = {dataInMem_hi_lo_hi_hi_lo_hi_3, dataInMem_hi_lo_hi_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_lo_hi_hi_hi_lo_3 = {dataInMem_hi_224, dataInMem_lo_96, dataInMem_hi_223, dataInMem_lo_95};
  wire [63:0]       dataInMem_hi_lo_hi_hi_hi_hi_3 = {dataInMem_hi_226, dataInMem_lo_98, dataInMem_hi_225, dataInMem_lo_97};
  wire [127:0]      dataInMem_hi_lo_hi_hi_hi_3 = {dataInMem_hi_lo_hi_hi_hi_hi_3, dataInMem_hi_lo_hi_hi_hi_lo_3};
  wire [255:0]      dataInMem_hi_lo_hi_hi_3 = {dataInMem_hi_lo_hi_hi_hi_3, dataInMem_hi_lo_hi_hi_lo_3};
  wire [511:0]      dataInMem_hi_lo_hi_3 = {dataInMem_hi_lo_hi_hi_3, dataInMem_hi_lo_hi_lo_3};
  wire [1023:0]     dataInMem_hi_lo_3 = {dataInMem_hi_lo_hi_3, dataInMem_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_lo_lo_lo_lo_3 = {dataInMem_hi_228, dataInMem_lo_100, dataInMem_hi_227, dataInMem_lo_99};
  wire [63:0]       dataInMem_hi_hi_lo_lo_lo_hi_3 = {dataInMem_hi_230, dataInMem_lo_102, dataInMem_hi_229, dataInMem_lo_101};
  wire [127:0]      dataInMem_hi_hi_lo_lo_lo_3 = {dataInMem_hi_hi_lo_lo_lo_hi_3, dataInMem_hi_hi_lo_lo_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_lo_lo_hi_lo_3 = {dataInMem_hi_232, dataInMem_lo_104, dataInMem_hi_231, dataInMem_lo_103};
  wire [63:0]       dataInMem_hi_hi_lo_lo_hi_hi_3 = {dataInMem_hi_234, dataInMem_lo_106, dataInMem_hi_233, dataInMem_lo_105};
  wire [127:0]      dataInMem_hi_hi_lo_lo_hi_3 = {dataInMem_hi_hi_lo_lo_hi_hi_3, dataInMem_hi_hi_lo_lo_hi_lo_3};
  wire [255:0]      dataInMem_hi_hi_lo_lo_3 = {dataInMem_hi_hi_lo_lo_hi_3, dataInMem_hi_hi_lo_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_lo_hi_lo_lo_3 = {dataInMem_hi_236, dataInMem_lo_108, dataInMem_hi_235, dataInMem_lo_107};
  wire [63:0]       dataInMem_hi_hi_lo_hi_lo_hi_3 = {dataInMem_hi_238, dataInMem_lo_110, dataInMem_hi_237, dataInMem_lo_109};
  wire [127:0]      dataInMem_hi_hi_lo_hi_lo_3 = {dataInMem_hi_hi_lo_hi_lo_hi_3, dataInMem_hi_hi_lo_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_lo_hi_hi_lo_3 = {dataInMem_hi_240, dataInMem_lo_112, dataInMem_hi_239, dataInMem_lo_111};
  wire [63:0]       dataInMem_hi_hi_lo_hi_hi_hi_3 = {dataInMem_hi_242, dataInMem_lo_114, dataInMem_hi_241, dataInMem_lo_113};
  wire [127:0]      dataInMem_hi_hi_lo_hi_hi_3 = {dataInMem_hi_hi_lo_hi_hi_hi_3, dataInMem_hi_hi_lo_hi_hi_lo_3};
  wire [255:0]      dataInMem_hi_hi_lo_hi_3 = {dataInMem_hi_hi_lo_hi_hi_3, dataInMem_hi_hi_lo_hi_lo_3};
  wire [511:0]      dataInMem_hi_hi_lo_3 = {dataInMem_hi_hi_lo_hi_3, dataInMem_hi_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_hi_lo_lo_lo_3 = {dataInMem_hi_244, dataInMem_lo_116, dataInMem_hi_243, dataInMem_lo_115};
  wire [63:0]       dataInMem_hi_hi_hi_lo_lo_hi_3 = {dataInMem_hi_246, dataInMem_lo_118, dataInMem_hi_245, dataInMem_lo_117};
  wire [127:0]      dataInMem_hi_hi_hi_lo_lo_3 = {dataInMem_hi_hi_hi_lo_lo_hi_3, dataInMem_hi_hi_hi_lo_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_hi_lo_hi_lo_3 = {dataInMem_hi_248, dataInMem_lo_120, dataInMem_hi_247, dataInMem_lo_119};
  wire [63:0]       dataInMem_hi_hi_hi_lo_hi_hi_3 = {dataInMem_hi_250, dataInMem_lo_122, dataInMem_hi_249, dataInMem_lo_121};
  wire [127:0]      dataInMem_hi_hi_hi_lo_hi_3 = {dataInMem_hi_hi_hi_lo_hi_hi_3, dataInMem_hi_hi_hi_lo_hi_lo_3};
  wire [255:0]      dataInMem_hi_hi_hi_lo_3 = {dataInMem_hi_hi_hi_lo_hi_3, dataInMem_hi_hi_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_hi_hi_lo_lo_3 = {dataInMem_hi_252, dataInMem_lo_124, dataInMem_hi_251, dataInMem_lo_123};
  wire [63:0]       dataInMem_hi_hi_hi_hi_lo_hi_3 = {dataInMem_hi_254, dataInMem_lo_126, dataInMem_hi_253, dataInMem_lo_125};
  wire [127:0]      dataInMem_hi_hi_hi_hi_lo_3 = {dataInMem_hi_hi_hi_hi_lo_hi_3, dataInMem_hi_hi_hi_hi_lo_lo_3};
  wire [63:0]       dataInMem_hi_hi_hi_hi_hi_lo_3 = {dataInMem_hi_256, dataInMem_lo_128, dataInMem_hi_255, dataInMem_lo_127};
  wire [63:0]       dataInMem_hi_hi_hi_hi_hi_hi_3 = {dataInMem_hi_258, dataInMem_lo_130, dataInMem_hi_257, dataInMem_lo_129};
  wire [127:0]      dataInMem_hi_hi_hi_hi_hi_3 = {dataInMem_hi_hi_hi_hi_hi_hi_3, dataInMem_hi_hi_hi_hi_hi_lo_3};
  wire [255:0]      dataInMem_hi_hi_hi_hi_3 = {dataInMem_hi_hi_hi_hi_hi_3, dataInMem_hi_hi_hi_hi_lo_3};
  wire [511:0]      dataInMem_hi_hi_hi_3 = {dataInMem_hi_hi_hi_hi_3, dataInMem_hi_hi_hi_lo_3};
  wire [1023:0]     dataInMem_hi_hi_3 = {dataInMem_hi_hi_hi_3, dataInMem_hi_hi_lo_3};
  wire [2047:0]     dataInMem_hi_259 = {dataInMem_hi_hi_3, dataInMem_hi_lo_3};
  wire [4095:0]     dataInMem_3 = {dataInMem_hi_259, dataInMem_lo_131};
  wire [1023:0]     regroupCacheLine_3_0 = dataInMem_3[1023:0];
  wire [1023:0]     regroupCacheLine_3_1 = dataInMem_3[2047:1024];
  wire [1023:0]     regroupCacheLine_3_2 = dataInMem_3[3071:2048];
  wire [1023:0]     regroupCacheLine_3_3 = dataInMem_3[4095:3072];
  wire [1023:0]     res_24 = regroupCacheLine_3_0;
  wire [1023:0]     res_25 = regroupCacheLine_3_1;
  wire [1023:0]     res_26 = regroupCacheLine_3_2;
  wire [1023:0]     res_27 = regroupCacheLine_3_3;
  wire [2047:0]     lo_lo_3 = {res_25, res_24};
  wire [2047:0]     lo_hi_3 = {res_27, res_26};
  wire [4095:0]     lo_3 = {lo_hi_3, lo_lo_3};
  wire [8191:0]     regroupLoadData_0_3 = {4096'h0, lo_3};
  wire [15:0]       _GEN_390 = {dataRegroupBySew_4_0, dataRegroupBySew_3_0};
  wire [15:0]       dataInMem_hi_hi_4;
  assign dataInMem_hi_hi_4 = _GEN_390;
  wire [15:0]       dataInMem_hi_lo_6;
  assign dataInMem_hi_lo_6 = _GEN_390;
  wire [23:0]       dataInMem_hi_260 = {dataInMem_hi_hi_4, dataRegroupBySew_2_0};
  wire [15:0]       _GEN_391 = {dataRegroupBySew_4_1, dataRegroupBySew_3_1};
  wire [15:0]       dataInMem_hi_hi_5;
  assign dataInMem_hi_hi_5 = _GEN_391;
  wire [15:0]       dataInMem_hi_lo_7;
  assign dataInMem_hi_lo_7 = _GEN_391;
  wire [23:0]       dataInMem_hi_261 = {dataInMem_hi_hi_5, dataRegroupBySew_2_1};
  wire [15:0]       _GEN_392 = {dataRegroupBySew_4_2, dataRegroupBySew_3_2};
  wire [15:0]       dataInMem_hi_hi_6;
  assign dataInMem_hi_hi_6 = _GEN_392;
  wire [15:0]       dataInMem_hi_lo_8;
  assign dataInMem_hi_lo_8 = _GEN_392;
  wire [23:0]       dataInMem_hi_262 = {dataInMem_hi_hi_6, dataRegroupBySew_2_2};
  wire [15:0]       _GEN_393 = {dataRegroupBySew_4_3, dataRegroupBySew_3_3};
  wire [15:0]       dataInMem_hi_hi_7;
  assign dataInMem_hi_hi_7 = _GEN_393;
  wire [15:0]       dataInMem_hi_lo_9;
  assign dataInMem_hi_lo_9 = _GEN_393;
  wire [23:0]       dataInMem_hi_263 = {dataInMem_hi_hi_7, dataRegroupBySew_2_3};
  wire [15:0]       _GEN_394 = {dataRegroupBySew_4_4, dataRegroupBySew_3_4};
  wire [15:0]       dataInMem_hi_hi_8;
  assign dataInMem_hi_hi_8 = _GEN_394;
  wire [15:0]       dataInMem_hi_lo_10;
  assign dataInMem_hi_lo_10 = _GEN_394;
  wire [23:0]       dataInMem_hi_264 = {dataInMem_hi_hi_8, dataRegroupBySew_2_4};
  wire [15:0]       _GEN_395 = {dataRegroupBySew_4_5, dataRegroupBySew_3_5};
  wire [15:0]       dataInMem_hi_hi_9;
  assign dataInMem_hi_hi_9 = _GEN_395;
  wire [15:0]       dataInMem_hi_lo_11;
  assign dataInMem_hi_lo_11 = _GEN_395;
  wire [23:0]       dataInMem_hi_265 = {dataInMem_hi_hi_9, dataRegroupBySew_2_5};
  wire [15:0]       _GEN_396 = {dataRegroupBySew_4_6, dataRegroupBySew_3_6};
  wire [15:0]       dataInMem_hi_hi_10;
  assign dataInMem_hi_hi_10 = _GEN_396;
  wire [15:0]       dataInMem_hi_lo_12;
  assign dataInMem_hi_lo_12 = _GEN_396;
  wire [23:0]       dataInMem_hi_266 = {dataInMem_hi_hi_10, dataRegroupBySew_2_6};
  wire [15:0]       _GEN_397 = {dataRegroupBySew_4_7, dataRegroupBySew_3_7};
  wire [15:0]       dataInMem_hi_hi_11;
  assign dataInMem_hi_hi_11 = _GEN_397;
  wire [15:0]       dataInMem_hi_lo_13;
  assign dataInMem_hi_lo_13 = _GEN_397;
  wire [23:0]       dataInMem_hi_267 = {dataInMem_hi_hi_11, dataRegroupBySew_2_7};
  wire [15:0]       _GEN_398 = {dataRegroupBySew_4_8, dataRegroupBySew_3_8};
  wire [15:0]       dataInMem_hi_hi_12;
  assign dataInMem_hi_hi_12 = _GEN_398;
  wire [15:0]       dataInMem_hi_lo_14;
  assign dataInMem_hi_lo_14 = _GEN_398;
  wire [23:0]       dataInMem_hi_268 = {dataInMem_hi_hi_12, dataRegroupBySew_2_8};
  wire [15:0]       _GEN_399 = {dataRegroupBySew_4_9, dataRegroupBySew_3_9};
  wire [15:0]       dataInMem_hi_hi_13;
  assign dataInMem_hi_hi_13 = _GEN_399;
  wire [15:0]       dataInMem_hi_lo_15;
  assign dataInMem_hi_lo_15 = _GEN_399;
  wire [23:0]       dataInMem_hi_269 = {dataInMem_hi_hi_13, dataRegroupBySew_2_9};
  wire [15:0]       _GEN_400 = {dataRegroupBySew_4_10, dataRegroupBySew_3_10};
  wire [15:0]       dataInMem_hi_hi_14;
  assign dataInMem_hi_hi_14 = _GEN_400;
  wire [15:0]       dataInMem_hi_lo_16;
  assign dataInMem_hi_lo_16 = _GEN_400;
  wire [23:0]       dataInMem_hi_270 = {dataInMem_hi_hi_14, dataRegroupBySew_2_10};
  wire [15:0]       _GEN_401 = {dataRegroupBySew_4_11, dataRegroupBySew_3_11};
  wire [15:0]       dataInMem_hi_hi_15;
  assign dataInMem_hi_hi_15 = _GEN_401;
  wire [15:0]       dataInMem_hi_lo_17;
  assign dataInMem_hi_lo_17 = _GEN_401;
  wire [23:0]       dataInMem_hi_271 = {dataInMem_hi_hi_15, dataRegroupBySew_2_11};
  wire [15:0]       _GEN_402 = {dataRegroupBySew_4_12, dataRegroupBySew_3_12};
  wire [15:0]       dataInMem_hi_hi_16;
  assign dataInMem_hi_hi_16 = _GEN_402;
  wire [15:0]       dataInMem_hi_lo_18;
  assign dataInMem_hi_lo_18 = _GEN_402;
  wire [23:0]       dataInMem_hi_272 = {dataInMem_hi_hi_16, dataRegroupBySew_2_12};
  wire [15:0]       _GEN_403 = {dataRegroupBySew_4_13, dataRegroupBySew_3_13};
  wire [15:0]       dataInMem_hi_hi_17;
  assign dataInMem_hi_hi_17 = _GEN_403;
  wire [15:0]       dataInMem_hi_lo_19;
  assign dataInMem_hi_lo_19 = _GEN_403;
  wire [23:0]       dataInMem_hi_273 = {dataInMem_hi_hi_17, dataRegroupBySew_2_13};
  wire [15:0]       _GEN_404 = {dataRegroupBySew_4_14, dataRegroupBySew_3_14};
  wire [15:0]       dataInMem_hi_hi_18;
  assign dataInMem_hi_hi_18 = _GEN_404;
  wire [15:0]       dataInMem_hi_lo_20;
  assign dataInMem_hi_lo_20 = _GEN_404;
  wire [23:0]       dataInMem_hi_274 = {dataInMem_hi_hi_18, dataRegroupBySew_2_14};
  wire [15:0]       _GEN_405 = {dataRegroupBySew_4_15, dataRegroupBySew_3_15};
  wire [15:0]       dataInMem_hi_hi_19;
  assign dataInMem_hi_hi_19 = _GEN_405;
  wire [15:0]       dataInMem_hi_lo_21;
  assign dataInMem_hi_lo_21 = _GEN_405;
  wire [23:0]       dataInMem_hi_275 = {dataInMem_hi_hi_19, dataRegroupBySew_2_15};
  wire [15:0]       _GEN_406 = {dataRegroupBySew_4_16, dataRegroupBySew_3_16};
  wire [15:0]       dataInMem_hi_hi_20;
  assign dataInMem_hi_hi_20 = _GEN_406;
  wire [15:0]       dataInMem_hi_lo_22;
  assign dataInMem_hi_lo_22 = _GEN_406;
  wire [23:0]       dataInMem_hi_276 = {dataInMem_hi_hi_20, dataRegroupBySew_2_16};
  wire [15:0]       _GEN_407 = {dataRegroupBySew_4_17, dataRegroupBySew_3_17};
  wire [15:0]       dataInMem_hi_hi_21;
  assign dataInMem_hi_hi_21 = _GEN_407;
  wire [15:0]       dataInMem_hi_lo_23;
  assign dataInMem_hi_lo_23 = _GEN_407;
  wire [23:0]       dataInMem_hi_277 = {dataInMem_hi_hi_21, dataRegroupBySew_2_17};
  wire [15:0]       _GEN_408 = {dataRegroupBySew_4_18, dataRegroupBySew_3_18};
  wire [15:0]       dataInMem_hi_hi_22;
  assign dataInMem_hi_hi_22 = _GEN_408;
  wire [15:0]       dataInMem_hi_lo_24;
  assign dataInMem_hi_lo_24 = _GEN_408;
  wire [23:0]       dataInMem_hi_278 = {dataInMem_hi_hi_22, dataRegroupBySew_2_18};
  wire [15:0]       _GEN_409 = {dataRegroupBySew_4_19, dataRegroupBySew_3_19};
  wire [15:0]       dataInMem_hi_hi_23;
  assign dataInMem_hi_hi_23 = _GEN_409;
  wire [15:0]       dataInMem_hi_lo_25;
  assign dataInMem_hi_lo_25 = _GEN_409;
  wire [23:0]       dataInMem_hi_279 = {dataInMem_hi_hi_23, dataRegroupBySew_2_19};
  wire [15:0]       _GEN_410 = {dataRegroupBySew_4_20, dataRegroupBySew_3_20};
  wire [15:0]       dataInMem_hi_hi_24;
  assign dataInMem_hi_hi_24 = _GEN_410;
  wire [15:0]       dataInMem_hi_lo_26;
  assign dataInMem_hi_lo_26 = _GEN_410;
  wire [23:0]       dataInMem_hi_280 = {dataInMem_hi_hi_24, dataRegroupBySew_2_20};
  wire [15:0]       _GEN_411 = {dataRegroupBySew_4_21, dataRegroupBySew_3_21};
  wire [15:0]       dataInMem_hi_hi_25;
  assign dataInMem_hi_hi_25 = _GEN_411;
  wire [15:0]       dataInMem_hi_lo_27;
  assign dataInMem_hi_lo_27 = _GEN_411;
  wire [23:0]       dataInMem_hi_281 = {dataInMem_hi_hi_25, dataRegroupBySew_2_21};
  wire [15:0]       _GEN_412 = {dataRegroupBySew_4_22, dataRegroupBySew_3_22};
  wire [15:0]       dataInMem_hi_hi_26;
  assign dataInMem_hi_hi_26 = _GEN_412;
  wire [15:0]       dataInMem_hi_lo_28;
  assign dataInMem_hi_lo_28 = _GEN_412;
  wire [23:0]       dataInMem_hi_282 = {dataInMem_hi_hi_26, dataRegroupBySew_2_22};
  wire [15:0]       _GEN_413 = {dataRegroupBySew_4_23, dataRegroupBySew_3_23};
  wire [15:0]       dataInMem_hi_hi_27;
  assign dataInMem_hi_hi_27 = _GEN_413;
  wire [15:0]       dataInMem_hi_lo_29;
  assign dataInMem_hi_lo_29 = _GEN_413;
  wire [23:0]       dataInMem_hi_283 = {dataInMem_hi_hi_27, dataRegroupBySew_2_23};
  wire [15:0]       _GEN_414 = {dataRegroupBySew_4_24, dataRegroupBySew_3_24};
  wire [15:0]       dataInMem_hi_hi_28;
  assign dataInMem_hi_hi_28 = _GEN_414;
  wire [15:0]       dataInMem_hi_lo_30;
  assign dataInMem_hi_lo_30 = _GEN_414;
  wire [23:0]       dataInMem_hi_284 = {dataInMem_hi_hi_28, dataRegroupBySew_2_24};
  wire [15:0]       _GEN_415 = {dataRegroupBySew_4_25, dataRegroupBySew_3_25};
  wire [15:0]       dataInMem_hi_hi_29;
  assign dataInMem_hi_hi_29 = _GEN_415;
  wire [15:0]       dataInMem_hi_lo_31;
  assign dataInMem_hi_lo_31 = _GEN_415;
  wire [23:0]       dataInMem_hi_285 = {dataInMem_hi_hi_29, dataRegroupBySew_2_25};
  wire [15:0]       _GEN_416 = {dataRegroupBySew_4_26, dataRegroupBySew_3_26};
  wire [15:0]       dataInMem_hi_hi_30;
  assign dataInMem_hi_hi_30 = _GEN_416;
  wire [15:0]       dataInMem_hi_lo_32;
  assign dataInMem_hi_lo_32 = _GEN_416;
  wire [23:0]       dataInMem_hi_286 = {dataInMem_hi_hi_30, dataRegroupBySew_2_26};
  wire [15:0]       _GEN_417 = {dataRegroupBySew_4_27, dataRegroupBySew_3_27};
  wire [15:0]       dataInMem_hi_hi_31;
  assign dataInMem_hi_hi_31 = _GEN_417;
  wire [15:0]       dataInMem_hi_lo_33;
  assign dataInMem_hi_lo_33 = _GEN_417;
  wire [23:0]       dataInMem_hi_287 = {dataInMem_hi_hi_31, dataRegroupBySew_2_27};
  wire [15:0]       _GEN_418 = {dataRegroupBySew_4_28, dataRegroupBySew_3_28};
  wire [15:0]       dataInMem_hi_hi_32;
  assign dataInMem_hi_hi_32 = _GEN_418;
  wire [15:0]       dataInMem_hi_lo_34;
  assign dataInMem_hi_lo_34 = _GEN_418;
  wire [23:0]       dataInMem_hi_288 = {dataInMem_hi_hi_32, dataRegroupBySew_2_28};
  wire [15:0]       _GEN_419 = {dataRegroupBySew_4_29, dataRegroupBySew_3_29};
  wire [15:0]       dataInMem_hi_hi_33;
  assign dataInMem_hi_hi_33 = _GEN_419;
  wire [15:0]       dataInMem_hi_lo_35;
  assign dataInMem_hi_lo_35 = _GEN_419;
  wire [23:0]       dataInMem_hi_289 = {dataInMem_hi_hi_33, dataRegroupBySew_2_29};
  wire [15:0]       _GEN_420 = {dataRegroupBySew_4_30, dataRegroupBySew_3_30};
  wire [15:0]       dataInMem_hi_hi_34;
  assign dataInMem_hi_hi_34 = _GEN_420;
  wire [15:0]       dataInMem_hi_lo_36;
  assign dataInMem_hi_lo_36 = _GEN_420;
  wire [23:0]       dataInMem_hi_290 = {dataInMem_hi_hi_34, dataRegroupBySew_2_30};
  wire [15:0]       _GEN_421 = {dataRegroupBySew_4_31, dataRegroupBySew_3_31};
  wire [15:0]       dataInMem_hi_hi_35;
  assign dataInMem_hi_hi_35 = _GEN_421;
  wire [15:0]       dataInMem_hi_lo_37;
  assign dataInMem_hi_lo_37 = _GEN_421;
  wire [23:0]       dataInMem_hi_291 = {dataInMem_hi_hi_35, dataRegroupBySew_2_31};
  wire [15:0]       _GEN_422 = {dataRegroupBySew_4_32, dataRegroupBySew_3_32};
  wire [15:0]       dataInMem_hi_hi_36;
  assign dataInMem_hi_hi_36 = _GEN_422;
  wire [15:0]       dataInMem_hi_lo_38;
  assign dataInMem_hi_lo_38 = _GEN_422;
  wire [23:0]       dataInMem_hi_292 = {dataInMem_hi_hi_36, dataRegroupBySew_2_32};
  wire [15:0]       _GEN_423 = {dataRegroupBySew_4_33, dataRegroupBySew_3_33};
  wire [15:0]       dataInMem_hi_hi_37;
  assign dataInMem_hi_hi_37 = _GEN_423;
  wire [15:0]       dataInMem_hi_lo_39;
  assign dataInMem_hi_lo_39 = _GEN_423;
  wire [23:0]       dataInMem_hi_293 = {dataInMem_hi_hi_37, dataRegroupBySew_2_33};
  wire [15:0]       _GEN_424 = {dataRegroupBySew_4_34, dataRegroupBySew_3_34};
  wire [15:0]       dataInMem_hi_hi_38;
  assign dataInMem_hi_hi_38 = _GEN_424;
  wire [15:0]       dataInMem_hi_lo_40;
  assign dataInMem_hi_lo_40 = _GEN_424;
  wire [23:0]       dataInMem_hi_294 = {dataInMem_hi_hi_38, dataRegroupBySew_2_34};
  wire [15:0]       _GEN_425 = {dataRegroupBySew_4_35, dataRegroupBySew_3_35};
  wire [15:0]       dataInMem_hi_hi_39;
  assign dataInMem_hi_hi_39 = _GEN_425;
  wire [15:0]       dataInMem_hi_lo_41;
  assign dataInMem_hi_lo_41 = _GEN_425;
  wire [23:0]       dataInMem_hi_295 = {dataInMem_hi_hi_39, dataRegroupBySew_2_35};
  wire [15:0]       _GEN_426 = {dataRegroupBySew_4_36, dataRegroupBySew_3_36};
  wire [15:0]       dataInMem_hi_hi_40;
  assign dataInMem_hi_hi_40 = _GEN_426;
  wire [15:0]       dataInMem_hi_lo_42;
  assign dataInMem_hi_lo_42 = _GEN_426;
  wire [23:0]       dataInMem_hi_296 = {dataInMem_hi_hi_40, dataRegroupBySew_2_36};
  wire [15:0]       _GEN_427 = {dataRegroupBySew_4_37, dataRegroupBySew_3_37};
  wire [15:0]       dataInMem_hi_hi_41;
  assign dataInMem_hi_hi_41 = _GEN_427;
  wire [15:0]       dataInMem_hi_lo_43;
  assign dataInMem_hi_lo_43 = _GEN_427;
  wire [23:0]       dataInMem_hi_297 = {dataInMem_hi_hi_41, dataRegroupBySew_2_37};
  wire [15:0]       _GEN_428 = {dataRegroupBySew_4_38, dataRegroupBySew_3_38};
  wire [15:0]       dataInMem_hi_hi_42;
  assign dataInMem_hi_hi_42 = _GEN_428;
  wire [15:0]       dataInMem_hi_lo_44;
  assign dataInMem_hi_lo_44 = _GEN_428;
  wire [23:0]       dataInMem_hi_298 = {dataInMem_hi_hi_42, dataRegroupBySew_2_38};
  wire [15:0]       _GEN_429 = {dataRegroupBySew_4_39, dataRegroupBySew_3_39};
  wire [15:0]       dataInMem_hi_hi_43;
  assign dataInMem_hi_hi_43 = _GEN_429;
  wire [15:0]       dataInMem_hi_lo_45;
  assign dataInMem_hi_lo_45 = _GEN_429;
  wire [23:0]       dataInMem_hi_299 = {dataInMem_hi_hi_43, dataRegroupBySew_2_39};
  wire [15:0]       _GEN_430 = {dataRegroupBySew_4_40, dataRegroupBySew_3_40};
  wire [15:0]       dataInMem_hi_hi_44;
  assign dataInMem_hi_hi_44 = _GEN_430;
  wire [15:0]       dataInMem_hi_lo_46;
  assign dataInMem_hi_lo_46 = _GEN_430;
  wire [23:0]       dataInMem_hi_300 = {dataInMem_hi_hi_44, dataRegroupBySew_2_40};
  wire [15:0]       _GEN_431 = {dataRegroupBySew_4_41, dataRegroupBySew_3_41};
  wire [15:0]       dataInMem_hi_hi_45;
  assign dataInMem_hi_hi_45 = _GEN_431;
  wire [15:0]       dataInMem_hi_lo_47;
  assign dataInMem_hi_lo_47 = _GEN_431;
  wire [23:0]       dataInMem_hi_301 = {dataInMem_hi_hi_45, dataRegroupBySew_2_41};
  wire [15:0]       _GEN_432 = {dataRegroupBySew_4_42, dataRegroupBySew_3_42};
  wire [15:0]       dataInMem_hi_hi_46;
  assign dataInMem_hi_hi_46 = _GEN_432;
  wire [15:0]       dataInMem_hi_lo_48;
  assign dataInMem_hi_lo_48 = _GEN_432;
  wire [23:0]       dataInMem_hi_302 = {dataInMem_hi_hi_46, dataRegroupBySew_2_42};
  wire [15:0]       _GEN_433 = {dataRegroupBySew_4_43, dataRegroupBySew_3_43};
  wire [15:0]       dataInMem_hi_hi_47;
  assign dataInMem_hi_hi_47 = _GEN_433;
  wire [15:0]       dataInMem_hi_lo_49;
  assign dataInMem_hi_lo_49 = _GEN_433;
  wire [23:0]       dataInMem_hi_303 = {dataInMem_hi_hi_47, dataRegroupBySew_2_43};
  wire [15:0]       _GEN_434 = {dataRegroupBySew_4_44, dataRegroupBySew_3_44};
  wire [15:0]       dataInMem_hi_hi_48;
  assign dataInMem_hi_hi_48 = _GEN_434;
  wire [15:0]       dataInMem_hi_lo_50;
  assign dataInMem_hi_lo_50 = _GEN_434;
  wire [23:0]       dataInMem_hi_304 = {dataInMem_hi_hi_48, dataRegroupBySew_2_44};
  wire [15:0]       _GEN_435 = {dataRegroupBySew_4_45, dataRegroupBySew_3_45};
  wire [15:0]       dataInMem_hi_hi_49;
  assign dataInMem_hi_hi_49 = _GEN_435;
  wire [15:0]       dataInMem_hi_lo_51;
  assign dataInMem_hi_lo_51 = _GEN_435;
  wire [23:0]       dataInMem_hi_305 = {dataInMem_hi_hi_49, dataRegroupBySew_2_45};
  wire [15:0]       _GEN_436 = {dataRegroupBySew_4_46, dataRegroupBySew_3_46};
  wire [15:0]       dataInMem_hi_hi_50;
  assign dataInMem_hi_hi_50 = _GEN_436;
  wire [15:0]       dataInMem_hi_lo_52;
  assign dataInMem_hi_lo_52 = _GEN_436;
  wire [23:0]       dataInMem_hi_306 = {dataInMem_hi_hi_50, dataRegroupBySew_2_46};
  wire [15:0]       _GEN_437 = {dataRegroupBySew_4_47, dataRegroupBySew_3_47};
  wire [15:0]       dataInMem_hi_hi_51;
  assign dataInMem_hi_hi_51 = _GEN_437;
  wire [15:0]       dataInMem_hi_lo_53;
  assign dataInMem_hi_lo_53 = _GEN_437;
  wire [23:0]       dataInMem_hi_307 = {dataInMem_hi_hi_51, dataRegroupBySew_2_47};
  wire [15:0]       _GEN_438 = {dataRegroupBySew_4_48, dataRegroupBySew_3_48};
  wire [15:0]       dataInMem_hi_hi_52;
  assign dataInMem_hi_hi_52 = _GEN_438;
  wire [15:0]       dataInMem_hi_lo_54;
  assign dataInMem_hi_lo_54 = _GEN_438;
  wire [23:0]       dataInMem_hi_308 = {dataInMem_hi_hi_52, dataRegroupBySew_2_48};
  wire [15:0]       _GEN_439 = {dataRegroupBySew_4_49, dataRegroupBySew_3_49};
  wire [15:0]       dataInMem_hi_hi_53;
  assign dataInMem_hi_hi_53 = _GEN_439;
  wire [15:0]       dataInMem_hi_lo_55;
  assign dataInMem_hi_lo_55 = _GEN_439;
  wire [23:0]       dataInMem_hi_309 = {dataInMem_hi_hi_53, dataRegroupBySew_2_49};
  wire [15:0]       _GEN_440 = {dataRegroupBySew_4_50, dataRegroupBySew_3_50};
  wire [15:0]       dataInMem_hi_hi_54;
  assign dataInMem_hi_hi_54 = _GEN_440;
  wire [15:0]       dataInMem_hi_lo_56;
  assign dataInMem_hi_lo_56 = _GEN_440;
  wire [23:0]       dataInMem_hi_310 = {dataInMem_hi_hi_54, dataRegroupBySew_2_50};
  wire [15:0]       _GEN_441 = {dataRegroupBySew_4_51, dataRegroupBySew_3_51};
  wire [15:0]       dataInMem_hi_hi_55;
  assign dataInMem_hi_hi_55 = _GEN_441;
  wire [15:0]       dataInMem_hi_lo_57;
  assign dataInMem_hi_lo_57 = _GEN_441;
  wire [23:0]       dataInMem_hi_311 = {dataInMem_hi_hi_55, dataRegroupBySew_2_51};
  wire [15:0]       _GEN_442 = {dataRegroupBySew_4_52, dataRegroupBySew_3_52};
  wire [15:0]       dataInMem_hi_hi_56;
  assign dataInMem_hi_hi_56 = _GEN_442;
  wire [15:0]       dataInMem_hi_lo_58;
  assign dataInMem_hi_lo_58 = _GEN_442;
  wire [23:0]       dataInMem_hi_312 = {dataInMem_hi_hi_56, dataRegroupBySew_2_52};
  wire [15:0]       _GEN_443 = {dataRegroupBySew_4_53, dataRegroupBySew_3_53};
  wire [15:0]       dataInMem_hi_hi_57;
  assign dataInMem_hi_hi_57 = _GEN_443;
  wire [15:0]       dataInMem_hi_lo_59;
  assign dataInMem_hi_lo_59 = _GEN_443;
  wire [23:0]       dataInMem_hi_313 = {dataInMem_hi_hi_57, dataRegroupBySew_2_53};
  wire [15:0]       _GEN_444 = {dataRegroupBySew_4_54, dataRegroupBySew_3_54};
  wire [15:0]       dataInMem_hi_hi_58;
  assign dataInMem_hi_hi_58 = _GEN_444;
  wire [15:0]       dataInMem_hi_lo_60;
  assign dataInMem_hi_lo_60 = _GEN_444;
  wire [23:0]       dataInMem_hi_314 = {dataInMem_hi_hi_58, dataRegroupBySew_2_54};
  wire [15:0]       _GEN_445 = {dataRegroupBySew_4_55, dataRegroupBySew_3_55};
  wire [15:0]       dataInMem_hi_hi_59;
  assign dataInMem_hi_hi_59 = _GEN_445;
  wire [15:0]       dataInMem_hi_lo_61;
  assign dataInMem_hi_lo_61 = _GEN_445;
  wire [23:0]       dataInMem_hi_315 = {dataInMem_hi_hi_59, dataRegroupBySew_2_55};
  wire [15:0]       _GEN_446 = {dataRegroupBySew_4_56, dataRegroupBySew_3_56};
  wire [15:0]       dataInMem_hi_hi_60;
  assign dataInMem_hi_hi_60 = _GEN_446;
  wire [15:0]       dataInMem_hi_lo_62;
  assign dataInMem_hi_lo_62 = _GEN_446;
  wire [23:0]       dataInMem_hi_316 = {dataInMem_hi_hi_60, dataRegroupBySew_2_56};
  wire [15:0]       _GEN_447 = {dataRegroupBySew_4_57, dataRegroupBySew_3_57};
  wire [15:0]       dataInMem_hi_hi_61;
  assign dataInMem_hi_hi_61 = _GEN_447;
  wire [15:0]       dataInMem_hi_lo_63;
  assign dataInMem_hi_lo_63 = _GEN_447;
  wire [23:0]       dataInMem_hi_317 = {dataInMem_hi_hi_61, dataRegroupBySew_2_57};
  wire [15:0]       _GEN_448 = {dataRegroupBySew_4_58, dataRegroupBySew_3_58};
  wire [15:0]       dataInMem_hi_hi_62;
  assign dataInMem_hi_hi_62 = _GEN_448;
  wire [15:0]       dataInMem_hi_lo_64;
  assign dataInMem_hi_lo_64 = _GEN_448;
  wire [23:0]       dataInMem_hi_318 = {dataInMem_hi_hi_62, dataRegroupBySew_2_58};
  wire [15:0]       _GEN_449 = {dataRegroupBySew_4_59, dataRegroupBySew_3_59};
  wire [15:0]       dataInMem_hi_hi_63;
  assign dataInMem_hi_hi_63 = _GEN_449;
  wire [15:0]       dataInMem_hi_lo_65;
  assign dataInMem_hi_lo_65 = _GEN_449;
  wire [23:0]       dataInMem_hi_319 = {dataInMem_hi_hi_63, dataRegroupBySew_2_59};
  wire [15:0]       _GEN_450 = {dataRegroupBySew_4_60, dataRegroupBySew_3_60};
  wire [15:0]       dataInMem_hi_hi_64;
  assign dataInMem_hi_hi_64 = _GEN_450;
  wire [15:0]       dataInMem_hi_lo_66;
  assign dataInMem_hi_lo_66 = _GEN_450;
  wire [23:0]       dataInMem_hi_320 = {dataInMem_hi_hi_64, dataRegroupBySew_2_60};
  wire [15:0]       _GEN_451 = {dataRegroupBySew_4_61, dataRegroupBySew_3_61};
  wire [15:0]       dataInMem_hi_hi_65;
  assign dataInMem_hi_hi_65 = _GEN_451;
  wire [15:0]       dataInMem_hi_lo_67;
  assign dataInMem_hi_lo_67 = _GEN_451;
  wire [23:0]       dataInMem_hi_321 = {dataInMem_hi_hi_65, dataRegroupBySew_2_61};
  wire [15:0]       _GEN_452 = {dataRegroupBySew_4_62, dataRegroupBySew_3_62};
  wire [15:0]       dataInMem_hi_hi_66;
  assign dataInMem_hi_hi_66 = _GEN_452;
  wire [15:0]       dataInMem_hi_lo_68;
  assign dataInMem_hi_lo_68 = _GEN_452;
  wire [23:0]       dataInMem_hi_322 = {dataInMem_hi_hi_66, dataRegroupBySew_2_62};
  wire [15:0]       _GEN_453 = {dataRegroupBySew_4_63, dataRegroupBySew_3_63};
  wire [15:0]       dataInMem_hi_hi_67;
  assign dataInMem_hi_hi_67 = _GEN_453;
  wire [15:0]       dataInMem_hi_lo_69;
  assign dataInMem_hi_lo_69 = _GEN_453;
  wire [23:0]       dataInMem_hi_323 = {dataInMem_hi_hi_67, dataRegroupBySew_2_63};
  wire [15:0]       _GEN_454 = {dataRegroupBySew_4_64, dataRegroupBySew_3_64};
  wire [15:0]       dataInMem_hi_hi_68;
  assign dataInMem_hi_hi_68 = _GEN_454;
  wire [15:0]       dataInMem_hi_lo_70;
  assign dataInMem_hi_lo_70 = _GEN_454;
  wire [23:0]       dataInMem_hi_324 = {dataInMem_hi_hi_68, dataRegroupBySew_2_64};
  wire [15:0]       _GEN_455 = {dataRegroupBySew_4_65, dataRegroupBySew_3_65};
  wire [15:0]       dataInMem_hi_hi_69;
  assign dataInMem_hi_hi_69 = _GEN_455;
  wire [15:0]       dataInMem_hi_lo_71;
  assign dataInMem_hi_lo_71 = _GEN_455;
  wire [23:0]       dataInMem_hi_325 = {dataInMem_hi_hi_69, dataRegroupBySew_2_65};
  wire [15:0]       _GEN_456 = {dataRegroupBySew_4_66, dataRegroupBySew_3_66};
  wire [15:0]       dataInMem_hi_hi_70;
  assign dataInMem_hi_hi_70 = _GEN_456;
  wire [15:0]       dataInMem_hi_lo_72;
  assign dataInMem_hi_lo_72 = _GEN_456;
  wire [23:0]       dataInMem_hi_326 = {dataInMem_hi_hi_70, dataRegroupBySew_2_66};
  wire [15:0]       _GEN_457 = {dataRegroupBySew_4_67, dataRegroupBySew_3_67};
  wire [15:0]       dataInMem_hi_hi_71;
  assign dataInMem_hi_hi_71 = _GEN_457;
  wire [15:0]       dataInMem_hi_lo_73;
  assign dataInMem_hi_lo_73 = _GEN_457;
  wire [23:0]       dataInMem_hi_327 = {dataInMem_hi_hi_71, dataRegroupBySew_2_67};
  wire [15:0]       _GEN_458 = {dataRegroupBySew_4_68, dataRegroupBySew_3_68};
  wire [15:0]       dataInMem_hi_hi_72;
  assign dataInMem_hi_hi_72 = _GEN_458;
  wire [15:0]       dataInMem_hi_lo_74;
  assign dataInMem_hi_lo_74 = _GEN_458;
  wire [23:0]       dataInMem_hi_328 = {dataInMem_hi_hi_72, dataRegroupBySew_2_68};
  wire [15:0]       _GEN_459 = {dataRegroupBySew_4_69, dataRegroupBySew_3_69};
  wire [15:0]       dataInMem_hi_hi_73;
  assign dataInMem_hi_hi_73 = _GEN_459;
  wire [15:0]       dataInMem_hi_lo_75;
  assign dataInMem_hi_lo_75 = _GEN_459;
  wire [23:0]       dataInMem_hi_329 = {dataInMem_hi_hi_73, dataRegroupBySew_2_69};
  wire [15:0]       _GEN_460 = {dataRegroupBySew_4_70, dataRegroupBySew_3_70};
  wire [15:0]       dataInMem_hi_hi_74;
  assign dataInMem_hi_hi_74 = _GEN_460;
  wire [15:0]       dataInMem_hi_lo_76;
  assign dataInMem_hi_lo_76 = _GEN_460;
  wire [23:0]       dataInMem_hi_330 = {dataInMem_hi_hi_74, dataRegroupBySew_2_70};
  wire [15:0]       _GEN_461 = {dataRegroupBySew_4_71, dataRegroupBySew_3_71};
  wire [15:0]       dataInMem_hi_hi_75;
  assign dataInMem_hi_hi_75 = _GEN_461;
  wire [15:0]       dataInMem_hi_lo_77;
  assign dataInMem_hi_lo_77 = _GEN_461;
  wire [23:0]       dataInMem_hi_331 = {dataInMem_hi_hi_75, dataRegroupBySew_2_71};
  wire [15:0]       _GEN_462 = {dataRegroupBySew_4_72, dataRegroupBySew_3_72};
  wire [15:0]       dataInMem_hi_hi_76;
  assign dataInMem_hi_hi_76 = _GEN_462;
  wire [15:0]       dataInMem_hi_lo_78;
  assign dataInMem_hi_lo_78 = _GEN_462;
  wire [23:0]       dataInMem_hi_332 = {dataInMem_hi_hi_76, dataRegroupBySew_2_72};
  wire [15:0]       _GEN_463 = {dataRegroupBySew_4_73, dataRegroupBySew_3_73};
  wire [15:0]       dataInMem_hi_hi_77;
  assign dataInMem_hi_hi_77 = _GEN_463;
  wire [15:0]       dataInMem_hi_lo_79;
  assign dataInMem_hi_lo_79 = _GEN_463;
  wire [23:0]       dataInMem_hi_333 = {dataInMem_hi_hi_77, dataRegroupBySew_2_73};
  wire [15:0]       _GEN_464 = {dataRegroupBySew_4_74, dataRegroupBySew_3_74};
  wire [15:0]       dataInMem_hi_hi_78;
  assign dataInMem_hi_hi_78 = _GEN_464;
  wire [15:0]       dataInMem_hi_lo_80;
  assign dataInMem_hi_lo_80 = _GEN_464;
  wire [23:0]       dataInMem_hi_334 = {dataInMem_hi_hi_78, dataRegroupBySew_2_74};
  wire [15:0]       _GEN_465 = {dataRegroupBySew_4_75, dataRegroupBySew_3_75};
  wire [15:0]       dataInMem_hi_hi_79;
  assign dataInMem_hi_hi_79 = _GEN_465;
  wire [15:0]       dataInMem_hi_lo_81;
  assign dataInMem_hi_lo_81 = _GEN_465;
  wire [23:0]       dataInMem_hi_335 = {dataInMem_hi_hi_79, dataRegroupBySew_2_75};
  wire [15:0]       _GEN_466 = {dataRegroupBySew_4_76, dataRegroupBySew_3_76};
  wire [15:0]       dataInMem_hi_hi_80;
  assign dataInMem_hi_hi_80 = _GEN_466;
  wire [15:0]       dataInMem_hi_lo_82;
  assign dataInMem_hi_lo_82 = _GEN_466;
  wire [23:0]       dataInMem_hi_336 = {dataInMem_hi_hi_80, dataRegroupBySew_2_76};
  wire [15:0]       _GEN_467 = {dataRegroupBySew_4_77, dataRegroupBySew_3_77};
  wire [15:0]       dataInMem_hi_hi_81;
  assign dataInMem_hi_hi_81 = _GEN_467;
  wire [15:0]       dataInMem_hi_lo_83;
  assign dataInMem_hi_lo_83 = _GEN_467;
  wire [23:0]       dataInMem_hi_337 = {dataInMem_hi_hi_81, dataRegroupBySew_2_77};
  wire [15:0]       _GEN_468 = {dataRegroupBySew_4_78, dataRegroupBySew_3_78};
  wire [15:0]       dataInMem_hi_hi_82;
  assign dataInMem_hi_hi_82 = _GEN_468;
  wire [15:0]       dataInMem_hi_lo_84;
  assign dataInMem_hi_lo_84 = _GEN_468;
  wire [23:0]       dataInMem_hi_338 = {dataInMem_hi_hi_82, dataRegroupBySew_2_78};
  wire [15:0]       _GEN_469 = {dataRegroupBySew_4_79, dataRegroupBySew_3_79};
  wire [15:0]       dataInMem_hi_hi_83;
  assign dataInMem_hi_hi_83 = _GEN_469;
  wire [15:0]       dataInMem_hi_lo_85;
  assign dataInMem_hi_lo_85 = _GEN_469;
  wire [23:0]       dataInMem_hi_339 = {dataInMem_hi_hi_83, dataRegroupBySew_2_79};
  wire [15:0]       _GEN_470 = {dataRegroupBySew_4_80, dataRegroupBySew_3_80};
  wire [15:0]       dataInMem_hi_hi_84;
  assign dataInMem_hi_hi_84 = _GEN_470;
  wire [15:0]       dataInMem_hi_lo_86;
  assign dataInMem_hi_lo_86 = _GEN_470;
  wire [23:0]       dataInMem_hi_340 = {dataInMem_hi_hi_84, dataRegroupBySew_2_80};
  wire [15:0]       _GEN_471 = {dataRegroupBySew_4_81, dataRegroupBySew_3_81};
  wire [15:0]       dataInMem_hi_hi_85;
  assign dataInMem_hi_hi_85 = _GEN_471;
  wire [15:0]       dataInMem_hi_lo_87;
  assign dataInMem_hi_lo_87 = _GEN_471;
  wire [23:0]       dataInMem_hi_341 = {dataInMem_hi_hi_85, dataRegroupBySew_2_81};
  wire [15:0]       _GEN_472 = {dataRegroupBySew_4_82, dataRegroupBySew_3_82};
  wire [15:0]       dataInMem_hi_hi_86;
  assign dataInMem_hi_hi_86 = _GEN_472;
  wire [15:0]       dataInMem_hi_lo_88;
  assign dataInMem_hi_lo_88 = _GEN_472;
  wire [23:0]       dataInMem_hi_342 = {dataInMem_hi_hi_86, dataRegroupBySew_2_82};
  wire [15:0]       _GEN_473 = {dataRegroupBySew_4_83, dataRegroupBySew_3_83};
  wire [15:0]       dataInMem_hi_hi_87;
  assign dataInMem_hi_hi_87 = _GEN_473;
  wire [15:0]       dataInMem_hi_lo_89;
  assign dataInMem_hi_lo_89 = _GEN_473;
  wire [23:0]       dataInMem_hi_343 = {dataInMem_hi_hi_87, dataRegroupBySew_2_83};
  wire [15:0]       _GEN_474 = {dataRegroupBySew_4_84, dataRegroupBySew_3_84};
  wire [15:0]       dataInMem_hi_hi_88;
  assign dataInMem_hi_hi_88 = _GEN_474;
  wire [15:0]       dataInMem_hi_lo_90;
  assign dataInMem_hi_lo_90 = _GEN_474;
  wire [23:0]       dataInMem_hi_344 = {dataInMem_hi_hi_88, dataRegroupBySew_2_84};
  wire [15:0]       _GEN_475 = {dataRegroupBySew_4_85, dataRegroupBySew_3_85};
  wire [15:0]       dataInMem_hi_hi_89;
  assign dataInMem_hi_hi_89 = _GEN_475;
  wire [15:0]       dataInMem_hi_lo_91;
  assign dataInMem_hi_lo_91 = _GEN_475;
  wire [23:0]       dataInMem_hi_345 = {dataInMem_hi_hi_89, dataRegroupBySew_2_85};
  wire [15:0]       _GEN_476 = {dataRegroupBySew_4_86, dataRegroupBySew_3_86};
  wire [15:0]       dataInMem_hi_hi_90;
  assign dataInMem_hi_hi_90 = _GEN_476;
  wire [15:0]       dataInMem_hi_lo_92;
  assign dataInMem_hi_lo_92 = _GEN_476;
  wire [23:0]       dataInMem_hi_346 = {dataInMem_hi_hi_90, dataRegroupBySew_2_86};
  wire [15:0]       _GEN_477 = {dataRegroupBySew_4_87, dataRegroupBySew_3_87};
  wire [15:0]       dataInMem_hi_hi_91;
  assign dataInMem_hi_hi_91 = _GEN_477;
  wire [15:0]       dataInMem_hi_lo_93;
  assign dataInMem_hi_lo_93 = _GEN_477;
  wire [23:0]       dataInMem_hi_347 = {dataInMem_hi_hi_91, dataRegroupBySew_2_87};
  wire [15:0]       _GEN_478 = {dataRegroupBySew_4_88, dataRegroupBySew_3_88};
  wire [15:0]       dataInMem_hi_hi_92;
  assign dataInMem_hi_hi_92 = _GEN_478;
  wire [15:0]       dataInMem_hi_lo_94;
  assign dataInMem_hi_lo_94 = _GEN_478;
  wire [23:0]       dataInMem_hi_348 = {dataInMem_hi_hi_92, dataRegroupBySew_2_88};
  wire [15:0]       _GEN_479 = {dataRegroupBySew_4_89, dataRegroupBySew_3_89};
  wire [15:0]       dataInMem_hi_hi_93;
  assign dataInMem_hi_hi_93 = _GEN_479;
  wire [15:0]       dataInMem_hi_lo_95;
  assign dataInMem_hi_lo_95 = _GEN_479;
  wire [23:0]       dataInMem_hi_349 = {dataInMem_hi_hi_93, dataRegroupBySew_2_89};
  wire [15:0]       _GEN_480 = {dataRegroupBySew_4_90, dataRegroupBySew_3_90};
  wire [15:0]       dataInMem_hi_hi_94;
  assign dataInMem_hi_hi_94 = _GEN_480;
  wire [15:0]       dataInMem_hi_lo_96;
  assign dataInMem_hi_lo_96 = _GEN_480;
  wire [23:0]       dataInMem_hi_350 = {dataInMem_hi_hi_94, dataRegroupBySew_2_90};
  wire [15:0]       _GEN_481 = {dataRegroupBySew_4_91, dataRegroupBySew_3_91};
  wire [15:0]       dataInMem_hi_hi_95;
  assign dataInMem_hi_hi_95 = _GEN_481;
  wire [15:0]       dataInMem_hi_lo_97;
  assign dataInMem_hi_lo_97 = _GEN_481;
  wire [23:0]       dataInMem_hi_351 = {dataInMem_hi_hi_95, dataRegroupBySew_2_91};
  wire [15:0]       _GEN_482 = {dataRegroupBySew_4_92, dataRegroupBySew_3_92};
  wire [15:0]       dataInMem_hi_hi_96;
  assign dataInMem_hi_hi_96 = _GEN_482;
  wire [15:0]       dataInMem_hi_lo_98;
  assign dataInMem_hi_lo_98 = _GEN_482;
  wire [23:0]       dataInMem_hi_352 = {dataInMem_hi_hi_96, dataRegroupBySew_2_92};
  wire [15:0]       _GEN_483 = {dataRegroupBySew_4_93, dataRegroupBySew_3_93};
  wire [15:0]       dataInMem_hi_hi_97;
  assign dataInMem_hi_hi_97 = _GEN_483;
  wire [15:0]       dataInMem_hi_lo_99;
  assign dataInMem_hi_lo_99 = _GEN_483;
  wire [23:0]       dataInMem_hi_353 = {dataInMem_hi_hi_97, dataRegroupBySew_2_93};
  wire [15:0]       _GEN_484 = {dataRegroupBySew_4_94, dataRegroupBySew_3_94};
  wire [15:0]       dataInMem_hi_hi_98;
  assign dataInMem_hi_hi_98 = _GEN_484;
  wire [15:0]       dataInMem_hi_lo_100;
  assign dataInMem_hi_lo_100 = _GEN_484;
  wire [23:0]       dataInMem_hi_354 = {dataInMem_hi_hi_98, dataRegroupBySew_2_94};
  wire [15:0]       _GEN_485 = {dataRegroupBySew_4_95, dataRegroupBySew_3_95};
  wire [15:0]       dataInMem_hi_hi_99;
  assign dataInMem_hi_hi_99 = _GEN_485;
  wire [15:0]       dataInMem_hi_lo_101;
  assign dataInMem_hi_lo_101 = _GEN_485;
  wire [23:0]       dataInMem_hi_355 = {dataInMem_hi_hi_99, dataRegroupBySew_2_95};
  wire [15:0]       _GEN_486 = {dataRegroupBySew_4_96, dataRegroupBySew_3_96};
  wire [15:0]       dataInMem_hi_hi_100;
  assign dataInMem_hi_hi_100 = _GEN_486;
  wire [15:0]       dataInMem_hi_lo_102;
  assign dataInMem_hi_lo_102 = _GEN_486;
  wire [23:0]       dataInMem_hi_356 = {dataInMem_hi_hi_100, dataRegroupBySew_2_96};
  wire [15:0]       _GEN_487 = {dataRegroupBySew_4_97, dataRegroupBySew_3_97};
  wire [15:0]       dataInMem_hi_hi_101;
  assign dataInMem_hi_hi_101 = _GEN_487;
  wire [15:0]       dataInMem_hi_lo_103;
  assign dataInMem_hi_lo_103 = _GEN_487;
  wire [23:0]       dataInMem_hi_357 = {dataInMem_hi_hi_101, dataRegroupBySew_2_97};
  wire [15:0]       _GEN_488 = {dataRegroupBySew_4_98, dataRegroupBySew_3_98};
  wire [15:0]       dataInMem_hi_hi_102;
  assign dataInMem_hi_hi_102 = _GEN_488;
  wire [15:0]       dataInMem_hi_lo_104;
  assign dataInMem_hi_lo_104 = _GEN_488;
  wire [23:0]       dataInMem_hi_358 = {dataInMem_hi_hi_102, dataRegroupBySew_2_98};
  wire [15:0]       _GEN_489 = {dataRegroupBySew_4_99, dataRegroupBySew_3_99};
  wire [15:0]       dataInMem_hi_hi_103;
  assign dataInMem_hi_hi_103 = _GEN_489;
  wire [15:0]       dataInMem_hi_lo_105;
  assign dataInMem_hi_lo_105 = _GEN_489;
  wire [23:0]       dataInMem_hi_359 = {dataInMem_hi_hi_103, dataRegroupBySew_2_99};
  wire [15:0]       _GEN_490 = {dataRegroupBySew_4_100, dataRegroupBySew_3_100};
  wire [15:0]       dataInMem_hi_hi_104;
  assign dataInMem_hi_hi_104 = _GEN_490;
  wire [15:0]       dataInMem_hi_lo_106;
  assign dataInMem_hi_lo_106 = _GEN_490;
  wire [23:0]       dataInMem_hi_360 = {dataInMem_hi_hi_104, dataRegroupBySew_2_100};
  wire [15:0]       _GEN_491 = {dataRegroupBySew_4_101, dataRegroupBySew_3_101};
  wire [15:0]       dataInMem_hi_hi_105;
  assign dataInMem_hi_hi_105 = _GEN_491;
  wire [15:0]       dataInMem_hi_lo_107;
  assign dataInMem_hi_lo_107 = _GEN_491;
  wire [23:0]       dataInMem_hi_361 = {dataInMem_hi_hi_105, dataRegroupBySew_2_101};
  wire [15:0]       _GEN_492 = {dataRegroupBySew_4_102, dataRegroupBySew_3_102};
  wire [15:0]       dataInMem_hi_hi_106;
  assign dataInMem_hi_hi_106 = _GEN_492;
  wire [15:0]       dataInMem_hi_lo_108;
  assign dataInMem_hi_lo_108 = _GEN_492;
  wire [23:0]       dataInMem_hi_362 = {dataInMem_hi_hi_106, dataRegroupBySew_2_102};
  wire [15:0]       _GEN_493 = {dataRegroupBySew_4_103, dataRegroupBySew_3_103};
  wire [15:0]       dataInMem_hi_hi_107;
  assign dataInMem_hi_hi_107 = _GEN_493;
  wire [15:0]       dataInMem_hi_lo_109;
  assign dataInMem_hi_lo_109 = _GEN_493;
  wire [23:0]       dataInMem_hi_363 = {dataInMem_hi_hi_107, dataRegroupBySew_2_103};
  wire [15:0]       _GEN_494 = {dataRegroupBySew_4_104, dataRegroupBySew_3_104};
  wire [15:0]       dataInMem_hi_hi_108;
  assign dataInMem_hi_hi_108 = _GEN_494;
  wire [15:0]       dataInMem_hi_lo_110;
  assign dataInMem_hi_lo_110 = _GEN_494;
  wire [23:0]       dataInMem_hi_364 = {dataInMem_hi_hi_108, dataRegroupBySew_2_104};
  wire [15:0]       _GEN_495 = {dataRegroupBySew_4_105, dataRegroupBySew_3_105};
  wire [15:0]       dataInMem_hi_hi_109;
  assign dataInMem_hi_hi_109 = _GEN_495;
  wire [15:0]       dataInMem_hi_lo_111;
  assign dataInMem_hi_lo_111 = _GEN_495;
  wire [23:0]       dataInMem_hi_365 = {dataInMem_hi_hi_109, dataRegroupBySew_2_105};
  wire [15:0]       _GEN_496 = {dataRegroupBySew_4_106, dataRegroupBySew_3_106};
  wire [15:0]       dataInMem_hi_hi_110;
  assign dataInMem_hi_hi_110 = _GEN_496;
  wire [15:0]       dataInMem_hi_lo_112;
  assign dataInMem_hi_lo_112 = _GEN_496;
  wire [23:0]       dataInMem_hi_366 = {dataInMem_hi_hi_110, dataRegroupBySew_2_106};
  wire [15:0]       _GEN_497 = {dataRegroupBySew_4_107, dataRegroupBySew_3_107};
  wire [15:0]       dataInMem_hi_hi_111;
  assign dataInMem_hi_hi_111 = _GEN_497;
  wire [15:0]       dataInMem_hi_lo_113;
  assign dataInMem_hi_lo_113 = _GEN_497;
  wire [23:0]       dataInMem_hi_367 = {dataInMem_hi_hi_111, dataRegroupBySew_2_107};
  wire [15:0]       _GEN_498 = {dataRegroupBySew_4_108, dataRegroupBySew_3_108};
  wire [15:0]       dataInMem_hi_hi_112;
  assign dataInMem_hi_hi_112 = _GEN_498;
  wire [15:0]       dataInMem_hi_lo_114;
  assign dataInMem_hi_lo_114 = _GEN_498;
  wire [23:0]       dataInMem_hi_368 = {dataInMem_hi_hi_112, dataRegroupBySew_2_108};
  wire [15:0]       _GEN_499 = {dataRegroupBySew_4_109, dataRegroupBySew_3_109};
  wire [15:0]       dataInMem_hi_hi_113;
  assign dataInMem_hi_hi_113 = _GEN_499;
  wire [15:0]       dataInMem_hi_lo_115;
  assign dataInMem_hi_lo_115 = _GEN_499;
  wire [23:0]       dataInMem_hi_369 = {dataInMem_hi_hi_113, dataRegroupBySew_2_109};
  wire [15:0]       _GEN_500 = {dataRegroupBySew_4_110, dataRegroupBySew_3_110};
  wire [15:0]       dataInMem_hi_hi_114;
  assign dataInMem_hi_hi_114 = _GEN_500;
  wire [15:0]       dataInMem_hi_lo_116;
  assign dataInMem_hi_lo_116 = _GEN_500;
  wire [23:0]       dataInMem_hi_370 = {dataInMem_hi_hi_114, dataRegroupBySew_2_110};
  wire [15:0]       _GEN_501 = {dataRegroupBySew_4_111, dataRegroupBySew_3_111};
  wire [15:0]       dataInMem_hi_hi_115;
  assign dataInMem_hi_hi_115 = _GEN_501;
  wire [15:0]       dataInMem_hi_lo_117;
  assign dataInMem_hi_lo_117 = _GEN_501;
  wire [23:0]       dataInMem_hi_371 = {dataInMem_hi_hi_115, dataRegroupBySew_2_111};
  wire [15:0]       _GEN_502 = {dataRegroupBySew_4_112, dataRegroupBySew_3_112};
  wire [15:0]       dataInMem_hi_hi_116;
  assign dataInMem_hi_hi_116 = _GEN_502;
  wire [15:0]       dataInMem_hi_lo_118;
  assign dataInMem_hi_lo_118 = _GEN_502;
  wire [23:0]       dataInMem_hi_372 = {dataInMem_hi_hi_116, dataRegroupBySew_2_112};
  wire [15:0]       _GEN_503 = {dataRegroupBySew_4_113, dataRegroupBySew_3_113};
  wire [15:0]       dataInMem_hi_hi_117;
  assign dataInMem_hi_hi_117 = _GEN_503;
  wire [15:0]       dataInMem_hi_lo_119;
  assign dataInMem_hi_lo_119 = _GEN_503;
  wire [23:0]       dataInMem_hi_373 = {dataInMem_hi_hi_117, dataRegroupBySew_2_113};
  wire [15:0]       _GEN_504 = {dataRegroupBySew_4_114, dataRegroupBySew_3_114};
  wire [15:0]       dataInMem_hi_hi_118;
  assign dataInMem_hi_hi_118 = _GEN_504;
  wire [15:0]       dataInMem_hi_lo_120;
  assign dataInMem_hi_lo_120 = _GEN_504;
  wire [23:0]       dataInMem_hi_374 = {dataInMem_hi_hi_118, dataRegroupBySew_2_114};
  wire [15:0]       _GEN_505 = {dataRegroupBySew_4_115, dataRegroupBySew_3_115};
  wire [15:0]       dataInMem_hi_hi_119;
  assign dataInMem_hi_hi_119 = _GEN_505;
  wire [15:0]       dataInMem_hi_lo_121;
  assign dataInMem_hi_lo_121 = _GEN_505;
  wire [23:0]       dataInMem_hi_375 = {dataInMem_hi_hi_119, dataRegroupBySew_2_115};
  wire [15:0]       _GEN_506 = {dataRegroupBySew_4_116, dataRegroupBySew_3_116};
  wire [15:0]       dataInMem_hi_hi_120;
  assign dataInMem_hi_hi_120 = _GEN_506;
  wire [15:0]       dataInMem_hi_lo_122;
  assign dataInMem_hi_lo_122 = _GEN_506;
  wire [23:0]       dataInMem_hi_376 = {dataInMem_hi_hi_120, dataRegroupBySew_2_116};
  wire [15:0]       _GEN_507 = {dataRegroupBySew_4_117, dataRegroupBySew_3_117};
  wire [15:0]       dataInMem_hi_hi_121;
  assign dataInMem_hi_hi_121 = _GEN_507;
  wire [15:0]       dataInMem_hi_lo_123;
  assign dataInMem_hi_lo_123 = _GEN_507;
  wire [23:0]       dataInMem_hi_377 = {dataInMem_hi_hi_121, dataRegroupBySew_2_117};
  wire [15:0]       _GEN_508 = {dataRegroupBySew_4_118, dataRegroupBySew_3_118};
  wire [15:0]       dataInMem_hi_hi_122;
  assign dataInMem_hi_hi_122 = _GEN_508;
  wire [15:0]       dataInMem_hi_lo_124;
  assign dataInMem_hi_lo_124 = _GEN_508;
  wire [23:0]       dataInMem_hi_378 = {dataInMem_hi_hi_122, dataRegroupBySew_2_118};
  wire [15:0]       _GEN_509 = {dataRegroupBySew_4_119, dataRegroupBySew_3_119};
  wire [15:0]       dataInMem_hi_hi_123;
  assign dataInMem_hi_hi_123 = _GEN_509;
  wire [15:0]       dataInMem_hi_lo_125;
  assign dataInMem_hi_lo_125 = _GEN_509;
  wire [23:0]       dataInMem_hi_379 = {dataInMem_hi_hi_123, dataRegroupBySew_2_119};
  wire [15:0]       _GEN_510 = {dataRegroupBySew_4_120, dataRegroupBySew_3_120};
  wire [15:0]       dataInMem_hi_hi_124;
  assign dataInMem_hi_hi_124 = _GEN_510;
  wire [15:0]       dataInMem_hi_lo_126;
  assign dataInMem_hi_lo_126 = _GEN_510;
  wire [23:0]       dataInMem_hi_380 = {dataInMem_hi_hi_124, dataRegroupBySew_2_120};
  wire [15:0]       _GEN_511 = {dataRegroupBySew_4_121, dataRegroupBySew_3_121};
  wire [15:0]       dataInMem_hi_hi_125;
  assign dataInMem_hi_hi_125 = _GEN_511;
  wire [15:0]       dataInMem_hi_lo_127;
  assign dataInMem_hi_lo_127 = _GEN_511;
  wire [23:0]       dataInMem_hi_381 = {dataInMem_hi_hi_125, dataRegroupBySew_2_121};
  wire [15:0]       _GEN_512 = {dataRegroupBySew_4_122, dataRegroupBySew_3_122};
  wire [15:0]       dataInMem_hi_hi_126;
  assign dataInMem_hi_hi_126 = _GEN_512;
  wire [15:0]       dataInMem_hi_lo_128;
  assign dataInMem_hi_lo_128 = _GEN_512;
  wire [23:0]       dataInMem_hi_382 = {dataInMem_hi_hi_126, dataRegroupBySew_2_122};
  wire [15:0]       _GEN_513 = {dataRegroupBySew_4_123, dataRegroupBySew_3_123};
  wire [15:0]       dataInMem_hi_hi_127;
  assign dataInMem_hi_hi_127 = _GEN_513;
  wire [15:0]       dataInMem_hi_lo_129;
  assign dataInMem_hi_lo_129 = _GEN_513;
  wire [23:0]       dataInMem_hi_383 = {dataInMem_hi_hi_127, dataRegroupBySew_2_123};
  wire [15:0]       _GEN_514 = {dataRegroupBySew_4_124, dataRegroupBySew_3_124};
  wire [15:0]       dataInMem_hi_hi_128;
  assign dataInMem_hi_hi_128 = _GEN_514;
  wire [15:0]       dataInMem_hi_lo_130;
  assign dataInMem_hi_lo_130 = _GEN_514;
  wire [23:0]       dataInMem_hi_384 = {dataInMem_hi_hi_128, dataRegroupBySew_2_124};
  wire [15:0]       _GEN_515 = {dataRegroupBySew_4_125, dataRegroupBySew_3_125};
  wire [15:0]       dataInMem_hi_hi_129;
  assign dataInMem_hi_hi_129 = _GEN_515;
  wire [15:0]       dataInMem_hi_lo_131;
  assign dataInMem_hi_lo_131 = _GEN_515;
  wire [23:0]       dataInMem_hi_385 = {dataInMem_hi_hi_129, dataRegroupBySew_2_125};
  wire [15:0]       _GEN_516 = {dataRegroupBySew_4_126, dataRegroupBySew_3_126};
  wire [15:0]       dataInMem_hi_hi_130;
  assign dataInMem_hi_hi_130 = _GEN_516;
  wire [15:0]       dataInMem_hi_lo_132;
  assign dataInMem_hi_lo_132 = _GEN_516;
  wire [23:0]       dataInMem_hi_386 = {dataInMem_hi_hi_130, dataRegroupBySew_2_126};
  wire [15:0]       _GEN_517 = {dataRegroupBySew_4_127, dataRegroupBySew_3_127};
  wire [15:0]       dataInMem_hi_hi_131;
  assign dataInMem_hi_hi_131 = _GEN_517;
  wire [15:0]       dataInMem_hi_lo_133;
  assign dataInMem_hi_lo_133 = _GEN_517;
  wire [23:0]       dataInMem_hi_387 = {dataInMem_hi_hi_131, dataRegroupBySew_2_127};
  wire [79:0]       dataInMem_lo_lo_lo_lo_lo_lo_4 = {dataInMem_hi_261, dataInMem_lo_133, dataInMem_hi_260, dataInMem_lo_132};
  wire [79:0]       dataInMem_lo_lo_lo_lo_lo_hi_4 = {dataInMem_hi_263, dataInMem_lo_135, dataInMem_hi_262, dataInMem_lo_134};
  wire [159:0]      dataInMem_lo_lo_lo_lo_lo_4 = {dataInMem_lo_lo_lo_lo_lo_hi_4, dataInMem_lo_lo_lo_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_lo_lo_lo_hi_lo_4 = {dataInMem_hi_265, dataInMem_lo_137, dataInMem_hi_264, dataInMem_lo_136};
  wire [79:0]       dataInMem_lo_lo_lo_lo_hi_hi_4 = {dataInMem_hi_267, dataInMem_lo_139, dataInMem_hi_266, dataInMem_lo_138};
  wire [159:0]      dataInMem_lo_lo_lo_lo_hi_4 = {dataInMem_lo_lo_lo_lo_hi_hi_4, dataInMem_lo_lo_lo_lo_hi_lo_4};
  wire [319:0]      dataInMem_lo_lo_lo_lo_4 = {dataInMem_lo_lo_lo_lo_hi_4, dataInMem_lo_lo_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_lo_lo_hi_lo_lo_4 = {dataInMem_hi_269, dataInMem_lo_141, dataInMem_hi_268, dataInMem_lo_140};
  wire [79:0]       dataInMem_lo_lo_lo_hi_lo_hi_4 = {dataInMem_hi_271, dataInMem_lo_143, dataInMem_hi_270, dataInMem_lo_142};
  wire [159:0]      dataInMem_lo_lo_lo_hi_lo_4 = {dataInMem_lo_lo_lo_hi_lo_hi_4, dataInMem_lo_lo_lo_hi_lo_lo_4};
  wire [79:0]       dataInMem_lo_lo_lo_hi_hi_lo_4 = {dataInMem_hi_273, dataInMem_lo_145, dataInMem_hi_272, dataInMem_lo_144};
  wire [79:0]       dataInMem_lo_lo_lo_hi_hi_hi_4 = {dataInMem_hi_275, dataInMem_lo_147, dataInMem_hi_274, dataInMem_lo_146};
  wire [159:0]      dataInMem_lo_lo_lo_hi_hi_4 = {dataInMem_lo_lo_lo_hi_hi_hi_4, dataInMem_lo_lo_lo_hi_hi_lo_4};
  wire [319:0]      dataInMem_lo_lo_lo_hi_4 = {dataInMem_lo_lo_lo_hi_hi_4, dataInMem_lo_lo_lo_hi_lo_4};
  wire [639:0]      dataInMem_lo_lo_lo_4 = {dataInMem_lo_lo_lo_hi_4, dataInMem_lo_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_lo_hi_lo_lo_lo_4 = {dataInMem_hi_277, dataInMem_lo_149, dataInMem_hi_276, dataInMem_lo_148};
  wire [79:0]       dataInMem_lo_lo_hi_lo_lo_hi_4 = {dataInMem_hi_279, dataInMem_lo_151, dataInMem_hi_278, dataInMem_lo_150};
  wire [159:0]      dataInMem_lo_lo_hi_lo_lo_4 = {dataInMem_lo_lo_hi_lo_lo_hi_4, dataInMem_lo_lo_hi_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_lo_hi_lo_hi_lo_4 = {dataInMem_hi_281, dataInMem_lo_153, dataInMem_hi_280, dataInMem_lo_152};
  wire [79:0]       dataInMem_lo_lo_hi_lo_hi_hi_4 = {dataInMem_hi_283, dataInMem_lo_155, dataInMem_hi_282, dataInMem_lo_154};
  wire [159:0]      dataInMem_lo_lo_hi_lo_hi_4 = {dataInMem_lo_lo_hi_lo_hi_hi_4, dataInMem_lo_lo_hi_lo_hi_lo_4};
  wire [319:0]      dataInMem_lo_lo_hi_lo_4 = {dataInMem_lo_lo_hi_lo_hi_4, dataInMem_lo_lo_hi_lo_lo_4};
  wire [79:0]       dataInMem_lo_lo_hi_hi_lo_lo_4 = {dataInMem_hi_285, dataInMem_lo_157, dataInMem_hi_284, dataInMem_lo_156};
  wire [79:0]       dataInMem_lo_lo_hi_hi_lo_hi_4 = {dataInMem_hi_287, dataInMem_lo_159, dataInMem_hi_286, dataInMem_lo_158};
  wire [159:0]      dataInMem_lo_lo_hi_hi_lo_4 = {dataInMem_lo_lo_hi_hi_lo_hi_4, dataInMem_lo_lo_hi_hi_lo_lo_4};
  wire [79:0]       dataInMem_lo_lo_hi_hi_hi_lo_4 = {dataInMem_hi_289, dataInMem_lo_161, dataInMem_hi_288, dataInMem_lo_160};
  wire [79:0]       dataInMem_lo_lo_hi_hi_hi_hi_4 = {dataInMem_hi_291, dataInMem_lo_163, dataInMem_hi_290, dataInMem_lo_162};
  wire [159:0]      dataInMem_lo_lo_hi_hi_hi_4 = {dataInMem_lo_lo_hi_hi_hi_hi_4, dataInMem_lo_lo_hi_hi_hi_lo_4};
  wire [319:0]      dataInMem_lo_lo_hi_hi_4 = {dataInMem_lo_lo_hi_hi_hi_4, dataInMem_lo_lo_hi_hi_lo_4};
  wire [639:0]      dataInMem_lo_lo_hi_4 = {dataInMem_lo_lo_hi_hi_4, dataInMem_lo_lo_hi_lo_4};
  wire [1279:0]     dataInMem_lo_lo_4 = {dataInMem_lo_lo_hi_4, dataInMem_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_lo_lo_lo_lo_4 = {dataInMem_hi_293, dataInMem_lo_165, dataInMem_hi_292, dataInMem_lo_164};
  wire [79:0]       dataInMem_lo_hi_lo_lo_lo_hi_4 = {dataInMem_hi_295, dataInMem_lo_167, dataInMem_hi_294, dataInMem_lo_166};
  wire [159:0]      dataInMem_lo_hi_lo_lo_lo_4 = {dataInMem_lo_hi_lo_lo_lo_hi_4, dataInMem_lo_hi_lo_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_lo_lo_hi_lo_4 = {dataInMem_hi_297, dataInMem_lo_169, dataInMem_hi_296, dataInMem_lo_168};
  wire [79:0]       dataInMem_lo_hi_lo_lo_hi_hi_4 = {dataInMem_hi_299, dataInMem_lo_171, dataInMem_hi_298, dataInMem_lo_170};
  wire [159:0]      dataInMem_lo_hi_lo_lo_hi_4 = {dataInMem_lo_hi_lo_lo_hi_hi_4, dataInMem_lo_hi_lo_lo_hi_lo_4};
  wire [319:0]      dataInMem_lo_hi_lo_lo_4 = {dataInMem_lo_hi_lo_lo_hi_4, dataInMem_lo_hi_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_lo_hi_lo_lo_4 = {dataInMem_hi_301, dataInMem_lo_173, dataInMem_hi_300, dataInMem_lo_172};
  wire [79:0]       dataInMem_lo_hi_lo_hi_lo_hi_4 = {dataInMem_hi_303, dataInMem_lo_175, dataInMem_hi_302, dataInMem_lo_174};
  wire [159:0]      dataInMem_lo_hi_lo_hi_lo_4 = {dataInMem_lo_hi_lo_hi_lo_hi_4, dataInMem_lo_hi_lo_hi_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_lo_hi_hi_lo_4 = {dataInMem_hi_305, dataInMem_lo_177, dataInMem_hi_304, dataInMem_lo_176};
  wire [79:0]       dataInMem_lo_hi_lo_hi_hi_hi_4 = {dataInMem_hi_307, dataInMem_lo_179, dataInMem_hi_306, dataInMem_lo_178};
  wire [159:0]      dataInMem_lo_hi_lo_hi_hi_4 = {dataInMem_lo_hi_lo_hi_hi_hi_4, dataInMem_lo_hi_lo_hi_hi_lo_4};
  wire [319:0]      dataInMem_lo_hi_lo_hi_4 = {dataInMem_lo_hi_lo_hi_hi_4, dataInMem_lo_hi_lo_hi_lo_4};
  wire [639:0]      dataInMem_lo_hi_lo_4 = {dataInMem_lo_hi_lo_hi_4, dataInMem_lo_hi_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_hi_lo_lo_lo_4 = {dataInMem_hi_309, dataInMem_lo_181, dataInMem_hi_308, dataInMem_lo_180};
  wire [79:0]       dataInMem_lo_hi_hi_lo_lo_hi_4 = {dataInMem_hi_311, dataInMem_lo_183, dataInMem_hi_310, dataInMem_lo_182};
  wire [159:0]      dataInMem_lo_hi_hi_lo_lo_4 = {dataInMem_lo_hi_hi_lo_lo_hi_4, dataInMem_lo_hi_hi_lo_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_hi_lo_hi_lo_4 = {dataInMem_hi_313, dataInMem_lo_185, dataInMem_hi_312, dataInMem_lo_184};
  wire [79:0]       dataInMem_lo_hi_hi_lo_hi_hi_4 = {dataInMem_hi_315, dataInMem_lo_187, dataInMem_hi_314, dataInMem_lo_186};
  wire [159:0]      dataInMem_lo_hi_hi_lo_hi_4 = {dataInMem_lo_hi_hi_lo_hi_hi_4, dataInMem_lo_hi_hi_lo_hi_lo_4};
  wire [319:0]      dataInMem_lo_hi_hi_lo_4 = {dataInMem_lo_hi_hi_lo_hi_4, dataInMem_lo_hi_hi_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_hi_hi_lo_lo_4 = {dataInMem_hi_317, dataInMem_lo_189, dataInMem_hi_316, dataInMem_lo_188};
  wire [79:0]       dataInMem_lo_hi_hi_hi_lo_hi_4 = {dataInMem_hi_319, dataInMem_lo_191, dataInMem_hi_318, dataInMem_lo_190};
  wire [159:0]      dataInMem_lo_hi_hi_hi_lo_4 = {dataInMem_lo_hi_hi_hi_lo_hi_4, dataInMem_lo_hi_hi_hi_lo_lo_4};
  wire [79:0]       dataInMem_lo_hi_hi_hi_hi_lo_4 = {dataInMem_hi_321, dataInMem_lo_193, dataInMem_hi_320, dataInMem_lo_192};
  wire [79:0]       dataInMem_lo_hi_hi_hi_hi_hi_4 = {dataInMem_hi_323, dataInMem_lo_195, dataInMem_hi_322, dataInMem_lo_194};
  wire [159:0]      dataInMem_lo_hi_hi_hi_hi_4 = {dataInMem_lo_hi_hi_hi_hi_hi_4, dataInMem_lo_hi_hi_hi_hi_lo_4};
  wire [319:0]      dataInMem_lo_hi_hi_hi_4 = {dataInMem_lo_hi_hi_hi_hi_4, dataInMem_lo_hi_hi_hi_lo_4};
  wire [639:0]      dataInMem_lo_hi_hi_4 = {dataInMem_lo_hi_hi_hi_4, dataInMem_lo_hi_hi_lo_4};
  wire [1279:0]     dataInMem_lo_hi_4 = {dataInMem_lo_hi_hi_4, dataInMem_lo_hi_lo_4};
  wire [2559:0]     dataInMem_lo_260 = {dataInMem_lo_hi_4, dataInMem_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_lo_lo_lo_lo_4 = {dataInMem_hi_325, dataInMem_lo_197, dataInMem_hi_324, dataInMem_lo_196};
  wire [79:0]       dataInMem_hi_lo_lo_lo_lo_hi_4 = {dataInMem_hi_327, dataInMem_lo_199, dataInMem_hi_326, dataInMem_lo_198};
  wire [159:0]      dataInMem_hi_lo_lo_lo_lo_4 = {dataInMem_hi_lo_lo_lo_lo_hi_4, dataInMem_hi_lo_lo_lo_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_lo_lo_hi_lo_4 = {dataInMem_hi_329, dataInMem_lo_201, dataInMem_hi_328, dataInMem_lo_200};
  wire [79:0]       dataInMem_hi_lo_lo_lo_hi_hi_4 = {dataInMem_hi_331, dataInMem_lo_203, dataInMem_hi_330, dataInMem_lo_202};
  wire [159:0]      dataInMem_hi_lo_lo_lo_hi_4 = {dataInMem_hi_lo_lo_lo_hi_hi_4, dataInMem_hi_lo_lo_lo_hi_lo_4};
  wire [319:0]      dataInMem_hi_lo_lo_lo_4 = {dataInMem_hi_lo_lo_lo_hi_4, dataInMem_hi_lo_lo_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_lo_hi_lo_lo_4 = {dataInMem_hi_333, dataInMem_lo_205, dataInMem_hi_332, dataInMem_lo_204};
  wire [79:0]       dataInMem_hi_lo_lo_hi_lo_hi_4 = {dataInMem_hi_335, dataInMem_lo_207, dataInMem_hi_334, dataInMem_lo_206};
  wire [159:0]      dataInMem_hi_lo_lo_hi_lo_4 = {dataInMem_hi_lo_lo_hi_lo_hi_4, dataInMem_hi_lo_lo_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_lo_hi_hi_lo_4 = {dataInMem_hi_337, dataInMem_lo_209, dataInMem_hi_336, dataInMem_lo_208};
  wire [79:0]       dataInMem_hi_lo_lo_hi_hi_hi_4 = {dataInMem_hi_339, dataInMem_lo_211, dataInMem_hi_338, dataInMem_lo_210};
  wire [159:0]      dataInMem_hi_lo_lo_hi_hi_4 = {dataInMem_hi_lo_lo_hi_hi_hi_4, dataInMem_hi_lo_lo_hi_hi_lo_4};
  wire [319:0]      dataInMem_hi_lo_lo_hi_4 = {dataInMem_hi_lo_lo_hi_hi_4, dataInMem_hi_lo_lo_hi_lo_4};
  wire [639:0]      dataInMem_hi_lo_lo_4 = {dataInMem_hi_lo_lo_hi_4, dataInMem_hi_lo_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_hi_lo_lo_lo_4 = {dataInMem_hi_341, dataInMem_lo_213, dataInMem_hi_340, dataInMem_lo_212};
  wire [79:0]       dataInMem_hi_lo_hi_lo_lo_hi_4 = {dataInMem_hi_343, dataInMem_lo_215, dataInMem_hi_342, dataInMem_lo_214};
  wire [159:0]      dataInMem_hi_lo_hi_lo_lo_4 = {dataInMem_hi_lo_hi_lo_lo_hi_4, dataInMem_hi_lo_hi_lo_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_hi_lo_hi_lo_4 = {dataInMem_hi_345, dataInMem_lo_217, dataInMem_hi_344, dataInMem_lo_216};
  wire [79:0]       dataInMem_hi_lo_hi_lo_hi_hi_4 = {dataInMem_hi_347, dataInMem_lo_219, dataInMem_hi_346, dataInMem_lo_218};
  wire [159:0]      dataInMem_hi_lo_hi_lo_hi_4 = {dataInMem_hi_lo_hi_lo_hi_hi_4, dataInMem_hi_lo_hi_lo_hi_lo_4};
  wire [319:0]      dataInMem_hi_lo_hi_lo_4 = {dataInMem_hi_lo_hi_lo_hi_4, dataInMem_hi_lo_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_hi_hi_lo_lo_4 = {dataInMem_hi_349, dataInMem_lo_221, dataInMem_hi_348, dataInMem_lo_220};
  wire [79:0]       dataInMem_hi_lo_hi_hi_lo_hi_4 = {dataInMem_hi_351, dataInMem_lo_223, dataInMem_hi_350, dataInMem_lo_222};
  wire [159:0]      dataInMem_hi_lo_hi_hi_lo_4 = {dataInMem_hi_lo_hi_hi_lo_hi_4, dataInMem_hi_lo_hi_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_lo_hi_hi_hi_lo_4 = {dataInMem_hi_353, dataInMem_lo_225, dataInMem_hi_352, dataInMem_lo_224};
  wire [79:0]       dataInMem_hi_lo_hi_hi_hi_hi_4 = {dataInMem_hi_355, dataInMem_lo_227, dataInMem_hi_354, dataInMem_lo_226};
  wire [159:0]      dataInMem_hi_lo_hi_hi_hi_4 = {dataInMem_hi_lo_hi_hi_hi_hi_4, dataInMem_hi_lo_hi_hi_hi_lo_4};
  wire [319:0]      dataInMem_hi_lo_hi_hi_4 = {dataInMem_hi_lo_hi_hi_hi_4, dataInMem_hi_lo_hi_hi_lo_4};
  wire [639:0]      dataInMem_hi_lo_hi_4 = {dataInMem_hi_lo_hi_hi_4, dataInMem_hi_lo_hi_lo_4};
  wire [1279:0]     dataInMem_hi_lo_4 = {dataInMem_hi_lo_hi_4, dataInMem_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_lo_lo_lo_lo_4 = {dataInMem_hi_357, dataInMem_lo_229, dataInMem_hi_356, dataInMem_lo_228};
  wire [79:0]       dataInMem_hi_hi_lo_lo_lo_hi_4 = {dataInMem_hi_359, dataInMem_lo_231, dataInMem_hi_358, dataInMem_lo_230};
  wire [159:0]      dataInMem_hi_hi_lo_lo_lo_4 = {dataInMem_hi_hi_lo_lo_lo_hi_4, dataInMem_hi_hi_lo_lo_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_lo_lo_hi_lo_4 = {dataInMem_hi_361, dataInMem_lo_233, dataInMem_hi_360, dataInMem_lo_232};
  wire [79:0]       dataInMem_hi_hi_lo_lo_hi_hi_4 = {dataInMem_hi_363, dataInMem_lo_235, dataInMem_hi_362, dataInMem_lo_234};
  wire [159:0]      dataInMem_hi_hi_lo_lo_hi_4 = {dataInMem_hi_hi_lo_lo_hi_hi_4, dataInMem_hi_hi_lo_lo_hi_lo_4};
  wire [319:0]      dataInMem_hi_hi_lo_lo_4 = {dataInMem_hi_hi_lo_lo_hi_4, dataInMem_hi_hi_lo_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_lo_hi_lo_lo_4 = {dataInMem_hi_365, dataInMem_lo_237, dataInMem_hi_364, dataInMem_lo_236};
  wire [79:0]       dataInMem_hi_hi_lo_hi_lo_hi_4 = {dataInMem_hi_367, dataInMem_lo_239, dataInMem_hi_366, dataInMem_lo_238};
  wire [159:0]      dataInMem_hi_hi_lo_hi_lo_4 = {dataInMem_hi_hi_lo_hi_lo_hi_4, dataInMem_hi_hi_lo_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_lo_hi_hi_lo_4 = {dataInMem_hi_369, dataInMem_lo_241, dataInMem_hi_368, dataInMem_lo_240};
  wire [79:0]       dataInMem_hi_hi_lo_hi_hi_hi_4 = {dataInMem_hi_371, dataInMem_lo_243, dataInMem_hi_370, dataInMem_lo_242};
  wire [159:0]      dataInMem_hi_hi_lo_hi_hi_4 = {dataInMem_hi_hi_lo_hi_hi_hi_4, dataInMem_hi_hi_lo_hi_hi_lo_4};
  wire [319:0]      dataInMem_hi_hi_lo_hi_4 = {dataInMem_hi_hi_lo_hi_hi_4, dataInMem_hi_hi_lo_hi_lo_4};
  wire [639:0]      dataInMem_hi_hi_lo_4 = {dataInMem_hi_hi_lo_hi_4, dataInMem_hi_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_hi_lo_lo_lo_4 = {dataInMem_hi_373, dataInMem_lo_245, dataInMem_hi_372, dataInMem_lo_244};
  wire [79:0]       dataInMem_hi_hi_hi_lo_lo_hi_4 = {dataInMem_hi_375, dataInMem_lo_247, dataInMem_hi_374, dataInMem_lo_246};
  wire [159:0]      dataInMem_hi_hi_hi_lo_lo_4 = {dataInMem_hi_hi_hi_lo_lo_hi_4, dataInMem_hi_hi_hi_lo_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_hi_lo_hi_lo_4 = {dataInMem_hi_377, dataInMem_lo_249, dataInMem_hi_376, dataInMem_lo_248};
  wire [79:0]       dataInMem_hi_hi_hi_lo_hi_hi_4 = {dataInMem_hi_379, dataInMem_lo_251, dataInMem_hi_378, dataInMem_lo_250};
  wire [159:0]      dataInMem_hi_hi_hi_lo_hi_4 = {dataInMem_hi_hi_hi_lo_hi_hi_4, dataInMem_hi_hi_hi_lo_hi_lo_4};
  wire [319:0]      dataInMem_hi_hi_hi_lo_4 = {dataInMem_hi_hi_hi_lo_hi_4, dataInMem_hi_hi_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_hi_hi_lo_lo_4 = {dataInMem_hi_381, dataInMem_lo_253, dataInMem_hi_380, dataInMem_lo_252};
  wire [79:0]       dataInMem_hi_hi_hi_hi_lo_hi_4 = {dataInMem_hi_383, dataInMem_lo_255, dataInMem_hi_382, dataInMem_lo_254};
  wire [159:0]      dataInMem_hi_hi_hi_hi_lo_4 = {dataInMem_hi_hi_hi_hi_lo_hi_4, dataInMem_hi_hi_hi_hi_lo_lo_4};
  wire [79:0]       dataInMem_hi_hi_hi_hi_hi_lo_4 = {dataInMem_hi_385, dataInMem_lo_257, dataInMem_hi_384, dataInMem_lo_256};
  wire [79:0]       dataInMem_hi_hi_hi_hi_hi_hi_4 = {dataInMem_hi_387, dataInMem_lo_259, dataInMem_hi_386, dataInMem_lo_258};
  wire [159:0]      dataInMem_hi_hi_hi_hi_hi_4 = {dataInMem_hi_hi_hi_hi_hi_hi_4, dataInMem_hi_hi_hi_hi_hi_lo_4};
  wire [319:0]      dataInMem_hi_hi_hi_hi_4 = {dataInMem_hi_hi_hi_hi_hi_4, dataInMem_hi_hi_hi_hi_lo_4};
  wire [639:0]      dataInMem_hi_hi_hi_4 = {dataInMem_hi_hi_hi_hi_4, dataInMem_hi_hi_hi_lo_4};
  wire [1279:0]     dataInMem_hi_hi_132 = {dataInMem_hi_hi_hi_4, dataInMem_hi_hi_lo_4};
  wire [2559:0]     dataInMem_hi_388 = {dataInMem_hi_hi_132, dataInMem_hi_lo_4};
  wire [5119:0]     dataInMem_4 = {dataInMem_hi_388, dataInMem_lo_260};
  wire [1023:0]     regroupCacheLine_4_0 = dataInMem_4[1023:0];
  wire [1023:0]     regroupCacheLine_4_1 = dataInMem_4[2047:1024];
  wire [1023:0]     regroupCacheLine_4_2 = dataInMem_4[3071:2048];
  wire [1023:0]     regroupCacheLine_4_3 = dataInMem_4[4095:3072];
  wire [1023:0]     regroupCacheLine_4_4 = dataInMem_4[5119:4096];
  wire [1023:0]     res_32 = regroupCacheLine_4_0;
  wire [1023:0]     res_33 = regroupCacheLine_4_1;
  wire [1023:0]     res_34 = regroupCacheLine_4_2;
  wire [1023:0]     res_35 = regroupCacheLine_4_3;
  wire [1023:0]     res_36 = regroupCacheLine_4_4;
  wire [2047:0]     lo_lo_4 = {res_33, res_32};
  wire [2047:0]     lo_hi_4 = {res_35, res_34};
  wire [4095:0]     lo_4 = {lo_hi_4, lo_lo_4};
  wire [2047:0]     hi_lo_4 = {1024'h0, res_36};
  wire [4095:0]     hi_4 = {2048'h0, hi_lo_4};
  wire [8191:0]     regroupLoadData_0_4 = {hi_4, lo_4};
  wire [23:0]       dataInMem_lo_261 = {dataInMem_lo_hi_5, dataRegroupBySew_0_0};
  wire [15:0]       _GEN_518 = {dataRegroupBySew_5_0, dataRegroupBySew_4_0};
  wire [15:0]       dataInMem_hi_hi_133;
  assign dataInMem_hi_hi_133 = _GEN_518;
  wire [15:0]       dataInMem_hi_lo_135;
  assign dataInMem_hi_lo_135 = _GEN_518;
  wire [23:0]       dataInMem_hi_389 = {dataInMem_hi_hi_133, dataRegroupBySew_3_0};
  wire [23:0]       dataInMem_lo_262 = {dataInMem_lo_hi_6, dataRegroupBySew_0_1};
  wire [15:0]       _GEN_519 = {dataRegroupBySew_5_1, dataRegroupBySew_4_1};
  wire [15:0]       dataInMem_hi_hi_134;
  assign dataInMem_hi_hi_134 = _GEN_519;
  wire [15:0]       dataInMem_hi_lo_136;
  assign dataInMem_hi_lo_136 = _GEN_519;
  wire [23:0]       dataInMem_hi_390 = {dataInMem_hi_hi_134, dataRegroupBySew_3_1};
  wire [23:0]       dataInMem_lo_263 = {dataInMem_lo_hi_7, dataRegroupBySew_0_2};
  wire [15:0]       _GEN_520 = {dataRegroupBySew_5_2, dataRegroupBySew_4_2};
  wire [15:0]       dataInMem_hi_hi_135;
  assign dataInMem_hi_hi_135 = _GEN_520;
  wire [15:0]       dataInMem_hi_lo_137;
  assign dataInMem_hi_lo_137 = _GEN_520;
  wire [23:0]       dataInMem_hi_391 = {dataInMem_hi_hi_135, dataRegroupBySew_3_2};
  wire [23:0]       dataInMem_lo_264 = {dataInMem_lo_hi_8, dataRegroupBySew_0_3};
  wire [15:0]       _GEN_521 = {dataRegroupBySew_5_3, dataRegroupBySew_4_3};
  wire [15:0]       dataInMem_hi_hi_136;
  assign dataInMem_hi_hi_136 = _GEN_521;
  wire [15:0]       dataInMem_hi_lo_138;
  assign dataInMem_hi_lo_138 = _GEN_521;
  wire [23:0]       dataInMem_hi_392 = {dataInMem_hi_hi_136, dataRegroupBySew_3_3};
  wire [23:0]       dataInMem_lo_265 = {dataInMem_lo_hi_9, dataRegroupBySew_0_4};
  wire [15:0]       _GEN_522 = {dataRegroupBySew_5_4, dataRegroupBySew_4_4};
  wire [15:0]       dataInMem_hi_hi_137;
  assign dataInMem_hi_hi_137 = _GEN_522;
  wire [15:0]       dataInMem_hi_lo_139;
  assign dataInMem_hi_lo_139 = _GEN_522;
  wire [23:0]       dataInMem_hi_393 = {dataInMem_hi_hi_137, dataRegroupBySew_3_4};
  wire [23:0]       dataInMem_lo_266 = {dataInMem_lo_hi_10, dataRegroupBySew_0_5};
  wire [15:0]       _GEN_523 = {dataRegroupBySew_5_5, dataRegroupBySew_4_5};
  wire [15:0]       dataInMem_hi_hi_138;
  assign dataInMem_hi_hi_138 = _GEN_523;
  wire [15:0]       dataInMem_hi_lo_140;
  assign dataInMem_hi_lo_140 = _GEN_523;
  wire [23:0]       dataInMem_hi_394 = {dataInMem_hi_hi_138, dataRegroupBySew_3_5};
  wire [23:0]       dataInMem_lo_267 = {dataInMem_lo_hi_11, dataRegroupBySew_0_6};
  wire [15:0]       _GEN_524 = {dataRegroupBySew_5_6, dataRegroupBySew_4_6};
  wire [15:0]       dataInMem_hi_hi_139;
  assign dataInMem_hi_hi_139 = _GEN_524;
  wire [15:0]       dataInMem_hi_lo_141;
  assign dataInMem_hi_lo_141 = _GEN_524;
  wire [23:0]       dataInMem_hi_395 = {dataInMem_hi_hi_139, dataRegroupBySew_3_6};
  wire [23:0]       dataInMem_lo_268 = {dataInMem_lo_hi_12, dataRegroupBySew_0_7};
  wire [15:0]       _GEN_525 = {dataRegroupBySew_5_7, dataRegroupBySew_4_7};
  wire [15:0]       dataInMem_hi_hi_140;
  assign dataInMem_hi_hi_140 = _GEN_525;
  wire [15:0]       dataInMem_hi_lo_142;
  assign dataInMem_hi_lo_142 = _GEN_525;
  wire [23:0]       dataInMem_hi_396 = {dataInMem_hi_hi_140, dataRegroupBySew_3_7};
  wire [23:0]       dataInMem_lo_269 = {dataInMem_lo_hi_13, dataRegroupBySew_0_8};
  wire [15:0]       _GEN_526 = {dataRegroupBySew_5_8, dataRegroupBySew_4_8};
  wire [15:0]       dataInMem_hi_hi_141;
  assign dataInMem_hi_hi_141 = _GEN_526;
  wire [15:0]       dataInMem_hi_lo_143;
  assign dataInMem_hi_lo_143 = _GEN_526;
  wire [23:0]       dataInMem_hi_397 = {dataInMem_hi_hi_141, dataRegroupBySew_3_8};
  wire [23:0]       dataInMem_lo_270 = {dataInMem_lo_hi_14, dataRegroupBySew_0_9};
  wire [15:0]       _GEN_527 = {dataRegroupBySew_5_9, dataRegroupBySew_4_9};
  wire [15:0]       dataInMem_hi_hi_142;
  assign dataInMem_hi_hi_142 = _GEN_527;
  wire [15:0]       dataInMem_hi_lo_144;
  assign dataInMem_hi_lo_144 = _GEN_527;
  wire [23:0]       dataInMem_hi_398 = {dataInMem_hi_hi_142, dataRegroupBySew_3_9};
  wire [23:0]       dataInMem_lo_271 = {dataInMem_lo_hi_15, dataRegroupBySew_0_10};
  wire [15:0]       _GEN_528 = {dataRegroupBySew_5_10, dataRegroupBySew_4_10};
  wire [15:0]       dataInMem_hi_hi_143;
  assign dataInMem_hi_hi_143 = _GEN_528;
  wire [15:0]       dataInMem_hi_lo_145;
  assign dataInMem_hi_lo_145 = _GEN_528;
  wire [23:0]       dataInMem_hi_399 = {dataInMem_hi_hi_143, dataRegroupBySew_3_10};
  wire [23:0]       dataInMem_lo_272 = {dataInMem_lo_hi_16, dataRegroupBySew_0_11};
  wire [15:0]       _GEN_529 = {dataRegroupBySew_5_11, dataRegroupBySew_4_11};
  wire [15:0]       dataInMem_hi_hi_144;
  assign dataInMem_hi_hi_144 = _GEN_529;
  wire [15:0]       dataInMem_hi_lo_146;
  assign dataInMem_hi_lo_146 = _GEN_529;
  wire [23:0]       dataInMem_hi_400 = {dataInMem_hi_hi_144, dataRegroupBySew_3_11};
  wire [23:0]       dataInMem_lo_273 = {dataInMem_lo_hi_17, dataRegroupBySew_0_12};
  wire [15:0]       _GEN_530 = {dataRegroupBySew_5_12, dataRegroupBySew_4_12};
  wire [15:0]       dataInMem_hi_hi_145;
  assign dataInMem_hi_hi_145 = _GEN_530;
  wire [15:0]       dataInMem_hi_lo_147;
  assign dataInMem_hi_lo_147 = _GEN_530;
  wire [23:0]       dataInMem_hi_401 = {dataInMem_hi_hi_145, dataRegroupBySew_3_12};
  wire [23:0]       dataInMem_lo_274 = {dataInMem_lo_hi_18, dataRegroupBySew_0_13};
  wire [15:0]       _GEN_531 = {dataRegroupBySew_5_13, dataRegroupBySew_4_13};
  wire [15:0]       dataInMem_hi_hi_146;
  assign dataInMem_hi_hi_146 = _GEN_531;
  wire [15:0]       dataInMem_hi_lo_148;
  assign dataInMem_hi_lo_148 = _GEN_531;
  wire [23:0]       dataInMem_hi_402 = {dataInMem_hi_hi_146, dataRegroupBySew_3_13};
  wire [23:0]       dataInMem_lo_275 = {dataInMem_lo_hi_19, dataRegroupBySew_0_14};
  wire [15:0]       _GEN_532 = {dataRegroupBySew_5_14, dataRegroupBySew_4_14};
  wire [15:0]       dataInMem_hi_hi_147;
  assign dataInMem_hi_hi_147 = _GEN_532;
  wire [15:0]       dataInMem_hi_lo_149;
  assign dataInMem_hi_lo_149 = _GEN_532;
  wire [23:0]       dataInMem_hi_403 = {dataInMem_hi_hi_147, dataRegroupBySew_3_14};
  wire [23:0]       dataInMem_lo_276 = {dataInMem_lo_hi_20, dataRegroupBySew_0_15};
  wire [15:0]       _GEN_533 = {dataRegroupBySew_5_15, dataRegroupBySew_4_15};
  wire [15:0]       dataInMem_hi_hi_148;
  assign dataInMem_hi_hi_148 = _GEN_533;
  wire [15:0]       dataInMem_hi_lo_150;
  assign dataInMem_hi_lo_150 = _GEN_533;
  wire [23:0]       dataInMem_hi_404 = {dataInMem_hi_hi_148, dataRegroupBySew_3_15};
  wire [23:0]       dataInMem_lo_277 = {dataInMem_lo_hi_21, dataRegroupBySew_0_16};
  wire [15:0]       _GEN_534 = {dataRegroupBySew_5_16, dataRegroupBySew_4_16};
  wire [15:0]       dataInMem_hi_hi_149;
  assign dataInMem_hi_hi_149 = _GEN_534;
  wire [15:0]       dataInMem_hi_lo_151;
  assign dataInMem_hi_lo_151 = _GEN_534;
  wire [23:0]       dataInMem_hi_405 = {dataInMem_hi_hi_149, dataRegroupBySew_3_16};
  wire [23:0]       dataInMem_lo_278 = {dataInMem_lo_hi_22, dataRegroupBySew_0_17};
  wire [15:0]       _GEN_535 = {dataRegroupBySew_5_17, dataRegroupBySew_4_17};
  wire [15:0]       dataInMem_hi_hi_150;
  assign dataInMem_hi_hi_150 = _GEN_535;
  wire [15:0]       dataInMem_hi_lo_152;
  assign dataInMem_hi_lo_152 = _GEN_535;
  wire [23:0]       dataInMem_hi_406 = {dataInMem_hi_hi_150, dataRegroupBySew_3_17};
  wire [23:0]       dataInMem_lo_279 = {dataInMem_lo_hi_23, dataRegroupBySew_0_18};
  wire [15:0]       _GEN_536 = {dataRegroupBySew_5_18, dataRegroupBySew_4_18};
  wire [15:0]       dataInMem_hi_hi_151;
  assign dataInMem_hi_hi_151 = _GEN_536;
  wire [15:0]       dataInMem_hi_lo_153;
  assign dataInMem_hi_lo_153 = _GEN_536;
  wire [23:0]       dataInMem_hi_407 = {dataInMem_hi_hi_151, dataRegroupBySew_3_18};
  wire [23:0]       dataInMem_lo_280 = {dataInMem_lo_hi_24, dataRegroupBySew_0_19};
  wire [15:0]       _GEN_537 = {dataRegroupBySew_5_19, dataRegroupBySew_4_19};
  wire [15:0]       dataInMem_hi_hi_152;
  assign dataInMem_hi_hi_152 = _GEN_537;
  wire [15:0]       dataInMem_hi_lo_154;
  assign dataInMem_hi_lo_154 = _GEN_537;
  wire [23:0]       dataInMem_hi_408 = {dataInMem_hi_hi_152, dataRegroupBySew_3_19};
  wire [23:0]       dataInMem_lo_281 = {dataInMem_lo_hi_25, dataRegroupBySew_0_20};
  wire [15:0]       _GEN_538 = {dataRegroupBySew_5_20, dataRegroupBySew_4_20};
  wire [15:0]       dataInMem_hi_hi_153;
  assign dataInMem_hi_hi_153 = _GEN_538;
  wire [15:0]       dataInMem_hi_lo_155;
  assign dataInMem_hi_lo_155 = _GEN_538;
  wire [23:0]       dataInMem_hi_409 = {dataInMem_hi_hi_153, dataRegroupBySew_3_20};
  wire [23:0]       dataInMem_lo_282 = {dataInMem_lo_hi_26, dataRegroupBySew_0_21};
  wire [15:0]       _GEN_539 = {dataRegroupBySew_5_21, dataRegroupBySew_4_21};
  wire [15:0]       dataInMem_hi_hi_154;
  assign dataInMem_hi_hi_154 = _GEN_539;
  wire [15:0]       dataInMem_hi_lo_156;
  assign dataInMem_hi_lo_156 = _GEN_539;
  wire [23:0]       dataInMem_hi_410 = {dataInMem_hi_hi_154, dataRegroupBySew_3_21};
  wire [23:0]       dataInMem_lo_283 = {dataInMem_lo_hi_27, dataRegroupBySew_0_22};
  wire [15:0]       _GEN_540 = {dataRegroupBySew_5_22, dataRegroupBySew_4_22};
  wire [15:0]       dataInMem_hi_hi_155;
  assign dataInMem_hi_hi_155 = _GEN_540;
  wire [15:0]       dataInMem_hi_lo_157;
  assign dataInMem_hi_lo_157 = _GEN_540;
  wire [23:0]       dataInMem_hi_411 = {dataInMem_hi_hi_155, dataRegroupBySew_3_22};
  wire [23:0]       dataInMem_lo_284 = {dataInMem_lo_hi_28, dataRegroupBySew_0_23};
  wire [15:0]       _GEN_541 = {dataRegroupBySew_5_23, dataRegroupBySew_4_23};
  wire [15:0]       dataInMem_hi_hi_156;
  assign dataInMem_hi_hi_156 = _GEN_541;
  wire [15:0]       dataInMem_hi_lo_158;
  assign dataInMem_hi_lo_158 = _GEN_541;
  wire [23:0]       dataInMem_hi_412 = {dataInMem_hi_hi_156, dataRegroupBySew_3_23};
  wire [23:0]       dataInMem_lo_285 = {dataInMem_lo_hi_29, dataRegroupBySew_0_24};
  wire [15:0]       _GEN_542 = {dataRegroupBySew_5_24, dataRegroupBySew_4_24};
  wire [15:0]       dataInMem_hi_hi_157;
  assign dataInMem_hi_hi_157 = _GEN_542;
  wire [15:0]       dataInMem_hi_lo_159;
  assign dataInMem_hi_lo_159 = _GEN_542;
  wire [23:0]       dataInMem_hi_413 = {dataInMem_hi_hi_157, dataRegroupBySew_3_24};
  wire [23:0]       dataInMem_lo_286 = {dataInMem_lo_hi_30, dataRegroupBySew_0_25};
  wire [15:0]       _GEN_543 = {dataRegroupBySew_5_25, dataRegroupBySew_4_25};
  wire [15:0]       dataInMem_hi_hi_158;
  assign dataInMem_hi_hi_158 = _GEN_543;
  wire [15:0]       dataInMem_hi_lo_160;
  assign dataInMem_hi_lo_160 = _GEN_543;
  wire [23:0]       dataInMem_hi_414 = {dataInMem_hi_hi_158, dataRegroupBySew_3_25};
  wire [23:0]       dataInMem_lo_287 = {dataInMem_lo_hi_31, dataRegroupBySew_0_26};
  wire [15:0]       _GEN_544 = {dataRegroupBySew_5_26, dataRegroupBySew_4_26};
  wire [15:0]       dataInMem_hi_hi_159;
  assign dataInMem_hi_hi_159 = _GEN_544;
  wire [15:0]       dataInMem_hi_lo_161;
  assign dataInMem_hi_lo_161 = _GEN_544;
  wire [23:0]       dataInMem_hi_415 = {dataInMem_hi_hi_159, dataRegroupBySew_3_26};
  wire [23:0]       dataInMem_lo_288 = {dataInMem_lo_hi_32, dataRegroupBySew_0_27};
  wire [15:0]       _GEN_545 = {dataRegroupBySew_5_27, dataRegroupBySew_4_27};
  wire [15:0]       dataInMem_hi_hi_160;
  assign dataInMem_hi_hi_160 = _GEN_545;
  wire [15:0]       dataInMem_hi_lo_162;
  assign dataInMem_hi_lo_162 = _GEN_545;
  wire [23:0]       dataInMem_hi_416 = {dataInMem_hi_hi_160, dataRegroupBySew_3_27};
  wire [23:0]       dataInMem_lo_289 = {dataInMem_lo_hi_33, dataRegroupBySew_0_28};
  wire [15:0]       _GEN_546 = {dataRegroupBySew_5_28, dataRegroupBySew_4_28};
  wire [15:0]       dataInMem_hi_hi_161;
  assign dataInMem_hi_hi_161 = _GEN_546;
  wire [15:0]       dataInMem_hi_lo_163;
  assign dataInMem_hi_lo_163 = _GEN_546;
  wire [23:0]       dataInMem_hi_417 = {dataInMem_hi_hi_161, dataRegroupBySew_3_28};
  wire [23:0]       dataInMem_lo_290 = {dataInMem_lo_hi_34, dataRegroupBySew_0_29};
  wire [15:0]       _GEN_547 = {dataRegroupBySew_5_29, dataRegroupBySew_4_29};
  wire [15:0]       dataInMem_hi_hi_162;
  assign dataInMem_hi_hi_162 = _GEN_547;
  wire [15:0]       dataInMem_hi_lo_164;
  assign dataInMem_hi_lo_164 = _GEN_547;
  wire [23:0]       dataInMem_hi_418 = {dataInMem_hi_hi_162, dataRegroupBySew_3_29};
  wire [23:0]       dataInMem_lo_291 = {dataInMem_lo_hi_35, dataRegroupBySew_0_30};
  wire [15:0]       _GEN_548 = {dataRegroupBySew_5_30, dataRegroupBySew_4_30};
  wire [15:0]       dataInMem_hi_hi_163;
  assign dataInMem_hi_hi_163 = _GEN_548;
  wire [15:0]       dataInMem_hi_lo_165;
  assign dataInMem_hi_lo_165 = _GEN_548;
  wire [23:0]       dataInMem_hi_419 = {dataInMem_hi_hi_163, dataRegroupBySew_3_30};
  wire [23:0]       dataInMem_lo_292 = {dataInMem_lo_hi_36, dataRegroupBySew_0_31};
  wire [15:0]       _GEN_549 = {dataRegroupBySew_5_31, dataRegroupBySew_4_31};
  wire [15:0]       dataInMem_hi_hi_164;
  assign dataInMem_hi_hi_164 = _GEN_549;
  wire [15:0]       dataInMem_hi_lo_166;
  assign dataInMem_hi_lo_166 = _GEN_549;
  wire [23:0]       dataInMem_hi_420 = {dataInMem_hi_hi_164, dataRegroupBySew_3_31};
  wire [23:0]       dataInMem_lo_293 = {dataInMem_lo_hi_37, dataRegroupBySew_0_32};
  wire [15:0]       _GEN_550 = {dataRegroupBySew_5_32, dataRegroupBySew_4_32};
  wire [15:0]       dataInMem_hi_hi_165;
  assign dataInMem_hi_hi_165 = _GEN_550;
  wire [15:0]       dataInMem_hi_lo_167;
  assign dataInMem_hi_lo_167 = _GEN_550;
  wire [23:0]       dataInMem_hi_421 = {dataInMem_hi_hi_165, dataRegroupBySew_3_32};
  wire [23:0]       dataInMem_lo_294 = {dataInMem_lo_hi_38, dataRegroupBySew_0_33};
  wire [15:0]       _GEN_551 = {dataRegroupBySew_5_33, dataRegroupBySew_4_33};
  wire [15:0]       dataInMem_hi_hi_166;
  assign dataInMem_hi_hi_166 = _GEN_551;
  wire [15:0]       dataInMem_hi_lo_168;
  assign dataInMem_hi_lo_168 = _GEN_551;
  wire [23:0]       dataInMem_hi_422 = {dataInMem_hi_hi_166, dataRegroupBySew_3_33};
  wire [23:0]       dataInMem_lo_295 = {dataInMem_lo_hi_39, dataRegroupBySew_0_34};
  wire [15:0]       _GEN_552 = {dataRegroupBySew_5_34, dataRegroupBySew_4_34};
  wire [15:0]       dataInMem_hi_hi_167;
  assign dataInMem_hi_hi_167 = _GEN_552;
  wire [15:0]       dataInMem_hi_lo_169;
  assign dataInMem_hi_lo_169 = _GEN_552;
  wire [23:0]       dataInMem_hi_423 = {dataInMem_hi_hi_167, dataRegroupBySew_3_34};
  wire [23:0]       dataInMem_lo_296 = {dataInMem_lo_hi_40, dataRegroupBySew_0_35};
  wire [15:0]       _GEN_553 = {dataRegroupBySew_5_35, dataRegroupBySew_4_35};
  wire [15:0]       dataInMem_hi_hi_168;
  assign dataInMem_hi_hi_168 = _GEN_553;
  wire [15:0]       dataInMem_hi_lo_170;
  assign dataInMem_hi_lo_170 = _GEN_553;
  wire [23:0]       dataInMem_hi_424 = {dataInMem_hi_hi_168, dataRegroupBySew_3_35};
  wire [23:0]       dataInMem_lo_297 = {dataInMem_lo_hi_41, dataRegroupBySew_0_36};
  wire [15:0]       _GEN_554 = {dataRegroupBySew_5_36, dataRegroupBySew_4_36};
  wire [15:0]       dataInMem_hi_hi_169;
  assign dataInMem_hi_hi_169 = _GEN_554;
  wire [15:0]       dataInMem_hi_lo_171;
  assign dataInMem_hi_lo_171 = _GEN_554;
  wire [23:0]       dataInMem_hi_425 = {dataInMem_hi_hi_169, dataRegroupBySew_3_36};
  wire [23:0]       dataInMem_lo_298 = {dataInMem_lo_hi_42, dataRegroupBySew_0_37};
  wire [15:0]       _GEN_555 = {dataRegroupBySew_5_37, dataRegroupBySew_4_37};
  wire [15:0]       dataInMem_hi_hi_170;
  assign dataInMem_hi_hi_170 = _GEN_555;
  wire [15:0]       dataInMem_hi_lo_172;
  assign dataInMem_hi_lo_172 = _GEN_555;
  wire [23:0]       dataInMem_hi_426 = {dataInMem_hi_hi_170, dataRegroupBySew_3_37};
  wire [23:0]       dataInMem_lo_299 = {dataInMem_lo_hi_43, dataRegroupBySew_0_38};
  wire [15:0]       _GEN_556 = {dataRegroupBySew_5_38, dataRegroupBySew_4_38};
  wire [15:0]       dataInMem_hi_hi_171;
  assign dataInMem_hi_hi_171 = _GEN_556;
  wire [15:0]       dataInMem_hi_lo_173;
  assign dataInMem_hi_lo_173 = _GEN_556;
  wire [23:0]       dataInMem_hi_427 = {dataInMem_hi_hi_171, dataRegroupBySew_3_38};
  wire [23:0]       dataInMem_lo_300 = {dataInMem_lo_hi_44, dataRegroupBySew_0_39};
  wire [15:0]       _GEN_557 = {dataRegroupBySew_5_39, dataRegroupBySew_4_39};
  wire [15:0]       dataInMem_hi_hi_172;
  assign dataInMem_hi_hi_172 = _GEN_557;
  wire [15:0]       dataInMem_hi_lo_174;
  assign dataInMem_hi_lo_174 = _GEN_557;
  wire [23:0]       dataInMem_hi_428 = {dataInMem_hi_hi_172, dataRegroupBySew_3_39};
  wire [23:0]       dataInMem_lo_301 = {dataInMem_lo_hi_45, dataRegroupBySew_0_40};
  wire [15:0]       _GEN_558 = {dataRegroupBySew_5_40, dataRegroupBySew_4_40};
  wire [15:0]       dataInMem_hi_hi_173;
  assign dataInMem_hi_hi_173 = _GEN_558;
  wire [15:0]       dataInMem_hi_lo_175;
  assign dataInMem_hi_lo_175 = _GEN_558;
  wire [23:0]       dataInMem_hi_429 = {dataInMem_hi_hi_173, dataRegroupBySew_3_40};
  wire [23:0]       dataInMem_lo_302 = {dataInMem_lo_hi_46, dataRegroupBySew_0_41};
  wire [15:0]       _GEN_559 = {dataRegroupBySew_5_41, dataRegroupBySew_4_41};
  wire [15:0]       dataInMem_hi_hi_174;
  assign dataInMem_hi_hi_174 = _GEN_559;
  wire [15:0]       dataInMem_hi_lo_176;
  assign dataInMem_hi_lo_176 = _GEN_559;
  wire [23:0]       dataInMem_hi_430 = {dataInMem_hi_hi_174, dataRegroupBySew_3_41};
  wire [23:0]       dataInMem_lo_303 = {dataInMem_lo_hi_47, dataRegroupBySew_0_42};
  wire [15:0]       _GEN_560 = {dataRegroupBySew_5_42, dataRegroupBySew_4_42};
  wire [15:0]       dataInMem_hi_hi_175;
  assign dataInMem_hi_hi_175 = _GEN_560;
  wire [15:0]       dataInMem_hi_lo_177;
  assign dataInMem_hi_lo_177 = _GEN_560;
  wire [23:0]       dataInMem_hi_431 = {dataInMem_hi_hi_175, dataRegroupBySew_3_42};
  wire [23:0]       dataInMem_lo_304 = {dataInMem_lo_hi_48, dataRegroupBySew_0_43};
  wire [15:0]       _GEN_561 = {dataRegroupBySew_5_43, dataRegroupBySew_4_43};
  wire [15:0]       dataInMem_hi_hi_176;
  assign dataInMem_hi_hi_176 = _GEN_561;
  wire [15:0]       dataInMem_hi_lo_178;
  assign dataInMem_hi_lo_178 = _GEN_561;
  wire [23:0]       dataInMem_hi_432 = {dataInMem_hi_hi_176, dataRegroupBySew_3_43};
  wire [23:0]       dataInMem_lo_305 = {dataInMem_lo_hi_49, dataRegroupBySew_0_44};
  wire [15:0]       _GEN_562 = {dataRegroupBySew_5_44, dataRegroupBySew_4_44};
  wire [15:0]       dataInMem_hi_hi_177;
  assign dataInMem_hi_hi_177 = _GEN_562;
  wire [15:0]       dataInMem_hi_lo_179;
  assign dataInMem_hi_lo_179 = _GEN_562;
  wire [23:0]       dataInMem_hi_433 = {dataInMem_hi_hi_177, dataRegroupBySew_3_44};
  wire [23:0]       dataInMem_lo_306 = {dataInMem_lo_hi_50, dataRegroupBySew_0_45};
  wire [15:0]       _GEN_563 = {dataRegroupBySew_5_45, dataRegroupBySew_4_45};
  wire [15:0]       dataInMem_hi_hi_178;
  assign dataInMem_hi_hi_178 = _GEN_563;
  wire [15:0]       dataInMem_hi_lo_180;
  assign dataInMem_hi_lo_180 = _GEN_563;
  wire [23:0]       dataInMem_hi_434 = {dataInMem_hi_hi_178, dataRegroupBySew_3_45};
  wire [23:0]       dataInMem_lo_307 = {dataInMem_lo_hi_51, dataRegroupBySew_0_46};
  wire [15:0]       _GEN_564 = {dataRegroupBySew_5_46, dataRegroupBySew_4_46};
  wire [15:0]       dataInMem_hi_hi_179;
  assign dataInMem_hi_hi_179 = _GEN_564;
  wire [15:0]       dataInMem_hi_lo_181;
  assign dataInMem_hi_lo_181 = _GEN_564;
  wire [23:0]       dataInMem_hi_435 = {dataInMem_hi_hi_179, dataRegroupBySew_3_46};
  wire [23:0]       dataInMem_lo_308 = {dataInMem_lo_hi_52, dataRegroupBySew_0_47};
  wire [15:0]       _GEN_565 = {dataRegroupBySew_5_47, dataRegroupBySew_4_47};
  wire [15:0]       dataInMem_hi_hi_180;
  assign dataInMem_hi_hi_180 = _GEN_565;
  wire [15:0]       dataInMem_hi_lo_182;
  assign dataInMem_hi_lo_182 = _GEN_565;
  wire [23:0]       dataInMem_hi_436 = {dataInMem_hi_hi_180, dataRegroupBySew_3_47};
  wire [23:0]       dataInMem_lo_309 = {dataInMem_lo_hi_53, dataRegroupBySew_0_48};
  wire [15:0]       _GEN_566 = {dataRegroupBySew_5_48, dataRegroupBySew_4_48};
  wire [15:0]       dataInMem_hi_hi_181;
  assign dataInMem_hi_hi_181 = _GEN_566;
  wire [15:0]       dataInMem_hi_lo_183;
  assign dataInMem_hi_lo_183 = _GEN_566;
  wire [23:0]       dataInMem_hi_437 = {dataInMem_hi_hi_181, dataRegroupBySew_3_48};
  wire [23:0]       dataInMem_lo_310 = {dataInMem_lo_hi_54, dataRegroupBySew_0_49};
  wire [15:0]       _GEN_567 = {dataRegroupBySew_5_49, dataRegroupBySew_4_49};
  wire [15:0]       dataInMem_hi_hi_182;
  assign dataInMem_hi_hi_182 = _GEN_567;
  wire [15:0]       dataInMem_hi_lo_184;
  assign dataInMem_hi_lo_184 = _GEN_567;
  wire [23:0]       dataInMem_hi_438 = {dataInMem_hi_hi_182, dataRegroupBySew_3_49};
  wire [23:0]       dataInMem_lo_311 = {dataInMem_lo_hi_55, dataRegroupBySew_0_50};
  wire [15:0]       _GEN_568 = {dataRegroupBySew_5_50, dataRegroupBySew_4_50};
  wire [15:0]       dataInMem_hi_hi_183;
  assign dataInMem_hi_hi_183 = _GEN_568;
  wire [15:0]       dataInMem_hi_lo_185;
  assign dataInMem_hi_lo_185 = _GEN_568;
  wire [23:0]       dataInMem_hi_439 = {dataInMem_hi_hi_183, dataRegroupBySew_3_50};
  wire [23:0]       dataInMem_lo_312 = {dataInMem_lo_hi_56, dataRegroupBySew_0_51};
  wire [15:0]       _GEN_569 = {dataRegroupBySew_5_51, dataRegroupBySew_4_51};
  wire [15:0]       dataInMem_hi_hi_184;
  assign dataInMem_hi_hi_184 = _GEN_569;
  wire [15:0]       dataInMem_hi_lo_186;
  assign dataInMem_hi_lo_186 = _GEN_569;
  wire [23:0]       dataInMem_hi_440 = {dataInMem_hi_hi_184, dataRegroupBySew_3_51};
  wire [23:0]       dataInMem_lo_313 = {dataInMem_lo_hi_57, dataRegroupBySew_0_52};
  wire [15:0]       _GEN_570 = {dataRegroupBySew_5_52, dataRegroupBySew_4_52};
  wire [15:0]       dataInMem_hi_hi_185;
  assign dataInMem_hi_hi_185 = _GEN_570;
  wire [15:0]       dataInMem_hi_lo_187;
  assign dataInMem_hi_lo_187 = _GEN_570;
  wire [23:0]       dataInMem_hi_441 = {dataInMem_hi_hi_185, dataRegroupBySew_3_52};
  wire [23:0]       dataInMem_lo_314 = {dataInMem_lo_hi_58, dataRegroupBySew_0_53};
  wire [15:0]       _GEN_571 = {dataRegroupBySew_5_53, dataRegroupBySew_4_53};
  wire [15:0]       dataInMem_hi_hi_186;
  assign dataInMem_hi_hi_186 = _GEN_571;
  wire [15:0]       dataInMem_hi_lo_188;
  assign dataInMem_hi_lo_188 = _GEN_571;
  wire [23:0]       dataInMem_hi_442 = {dataInMem_hi_hi_186, dataRegroupBySew_3_53};
  wire [23:0]       dataInMem_lo_315 = {dataInMem_lo_hi_59, dataRegroupBySew_0_54};
  wire [15:0]       _GEN_572 = {dataRegroupBySew_5_54, dataRegroupBySew_4_54};
  wire [15:0]       dataInMem_hi_hi_187;
  assign dataInMem_hi_hi_187 = _GEN_572;
  wire [15:0]       dataInMem_hi_lo_189;
  assign dataInMem_hi_lo_189 = _GEN_572;
  wire [23:0]       dataInMem_hi_443 = {dataInMem_hi_hi_187, dataRegroupBySew_3_54};
  wire [23:0]       dataInMem_lo_316 = {dataInMem_lo_hi_60, dataRegroupBySew_0_55};
  wire [15:0]       _GEN_573 = {dataRegroupBySew_5_55, dataRegroupBySew_4_55};
  wire [15:0]       dataInMem_hi_hi_188;
  assign dataInMem_hi_hi_188 = _GEN_573;
  wire [15:0]       dataInMem_hi_lo_190;
  assign dataInMem_hi_lo_190 = _GEN_573;
  wire [23:0]       dataInMem_hi_444 = {dataInMem_hi_hi_188, dataRegroupBySew_3_55};
  wire [23:0]       dataInMem_lo_317 = {dataInMem_lo_hi_61, dataRegroupBySew_0_56};
  wire [15:0]       _GEN_574 = {dataRegroupBySew_5_56, dataRegroupBySew_4_56};
  wire [15:0]       dataInMem_hi_hi_189;
  assign dataInMem_hi_hi_189 = _GEN_574;
  wire [15:0]       dataInMem_hi_lo_191;
  assign dataInMem_hi_lo_191 = _GEN_574;
  wire [23:0]       dataInMem_hi_445 = {dataInMem_hi_hi_189, dataRegroupBySew_3_56};
  wire [23:0]       dataInMem_lo_318 = {dataInMem_lo_hi_62, dataRegroupBySew_0_57};
  wire [15:0]       _GEN_575 = {dataRegroupBySew_5_57, dataRegroupBySew_4_57};
  wire [15:0]       dataInMem_hi_hi_190;
  assign dataInMem_hi_hi_190 = _GEN_575;
  wire [15:0]       dataInMem_hi_lo_192;
  assign dataInMem_hi_lo_192 = _GEN_575;
  wire [23:0]       dataInMem_hi_446 = {dataInMem_hi_hi_190, dataRegroupBySew_3_57};
  wire [23:0]       dataInMem_lo_319 = {dataInMem_lo_hi_63, dataRegroupBySew_0_58};
  wire [15:0]       _GEN_576 = {dataRegroupBySew_5_58, dataRegroupBySew_4_58};
  wire [15:0]       dataInMem_hi_hi_191;
  assign dataInMem_hi_hi_191 = _GEN_576;
  wire [15:0]       dataInMem_hi_lo_193;
  assign dataInMem_hi_lo_193 = _GEN_576;
  wire [23:0]       dataInMem_hi_447 = {dataInMem_hi_hi_191, dataRegroupBySew_3_58};
  wire [23:0]       dataInMem_lo_320 = {dataInMem_lo_hi_64, dataRegroupBySew_0_59};
  wire [15:0]       _GEN_577 = {dataRegroupBySew_5_59, dataRegroupBySew_4_59};
  wire [15:0]       dataInMem_hi_hi_192;
  assign dataInMem_hi_hi_192 = _GEN_577;
  wire [15:0]       dataInMem_hi_lo_194;
  assign dataInMem_hi_lo_194 = _GEN_577;
  wire [23:0]       dataInMem_hi_448 = {dataInMem_hi_hi_192, dataRegroupBySew_3_59};
  wire [23:0]       dataInMem_lo_321 = {dataInMem_lo_hi_65, dataRegroupBySew_0_60};
  wire [15:0]       _GEN_578 = {dataRegroupBySew_5_60, dataRegroupBySew_4_60};
  wire [15:0]       dataInMem_hi_hi_193;
  assign dataInMem_hi_hi_193 = _GEN_578;
  wire [15:0]       dataInMem_hi_lo_195;
  assign dataInMem_hi_lo_195 = _GEN_578;
  wire [23:0]       dataInMem_hi_449 = {dataInMem_hi_hi_193, dataRegroupBySew_3_60};
  wire [23:0]       dataInMem_lo_322 = {dataInMem_lo_hi_66, dataRegroupBySew_0_61};
  wire [15:0]       _GEN_579 = {dataRegroupBySew_5_61, dataRegroupBySew_4_61};
  wire [15:0]       dataInMem_hi_hi_194;
  assign dataInMem_hi_hi_194 = _GEN_579;
  wire [15:0]       dataInMem_hi_lo_196;
  assign dataInMem_hi_lo_196 = _GEN_579;
  wire [23:0]       dataInMem_hi_450 = {dataInMem_hi_hi_194, dataRegroupBySew_3_61};
  wire [23:0]       dataInMem_lo_323 = {dataInMem_lo_hi_67, dataRegroupBySew_0_62};
  wire [15:0]       _GEN_580 = {dataRegroupBySew_5_62, dataRegroupBySew_4_62};
  wire [15:0]       dataInMem_hi_hi_195;
  assign dataInMem_hi_hi_195 = _GEN_580;
  wire [15:0]       dataInMem_hi_lo_197;
  assign dataInMem_hi_lo_197 = _GEN_580;
  wire [23:0]       dataInMem_hi_451 = {dataInMem_hi_hi_195, dataRegroupBySew_3_62};
  wire [23:0]       dataInMem_lo_324 = {dataInMem_lo_hi_68, dataRegroupBySew_0_63};
  wire [15:0]       _GEN_581 = {dataRegroupBySew_5_63, dataRegroupBySew_4_63};
  wire [15:0]       dataInMem_hi_hi_196;
  assign dataInMem_hi_hi_196 = _GEN_581;
  wire [15:0]       dataInMem_hi_lo_198;
  assign dataInMem_hi_lo_198 = _GEN_581;
  wire [23:0]       dataInMem_hi_452 = {dataInMem_hi_hi_196, dataRegroupBySew_3_63};
  wire [23:0]       dataInMem_lo_325 = {dataInMem_lo_hi_69, dataRegroupBySew_0_64};
  wire [15:0]       _GEN_582 = {dataRegroupBySew_5_64, dataRegroupBySew_4_64};
  wire [15:0]       dataInMem_hi_hi_197;
  assign dataInMem_hi_hi_197 = _GEN_582;
  wire [15:0]       dataInMem_hi_lo_199;
  assign dataInMem_hi_lo_199 = _GEN_582;
  wire [23:0]       dataInMem_hi_453 = {dataInMem_hi_hi_197, dataRegroupBySew_3_64};
  wire [23:0]       dataInMem_lo_326 = {dataInMem_lo_hi_70, dataRegroupBySew_0_65};
  wire [15:0]       _GEN_583 = {dataRegroupBySew_5_65, dataRegroupBySew_4_65};
  wire [15:0]       dataInMem_hi_hi_198;
  assign dataInMem_hi_hi_198 = _GEN_583;
  wire [15:0]       dataInMem_hi_lo_200;
  assign dataInMem_hi_lo_200 = _GEN_583;
  wire [23:0]       dataInMem_hi_454 = {dataInMem_hi_hi_198, dataRegroupBySew_3_65};
  wire [23:0]       dataInMem_lo_327 = {dataInMem_lo_hi_71, dataRegroupBySew_0_66};
  wire [15:0]       _GEN_584 = {dataRegroupBySew_5_66, dataRegroupBySew_4_66};
  wire [15:0]       dataInMem_hi_hi_199;
  assign dataInMem_hi_hi_199 = _GEN_584;
  wire [15:0]       dataInMem_hi_lo_201;
  assign dataInMem_hi_lo_201 = _GEN_584;
  wire [23:0]       dataInMem_hi_455 = {dataInMem_hi_hi_199, dataRegroupBySew_3_66};
  wire [23:0]       dataInMem_lo_328 = {dataInMem_lo_hi_72, dataRegroupBySew_0_67};
  wire [15:0]       _GEN_585 = {dataRegroupBySew_5_67, dataRegroupBySew_4_67};
  wire [15:0]       dataInMem_hi_hi_200;
  assign dataInMem_hi_hi_200 = _GEN_585;
  wire [15:0]       dataInMem_hi_lo_202;
  assign dataInMem_hi_lo_202 = _GEN_585;
  wire [23:0]       dataInMem_hi_456 = {dataInMem_hi_hi_200, dataRegroupBySew_3_67};
  wire [23:0]       dataInMem_lo_329 = {dataInMem_lo_hi_73, dataRegroupBySew_0_68};
  wire [15:0]       _GEN_586 = {dataRegroupBySew_5_68, dataRegroupBySew_4_68};
  wire [15:0]       dataInMem_hi_hi_201;
  assign dataInMem_hi_hi_201 = _GEN_586;
  wire [15:0]       dataInMem_hi_lo_203;
  assign dataInMem_hi_lo_203 = _GEN_586;
  wire [23:0]       dataInMem_hi_457 = {dataInMem_hi_hi_201, dataRegroupBySew_3_68};
  wire [23:0]       dataInMem_lo_330 = {dataInMem_lo_hi_74, dataRegroupBySew_0_69};
  wire [15:0]       _GEN_587 = {dataRegroupBySew_5_69, dataRegroupBySew_4_69};
  wire [15:0]       dataInMem_hi_hi_202;
  assign dataInMem_hi_hi_202 = _GEN_587;
  wire [15:0]       dataInMem_hi_lo_204;
  assign dataInMem_hi_lo_204 = _GEN_587;
  wire [23:0]       dataInMem_hi_458 = {dataInMem_hi_hi_202, dataRegroupBySew_3_69};
  wire [23:0]       dataInMem_lo_331 = {dataInMem_lo_hi_75, dataRegroupBySew_0_70};
  wire [15:0]       _GEN_588 = {dataRegroupBySew_5_70, dataRegroupBySew_4_70};
  wire [15:0]       dataInMem_hi_hi_203;
  assign dataInMem_hi_hi_203 = _GEN_588;
  wire [15:0]       dataInMem_hi_lo_205;
  assign dataInMem_hi_lo_205 = _GEN_588;
  wire [23:0]       dataInMem_hi_459 = {dataInMem_hi_hi_203, dataRegroupBySew_3_70};
  wire [23:0]       dataInMem_lo_332 = {dataInMem_lo_hi_76, dataRegroupBySew_0_71};
  wire [15:0]       _GEN_589 = {dataRegroupBySew_5_71, dataRegroupBySew_4_71};
  wire [15:0]       dataInMem_hi_hi_204;
  assign dataInMem_hi_hi_204 = _GEN_589;
  wire [15:0]       dataInMem_hi_lo_206;
  assign dataInMem_hi_lo_206 = _GEN_589;
  wire [23:0]       dataInMem_hi_460 = {dataInMem_hi_hi_204, dataRegroupBySew_3_71};
  wire [23:0]       dataInMem_lo_333 = {dataInMem_lo_hi_77, dataRegroupBySew_0_72};
  wire [15:0]       _GEN_590 = {dataRegroupBySew_5_72, dataRegroupBySew_4_72};
  wire [15:0]       dataInMem_hi_hi_205;
  assign dataInMem_hi_hi_205 = _GEN_590;
  wire [15:0]       dataInMem_hi_lo_207;
  assign dataInMem_hi_lo_207 = _GEN_590;
  wire [23:0]       dataInMem_hi_461 = {dataInMem_hi_hi_205, dataRegroupBySew_3_72};
  wire [23:0]       dataInMem_lo_334 = {dataInMem_lo_hi_78, dataRegroupBySew_0_73};
  wire [15:0]       _GEN_591 = {dataRegroupBySew_5_73, dataRegroupBySew_4_73};
  wire [15:0]       dataInMem_hi_hi_206;
  assign dataInMem_hi_hi_206 = _GEN_591;
  wire [15:0]       dataInMem_hi_lo_208;
  assign dataInMem_hi_lo_208 = _GEN_591;
  wire [23:0]       dataInMem_hi_462 = {dataInMem_hi_hi_206, dataRegroupBySew_3_73};
  wire [23:0]       dataInMem_lo_335 = {dataInMem_lo_hi_79, dataRegroupBySew_0_74};
  wire [15:0]       _GEN_592 = {dataRegroupBySew_5_74, dataRegroupBySew_4_74};
  wire [15:0]       dataInMem_hi_hi_207;
  assign dataInMem_hi_hi_207 = _GEN_592;
  wire [15:0]       dataInMem_hi_lo_209;
  assign dataInMem_hi_lo_209 = _GEN_592;
  wire [23:0]       dataInMem_hi_463 = {dataInMem_hi_hi_207, dataRegroupBySew_3_74};
  wire [23:0]       dataInMem_lo_336 = {dataInMem_lo_hi_80, dataRegroupBySew_0_75};
  wire [15:0]       _GEN_593 = {dataRegroupBySew_5_75, dataRegroupBySew_4_75};
  wire [15:0]       dataInMem_hi_hi_208;
  assign dataInMem_hi_hi_208 = _GEN_593;
  wire [15:0]       dataInMem_hi_lo_210;
  assign dataInMem_hi_lo_210 = _GEN_593;
  wire [23:0]       dataInMem_hi_464 = {dataInMem_hi_hi_208, dataRegroupBySew_3_75};
  wire [23:0]       dataInMem_lo_337 = {dataInMem_lo_hi_81, dataRegroupBySew_0_76};
  wire [15:0]       _GEN_594 = {dataRegroupBySew_5_76, dataRegroupBySew_4_76};
  wire [15:0]       dataInMem_hi_hi_209;
  assign dataInMem_hi_hi_209 = _GEN_594;
  wire [15:0]       dataInMem_hi_lo_211;
  assign dataInMem_hi_lo_211 = _GEN_594;
  wire [23:0]       dataInMem_hi_465 = {dataInMem_hi_hi_209, dataRegroupBySew_3_76};
  wire [23:0]       dataInMem_lo_338 = {dataInMem_lo_hi_82, dataRegroupBySew_0_77};
  wire [15:0]       _GEN_595 = {dataRegroupBySew_5_77, dataRegroupBySew_4_77};
  wire [15:0]       dataInMem_hi_hi_210;
  assign dataInMem_hi_hi_210 = _GEN_595;
  wire [15:0]       dataInMem_hi_lo_212;
  assign dataInMem_hi_lo_212 = _GEN_595;
  wire [23:0]       dataInMem_hi_466 = {dataInMem_hi_hi_210, dataRegroupBySew_3_77};
  wire [23:0]       dataInMem_lo_339 = {dataInMem_lo_hi_83, dataRegroupBySew_0_78};
  wire [15:0]       _GEN_596 = {dataRegroupBySew_5_78, dataRegroupBySew_4_78};
  wire [15:0]       dataInMem_hi_hi_211;
  assign dataInMem_hi_hi_211 = _GEN_596;
  wire [15:0]       dataInMem_hi_lo_213;
  assign dataInMem_hi_lo_213 = _GEN_596;
  wire [23:0]       dataInMem_hi_467 = {dataInMem_hi_hi_211, dataRegroupBySew_3_78};
  wire [23:0]       dataInMem_lo_340 = {dataInMem_lo_hi_84, dataRegroupBySew_0_79};
  wire [15:0]       _GEN_597 = {dataRegroupBySew_5_79, dataRegroupBySew_4_79};
  wire [15:0]       dataInMem_hi_hi_212;
  assign dataInMem_hi_hi_212 = _GEN_597;
  wire [15:0]       dataInMem_hi_lo_214;
  assign dataInMem_hi_lo_214 = _GEN_597;
  wire [23:0]       dataInMem_hi_468 = {dataInMem_hi_hi_212, dataRegroupBySew_3_79};
  wire [23:0]       dataInMem_lo_341 = {dataInMem_lo_hi_85, dataRegroupBySew_0_80};
  wire [15:0]       _GEN_598 = {dataRegroupBySew_5_80, dataRegroupBySew_4_80};
  wire [15:0]       dataInMem_hi_hi_213;
  assign dataInMem_hi_hi_213 = _GEN_598;
  wire [15:0]       dataInMem_hi_lo_215;
  assign dataInMem_hi_lo_215 = _GEN_598;
  wire [23:0]       dataInMem_hi_469 = {dataInMem_hi_hi_213, dataRegroupBySew_3_80};
  wire [23:0]       dataInMem_lo_342 = {dataInMem_lo_hi_86, dataRegroupBySew_0_81};
  wire [15:0]       _GEN_599 = {dataRegroupBySew_5_81, dataRegroupBySew_4_81};
  wire [15:0]       dataInMem_hi_hi_214;
  assign dataInMem_hi_hi_214 = _GEN_599;
  wire [15:0]       dataInMem_hi_lo_216;
  assign dataInMem_hi_lo_216 = _GEN_599;
  wire [23:0]       dataInMem_hi_470 = {dataInMem_hi_hi_214, dataRegroupBySew_3_81};
  wire [23:0]       dataInMem_lo_343 = {dataInMem_lo_hi_87, dataRegroupBySew_0_82};
  wire [15:0]       _GEN_600 = {dataRegroupBySew_5_82, dataRegroupBySew_4_82};
  wire [15:0]       dataInMem_hi_hi_215;
  assign dataInMem_hi_hi_215 = _GEN_600;
  wire [15:0]       dataInMem_hi_lo_217;
  assign dataInMem_hi_lo_217 = _GEN_600;
  wire [23:0]       dataInMem_hi_471 = {dataInMem_hi_hi_215, dataRegroupBySew_3_82};
  wire [23:0]       dataInMem_lo_344 = {dataInMem_lo_hi_88, dataRegroupBySew_0_83};
  wire [15:0]       _GEN_601 = {dataRegroupBySew_5_83, dataRegroupBySew_4_83};
  wire [15:0]       dataInMem_hi_hi_216;
  assign dataInMem_hi_hi_216 = _GEN_601;
  wire [15:0]       dataInMem_hi_lo_218;
  assign dataInMem_hi_lo_218 = _GEN_601;
  wire [23:0]       dataInMem_hi_472 = {dataInMem_hi_hi_216, dataRegroupBySew_3_83};
  wire [23:0]       dataInMem_lo_345 = {dataInMem_lo_hi_89, dataRegroupBySew_0_84};
  wire [15:0]       _GEN_602 = {dataRegroupBySew_5_84, dataRegroupBySew_4_84};
  wire [15:0]       dataInMem_hi_hi_217;
  assign dataInMem_hi_hi_217 = _GEN_602;
  wire [15:0]       dataInMem_hi_lo_219;
  assign dataInMem_hi_lo_219 = _GEN_602;
  wire [23:0]       dataInMem_hi_473 = {dataInMem_hi_hi_217, dataRegroupBySew_3_84};
  wire [23:0]       dataInMem_lo_346 = {dataInMem_lo_hi_90, dataRegroupBySew_0_85};
  wire [15:0]       _GEN_603 = {dataRegroupBySew_5_85, dataRegroupBySew_4_85};
  wire [15:0]       dataInMem_hi_hi_218;
  assign dataInMem_hi_hi_218 = _GEN_603;
  wire [15:0]       dataInMem_hi_lo_220;
  assign dataInMem_hi_lo_220 = _GEN_603;
  wire [23:0]       dataInMem_hi_474 = {dataInMem_hi_hi_218, dataRegroupBySew_3_85};
  wire [23:0]       dataInMem_lo_347 = {dataInMem_lo_hi_91, dataRegroupBySew_0_86};
  wire [15:0]       _GEN_604 = {dataRegroupBySew_5_86, dataRegroupBySew_4_86};
  wire [15:0]       dataInMem_hi_hi_219;
  assign dataInMem_hi_hi_219 = _GEN_604;
  wire [15:0]       dataInMem_hi_lo_221;
  assign dataInMem_hi_lo_221 = _GEN_604;
  wire [23:0]       dataInMem_hi_475 = {dataInMem_hi_hi_219, dataRegroupBySew_3_86};
  wire [23:0]       dataInMem_lo_348 = {dataInMem_lo_hi_92, dataRegroupBySew_0_87};
  wire [15:0]       _GEN_605 = {dataRegroupBySew_5_87, dataRegroupBySew_4_87};
  wire [15:0]       dataInMem_hi_hi_220;
  assign dataInMem_hi_hi_220 = _GEN_605;
  wire [15:0]       dataInMem_hi_lo_222;
  assign dataInMem_hi_lo_222 = _GEN_605;
  wire [23:0]       dataInMem_hi_476 = {dataInMem_hi_hi_220, dataRegroupBySew_3_87};
  wire [23:0]       dataInMem_lo_349 = {dataInMem_lo_hi_93, dataRegroupBySew_0_88};
  wire [15:0]       _GEN_606 = {dataRegroupBySew_5_88, dataRegroupBySew_4_88};
  wire [15:0]       dataInMem_hi_hi_221;
  assign dataInMem_hi_hi_221 = _GEN_606;
  wire [15:0]       dataInMem_hi_lo_223;
  assign dataInMem_hi_lo_223 = _GEN_606;
  wire [23:0]       dataInMem_hi_477 = {dataInMem_hi_hi_221, dataRegroupBySew_3_88};
  wire [23:0]       dataInMem_lo_350 = {dataInMem_lo_hi_94, dataRegroupBySew_0_89};
  wire [15:0]       _GEN_607 = {dataRegroupBySew_5_89, dataRegroupBySew_4_89};
  wire [15:0]       dataInMem_hi_hi_222;
  assign dataInMem_hi_hi_222 = _GEN_607;
  wire [15:0]       dataInMem_hi_lo_224;
  assign dataInMem_hi_lo_224 = _GEN_607;
  wire [23:0]       dataInMem_hi_478 = {dataInMem_hi_hi_222, dataRegroupBySew_3_89};
  wire [23:0]       dataInMem_lo_351 = {dataInMem_lo_hi_95, dataRegroupBySew_0_90};
  wire [15:0]       _GEN_608 = {dataRegroupBySew_5_90, dataRegroupBySew_4_90};
  wire [15:0]       dataInMem_hi_hi_223;
  assign dataInMem_hi_hi_223 = _GEN_608;
  wire [15:0]       dataInMem_hi_lo_225;
  assign dataInMem_hi_lo_225 = _GEN_608;
  wire [23:0]       dataInMem_hi_479 = {dataInMem_hi_hi_223, dataRegroupBySew_3_90};
  wire [23:0]       dataInMem_lo_352 = {dataInMem_lo_hi_96, dataRegroupBySew_0_91};
  wire [15:0]       _GEN_609 = {dataRegroupBySew_5_91, dataRegroupBySew_4_91};
  wire [15:0]       dataInMem_hi_hi_224;
  assign dataInMem_hi_hi_224 = _GEN_609;
  wire [15:0]       dataInMem_hi_lo_226;
  assign dataInMem_hi_lo_226 = _GEN_609;
  wire [23:0]       dataInMem_hi_480 = {dataInMem_hi_hi_224, dataRegroupBySew_3_91};
  wire [23:0]       dataInMem_lo_353 = {dataInMem_lo_hi_97, dataRegroupBySew_0_92};
  wire [15:0]       _GEN_610 = {dataRegroupBySew_5_92, dataRegroupBySew_4_92};
  wire [15:0]       dataInMem_hi_hi_225;
  assign dataInMem_hi_hi_225 = _GEN_610;
  wire [15:0]       dataInMem_hi_lo_227;
  assign dataInMem_hi_lo_227 = _GEN_610;
  wire [23:0]       dataInMem_hi_481 = {dataInMem_hi_hi_225, dataRegroupBySew_3_92};
  wire [23:0]       dataInMem_lo_354 = {dataInMem_lo_hi_98, dataRegroupBySew_0_93};
  wire [15:0]       _GEN_611 = {dataRegroupBySew_5_93, dataRegroupBySew_4_93};
  wire [15:0]       dataInMem_hi_hi_226;
  assign dataInMem_hi_hi_226 = _GEN_611;
  wire [15:0]       dataInMem_hi_lo_228;
  assign dataInMem_hi_lo_228 = _GEN_611;
  wire [23:0]       dataInMem_hi_482 = {dataInMem_hi_hi_226, dataRegroupBySew_3_93};
  wire [23:0]       dataInMem_lo_355 = {dataInMem_lo_hi_99, dataRegroupBySew_0_94};
  wire [15:0]       _GEN_612 = {dataRegroupBySew_5_94, dataRegroupBySew_4_94};
  wire [15:0]       dataInMem_hi_hi_227;
  assign dataInMem_hi_hi_227 = _GEN_612;
  wire [15:0]       dataInMem_hi_lo_229;
  assign dataInMem_hi_lo_229 = _GEN_612;
  wire [23:0]       dataInMem_hi_483 = {dataInMem_hi_hi_227, dataRegroupBySew_3_94};
  wire [23:0]       dataInMem_lo_356 = {dataInMem_lo_hi_100, dataRegroupBySew_0_95};
  wire [15:0]       _GEN_613 = {dataRegroupBySew_5_95, dataRegroupBySew_4_95};
  wire [15:0]       dataInMem_hi_hi_228;
  assign dataInMem_hi_hi_228 = _GEN_613;
  wire [15:0]       dataInMem_hi_lo_230;
  assign dataInMem_hi_lo_230 = _GEN_613;
  wire [23:0]       dataInMem_hi_484 = {dataInMem_hi_hi_228, dataRegroupBySew_3_95};
  wire [23:0]       dataInMem_lo_357 = {dataInMem_lo_hi_101, dataRegroupBySew_0_96};
  wire [15:0]       _GEN_614 = {dataRegroupBySew_5_96, dataRegroupBySew_4_96};
  wire [15:0]       dataInMem_hi_hi_229;
  assign dataInMem_hi_hi_229 = _GEN_614;
  wire [15:0]       dataInMem_hi_lo_231;
  assign dataInMem_hi_lo_231 = _GEN_614;
  wire [23:0]       dataInMem_hi_485 = {dataInMem_hi_hi_229, dataRegroupBySew_3_96};
  wire [23:0]       dataInMem_lo_358 = {dataInMem_lo_hi_102, dataRegroupBySew_0_97};
  wire [15:0]       _GEN_615 = {dataRegroupBySew_5_97, dataRegroupBySew_4_97};
  wire [15:0]       dataInMem_hi_hi_230;
  assign dataInMem_hi_hi_230 = _GEN_615;
  wire [15:0]       dataInMem_hi_lo_232;
  assign dataInMem_hi_lo_232 = _GEN_615;
  wire [23:0]       dataInMem_hi_486 = {dataInMem_hi_hi_230, dataRegroupBySew_3_97};
  wire [23:0]       dataInMem_lo_359 = {dataInMem_lo_hi_103, dataRegroupBySew_0_98};
  wire [15:0]       _GEN_616 = {dataRegroupBySew_5_98, dataRegroupBySew_4_98};
  wire [15:0]       dataInMem_hi_hi_231;
  assign dataInMem_hi_hi_231 = _GEN_616;
  wire [15:0]       dataInMem_hi_lo_233;
  assign dataInMem_hi_lo_233 = _GEN_616;
  wire [23:0]       dataInMem_hi_487 = {dataInMem_hi_hi_231, dataRegroupBySew_3_98};
  wire [23:0]       dataInMem_lo_360 = {dataInMem_lo_hi_104, dataRegroupBySew_0_99};
  wire [15:0]       _GEN_617 = {dataRegroupBySew_5_99, dataRegroupBySew_4_99};
  wire [15:0]       dataInMem_hi_hi_232;
  assign dataInMem_hi_hi_232 = _GEN_617;
  wire [15:0]       dataInMem_hi_lo_234;
  assign dataInMem_hi_lo_234 = _GEN_617;
  wire [23:0]       dataInMem_hi_488 = {dataInMem_hi_hi_232, dataRegroupBySew_3_99};
  wire [23:0]       dataInMem_lo_361 = {dataInMem_lo_hi_105, dataRegroupBySew_0_100};
  wire [15:0]       _GEN_618 = {dataRegroupBySew_5_100, dataRegroupBySew_4_100};
  wire [15:0]       dataInMem_hi_hi_233;
  assign dataInMem_hi_hi_233 = _GEN_618;
  wire [15:0]       dataInMem_hi_lo_235;
  assign dataInMem_hi_lo_235 = _GEN_618;
  wire [23:0]       dataInMem_hi_489 = {dataInMem_hi_hi_233, dataRegroupBySew_3_100};
  wire [23:0]       dataInMem_lo_362 = {dataInMem_lo_hi_106, dataRegroupBySew_0_101};
  wire [15:0]       _GEN_619 = {dataRegroupBySew_5_101, dataRegroupBySew_4_101};
  wire [15:0]       dataInMem_hi_hi_234;
  assign dataInMem_hi_hi_234 = _GEN_619;
  wire [15:0]       dataInMem_hi_lo_236;
  assign dataInMem_hi_lo_236 = _GEN_619;
  wire [23:0]       dataInMem_hi_490 = {dataInMem_hi_hi_234, dataRegroupBySew_3_101};
  wire [23:0]       dataInMem_lo_363 = {dataInMem_lo_hi_107, dataRegroupBySew_0_102};
  wire [15:0]       _GEN_620 = {dataRegroupBySew_5_102, dataRegroupBySew_4_102};
  wire [15:0]       dataInMem_hi_hi_235;
  assign dataInMem_hi_hi_235 = _GEN_620;
  wire [15:0]       dataInMem_hi_lo_237;
  assign dataInMem_hi_lo_237 = _GEN_620;
  wire [23:0]       dataInMem_hi_491 = {dataInMem_hi_hi_235, dataRegroupBySew_3_102};
  wire [23:0]       dataInMem_lo_364 = {dataInMem_lo_hi_108, dataRegroupBySew_0_103};
  wire [15:0]       _GEN_621 = {dataRegroupBySew_5_103, dataRegroupBySew_4_103};
  wire [15:0]       dataInMem_hi_hi_236;
  assign dataInMem_hi_hi_236 = _GEN_621;
  wire [15:0]       dataInMem_hi_lo_238;
  assign dataInMem_hi_lo_238 = _GEN_621;
  wire [23:0]       dataInMem_hi_492 = {dataInMem_hi_hi_236, dataRegroupBySew_3_103};
  wire [23:0]       dataInMem_lo_365 = {dataInMem_lo_hi_109, dataRegroupBySew_0_104};
  wire [15:0]       _GEN_622 = {dataRegroupBySew_5_104, dataRegroupBySew_4_104};
  wire [15:0]       dataInMem_hi_hi_237;
  assign dataInMem_hi_hi_237 = _GEN_622;
  wire [15:0]       dataInMem_hi_lo_239;
  assign dataInMem_hi_lo_239 = _GEN_622;
  wire [23:0]       dataInMem_hi_493 = {dataInMem_hi_hi_237, dataRegroupBySew_3_104};
  wire [23:0]       dataInMem_lo_366 = {dataInMem_lo_hi_110, dataRegroupBySew_0_105};
  wire [15:0]       _GEN_623 = {dataRegroupBySew_5_105, dataRegroupBySew_4_105};
  wire [15:0]       dataInMem_hi_hi_238;
  assign dataInMem_hi_hi_238 = _GEN_623;
  wire [15:0]       dataInMem_hi_lo_240;
  assign dataInMem_hi_lo_240 = _GEN_623;
  wire [23:0]       dataInMem_hi_494 = {dataInMem_hi_hi_238, dataRegroupBySew_3_105};
  wire [23:0]       dataInMem_lo_367 = {dataInMem_lo_hi_111, dataRegroupBySew_0_106};
  wire [15:0]       _GEN_624 = {dataRegroupBySew_5_106, dataRegroupBySew_4_106};
  wire [15:0]       dataInMem_hi_hi_239;
  assign dataInMem_hi_hi_239 = _GEN_624;
  wire [15:0]       dataInMem_hi_lo_241;
  assign dataInMem_hi_lo_241 = _GEN_624;
  wire [23:0]       dataInMem_hi_495 = {dataInMem_hi_hi_239, dataRegroupBySew_3_106};
  wire [23:0]       dataInMem_lo_368 = {dataInMem_lo_hi_112, dataRegroupBySew_0_107};
  wire [15:0]       _GEN_625 = {dataRegroupBySew_5_107, dataRegroupBySew_4_107};
  wire [15:0]       dataInMem_hi_hi_240;
  assign dataInMem_hi_hi_240 = _GEN_625;
  wire [15:0]       dataInMem_hi_lo_242;
  assign dataInMem_hi_lo_242 = _GEN_625;
  wire [23:0]       dataInMem_hi_496 = {dataInMem_hi_hi_240, dataRegroupBySew_3_107};
  wire [23:0]       dataInMem_lo_369 = {dataInMem_lo_hi_113, dataRegroupBySew_0_108};
  wire [15:0]       _GEN_626 = {dataRegroupBySew_5_108, dataRegroupBySew_4_108};
  wire [15:0]       dataInMem_hi_hi_241;
  assign dataInMem_hi_hi_241 = _GEN_626;
  wire [15:0]       dataInMem_hi_lo_243;
  assign dataInMem_hi_lo_243 = _GEN_626;
  wire [23:0]       dataInMem_hi_497 = {dataInMem_hi_hi_241, dataRegroupBySew_3_108};
  wire [23:0]       dataInMem_lo_370 = {dataInMem_lo_hi_114, dataRegroupBySew_0_109};
  wire [15:0]       _GEN_627 = {dataRegroupBySew_5_109, dataRegroupBySew_4_109};
  wire [15:0]       dataInMem_hi_hi_242;
  assign dataInMem_hi_hi_242 = _GEN_627;
  wire [15:0]       dataInMem_hi_lo_244;
  assign dataInMem_hi_lo_244 = _GEN_627;
  wire [23:0]       dataInMem_hi_498 = {dataInMem_hi_hi_242, dataRegroupBySew_3_109};
  wire [23:0]       dataInMem_lo_371 = {dataInMem_lo_hi_115, dataRegroupBySew_0_110};
  wire [15:0]       _GEN_628 = {dataRegroupBySew_5_110, dataRegroupBySew_4_110};
  wire [15:0]       dataInMem_hi_hi_243;
  assign dataInMem_hi_hi_243 = _GEN_628;
  wire [15:0]       dataInMem_hi_lo_245;
  assign dataInMem_hi_lo_245 = _GEN_628;
  wire [23:0]       dataInMem_hi_499 = {dataInMem_hi_hi_243, dataRegroupBySew_3_110};
  wire [23:0]       dataInMem_lo_372 = {dataInMem_lo_hi_116, dataRegroupBySew_0_111};
  wire [15:0]       _GEN_629 = {dataRegroupBySew_5_111, dataRegroupBySew_4_111};
  wire [15:0]       dataInMem_hi_hi_244;
  assign dataInMem_hi_hi_244 = _GEN_629;
  wire [15:0]       dataInMem_hi_lo_246;
  assign dataInMem_hi_lo_246 = _GEN_629;
  wire [23:0]       dataInMem_hi_500 = {dataInMem_hi_hi_244, dataRegroupBySew_3_111};
  wire [23:0]       dataInMem_lo_373 = {dataInMem_lo_hi_117, dataRegroupBySew_0_112};
  wire [15:0]       _GEN_630 = {dataRegroupBySew_5_112, dataRegroupBySew_4_112};
  wire [15:0]       dataInMem_hi_hi_245;
  assign dataInMem_hi_hi_245 = _GEN_630;
  wire [15:0]       dataInMem_hi_lo_247;
  assign dataInMem_hi_lo_247 = _GEN_630;
  wire [23:0]       dataInMem_hi_501 = {dataInMem_hi_hi_245, dataRegroupBySew_3_112};
  wire [23:0]       dataInMem_lo_374 = {dataInMem_lo_hi_118, dataRegroupBySew_0_113};
  wire [15:0]       _GEN_631 = {dataRegroupBySew_5_113, dataRegroupBySew_4_113};
  wire [15:0]       dataInMem_hi_hi_246;
  assign dataInMem_hi_hi_246 = _GEN_631;
  wire [15:0]       dataInMem_hi_lo_248;
  assign dataInMem_hi_lo_248 = _GEN_631;
  wire [23:0]       dataInMem_hi_502 = {dataInMem_hi_hi_246, dataRegroupBySew_3_113};
  wire [23:0]       dataInMem_lo_375 = {dataInMem_lo_hi_119, dataRegroupBySew_0_114};
  wire [15:0]       _GEN_632 = {dataRegroupBySew_5_114, dataRegroupBySew_4_114};
  wire [15:0]       dataInMem_hi_hi_247;
  assign dataInMem_hi_hi_247 = _GEN_632;
  wire [15:0]       dataInMem_hi_lo_249;
  assign dataInMem_hi_lo_249 = _GEN_632;
  wire [23:0]       dataInMem_hi_503 = {dataInMem_hi_hi_247, dataRegroupBySew_3_114};
  wire [23:0]       dataInMem_lo_376 = {dataInMem_lo_hi_120, dataRegroupBySew_0_115};
  wire [15:0]       _GEN_633 = {dataRegroupBySew_5_115, dataRegroupBySew_4_115};
  wire [15:0]       dataInMem_hi_hi_248;
  assign dataInMem_hi_hi_248 = _GEN_633;
  wire [15:0]       dataInMem_hi_lo_250;
  assign dataInMem_hi_lo_250 = _GEN_633;
  wire [23:0]       dataInMem_hi_504 = {dataInMem_hi_hi_248, dataRegroupBySew_3_115};
  wire [23:0]       dataInMem_lo_377 = {dataInMem_lo_hi_121, dataRegroupBySew_0_116};
  wire [15:0]       _GEN_634 = {dataRegroupBySew_5_116, dataRegroupBySew_4_116};
  wire [15:0]       dataInMem_hi_hi_249;
  assign dataInMem_hi_hi_249 = _GEN_634;
  wire [15:0]       dataInMem_hi_lo_251;
  assign dataInMem_hi_lo_251 = _GEN_634;
  wire [23:0]       dataInMem_hi_505 = {dataInMem_hi_hi_249, dataRegroupBySew_3_116};
  wire [23:0]       dataInMem_lo_378 = {dataInMem_lo_hi_122, dataRegroupBySew_0_117};
  wire [15:0]       _GEN_635 = {dataRegroupBySew_5_117, dataRegroupBySew_4_117};
  wire [15:0]       dataInMem_hi_hi_250;
  assign dataInMem_hi_hi_250 = _GEN_635;
  wire [15:0]       dataInMem_hi_lo_252;
  assign dataInMem_hi_lo_252 = _GEN_635;
  wire [23:0]       dataInMem_hi_506 = {dataInMem_hi_hi_250, dataRegroupBySew_3_117};
  wire [23:0]       dataInMem_lo_379 = {dataInMem_lo_hi_123, dataRegroupBySew_0_118};
  wire [15:0]       _GEN_636 = {dataRegroupBySew_5_118, dataRegroupBySew_4_118};
  wire [15:0]       dataInMem_hi_hi_251;
  assign dataInMem_hi_hi_251 = _GEN_636;
  wire [15:0]       dataInMem_hi_lo_253;
  assign dataInMem_hi_lo_253 = _GEN_636;
  wire [23:0]       dataInMem_hi_507 = {dataInMem_hi_hi_251, dataRegroupBySew_3_118};
  wire [23:0]       dataInMem_lo_380 = {dataInMem_lo_hi_124, dataRegroupBySew_0_119};
  wire [15:0]       _GEN_637 = {dataRegroupBySew_5_119, dataRegroupBySew_4_119};
  wire [15:0]       dataInMem_hi_hi_252;
  assign dataInMem_hi_hi_252 = _GEN_637;
  wire [15:0]       dataInMem_hi_lo_254;
  assign dataInMem_hi_lo_254 = _GEN_637;
  wire [23:0]       dataInMem_hi_508 = {dataInMem_hi_hi_252, dataRegroupBySew_3_119};
  wire [23:0]       dataInMem_lo_381 = {dataInMem_lo_hi_125, dataRegroupBySew_0_120};
  wire [15:0]       _GEN_638 = {dataRegroupBySew_5_120, dataRegroupBySew_4_120};
  wire [15:0]       dataInMem_hi_hi_253;
  assign dataInMem_hi_hi_253 = _GEN_638;
  wire [15:0]       dataInMem_hi_lo_255;
  assign dataInMem_hi_lo_255 = _GEN_638;
  wire [23:0]       dataInMem_hi_509 = {dataInMem_hi_hi_253, dataRegroupBySew_3_120};
  wire [23:0]       dataInMem_lo_382 = {dataInMem_lo_hi_126, dataRegroupBySew_0_121};
  wire [15:0]       _GEN_639 = {dataRegroupBySew_5_121, dataRegroupBySew_4_121};
  wire [15:0]       dataInMem_hi_hi_254;
  assign dataInMem_hi_hi_254 = _GEN_639;
  wire [15:0]       dataInMem_hi_lo_256;
  assign dataInMem_hi_lo_256 = _GEN_639;
  wire [23:0]       dataInMem_hi_510 = {dataInMem_hi_hi_254, dataRegroupBySew_3_121};
  wire [23:0]       dataInMem_lo_383 = {dataInMem_lo_hi_127, dataRegroupBySew_0_122};
  wire [15:0]       _GEN_640 = {dataRegroupBySew_5_122, dataRegroupBySew_4_122};
  wire [15:0]       dataInMem_hi_hi_255;
  assign dataInMem_hi_hi_255 = _GEN_640;
  wire [15:0]       dataInMem_hi_lo_257;
  assign dataInMem_hi_lo_257 = _GEN_640;
  wire [23:0]       dataInMem_hi_511 = {dataInMem_hi_hi_255, dataRegroupBySew_3_122};
  wire [23:0]       dataInMem_lo_384 = {dataInMem_lo_hi_128, dataRegroupBySew_0_123};
  wire [15:0]       _GEN_641 = {dataRegroupBySew_5_123, dataRegroupBySew_4_123};
  wire [15:0]       dataInMem_hi_hi_256;
  assign dataInMem_hi_hi_256 = _GEN_641;
  wire [15:0]       dataInMem_hi_lo_258;
  assign dataInMem_hi_lo_258 = _GEN_641;
  wire [23:0]       dataInMem_hi_512 = {dataInMem_hi_hi_256, dataRegroupBySew_3_123};
  wire [23:0]       dataInMem_lo_385 = {dataInMem_lo_hi_129, dataRegroupBySew_0_124};
  wire [15:0]       _GEN_642 = {dataRegroupBySew_5_124, dataRegroupBySew_4_124};
  wire [15:0]       dataInMem_hi_hi_257;
  assign dataInMem_hi_hi_257 = _GEN_642;
  wire [15:0]       dataInMem_hi_lo_259;
  assign dataInMem_hi_lo_259 = _GEN_642;
  wire [23:0]       dataInMem_hi_513 = {dataInMem_hi_hi_257, dataRegroupBySew_3_124};
  wire [23:0]       dataInMem_lo_386 = {dataInMem_lo_hi_130, dataRegroupBySew_0_125};
  wire [15:0]       _GEN_643 = {dataRegroupBySew_5_125, dataRegroupBySew_4_125};
  wire [15:0]       dataInMem_hi_hi_258;
  assign dataInMem_hi_hi_258 = _GEN_643;
  wire [15:0]       dataInMem_hi_lo_260;
  assign dataInMem_hi_lo_260 = _GEN_643;
  wire [23:0]       dataInMem_hi_514 = {dataInMem_hi_hi_258, dataRegroupBySew_3_125};
  wire [23:0]       dataInMem_lo_387 = {dataInMem_lo_hi_131, dataRegroupBySew_0_126};
  wire [15:0]       _GEN_644 = {dataRegroupBySew_5_126, dataRegroupBySew_4_126};
  wire [15:0]       dataInMem_hi_hi_259;
  assign dataInMem_hi_hi_259 = _GEN_644;
  wire [15:0]       dataInMem_hi_lo_261;
  assign dataInMem_hi_lo_261 = _GEN_644;
  wire [23:0]       dataInMem_hi_515 = {dataInMem_hi_hi_259, dataRegroupBySew_3_126};
  wire [23:0]       dataInMem_lo_388 = {dataInMem_lo_hi_132, dataRegroupBySew_0_127};
  wire [15:0]       _GEN_645 = {dataRegroupBySew_5_127, dataRegroupBySew_4_127};
  wire [15:0]       dataInMem_hi_hi_260;
  assign dataInMem_hi_hi_260 = _GEN_645;
  wire [15:0]       dataInMem_hi_lo_262;
  assign dataInMem_hi_lo_262 = _GEN_645;
  wire [23:0]       dataInMem_hi_516 = {dataInMem_hi_hi_260, dataRegroupBySew_3_127};
  wire [95:0]       dataInMem_lo_lo_lo_lo_lo_lo_5 = {dataInMem_hi_390, dataInMem_lo_262, dataInMem_hi_389, dataInMem_lo_261};
  wire [95:0]       dataInMem_lo_lo_lo_lo_lo_hi_5 = {dataInMem_hi_392, dataInMem_lo_264, dataInMem_hi_391, dataInMem_lo_263};
  wire [191:0]      dataInMem_lo_lo_lo_lo_lo_5 = {dataInMem_lo_lo_lo_lo_lo_hi_5, dataInMem_lo_lo_lo_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_lo_lo_lo_hi_lo_5 = {dataInMem_hi_394, dataInMem_lo_266, dataInMem_hi_393, dataInMem_lo_265};
  wire [95:0]       dataInMem_lo_lo_lo_lo_hi_hi_5 = {dataInMem_hi_396, dataInMem_lo_268, dataInMem_hi_395, dataInMem_lo_267};
  wire [191:0]      dataInMem_lo_lo_lo_lo_hi_5 = {dataInMem_lo_lo_lo_lo_hi_hi_5, dataInMem_lo_lo_lo_lo_hi_lo_5};
  wire [383:0]      dataInMem_lo_lo_lo_lo_5 = {dataInMem_lo_lo_lo_lo_hi_5, dataInMem_lo_lo_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_lo_lo_hi_lo_lo_5 = {dataInMem_hi_398, dataInMem_lo_270, dataInMem_hi_397, dataInMem_lo_269};
  wire [95:0]       dataInMem_lo_lo_lo_hi_lo_hi_5 = {dataInMem_hi_400, dataInMem_lo_272, dataInMem_hi_399, dataInMem_lo_271};
  wire [191:0]      dataInMem_lo_lo_lo_hi_lo_5 = {dataInMem_lo_lo_lo_hi_lo_hi_5, dataInMem_lo_lo_lo_hi_lo_lo_5};
  wire [95:0]       dataInMem_lo_lo_lo_hi_hi_lo_5 = {dataInMem_hi_402, dataInMem_lo_274, dataInMem_hi_401, dataInMem_lo_273};
  wire [95:0]       dataInMem_lo_lo_lo_hi_hi_hi_5 = {dataInMem_hi_404, dataInMem_lo_276, dataInMem_hi_403, dataInMem_lo_275};
  wire [191:0]      dataInMem_lo_lo_lo_hi_hi_5 = {dataInMem_lo_lo_lo_hi_hi_hi_5, dataInMem_lo_lo_lo_hi_hi_lo_5};
  wire [383:0]      dataInMem_lo_lo_lo_hi_5 = {dataInMem_lo_lo_lo_hi_hi_5, dataInMem_lo_lo_lo_hi_lo_5};
  wire [767:0]      dataInMem_lo_lo_lo_5 = {dataInMem_lo_lo_lo_hi_5, dataInMem_lo_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_lo_hi_lo_lo_lo_5 = {dataInMem_hi_406, dataInMem_lo_278, dataInMem_hi_405, dataInMem_lo_277};
  wire [95:0]       dataInMem_lo_lo_hi_lo_lo_hi_5 = {dataInMem_hi_408, dataInMem_lo_280, dataInMem_hi_407, dataInMem_lo_279};
  wire [191:0]      dataInMem_lo_lo_hi_lo_lo_5 = {dataInMem_lo_lo_hi_lo_lo_hi_5, dataInMem_lo_lo_hi_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_lo_hi_lo_hi_lo_5 = {dataInMem_hi_410, dataInMem_lo_282, dataInMem_hi_409, dataInMem_lo_281};
  wire [95:0]       dataInMem_lo_lo_hi_lo_hi_hi_5 = {dataInMem_hi_412, dataInMem_lo_284, dataInMem_hi_411, dataInMem_lo_283};
  wire [191:0]      dataInMem_lo_lo_hi_lo_hi_5 = {dataInMem_lo_lo_hi_lo_hi_hi_5, dataInMem_lo_lo_hi_lo_hi_lo_5};
  wire [383:0]      dataInMem_lo_lo_hi_lo_5 = {dataInMem_lo_lo_hi_lo_hi_5, dataInMem_lo_lo_hi_lo_lo_5};
  wire [95:0]       dataInMem_lo_lo_hi_hi_lo_lo_5 = {dataInMem_hi_414, dataInMem_lo_286, dataInMem_hi_413, dataInMem_lo_285};
  wire [95:0]       dataInMem_lo_lo_hi_hi_lo_hi_5 = {dataInMem_hi_416, dataInMem_lo_288, dataInMem_hi_415, dataInMem_lo_287};
  wire [191:0]      dataInMem_lo_lo_hi_hi_lo_5 = {dataInMem_lo_lo_hi_hi_lo_hi_5, dataInMem_lo_lo_hi_hi_lo_lo_5};
  wire [95:0]       dataInMem_lo_lo_hi_hi_hi_lo_5 = {dataInMem_hi_418, dataInMem_lo_290, dataInMem_hi_417, dataInMem_lo_289};
  wire [95:0]       dataInMem_lo_lo_hi_hi_hi_hi_5 = {dataInMem_hi_420, dataInMem_lo_292, dataInMem_hi_419, dataInMem_lo_291};
  wire [191:0]      dataInMem_lo_lo_hi_hi_hi_5 = {dataInMem_lo_lo_hi_hi_hi_hi_5, dataInMem_lo_lo_hi_hi_hi_lo_5};
  wire [383:0]      dataInMem_lo_lo_hi_hi_5 = {dataInMem_lo_lo_hi_hi_hi_5, dataInMem_lo_lo_hi_hi_lo_5};
  wire [767:0]      dataInMem_lo_lo_hi_5 = {dataInMem_lo_lo_hi_hi_5, dataInMem_lo_lo_hi_lo_5};
  wire [1535:0]     dataInMem_lo_lo_5 = {dataInMem_lo_lo_hi_5, dataInMem_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_lo_lo_lo_lo_5 = {dataInMem_hi_422, dataInMem_lo_294, dataInMem_hi_421, dataInMem_lo_293};
  wire [95:0]       dataInMem_lo_hi_lo_lo_lo_hi_5 = {dataInMem_hi_424, dataInMem_lo_296, dataInMem_hi_423, dataInMem_lo_295};
  wire [191:0]      dataInMem_lo_hi_lo_lo_lo_5 = {dataInMem_lo_hi_lo_lo_lo_hi_5, dataInMem_lo_hi_lo_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_lo_lo_hi_lo_5 = {dataInMem_hi_426, dataInMem_lo_298, dataInMem_hi_425, dataInMem_lo_297};
  wire [95:0]       dataInMem_lo_hi_lo_lo_hi_hi_5 = {dataInMem_hi_428, dataInMem_lo_300, dataInMem_hi_427, dataInMem_lo_299};
  wire [191:0]      dataInMem_lo_hi_lo_lo_hi_5 = {dataInMem_lo_hi_lo_lo_hi_hi_5, dataInMem_lo_hi_lo_lo_hi_lo_5};
  wire [383:0]      dataInMem_lo_hi_lo_lo_5 = {dataInMem_lo_hi_lo_lo_hi_5, dataInMem_lo_hi_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_lo_hi_lo_lo_5 = {dataInMem_hi_430, dataInMem_lo_302, dataInMem_hi_429, dataInMem_lo_301};
  wire [95:0]       dataInMem_lo_hi_lo_hi_lo_hi_5 = {dataInMem_hi_432, dataInMem_lo_304, dataInMem_hi_431, dataInMem_lo_303};
  wire [191:0]      dataInMem_lo_hi_lo_hi_lo_5 = {dataInMem_lo_hi_lo_hi_lo_hi_5, dataInMem_lo_hi_lo_hi_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_lo_hi_hi_lo_5 = {dataInMem_hi_434, dataInMem_lo_306, dataInMem_hi_433, dataInMem_lo_305};
  wire [95:0]       dataInMem_lo_hi_lo_hi_hi_hi_5 = {dataInMem_hi_436, dataInMem_lo_308, dataInMem_hi_435, dataInMem_lo_307};
  wire [191:0]      dataInMem_lo_hi_lo_hi_hi_5 = {dataInMem_lo_hi_lo_hi_hi_hi_5, dataInMem_lo_hi_lo_hi_hi_lo_5};
  wire [383:0]      dataInMem_lo_hi_lo_hi_5 = {dataInMem_lo_hi_lo_hi_hi_5, dataInMem_lo_hi_lo_hi_lo_5};
  wire [767:0]      dataInMem_lo_hi_lo_5 = {dataInMem_lo_hi_lo_hi_5, dataInMem_lo_hi_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_hi_lo_lo_lo_5 = {dataInMem_hi_438, dataInMem_lo_310, dataInMem_hi_437, dataInMem_lo_309};
  wire [95:0]       dataInMem_lo_hi_hi_lo_lo_hi_5 = {dataInMem_hi_440, dataInMem_lo_312, dataInMem_hi_439, dataInMem_lo_311};
  wire [191:0]      dataInMem_lo_hi_hi_lo_lo_5 = {dataInMem_lo_hi_hi_lo_lo_hi_5, dataInMem_lo_hi_hi_lo_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_hi_lo_hi_lo_5 = {dataInMem_hi_442, dataInMem_lo_314, dataInMem_hi_441, dataInMem_lo_313};
  wire [95:0]       dataInMem_lo_hi_hi_lo_hi_hi_5 = {dataInMem_hi_444, dataInMem_lo_316, dataInMem_hi_443, dataInMem_lo_315};
  wire [191:0]      dataInMem_lo_hi_hi_lo_hi_5 = {dataInMem_lo_hi_hi_lo_hi_hi_5, dataInMem_lo_hi_hi_lo_hi_lo_5};
  wire [383:0]      dataInMem_lo_hi_hi_lo_5 = {dataInMem_lo_hi_hi_lo_hi_5, dataInMem_lo_hi_hi_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_hi_hi_lo_lo_5 = {dataInMem_hi_446, dataInMem_lo_318, dataInMem_hi_445, dataInMem_lo_317};
  wire [95:0]       dataInMem_lo_hi_hi_hi_lo_hi_5 = {dataInMem_hi_448, dataInMem_lo_320, dataInMem_hi_447, dataInMem_lo_319};
  wire [191:0]      dataInMem_lo_hi_hi_hi_lo_5 = {dataInMem_lo_hi_hi_hi_lo_hi_5, dataInMem_lo_hi_hi_hi_lo_lo_5};
  wire [95:0]       dataInMem_lo_hi_hi_hi_hi_lo_5 = {dataInMem_hi_450, dataInMem_lo_322, dataInMem_hi_449, dataInMem_lo_321};
  wire [95:0]       dataInMem_lo_hi_hi_hi_hi_hi_5 = {dataInMem_hi_452, dataInMem_lo_324, dataInMem_hi_451, dataInMem_lo_323};
  wire [191:0]      dataInMem_lo_hi_hi_hi_hi_5 = {dataInMem_lo_hi_hi_hi_hi_hi_5, dataInMem_lo_hi_hi_hi_hi_lo_5};
  wire [383:0]      dataInMem_lo_hi_hi_hi_5 = {dataInMem_lo_hi_hi_hi_hi_5, dataInMem_lo_hi_hi_hi_lo_5};
  wire [767:0]      dataInMem_lo_hi_hi_5 = {dataInMem_lo_hi_hi_hi_5, dataInMem_lo_hi_hi_lo_5};
  wire [1535:0]     dataInMem_lo_hi_133 = {dataInMem_lo_hi_hi_5, dataInMem_lo_hi_lo_5};
  wire [3071:0]     dataInMem_lo_389 = {dataInMem_lo_hi_133, dataInMem_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_lo_lo_lo_lo_5 = {dataInMem_hi_454, dataInMem_lo_326, dataInMem_hi_453, dataInMem_lo_325};
  wire [95:0]       dataInMem_hi_lo_lo_lo_lo_hi_5 = {dataInMem_hi_456, dataInMem_lo_328, dataInMem_hi_455, dataInMem_lo_327};
  wire [191:0]      dataInMem_hi_lo_lo_lo_lo_5 = {dataInMem_hi_lo_lo_lo_lo_hi_5, dataInMem_hi_lo_lo_lo_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_lo_lo_hi_lo_5 = {dataInMem_hi_458, dataInMem_lo_330, dataInMem_hi_457, dataInMem_lo_329};
  wire [95:0]       dataInMem_hi_lo_lo_lo_hi_hi_5 = {dataInMem_hi_460, dataInMem_lo_332, dataInMem_hi_459, dataInMem_lo_331};
  wire [191:0]      dataInMem_hi_lo_lo_lo_hi_5 = {dataInMem_hi_lo_lo_lo_hi_hi_5, dataInMem_hi_lo_lo_lo_hi_lo_5};
  wire [383:0]      dataInMem_hi_lo_lo_lo_5 = {dataInMem_hi_lo_lo_lo_hi_5, dataInMem_hi_lo_lo_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_lo_hi_lo_lo_5 = {dataInMem_hi_462, dataInMem_lo_334, dataInMem_hi_461, dataInMem_lo_333};
  wire [95:0]       dataInMem_hi_lo_lo_hi_lo_hi_5 = {dataInMem_hi_464, dataInMem_lo_336, dataInMem_hi_463, dataInMem_lo_335};
  wire [191:0]      dataInMem_hi_lo_lo_hi_lo_5 = {dataInMem_hi_lo_lo_hi_lo_hi_5, dataInMem_hi_lo_lo_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_lo_hi_hi_lo_5 = {dataInMem_hi_466, dataInMem_lo_338, dataInMem_hi_465, dataInMem_lo_337};
  wire [95:0]       dataInMem_hi_lo_lo_hi_hi_hi_5 = {dataInMem_hi_468, dataInMem_lo_340, dataInMem_hi_467, dataInMem_lo_339};
  wire [191:0]      dataInMem_hi_lo_lo_hi_hi_5 = {dataInMem_hi_lo_lo_hi_hi_hi_5, dataInMem_hi_lo_lo_hi_hi_lo_5};
  wire [383:0]      dataInMem_hi_lo_lo_hi_5 = {dataInMem_hi_lo_lo_hi_hi_5, dataInMem_hi_lo_lo_hi_lo_5};
  wire [767:0]      dataInMem_hi_lo_lo_5 = {dataInMem_hi_lo_lo_hi_5, dataInMem_hi_lo_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_hi_lo_lo_lo_5 = {dataInMem_hi_470, dataInMem_lo_342, dataInMem_hi_469, dataInMem_lo_341};
  wire [95:0]       dataInMem_hi_lo_hi_lo_lo_hi_5 = {dataInMem_hi_472, dataInMem_lo_344, dataInMem_hi_471, dataInMem_lo_343};
  wire [191:0]      dataInMem_hi_lo_hi_lo_lo_5 = {dataInMem_hi_lo_hi_lo_lo_hi_5, dataInMem_hi_lo_hi_lo_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_hi_lo_hi_lo_5 = {dataInMem_hi_474, dataInMem_lo_346, dataInMem_hi_473, dataInMem_lo_345};
  wire [95:0]       dataInMem_hi_lo_hi_lo_hi_hi_5 = {dataInMem_hi_476, dataInMem_lo_348, dataInMem_hi_475, dataInMem_lo_347};
  wire [191:0]      dataInMem_hi_lo_hi_lo_hi_5 = {dataInMem_hi_lo_hi_lo_hi_hi_5, dataInMem_hi_lo_hi_lo_hi_lo_5};
  wire [383:0]      dataInMem_hi_lo_hi_lo_5 = {dataInMem_hi_lo_hi_lo_hi_5, dataInMem_hi_lo_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_hi_hi_lo_lo_5 = {dataInMem_hi_478, dataInMem_lo_350, dataInMem_hi_477, dataInMem_lo_349};
  wire [95:0]       dataInMem_hi_lo_hi_hi_lo_hi_5 = {dataInMem_hi_480, dataInMem_lo_352, dataInMem_hi_479, dataInMem_lo_351};
  wire [191:0]      dataInMem_hi_lo_hi_hi_lo_5 = {dataInMem_hi_lo_hi_hi_lo_hi_5, dataInMem_hi_lo_hi_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_lo_hi_hi_hi_lo_5 = {dataInMem_hi_482, dataInMem_lo_354, dataInMem_hi_481, dataInMem_lo_353};
  wire [95:0]       dataInMem_hi_lo_hi_hi_hi_hi_5 = {dataInMem_hi_484, dataInMem_lo_356, dataInMem_hi_483, dataInMem_lo_355};
  wire [191:0]      dataInMem_hi_lo_hi_hi_hi_5 = {dataInMem_hi_lo_hi_hi_hi_hi_5, dataInMem_hi_lo_hi_hi_hi_lo_5};
  wire [383:0]      dataInMem_hi_lo_hi_hi_5 = {dataInMem_hi_lo_hi_hi_hi_5, dataInMem_hi_lo_hi_hi_lo_5};
  wire [767:0]      dataInMem_hi_lo_hi_5 = {dataInMem_hi_lo_hi_hi_5, dataInMem_hi_lo_hi_lo_5};
  wire [1535:0]     dataInMem_hi_lo_5 = {dataInMem_hi_lo_hi_5, dataInMem_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_lo_lo_lo_lo_5 = {dataInMem_hi_486, dataInMem_lo_358, dataInMem_hi_485, dataInMem_lo_357};
  wire [95:0]       dataInMem_hi_hi_lo_lo_lo_hi_5 = {dataInMem_hi_488, dataInMem_lo_360, dataInMem_hi_487, dataInMem_lo_359};
  wire [191:0]      dataInMem_hi_hi_lo_lo_lo_5 = {dataInMem_hi_hi_lo_lo_lo_hi_5, dataInMem_hi_hi_lo_lo_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_lo_lo_hi_lo_5 = {dataInMem_hi_490, dataInMem_lo_362, dataInMem_hi_489, dataInMem_lo_361};
  wire [95:0]       dataInMem_hi_hi_lo_lo_hi_hi_5 = {dataInMem_hi_492, dataInMem_lo_364, dataInMem_hi_491, dataInMem_lo_363};
  wire [191:0]      dataInMem_hi_hi_lo_lo_hi_5 = {dataInMem_hi_hi_lo_lo_hi_hi_5, dataInMem_hi_hi_lo_lo_hi_lo_5};
  wire [383:0]      dataInMem_hi_hi_lo_lo_5 = {dataInMem_hi_hi_lo_lo_hi_5, dataInMem_hi_hi_lo_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_lo_hi_lo_lo_5 = {dataInMem_hi_494, dataInMem_lo_366, dataInMem_hi_493, dataInMem_lo_365};
  wire [95:0]       dataInMem_hi_hi_lo_hi_lo_hi_5 = {dataInMem_hi_496, dataInMem_lo_368, dataInMem_hi_495, dataInMem_lo_367};
  wire [191:0]      dataInMem_hi_hi_lo_hi_lo_5 = {dataInMem_hi_hi_lo_hi_lo_hi_5, dataInMem_hi_hi_lo_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_lo_hi_hi_lo_5 = {dataInMem_hi_498, dataInMem_lo_370, dataInMem_hi_497, dataInMem_lo_369};
  wire [95:0]       dataInMem_hi_hi_lo_hi_hi_hi_5 = {dataInMem_hi_500, dataInMem_lo_372, dataInMem_hi_499, dataInMem_lo_371};
  wire [191:0]      dataInMem_hi_hi_lo_hi_hi_5 = {dataInMem_hi_hi_lo_hi_hi_hi_5, dataInMem_hi_hi_lo_hi_hi_lo_5};
  wire [383:0]      dataInMem_hi_hi_lo_hi_5 = {dataInMem_hi_hi_lo_hi_hi_5, dataInMem_hi_hi_lo_hi_lo_5};
  wire [767:0]      dataInMem_hi_hi_lo_5 = {dataInMem_hi_hi_lo_hi_5, dataInMem_hi_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_hi_lo_lo_lo_5 = {dataInMem_hi_502, dataInMem_lo_374, dataInMem_hi_501, dataInMem_lo_373};
  wire [95:0]       dataInMem_hi_hi_hi_lo_lo_hi_5 = {dataInMem_hi_504, dataInMem_lo_376, dataInMem_hi_503, dataInMem_lo_375};
  wire [191:0]      dataInMem_hi_hi_hi_lo_lo_5 = {dataInMem_hi_hi_hi_lo_lo_hi_5, dataInMem_hi_hi_hi_lo_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_hi_lo_hi_lo_5 = {dataInMem_hi_506, dataInMem_lo_378, dataInMem_hi_505, dataInMem_lo_377};
  wire [95:0]       dataInMem_hi_hi_hi_lo_hi_hi_5 = {dataInMem_hi_508, dataInMem_lo_380, dataInMem_hi_507, dataInMem_lo_379};
  wire [191:0]      dataInMem_hi_hi_hi_lo_hi_5 = {dataInMem_hi_hi_hi_lo_hi_hi_5, dataInMem_hi_hi_hi_lo_hi_lo_5};
  wire [383:0]      dataInMem_hi_hi_hi_lo_5 = {dataInMem_hi_hi_hi_lo_hi_5, dataInMem_hi_hi_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_hi_hi_lo_lo_5 = {dataInMem_hi_510, dataInMem_lo_382, dataInMem_hi_509, dataInMem_lo_381};
  wire [95:0]       dataInMem_hi_hi_hi_hi_lo_hi_5 = {dataInMem_hi_512, dataInMem_lo_384, dataInMem_hi_511, dataInMem_lo_383};
  wire [191:0]      dataInMem_hi_hi_hi_hi_lo_5 = {dataInMem_hi_hi_hi_hi_lo_hi_5, dataInMem_hi_hi_hi_hi_lo_lo_5};
  wire [95:0]       dataInMem_hi_hi_hi_hi_hi_lo_5 = {dataInMem_hi_514, dataInMem_lo_386, dataInMem_hi_513, dataInMem_lo_385};
  wire [95:0]       dataInMem_hi_hi_hi_hi_hi_hi_5 = {dataInMem_hi_516, dataInMem_lo_388, dataInMem_hi_515, dataInMem_lo_387};
  wire [191:0]      dataInMem_hi_hi_hi_hi_hi_5 = {dataInMem_hi_hi_hi_hi_hi_hi_5, dataInMem_hi_hi_hi_hi_hi_lo_5};
  wire [383:0]      dataInMem_hi_hi_hi_hi_5 = {dataInMem_hi_hi_hi_hi_hi_5, dataInMem_hi_hi_hi_hi_lo_5};
  wire [767:0]      dataInMem_hi_hi_hi_5 = {dataInMem_hi_hi_hi_hi_5, dataInMem_hi_hi_hi_lo_5};
  wire [1535:0]     dataInMem_hi_hi_261 = {dataInMem_hi_hi_hi_5, dataInMem_hi_hi_lo_5};
  wire [3071:0]     dataInMem_hi_517 = {dataInMem_hi_hi_261, dataInMem_hi_lo_5};
  wire [6143:0]     dataInMem_5 = {dataInMem_hi_517, dataInMem_lo_389};
  wire [1023:0]     regroupCacheLine_5_0 = dataInMem_5[1023:0];
  wire [1023:0]     regroupCacheLine_5_1 = dataInMem_5[2047:1024];
  wire [1023:0]     regroupCacheLine_5_2 = dataInMem_5[3071:2048];
  wire [1023:0]     regroupCacheLine_5_3 = dataInMem_5[4095:3072];
  wire [1023:0]     regroupCacheLine_5_4 = dataInMem_5[5119:4096];
  wire [1023:0]     regroupCacheLine_5_5 = dataInMem_5[6143:5120];
  wire [1023:0]     res_40 = regroupCacheLine_5_0;
  wire [1023:0]     res_41 = regroupCacheLine_5_1;
  wire [1023:0]     res_42 = regroupCacheLine_5_2;
  wire [1023:0]     res_43 = regroupCacheLine_5_3;
  wire [1023:0]     res_44 = regroupCacheLine_5_4;
  wire [1023:0]     res_45 = regroupCacheLine_5_5;
  wire [2047:0]     lo_lo_5 = {res_41, res_40};
  wire [2047:0]     lo_hi_5 = {res_43, res_42};
  wire [4095:0]     lo_5 = {lo_hi_5, lo_lo_5};
  wire [2047:0]     hi_lo_5 = {res_45, res_44};
  wire [4095:0]     hi_5 = {2048'h0, hi_lo_5};
  wire [8191:0]     regroupLoadData_0_5 = {hi_5, lo_5};
  wire [23:0]       dataInMem_lo_390 = {dataInMem_lo_hi_134, dataRegroupBySew_0_0};
  wire [15:0]       dataInMem_hi_hi_262 = {dataRegroupBySew_6_0, dataRegroupBySew_5_0};
  wire [31:0]       dataInMem_hi_518 = {dataInMem_hi_hi_262, dataInMem_hi_lo_6};
  wire [23:0]       dataInMem_lo_391 = {dataInMem_lo_hi_135, dataRegroupBySew_0_1};
  wire [15:0]       dataInMem_hi_hi_263 = {dataRegroupBySew_6_1, dataRegroupBySew_5_1};
  wire [31:0]       dataInMem_hi_519 = {dataInMem_hi_hi_263, dataInMem_hi_lo_7};
  wire [23:0]       dataInMem_lo_392 = {dataInMem_lo_hi_136, dataRegroupBySew_0_2};
  wire [15:0]       dataInMem_hi_hi_264 = {dataRegroupBySew_6_2, dataRegroupBySew_5_2};
  wire [31:0]       dataInMem_hi_520 = {dataInMem_hi_hi_264, dataInMem_hi_lo_8};
  wire [23:0]       dataInMem_lo_393 = {dataInMem_lo_hi_137, dataRegroupBySew_0_3};
  wire [15:0]       dataInMem_hi_hi_265 = {dataRegroupBySew_6_3, dataRegroupBySew_5_3};
  wire [31:0]       dataInMem_hi_521 = {dataInMem_hi_hi_265, dataInMem_hi_lo_9};
  wire [23:0]       dataInMem_lo_394 = {dataInMem_lo_hi_138, dataRegroupBySew_0_4};
  wire [15:0]       dataInMem_hi_hi_266 = {dataRegroupBySew_6_4, dataRegroupBySew_5_4};
  wire [31:0]       dataInMem_hi_522 = {dataInMem_hi_hi_266, dataInMem_hi_lo_10};
  wire [23:0]       dataInMem_lo_395 = {dataInMem_lo_hi_139, dataRegroupBySew_0_5};
  wire [15:0]       dataInMem_hi_hi_267 = {dataRegroupBySew_6_5, dataRegroupBySew_5_5};
  wire [31:0]       dataInMem_hi_523 = {dataInMem_hi_hi_267, dataInMem_hi_lo_11};
  wire [23:0]       dataInMem_lo_396 = {dataInMem_lo_hi_140, dataRegroupBySew_0_6};
  wire [15:0]       dataInMem_hi_hi_268 = {dataRegroupBySew_6_6, dataRegroupBySew_5_6};
  wire [31:0]       dataInMem_hi_524 = {dataInMem_hi_hi_268, dataInMem_hi_lo_12};
  wire [23:0]       dataInMem_lo_397 = {dataInMem_lo_hi_141, dataRegroupBySew_0_7};
  wire [15:0]       dataInMem_hi_hi_269 = {dataRegroupBySew_6_7, dataRegroupBySew_5_7};
  wire [31:0]       dataInMem_hi_525 = {dataInMem_hi_hi_269, dataInMem_hi_lo_13};
  wire [23:0]       dataInMem_lo_398 = {dataInMem_lo_hi_142, dataRegroupBySew_0_8};
  wire [15:0]       dataInMem_hi_hi_270 = {dataRegroupBySew_6_8, dataRegroupBySew_5_8};
  wire [31:0]       dataInMem_hi_526 = {dataInMem_hi_hi_270, dataInMem_hi_lo_14};
  wire [23:0]       dataInMem_lo_399 = {dataInMem_lo_hi_143, dataRegroupBySew_0_9};
  wire [15:0]       dataInMem_hi_hi_271 = {dataRegroupBySew_6_9, dataRegroupBySew_5_9};
  wire [31:0]       dataInMem_hi_527 = {dataInMem_hi_hi_271, dataInMem_hi_lo_15};
  wire [23:0]       dataInMem_lo_400 = {dataInMem_lo_hi_144, dataRegroupBySew_0_10};
  wire [15:0]       dataInMem_hi_hi_272 = {dataRegroupBySew_6_10, dataRegroupBySew_5_10};
  wire [31:0]       dataInMem_hi_528 = {dataInMem_hi_hi_272, dataInMem_hi_lo_16};
  wire [23:0]       dataInMem_lo_401 = {dataInMem_lo_hi_145, dataRegroupBySew_0_11};
  wire [15:0]       dataInMem_hi_hi_273 = {dataRegroupBySew_6_11, dataRegroupBySew_5_11};
  wire [31:0]       dataInMem_hi_529 = {dataInMem_hi_hi_273, dataInMem_hi_lo_17};
  wire [23:0]       dataInMem_lo_402 = {dataInMem_lo_hi_146, dataRegroupBySew_0_12};
  wire [15:0]       dataInMem_hi_hi_274 = {dataRegroupBySew_6_12, dataRegroupBySew_5_12};
  wire [31:0]       dataInMem_hi_530 = {dataInMem_hi_hi_274, dataInMem_hi_lo_18};
  wire [23:0]       dataInMem_lo_403 = {dataInMem_lo_hi_147, dataRegroupBySew_0_13};
  wire [15:0]       dataInMem_hi_hi_275 = {dataRegroupBySew_6_13, dataRegroupBySew_5_13};
  wire [31:0]       dataInMem_hi_531 = {dataInMem_hi_hi_275, dataInMem_hi_lo_19};
  wire [23:0]       dataInMem_lo_404 = {dataInMem_lo_hi_148, dataRegroupBySew_0_14};
  wire [15:0]       dataInMem_hi_hi_276 = {dataRegroupBySew_6_14, dataRegroupBySew_5_14};
  wire [31:0]       dataInMem_hi_532 = {dataInMem_hi_hi_276, dataInMem_hi_lo_20};
  wire [23:0]       dataInMem_lo_405 = {dataInMem_lo_hi_149, dataRegroupBySew_0_15};
  wire [15:0]       dataInMem_hi_hi_277 = {dataRegroupBySew_6_15, dataRegroupBySew_5_15};
  wire [31:0]       dataInMem_hi_533 = {dataInMem_hi_hi_277, dataInMem_hi_lo_21};
  wire [23:0]       dataInMem_lo_406 = {dataInMem_lo_hi_150, dataRegroupBySew_0_16};
  wire [15:0]       dataInMem_hi_hi_278 = {dataRegroupBySew_6_16, dataRegroupBySew_5_16};
  wire [31:0]       dataInMem_hi_534 = {dataInMem_hi_hi_278, dataInMem_hi_lo_22};
  wire [23:0]       dataInMem_lo_407 = {dataInMem_lo_hi_151, dataRegroupBySew_0_17};
  wire [15:0]       dataInMem_hi_hi_279 = {dataRegroupBySew_6_17, dataRegroupBySew_5_17};
  wire [31:0]       dataInMem_hi_535 = {dataInMem_hi_hi_279, dataInMem_hi_lo_23};
  wire [23:0]       dataInMem_lo_408 = {dataInMem_lo_hi_152, dataRegroupBySew_0_18};
  wire [15:0]       dataInMem_hi_hi_280 = {dataRegroupBySew_6_18, dataRegroupBySew_5_18};
  wire [31:0]       dataInMem_hi_536 = {dataInMem_hi_hi_280, dataInMem_hi_lo_24};
  wire [23:0]       dataInMem_lo_409 = {dataInMem_lo_hi_153, dataRegroupBySew_0_19};
  wire [15:0]       dataInMem_hi_hi_281 = {dataRegroupBySew_6_19, dataRegroupBySew_5_19};
  wire [31:0]       dataInMem_hi_537 = {dataInMem_hi_hi_281, dataInMem_hi_lo_25};
  wire [23:0]       dataInMem_lo_410 = {dataInMem_lo_hi_154, dataRegroupBySew_0_20};
  wire [15:0]       dataInMem_hi_hi_282 = {dataRegroupBySew_6_20, dataRegroupBySew_5_20};
  wire [31:0]       dataInMem_hi_538 = {dataInMem_hi_hi_282, dataInMem_hi_lo_26};
  wire [23:0]       dataInMem_lo_411 = {dataInMem_lo_hi_155, dataRegroupBySew_0_21};
  wire [15:0]       dataInMem_hi_hi_283 = {dataRegroupBySew_6_21, dataRegroupBySew_5_21};
  wire [31:0]       dataInMem_hi_539 = {dataInMem_hi_hi_283, dataInMem_hi_lo_27};
  wire [23:0]       dataInMem_lo_412 = {dataInMem_lo_hi_156, dataRegroupBySew_0_22};
  wire [15:0]       dataInMem_hi_hi_284 = {dataRegroupBySew_6_22, dataRegroupBySew_5_22};
  wire [31:0]       dataInMem_hi_540 = {dataInMem_hi_hi_284, dataInMem_hi_lo_28};
  wire [23:0]       dataInMem_lo_413 = {dataInMem_lo_hi_157, dataRegroupBySew_0_23};
  wire [15:0]       dataInMem_hi_hi_285 = {dataRegroupBySew_6_23, dataRegroupBySew_5_23};
  wire [31:0]       dataInMem_hi_541 = {dataInMem_hi_hi_285, dataInMem_hi_lo_29};
  wire [23:0]       dataInMem_lo_414 = {dataInMem_lo_hi_158, dataRegroupBySew_0_24};
  wire [15:0]       dataInMem_hi_hi_286 = {dataRegroupBySew_6_24, dataRegroupBySew_5_24};
  wire [31:0]       dataInMem_hi_542 = {dataInMem_hi_hi_286, dataInMem_hi_lo_30};
  wire [23:0]       dataInMem_lo_415 = {dataInMem_lo_hi_159, dataRegroupBySew_0_25};
  wire [15:0]       dataInMem_hi_hi_287 = {dataRegroupBySew_6_25, dataRegroupBySew_5_25};
  wire [31:0]       dataInMem_hi_543 = {dataInMem_hi_hi_287, dataInMem_hi_lo_31};
  wire [23:0]       dataInMem_lo_416 = {dataInMem_lo_hi_160, dataRegroupBySew_0_26};
  wire [15:0]       dataInMem_hi_hi_288 = {dataRegroupBySew_6_26, dataRegroupBySew_5_26};
  wire [31:0]       dataInMem_hi_544 = {dataInMem_hi_hi_288, dataInMem_hi_lo_32};
  wire [23:0]       dataInMem_lo_417 = {dataInMem_lo_hi_161, dataRegroupBySew_0_27};
  wire [15:0]       dataInMem_hi_hi_289 = {dataRegroupBySew_6_27, dataRegroupBySew_5_27};
  wire [31:0]       dataInMem_hi_545 = {dataInMem_hi_hi_289, dataInMem_hi_lo_33};
  wire [23:0]       dataInMem_lo_418 = {dataInMem_lo_hi_162, dataRegroupBySew_0_28};
  wire [15:0]       dataInMem_hi_hi_290 = {dataRegroupBySew_6_28, dataRegroupBySew_5_28};
  wire [31:0]       dataInMem_hi_546 = {dataInMem_hi_hi_290, dataInMem_hi_lo_34};
  wire [23:0]       dataInMem_lo_419 = {dataInMem_lo_hi_163, dataRegroupBySew_0_29};
  wire [15:0]       dataInMem_hi_hi_291 = {dataRegroupBySew_6_29, dataRegroupBySew_5_29};
  wire [31:0]       dataInMem_hi_547 = {dataInMem_hi_hi_291, dataInMem_hi_lo_35};
  wire [23:0]       dataInMem_lo_420 = {dataInMem_lo_hi_164, dataRegroupBySew_0_30};
  wire [15:0]       dataInMem_hi_hi_292 = {dataRegroupBySew_6_30, dataRegroupBySew_5_30};
  wire [31:0]       dataInMem_hi_548 = {dataInMem_hi_hi_292, dataInMem_hi_lo_36};
  wire [23:0]       dataInMem_lo_421 = {dataInMem_lo_hi_165, dataRegroupBySew_0_31};
  wire [15:0]       dataInMem_hi_hi_293 = {dataRegroupBySew_6_31, dataRegroupBySew_5_31};
  wire [31:0]       dataInMem_hi_549 = {dataInMem_hi_hi_293, dataInMem_hi_lo_37};
  wire [23:0]       dataInMem_lo_422 = {dataInMem_lo_hi_166, dataRegroupBySew_0_32};
  wire [15:0]       dataInMem_hi_hi_294 = {dataRegroupBySew_6_32, dataRegroupBySew_5_32};
  wire [31:0]       dataInMem_hi_550 = {dataInMem_hi_hi_294, dataInMem_hi_lo_38};
  wire [23:0]       dataInMem_lo_423 = {dataInMem_lo_hi_167, dataRegroupBySew_0_33};
  wire [15:0]       dataInMem_hi_hi_295 = {dataRegroupBySew_6_33, dataRegroupBySew_5_33};
  wire [31:0]       dataInMem_hi_551 = {dataInMem_hi_hi_295, dataInMem_hi_lo_39};
  wire [23:0]       dataInMem_lo_424 = {dataInMem_lo_hi_168, dataRegroupBySew_0_34};
  wire [15:0]       dataInMem_hi_hi_296 = {dataRegroupBySew_6_34, dataRegroupBySew_5_34};
  wire [31:0]       dataInMem_hi_552 = {dataInMem_hi_hi_296, dataInMem_hi_lo_40};
  wire [23:0]       dataInMem_lo_425 = {dataInMem_lo_hi_169, dataRegroupBySew_0_35};
  wire [15:0]       dataInMem_hi_hi_297 = {dataRegroupBySew_6_35, dataRegroupBySew_5_35};
  wire [31:0]       dataInMem_hi_553 = {dataInMem_hi_hi_297, dataInMem_hi_lo_41};
  wire [23:0]       dataInMem_lo_426 = {dataInMem_lo_hi_170, dataRegroupBySew_0_36};
  wire [15:0]       dataInMem_hi_hi_298 = {dataRegroupBySew_6_36, dataRegroupBySew_5_36};
  wire [31:0]       dataInMem_hi_554 = {dataInMem_hi_hi_298, dataInMem_hi_lo_42};
  wire [23:0]       dataInMem_lo_427 = {dataInMem_lo_hi_171, dataRegroupBySew_0_37};
  wire [15:0]       dataInMem_hi_hi_299 = {dataRegroupBySew_6_37, dataRegroupBySew_5_37};
  wire [31:0]       dataInMem_hi_555 = {dataInMem_hi_hi_299, dataInMem_hi_lo_43};
  wire [23:0]       dataInMem_lo_428 = {dataInMem_lo_hi_172, dataRegroupBySew_0_38};
  wire [15:0]       dataInMem_hi_hi_300 = {dataRegroupBySew_6_38, dataRegroupBySew_5_38};
  wire [31:0]       dataInMem_hi_556 = {dataInMem_hi_hi_300, dataInMem_hi_lo_44};
  wire [23:0]       dataInMem_lo_429 = {dataInMem_lo_hi_173, dataRegroupBySew_0_39};
  wire [15:0]       dataInMem_hi_hi_301 = {dataRegroupBySew_6_39, dataRegroupBySew_5_39};
  wire [31:0]       dataInMem_hi_557 = {dataInMem_hi_hi_301, dataInMem_hi_lo_45};
  wire [23:0]       dataInMem_lo_430 = {dataInMem_lo_hi_174, dataRegroupBySew_0_40};
  wire [15:0]       dataInMem_hi_hi_302 = {dataRegroupBySew_6_40, dataRegroupBySew_5_40};
  wire [31:0]       dataInMem_hi_558 = {dataInMem_hi_hi_302, dataInMem_hi_lo_46};
  wire [23:0]       dataInMem_lo_431 = {dataInMem_lo_hi_175, dataRegroupBySew_0_41};
  wire [15:0]       dataInMem_hi_hi_303 = {dataRegroupBySew_6_41, dataRegroupBySew_5_41};
  wire [31:0]       dataInMem_hi_559 = {dataInMem_hi_hi_303, dataInMem_hi_lo_47};
  wire [23:0]       dataInMem_lo_432 = {dataInMem_lo_hi_176, dataRegroupBySew_0_42};
  wire [15:0]       dataInMem_hi_hi_304 = {dataRegroupBySew_6_42, dataRegroupBySew_5_42};
  wire [31:0]       dataInMem_hi_560 = {dataInMem_hi_hi_304, dataInMem_hi_lo_48};
  wire [23:0]       dataInMem_lo_433 = {dataInMem_lo_hi_177, dataRegroupBySew_0_43};
  wire [15:0]       dataInMem_hi_hi_305 = {dataRegroupBySew_6_43, dataRegroupBySew_5_43};
  wire [31:0]       dataInMem_hi_561 = {dataInMem_hi_hi_305, dataInMem_hi_lo_49};
  wire [23:0]       dataInMem_lo_434 = {dataInMem_lo_hi_178, dataRegroupBySew_0_44};
  wire [15:0]       dataInMem_hi_hi_306 = {dataRegroupBySew_6_44, dataRegroupBySew_5_44};
  wire [31:0]       dataInMem_hi_562 = {dataInMem_hi_hi_306, dataInMem_hi_lo_50};
  wire [23:0]       dataInMem_lo_435 = {dataInMem_lo_hi_179, dataRegroupBySew_0_45};
  wire [15:0]       dataInMem_hi_hi_307 = {dataRegroupBySew_6_45, dataRegroupBySew_5_45};
  wire [31:0]       dataInMem_hi_563 = {dataInMem_hi_hi_307, dataInMem_hi_lo_51};
  wire [23:0]       dataInMem_lo_436 = {dataInMem_lo_hi_180, dataRegroupBySew_0_46};
  wire [15:0]       dataInMem_hi_hi_308 = {dataRegroupBySew_6_46, dataRegroupBySew_5_46};
  wire [31:0]       dataInMem_hi_564 = {dataInMem_hi_hi_308, dataInMem_hi_lo_52};
  wire [23:0]       dataInMem_lo_437 = {dataInMem_lo_hi_181, dataRegroupBySew_0_47};
  wire [15:0]       dataInMem_hi_hi_309 = {dataRegroupBySew_6_47, dataRegroupBySew_5_47};
  wire [31:0]       dataInMem_hi_565 = {dataInMem_hi_hi_309, dataInMem_hi_lo_53};
  wire [23:0]       dataInMem_lo_438 = {dataInMem_lo_hi_182, dataRegroupBySew_0_48};
  wire [15:0]       dataInMem_hi_hi_310 = {dataRegroupBySew_6_48, dataRegroupBySew_5_48};
  wire [31:0]       dataInMem_hi_566 = {dataInMem_hi_hi_310, dataInMem_hi_lo_54};
  wire [23:0]       dataInMem_lo_439 = {dataInMem_lo_hi_183, dataRegroupBySew_0_49};
  wire [15:0]       dataInMem_hi_hi_311 = {dataRegroupBySew_6_49, dataRegroupBySew_5_49};
  wire [31:0]       dataInMem_hi_567 = {dataInMem_hi_hi_311, dataInMem_hi_lo_55};
  wire [23:0]       dataInMem_lo_440 = {dataInMem_lo_hi_184, dataRegroupBySew_0_50};
  wire [15:0]       dataInMem_hi_hi_312 = {dataRegroupBySew_6_50, dataRegroupBySew_5_50};
  wire [31:0]       dataInMem_hi_568 = {dataInMem_hi_hi_312, dataInMem_hi_lo_56};
  wire [23:0]       dataInMem_lo_441 = {dataInMem_lo_hi_185, dataRegroupBySew_0_51};
  wire [15:0]       dataInMem_hi_hi_313 = {dataRegroupBySew_6_51, dataRegroupBySew_5_51};
  wire [31:0]       dataInMem_hi_569 = {dataInMem_hi_hi_313, dataInMem_hi_lo_57};
  wire [23:0]       dataInMem_lo_442 = {dataInMem_lo_hi_186, dataRegroupBySew_0_52};
  wire [15:0]       dataInMem_hi_hi_314 = {dataRegroupBySew_6_52, dataRegroupBySew_5_52};
  wire [31:0]       dataInMem_hi_570 = {dataInMem_hi_hi_314, dataInMem_hi_lo_58};
  wire [23:0]       dataInMem_lo_443 = {dataInMem_lo_hi_187, dataRegroupBySew_0_53};
  wire [15:0]       dataInMem_hi_hi_315 = {dataRegroupBySew_6_53, dataRegroupBySew_5_53};
  wire [31:0]       dataInMem_hi_571 = {dataInMem_hi_hi_315, dataInMem_hi_lo_59};
  wire [23:0]       dataInMem_lo_444 = {dataInMem_lo_hi_188, dataRegroupBySew_0_54};
  wire [15:0]       dataInMem_hi_hi_316 = {dataRegroupBySew_6_54, dataRegroupBySew_5_54};
  wire [31:0]       dataInMem_hi_572 = {dataInMem_hi_hi_316, dataInMem_hi_lo_60};
  wire [23:0]       dataInMem_lo_445 = {dataInMem_lo_hi_189, dataRegroupBySew_0_55};
  wire [15:0]       dataInMem_hi_hi_317 = {dataRegroupBySew_6_55, dataRegroupBySew_5_55};
  wire [31:0]       dataInMem_hi_573 = {dataInMem_hi_hi_317, dataInMem_hi_lo_61};
  wire [23:0]       dataInMem_lo_446 = {dataInMem_lo_hi_190, dataRegroupBySew_0_56};
  wire [15:0]       dataInMem_hi_hi_318 = {dataRegroupBySew_6_56, dataRegroupBySew_5_56};
  wire [31:0]       dataInMem_hi_574 = {dataInMem_hi_hi_318, dataInMem_hi_lo_62};
  wire [23:0]       dataInMem_lo_447 = {dataInMem_lo_hi_191, dataRegroupBySew_0_57};
  wire [15:0]       dataInMem_hi_hi_319 = {dataRegroupBySew_6_57, dataRegroupBySew_5_57};
  wire [31:0]       dataInMem_hi_575 = {dataInMem_hi_hi_319, dataInMem_hi_lo_63};
  wire [23:0]       dataInMem_lo_448 = {dataInMem_lo_hi_192, dataRegroupBySew_0_58};
  wire [15:0]       dataInMem_hi_hi_320 = {dataRegroupBySew_6_58, dataRegroupBySew_5_58};
  wire [31:0]       dataInMem_hi_576 = {dataInMem_hi_hi_320, dataInMem_hi_lo_64};
  wire [23:0]       dataInMem_lo_449 = {dataInMem_lo_hi_193, dataRegroupBySew_0_59};
  wire [15:0]       dataInMem_hi_hi_321 = {dataRegroupBySew_6_59, dataRegroupBySew_5_59};
  wire [31:0]       dataInMem_hi_577 = {dataInMem_hi_hi_321, dataInMem_hi_lo_65};
  wire [23:0]       dataInMem_lo_450 = {dataInMem_lo_hi_194, dataRegroupBySew_0_60};
  wire [15:0]       dataInMem_hi_hi_322 = {dataRegroupBySew_6_60, dataRegroupBySew_5_60};
  wire [31:0]       dataInMem_hi_578 = {dataInMem_hi_hi_322, dataInMem_hi_lo_66};
  wire [23:0]       dataInMem_lo_451 = {dataInMem_lo_hi_195, dataRegroupBySew_0_61};
  wire [15:0]       dataInMem_hi_hi_323 = {dataRegroupBySew_6_61, dataRegroupBySew_5_61};
  wire [31:0]       dataInMem_hi_579 = {dataInMem_hi_hi_323, dataInMem_hi_lo_67};
  wire [23:0]       dataInMem_lo_452 = {dataInMem_lo_hi_196, dataRegroupBySew_0_62};
  wire [15:0]       dataInMem_hi_hi_324 = {dataRegroupBySew_6_62, dataRegroupBySew_5_62};
  wire [31:0]       dataInMem_hi_580 = {dataInMem_hi_hi_324, dataInMem_hi_lo_68};
  wire [23:0]       dataInMem_lo_453 = {dataInMem_lo_hi_197, dataRegroupBySew_0_63};
  wire [15:0]       dataInMem_hi_hi_325 = {dataRegroupBySew_6_63, dataRegroupBySew_5_63};
  wire [31:0]       dataInMem_hi_581 = {dataInMem_hi_hi_325, dataInMem_hi_lo_69};
  wire [23:0]       dataInMem_lo_454 = {dataInMem_lo_hi_198, dataRegroupBySew_0_64};
  wire [15:0]       dataInMem_hi_hi_326 = {dataRegroupBySew_6_64, dataRegroupBySew_5_64};
  wire [31:0]       dataInMem_hi_582 = {dataInMem_hi_hi_326, dataInMem_hi_lo_70};
  wire [23:0]       dataInMem_lo_455 = {dataInMem_lo_hi_199, dataRegroupBySew_0_65};
  wire [15:0]       dataInMem_hi_hi_327 = {dataRegroupBySew_6_65, dataRegroupBySew_5_65};
  wire [31:0]       dataInMem_hi_583 = {dataInMem_hi_hi_327, dataInMem_hi_lo_71};
  wire [23:0]       dataInMem_lo_456 = {dataInMem_lo_hi_200, dataRegroupBySew_0_66};
  wire [15:0]       dataInMem_hi_hi_328 = {dataRegroupBySew_6_66, dataRegroupBySew_5_66};
  wire [31:0]       dataInMem_hi_584 = {dataInMem_hi_hi_328, dataInMem_hi_lo_72};
  wire [23:0]       dataInMem_lo_457 = {dataInMem_lo_hi_201, dataRegroupBySew_0_67};
  wire [15:0]       dataInMem_hi_hi_329 = {dataRegroupBySew_6_67, dataRegroupBySew_5_67};
  wire [31:0]       dataInMem_hi_585 = {dataInMem_hi_hi_329, dataInMem_hi_lo_73};
  wire [23:0]       dataInMem_lo_458 = {dataInMem_lo_hi_202, dataRegroupBySew_0_68};
  wire [15:0]       dataInMem_hi_hi_330 = {dataRegroupBySew_6_68, dataRegroupBySew_5_68};
  wire [31:0]       dataInMem_hi_586 = {dataInMem_hi_hi_330, dataInMem_hi_lo_74};
  wire [23:0]       dataInMem_lo_459 = {dataInMem_lo_hi_203, dataRegroupBySew_0_69};
  wire [15:0]       dataInMem_hi_hi_331 = {dataRegroupBySew_6_69, dataRegroupBySew_5_69};
  wire [31:0]       dataInMem_hi_587 = {dataInMem_hi_hi_331, dataInMem_hi_lo_75};
  wire [23:0]       dataInMem_lo_460 = {dataInMem_lo_hi_204, dataRegroupBySew_0_70};
  wire [15:0]       dataInMem_hi_hi_332 = {dataRegroupBySew_6_70, dataRegroupBySew_5_70};
  wire [31:0]       dataInMem_hi_588 = {dataInMem_hi_hi_332, dataInMem_hi_lo_76};
  wire [23:0]       dataInMem_lo_461 = {dataInMem_lo_hi_205, dataRegroupBySew_0_71};
  wire [15:0]       dataInMem_hi_hi_333 = {dataRegroupBySew_6_71, dataRegroupBySew_5_71};
  wire [31:0]       dataInMem_hi_589 = {dataInMem_hi_hi_333, dataInMem_hi_lo_77};
  wire [23:0]       dataInMem_lo_462 = {dataInMem_lo_hi_206, dataRegroupBySew_0_72};
  wire [15:0]       dataInMem_hi_hi_334 = {dataRegroupBySew_6_72, dataRegroupBySew_5_72};
  wire [31:0]       dataInMem_hi_590 = {dataInMem_hi_hi_334, dataInMem_hi_lo_78};
  wire [23:0]       dataInMem_lo_463 = {dataInMem_lo_hi_207, dataRegroupBySew_0_73};
  wire [15:0]       dataInMem_hi_hi_335 = {dataRegroupBySew_6_73, dataRegroupBySew_5_73};
  wire [31:0]       dataInMem_hi_591 = {dataInMem_hi_hi_335, dataInMem_hi_lo_79};
  wire [23:0]       dataInMem_lo_464 = {dataInMem_lo_hi_208, dataRegroupBySew_0_74};
  wire [15:0]       dataInMem_hi_hi_336 = {dataRegroupBySew_6_74, dataRegroupBySew_5_74};
  wire [31:0]       dataInMem_hi_592 = {dataInMem_hi_hi_336, dataInMem_hi_lo_80};
  wire [23:0]       dataInMem_lo_465 = {dataInMem_lo_hi_209, dataRegroupBySew_0_75};
  wire [15:0]       dataInMem_hi_hi_337 = {dataRegroupBySew_6_75, dataRegroupBySew_5_75};
  wire [31:0]       dataInMem_hi_593 = {dataInMem_hi_hi_337, dataInMem_hi_lo_81};
  wire [23:0]       dataInMem_lo_466 = {dataInMem_lo_hi_210, dataRegroupBySew_0_76};
  wire [15:0]       dataInMem_hi_hi_338 = {dataRegroupBySew_6_76, dataRegroupBySew_5_76};
  wire [31:0]       dataInMem_hi_594 = {dataInMem_hi_hi_338, dataInMem_hi_lo_82};
  wire [23:0]       dataInMem_lo_467 = {dataInMem_lo_hi_211, dataRegroupBySew_0_77};
  wire [15:0]       dataInMem_hi_hi_339 = {dataRegroupBySew_6_77, dataRegroupBySew_5_77};
  wire [31:0]       dataInMem_hi_595 = {dataInMem_hi_hi_339, dataInMem_hi_lo_83};
  wire [23:0]       dataInMem_lo_468 = {dataInMem_lo_hi_212, dataRegroupBySew_0_78};
  wire [15:0]       dataInMem_hi_hi_340 = {dataRegroupBySew_6_78, dataRegroupBySew_5_78};
  wire [31:0]       dataInMem_hi_596 = {dataInMem_hi_hi_340, dataInMem_hi_lo_84};
  wire [23:0]       dataInMem_lo_469 = {dataInMem_lo_hi_213, dataRegroupBySew_0_79};
  wire [15:0]       dataInMem_hi_hi_341 = {dataRegroupBySew_6_79, dataRegroupBySew_5_79};
  wire [31:0]       dataInMem_hi_597 = {dataInMem_hi_hi_341, dataInMem_hi_lo_85};
  wire [23:0]       dataInMem_lo_470 = {dataInMem_lo_hi_214, dataRegroupBySew_0_80};
  wire [15:0]       dataInMem_hi_hi_342 = {dataRegroupBySew_6_80, dataRegroupBySew_5_80};
  wire [31:0]       dataInMem_hi_598 = {dataInMem_hi_hi_342, dataInMem_hi_lo_86};
  wire [23:0]       dataInMem_lo_471 = {dataInMem_lo_hi_215, dataRegroupBySew_0_81};
  wire [15:0]       dataInMem_hi_hi_343 = {dataRegroupBySew_6_81, dataRegroupBySew_5_81};
  wire [31:0]       dataInMem_hi_599 = {dataInMem_hi_hi_343, dataInMem_hi_lo_87};
  wire [23:0]       dataInMem_lo_472 = {dataInMem_lo_hi_216, dataRegroupBySew_0_82};
  wire [15:0]       dataInMem_hi_hi_344 = {dataRegroupBySew_6_82, dataRegroupBySew_5_82};
  wire [31:0]       dataInMem_hi_600 = {dataInMem_hi_hi_344, dataInMem_hi_lo_88};
  wire [23:0]       dataInMem_lo_473 = {dataInMem_lo_hi_217, dataRegroupBySew_0_83};
  wire [15:0]       dataInMem_hi_hi_345 = {dataRegroupBySew_6_83, dataRegroupBySew_5_83};
  wire [31:0]       dataInMem_hi_601 = {dataInMem_hi_hi_345, dataInMem_hi_lo_89};
  wire [23:0]       dataInMem_lo_474 = {dataInMem_lo_hi_218, dataRegroupBySew_0_84};
  wire [15:0]       dataInMem_hi_hi_346 = {dataRegroupBySew_6_84, dataRegroupBySew_5_84};
  wire [31:0]       dataInMem_hi_602 = {dataInMem_hi_hi_346, dataInMem_hi_lo_90};
  wire [23:0]       dataInMem_lo_475 = {dataInMem_lo_hi_219, dataRegroupBySew_0_85};
  wire [15:0]       dataInMem_hi_hi_347 = {dataRegroupBySew_6_85, dataRegroupBySew_5_85};
  wire [31:0]       dataInMem_hi_603 = {dataInMem_hi_hi_347, dataInMem_hi_lo_91};
  wire [23:0]       dataInMem_lo_476 = {dataInMem_lo_hi_220, dataRegroupBySew_0_86};
  wire [15:0]       dataInMem_hi_hi_348 = {dataRegroupBySew_6_86, dataRegroupBySew_5_86};
  wire [31:0]       dataInMem_hi_604 = {dataInMem_hi_hi_348, dataInMem_hi_lo_92};
  wire [23:0]       dataInMem_lo_477 = {dataInMem_lo_hi_221, dataRegroupBySew_0_87};
  wire [15:0]       dataInMem_hi_hi_349 = {dataRegroupBySew_6_87, dataRegroupBySew_5_87};
  wire [31:0]       dataInMem_hi_605 = {dataInMem_hi_hi_349, dataInMem_hi_lo_93};
  wire [23:0]       dataInMem_lo_478 = {dataInMem_lo_hi_222, dataRegroupBySew_0_88};
  wire [15:0]       dataInMem_hi_hi_350 = {dataRegroupBySew_6_88, dataRegroupBySew_5_88};
  wire [31:0]       dataInMem_hi_606 = {dataInMem_hi_hi_350, dataInMem_hi_lo_94};
  wire [23:0]       dataInMem_lo_479 = {dataInMem_lo_hi_223, dataRegroupBySew_0_89};
  wire [15:0]       dataInMem_hi_hi_351 = {dataRegroupBySew_6_89, dataRegroupBySew_5_89};
  wire [31:0]       dataInMem_hi_607 = {dataInMem_hi_hi_351, dataInMem_hi_lo_95};
  wire [23:0]       dataInMem_lo_480 = {dataInMem_lo_hi_224, dataRegroupBySew_0_90};
  wire [15:0]       dataInMem_hi_hi_352 = {dataRegroupBySew_6_90, dataRegroupBySew_5_90};
  wire [31:0]       dataInMem_hi_608 = {dataInMem_hi_hi_352, dataInMem_hi_lo_96};
  wire [23:0]       dataInMem_lo_481 = {dataInMem_lo_hi_225, dataRegroupBySew_0_91};
  wire [15:0]       dataInMem_hi_hi_353 = {dataRegroupBySew_6_91, dataRegroupBySew_5_91};
  wire [31:0]       dataInMem_hi_609 = {dataInMem_hi_hi_353, dataInMem_hi_lo_97};
  wire [23:0]       dataInMem_lo_482 = {dataInMem_lo_hi_226, dataRegroupBySew_0_92};
  wire [15:0]       dataInMem_hi_hi_354 = {dataRegroupBySew_6_92, dataRegroupBySew_5_92};
  wire [31:0]       dataInMem_hi_610 = {dataInMem_hi_hi_354, dataInMem_hi_lo_98};
  wire [23:0]       dataInMem_lo_483 = {dataInMem_lo_hi_227, dataRegroupBySew_0_93};
  wire [15:0]       dataInMem_hi_hi_355 = {dataRegroupBySew_6_93, dataRegroupBySew_5_93};
  wire [31:0]       dataInMem_hi_611 = {dataInMem_hi_hi_355, dataInMem_hi_lo_99};
  wire [23:0]       dataInMem_lo_484 = {dataInMem_lo_hi_228, dataRegroupBySew_0_94};
  wire [15:0]       dataInMem_hi_hi_356 = {dataRegroupBySew_6_94, dataRegroupBySew_5_94};
  wire [31:0]       dataInMem_hi_612 = {dataInMem_hi_hi_356, dataInMem_hi_lo_100};
  wire [23:0]       dataInMem_lo_485 = {dataInMem_lo_hi_229, dataRegroupBySew_0_95};
  wire [15:0]       dataInMem_hi_hi_357 = {dataRegroupBySew_6_95, dataRegroupBySew_5_95};
  wire [31:0]       dataInMem_hi_613 = {dataInMem_hi_hi_357, dataInMem_hi_lo_101};
  wire [23:0]       dataInMem_lo_486 = {dataInMem_lo_hi_230, dataRegroupBySew_0_96};
  wire [15:0]       dataInMem_hi_hi_358 = {dataRegroupBySew_6_96, dataRegroupBySew_5_96};
  wire [31:0]       dataInMem_hi_614 = {dataInMem_hi_hi_358, dataInMem_hi_lo_102};
  wire [23:0]       dataInMem_lo_487 = {dataInMem_lo_hi_231, dataRegroupBySew_0_97};
  wire [15:0]       dataInMem_hi_hi_359 = {dataRegroupBySew_6_97, dataRegroupBySew_5_97};
  wire [31:0]       dataInMem_hi_615 = {dataInMem_hi_hi_359, dataInMem_hi_lo_103};
  wire [23:0]       dataInMem_lo_488 = {dataInMem_lo_hi_232, dataRegroupBySew_0_98};
  wire [15:0]       dataInMem_hi_hi_360 = {dataRegroupBySew_6_98, dataRegroupBySew_5_98};
  wire [31:0]       dataInMem_hi_616 = {dataInMem_hi_hi_360, dataInMem_hi_lo_104};
  wire [23:0]       dataInMem_lo_489 = {dataInMem_lo_hi_233, dataRegroupBySew_0_99};
  wire [15:0]       dataInMem_hi_hi_361 = {dataRegroupBySew_6_99, dataRegroupBySew_5_99};
  wire [31:0]       dataInMem_hi_617 = {dataInMem_hi_hi_361, dataInMem_hi_lo_105};
  wire [23:0]       dataInMem_lo_490 = {dataInMem_lo_hi_234, dataRegroupBySew_0_100};
  wire [15:0]       dataInMem_hi_hi_362 = {dataRegroupBySew_6_100, dataRegroupBySew_5_100};
  wire [31:0]       dataInMem_hi_618 = {dataInMem_hi_hi_362, dataInMem_hi_lo_106};
  wire [23:0]       dataInMem_lo_491 = {dataInMem_lo_hi_235, dataRegroupBySew_0_101};
  wire [15:0]       dataInMem_hi_hi_363 = {dataRegroupBySew_6_101, dataRegroupBySew_5_101};
  wire [31:0]       dataInMem_hi_619 = {dataInMem_hi_hi_363, dataInMem_hi_lo_107};
  wire [23:0]       dataInMem_lo_492 = {dataInMem_lo_hi_236, dataRegroupBySew_0_102};
  wire [15:0]       dataInMem_hi_hi_364 = {dataRegroupBySew_6_102, dataRegroupBySew_5_102};
  wire [31:0]       dataInMem_hi_620 = {dataInMem_hi_hi_364, dataInMem_hi_lo_108};
  wire [23:0]       dataInMem_lo_493 = {dataInMem_lo_hi_237, dataRegroupBySew_0_103};
  wire [15:0]       dataInMem_hi_hi_365 = {dataRegroupBySew_6_103, dataRegroupBySew_5_103};
  wire [31:0]       dataInMem_hi_621 = {dataInMem_hi_hi_365, dataInMem_hi_lo_109};
  wire [23:0]       dataInMem_lo_494 = {dataInMem_lo_hi_238, dataRegroupBySew_0_104};
  wire [15:0]       dataInMem_hi_hi_366 = {dataRegroupBySew_6_104, dataRegroupBySew_5_104};
  wire [31:0]       dataInMem_hi_622 = {dataInMem_hi_hi_366, dataInMem_hi_lo_110};
  wire [23:0]       dataInMem_lo_495 = {dataInMem_lo_hi_239, dataRegroupBySew_0_105};
  wire [15:0]       dataInMem_hi_hi_367 = {dataRegroupBySew_6_105, dataRegroupBySew_5_105};
  wire [31:0]       dataInMem_hi_623 = {dataInMem_hi_hi_367, dataInMem_hi_lo_111};
  wire [23:0]       dataInMem_lo_496 = {dataInMem_lo_hi_240, dataRegroupBySew_0_106};
  wire [15:0]       dataInMem_hi_hi_368 = {dataRegroupBySew_6_106, dataRegroupBySew_5_106};
  wire [31:0]       dataInMem_hi_624 = {dataInMem_hi_hi_368, dataInMem_hi_lo_112};
  wire [23:0]       dataInMem_lo_497 = {dataInMem_lo_hi_241, dataRegroupBySew_0_107};
  wire [15:0]       dataInMem_hi_hi_369 = {dataRegroupBySew_6_107, dataRegroupBySew_5_107};
  wire [31:0]       dataInMem_hi_625 = {dataInMem_hi_hi_369, dataInMem_hi_lo_113};
  wire [23:0]       dataInMem_lo_498 = {dataInMem_lo_hi_242, dataRegroupBySew_0_108};
  wire [15:0]       dataInMem_hi_hi_370 = {dataRegroupBySew_6_108, dataRegroupBySew_5_108};
  wire [31:0]       dataInMem_hi_626 = {dataInMem_hi_hi_370, dataInMem_hi_lo_114};
  wire [23:0]       dataInMem_lo_499 = {dataInMem_lo_hi_243, dataRegroupBySew_0_109};
  wire [15:0]       dataInMem_hi_hi_371 = {dataRegroupBySew_6_109, dataRegroupBySew_5_109};
  wire [31:0]       dataInMem_hi_627 = {dataInMem_hi_hi_371, dataInMem_hi_lo_115};
  wire [23:0]       dataInMem_lo_500 = {dataInMem_lo_hi_244, dataRegroupBySew_0_110};
  wire [15:0]       dataInMem_hi_hi_372 = {dataRegroupBySew_6_110, dataRegroupBySew_5_110};
  wire [31:0]       dataInMem_hi_628 = {dataInMem_hi_hi_372, dataInMem_hi_lo_116};
  wire [23:0]       dataInMem_lo_501 = {dataInMem_lo_hi_245, dataRegroupBySew_0_111};
  wire [15:0]       dataInMem_hi_hi_373 = {dataRegroupBySew_6_111, dataRegroupBySew_5_111};
  wire [31:0]       dataInMem_hi_629 = {dataInMem_hi_hi_373, dataInMem_hi_lo_117};
  wire [23:0]       dataInMem_lo_502 = {dataInMem_lo_hi_246, dataRegroupBySew_0_112};
  wire [15:0]       dataInMem_hi_hi_374 = {dataRegroupBySew_6_112, dataRegroupBySew_5_112};
  wire [31:0]       dataInMem_hi_630 = {dataInMem_hi_hi_374, dataInMem_hi_lo_118};
  wire [23:0]       dataInMem_lo_503 = {dataInMem_lo_hi_247, dataRegroupBySew_0_113};
  wire [15:0]       dataInMem_hi_hi_375 = {dataRegroupBySew_6_113, dataRegroupBySew_5_113};
  wire [31:0]       dataInMem_hi_631 = {dataInMem_hi_hi_375, dataInMem_hi_lo_119};
  wire [23:0]       dataInMem_lo_504 = {dataInMem_lo_hi_248, dataRegroupBySew_0_114};
  wire [15:0]       dataInMem_hi_hi_376 = {dataRegroupBySew_6_114, dataRegroupBySew_5_114};
  wire [31:0]       dataInMem_hi_632 = {dataInMem_hi_hi_376, dataInMem_hi_lo_120};
  wire [23:0]       dataInMem_lo_505 = {dataInMem_lo_hi_249, dataRegroupBySew_0_115};
  wire [15:0]       dataInMem_hi_hi_377 = {dataRegroupBySew_6_115, dataRegroupBySew_5_115};
  wire [31:0]       dataInMem_hi_633 = {dataInMem_hi_hi_377, dataInMem_hi_lo_121};
  wire [23:0]       dataInMem_lo_506 = {dataInMem_lo_hi_250, dataRegroupBySew_0_116};
  wire [15:0]       dataInMem_hi_hi_378 = {dataRegroupBySew_6_116, dataRegroupBySew_5_116};
  wire [31:0]       dataInMem_hi_634 = {dataInMem_hi_hi_378, dataInMem_hi_lo_122};
  wire [23:0]       dataInMem_lo_507 = {dataInMem_lo_hi_251, dataRegroupBySew_0_117};
  wire [15:0]       dataInMem_hi_hi_379 = {dataRegroupBySew_6_117, dataRegroupBySew_5_117};
  wire [31:0]       dataInMem_hi_635 = {dataInMem_hi_hi_379, dataInMem_hi_lo_123};
  wire [23:0]       dataInMem_lo_508 = {dataInMem_lo_hi_252, dataRegroupBySew_0_118};
  wire [15:0]       dataInMem_hi_hi_380 = {dataRegroupBySew_6_118, dataRegroupBySew_5_118};
  wire [31:0]       dataInMem_hi_636 = {dataInMem_hi_hi_380, dataInMem_hi_lo_124};
  wire [23:0]       dataInMem_lo_509 = {dataInMem_lo_hi_253, dataRegroupBySew_0_119};
  wire [15:0]       dataInMem_hi_hi_381 = {dataRegroupBySew_6_119, dataRegroupBySew_5_119};
  wire [31:0]       dataInMem_hi_637 = {dataInMem_hi_hi_381, dataInMem_hi_lo_125};
  wire [23:0]       dataInMem_lo_510 = {dataInMem_lo_hi_254, dataRegroupBySew_0_120};
  wire [15:0]       dataInMem_hi_hi_382 = {dataRegroupBySew_6_120, dataRegroupBySew_5_120};
  wire [31:0]       dataInMem_hi_638 = {dataInMem_hi_hi_382, dataInMem_hi_lo_126};
  wire [23:0]       dataInMem_lo_511 = {dataInMem_lo_hi_255, dataRegroupBySew_0_121};
  wire [15:0]       dataInMem_hi_hi_383 = {dataRegroupBySew_6_121, dataRegroupBySew_5_121};
  wire [31:0]       dataInMem_hi_639 = {dataInMem_hi_hi_383, dataInMem_hi_lo_127};
  wire [23:0]       dataInMem_lo_512 = {dataInMem_lo_hi_256, dataRegroupBySew_0_122};
  wire [15:0]       dataInMem_hi_hi_384 = {dataRegroupBySew_6_122, dataRegroupBySew_5_122};
  wire [31:0]       dataInMem_hi_640 = {dataInMem_hi_hi_384, dataInMem_hi_lo_128};
  wire [23:0]       dataInMem_lo_513 = {dataInMem_lo_hi_257, dataRegroupBySew_0_123};
  wire [15:0]       dataInMem_hi_hi_385 = {dataRegroupBySew_6_123, dataRegroupBySew_5_123};
  wire [31:0]       dataInMem_hi_641 = {dataInMem_hi_hi_385, dataInMem_hi_lo_129};
  wire [23:0]       dataInMem_lo_514 = {dataInMem_lo_hi_258, dataRegroupBySew_0_124};
  wire [15:0]       dataInMem_hi_hi_386 = {dataRegroupBySew_6_124, dataRegroupBySew_5_124};
  wire [31:0]       dataInMem_hi_642 = {dataInMem_hi_hi_386, dataInMem_hi_lo_130};
  wire [23:0]       dataInMem_lo_515 = {dataInMem_lo_hi_259, dataRegroupBySew_0_125};
  wire [15:0]       dataInMem_hi_hi_387 = {dataRegroupBySew_6_125, dataRegroupBySew_5_125};
  wire [31:0]       dataInMem_hi_643 = {dataInMem_hi_hi_387, dataInMem_hi_lo_131};
  wire [23:0]       dataInMem_lo_516 = {dataInMem_lo_hi_260, dataRegroupBySew_0_126};
  wire [15:0]       dataInMem_hi_hi_388 = {dataRegroupBySew_6_126, dataRegroupBySew_5_126};
  wire [31:0]       dataInMem_hi_644 = {dataInMem_hi_hi_388, dataInMem_hi_lo_132};
  wire [23:0]       dataInMem_lo_517 = {dataInMem_lo_hi_261, dataRegroupBySew_0_127};
  wire [15:0]       dataInMem_hi_hi_389 = {dataRegroupBySew_6_127, dataRegroupBySew_5_127};
  wire [31:0]       dataInMem_hi_645 = {dataInMem_hi_hi_389, dataInMem_hi_lo_133};
  wire [111:0]      dataInMem_lo_lo_lo_lo_lo_lo_6 = {dataInMem_hi_519, dataInMem_lo_391, dataInMem_hi_518, dataInMem_lo_390};
  wire [111:0]      dataInMem_lo_lo_lo_lo_lo_hi_6 = {dataInMem_hi_521, dataInMem_lo_393, dataInMem_hi_520, dataInMem_lo_392};
  wire [223:0]      dataInMem_lo_lo_lo_lo_lo_6 = {dataInMem_lo_lo_lo_lo_lo_hi_6, dataInMem_lo_lo_lo_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_lo_lo_lo_hi_lo_6 = {dataInMem_hi_523, dataInMem_lo_395, dataInMem_hi_522, dataInMem_lo_394};
  wire [111:0]      dataInMem_lo_lo_lo_lo_hi_hi_6 = {dataInMem_hi_525, dataInMem_lo_397, dataInMem_hi_524, dataInMem_lo_396};
  wire [223:0]      dataInMem_lo_lo_lo_lo_hi_6 = {dataInMem_lo_lo_lo_lo_hi_hi_6, dataInMem_lo_lo_lo_lo_hi_lo_6};
  wire [447:0]      dataInMem_lo_lo_lo_lo_6 = {dataInMem_lo_lo_lo_lo_hi_6, dataInMem_lo_lo_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_lo_lo_hi_lo_lo_6 = {dataInMem_hi_527, dataInMem_lo_399, dataInMem_hi_526, dataInMem_lo_398};
  wire [111:0]      dataInMem_lo_lo_lo_hi_lo_hi_6 = {dataInMem_hi_529, dataInMem_lo_401, dataInMem_hi_528, dataInMem_lo_400};
  wire [223:0]      dataInMem_lo_lo_lo_hi_lo_6 = {dataInMem_lo_lo_lo_hi_lo_hi_6, dataInMem_lo_lo_lo_hi_lo_lo_6};
  wire [111:0]      dataInMem_lo_lo_lo_hi_hi_lo_6 = {dataInMem_hi_531, dataInMem_lo_403, dataInMem_hi_530, dataInMem_lo_402};
  wire [111:0]      dataInMem_lo_lo_lo_hi_hi_hi_6 = {dataInMem_hi_533, dataInMem_lo_405, dataInMem_hi_532, dataInMem_lo_404};
  wire [223:0]      dataInMem_lo_lo_lo_hi_hi_6 = {dataInMem_lo_lo_lo_hi_hi_hi_6, dataInMem_lo_lo_lo_hi_hi_lo_6};
  wire [447:0]      dataInMem_lo_lo_lo_hi_6 = {dataInMem_lo_lo_lo_hi_hi_6, dataInMem_lo_lo_lo_hi_lo_6};
  wire [895:0]      dataInMem_lo_lo_lo_6 = {dataInMem_lo_lo_lo_hi_6, dataInMem_lo_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_lo_hi_lo_lo_lo_6 = {dataInMem_hi_535, dataInMem_lo_407, dataInMem_hi_534, dataInMem_lo_406};
  wire [111:0]      dataInMem_lo_lo_hi_lo_lo_hi_6 = {dataInMem_hi_537, dataInMem_lo_409, dataInMem_hi_536, dataInMem_lo_408};
  wire [223:0]      dataInMem_lo_lo_hi_lo_lo_6 = {dataInMem_lo_lo_hi_lo_lo_hi_6, dataInMem_lo_lo_hi_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_lo_hi_lo_hi_lo_6 = {dataInMem_hi_539, dataInMem_lo_411, dataInMem_hi_538, dataInMem_lo_410};
  wire [111:0]      dataInMem_lo_lo_hi_lo_hi_hi_6 = {dataInMem_hi_541, dataInMem_lo_413, dataInMem_hi_540, dataInMem_lo_412};
  wire [223:0]      dataInMem_lo_lo_hi_lo_hi_6 = {dataInMem_lo_lo_hi_lo_hi_hi_6, dataInMem_lo_lo_hi_lo_hi_lo_6};
  wire [447:0]      dataInMem_lo_lo_hi_lo_6 = {dataInMem_lo_lo_hi_lo_hi_6, dataInMem_lo_lo_hi_lo_lo_6};
  wire [111:0]      dataInMem_lo_lo_hi_hi_lo_lo_6 = {dataInMem_hi_543, dataInMem_lo_415, dataInMem_hi_542, dataInMem_lo_414};
  wire [111:0]      dataInMem_lo_lo_hi_hi_lo_hi_6 = {dataInMem_hi_545, dataInMem_lo_417, dataInMem_hi_544, dataInMem_lo_416};
  wire [223:0]      dataInMem_lo_lo_hi_hi_lo_6 = {dataInMem_lo_lo_hi_hi_lo_hi_6, dataInMem_lo_lo_hi_hi_lo_lo_6};
  wire [111:0]      dataInMem_lo_lo_hi_hi_hi_lo_6 = {dataInMem_hi_547, dataInMem_lo_419, dataInMem_hi_546, dataInMem_lo_418};
  wire [111:0]      dataInMem_lo_lo_hi_hi_hi_hi_6 = {dataInMem_hi_549, dataInMem_lo_421, dataInMem_hi_548, dataInMem_lo_420};
  wire [223:0]      dataInMem_lo_lo_hi_hi_hi_6 = {dataInMem_lo_lo_hi_hi_hi_hi_6, dataInMem_lo_lo_hi_hi_hi_lo_6};
  wire [447:0]      dataInMem_lo_lo_hi_hi_6 = {dataInMem_lo_lo_hi_hi_hi_6, dataInMem_lo_lo_hi_hi_lo_6};
  wire [895:0]      dataInMem_lo_lo_hi_6 = {dataInMem_lo_lo_hi_hi_6, dataInMem_lo_lo_hi_lo_6};
  wire [1791:0]     dataInMem_lo_lo_6 = {dataInMem_lo_lo_hi_6, dataInMem_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_lo_lo_lo_lo_6 = {dataInMem_hi_551, dataInMem_lo_423, dataInMem_hi_550, dataInMem_lo_422};
  wire [111:0]      dataInMem_lo_hi_lo_lo_lo_hi_6 = {dataInMem_hi_553, dataInMem_lo_425, dataInMem_hi_552, dataInMem_lo_424};
  wire [223:0]      dataInMem_lo_hi_lo_lo_lo_6 = {dataInMem_lo_hi_lo_lo_lo_hi_6, dataInMem_lo_hi_lo_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_lo_lo_hi_lo_6 = {dataInMem_hi_555, dataInMem_lo_427, dataInMem_hi_554, dataInMem_lo_426};
  wire [111:0]      dataInMem_lo_hi_lo_lo_hi_hi_6 = {dataInMem_hi_557, dataInMem_lo_429, dataInMem_hi_556, dataInMem_lo_428};
  wire [223:0]      dataInMem_lo_hi_lo_lo_hi_6 = {dataInMem_lo_hi_lo_lo_hi_hi_6, dataInMem_lo_hi_lo_lo_hi_lo_6};
  wire [447:0]      dataInMem_lo_hi_lo_lo_6 = {dataInMem_lo_hi_lo_lo_hi_6, dataInMem_lo_hi_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_lo_hi_lo_lo_6 = {dataInMem_hi_559, dataInMem_lo_431, dataInMem_hi_558, dataInMem_lo_430};
  wire [111:0]      dataInMem_lo_hi_lo_hi_lo_hi_6 = {dataInMem_hi_561, dataInMem_lo_433, dataInMem_hi_560, dataInMem_lo_432};
  wire [223:0]      dataInMem_lo_hi_lo_hi_lo_6 = {dataInMem_lo_hi_lo_hi_lo_hi_6, dataInMem_lo_hi_lo_hi_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_lo_hi_hi_lo_6 = {dataInMem_hi_563, dataInMem_lo_435, dataInMem_hi_562, dataInMem_lo_434};
  wire [111:0]      dataInMem_lo_hi_lo_hi_hi_hi_6 = {dataInMem_hi_565, dataInMem_lo_437, dataInMem_hi_564, dataInMem_lo_436};
  wire [223:0]      dataInMem_lo_hi_lo_hi_hi_6 = {dataInMem_lo_hi_lo_hi_hi_hi_6, dataInMem_lo_hi_lo_hi_hi_lo_6};
  wire [447:0]      dataInMem_lo_hi_lo_hi_6 = {dataInMem_lo_hi_lo_hi_hi_6, dataInMem_lo_hi_lo_hi_lo_6};
  wire [895:0]      dataInMem_lo_hi_lo_6 = {dataInMem_lo_hi_lo_hi_6, dataInMem_lo_hi_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_hi_lo_lo_lo_6 = {dataInMem_hi_567, dataInMem_lo_439, dataInMem_hi_566, dataInMem_lo_438};
  wire [111:0]      dataInMem_lo_hi_hi_lo_lo_hi_6 = {dataInMem_hi_569, dataInMem_lo_441, dataInMem_hi_568, dataInMem_lo_440};
  wire [223:0]      dataInMem_lo_hi_hi_lo_lo_6 = {dataInMem_lo_hi_hi_lo_lo_hi_6, dataInMem_lo_hi_hi_lo_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_hi_lo_hi_lo_6 = {dataInMem_hi_571, dataInMem_lo_443, dataInMem_hi_570, dataInMem_lo_442};
  wire [111:0]      dataInMem_lo_hi_hi_lo_hi_hi_6 = {dataInMem_hi_573, dataInMem_lo_445, dataInMem_hi_572, dataInMem_lo_444};
  wire [223:0]      dataInMem_lo_hi_hi_lo_hi_6 = {dataInMem_lo_hi_hi_lo_hi_hi_6, dataInMem_lo_hi_hi_lo_hi_lo_6};
  wire [447:0]      dataInMem_lo_hi_hi_lo_6 = {dataInMem_lo_hi_hi_lo_hi_6, dataInMem_lo_hi_hi_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_hi_hi_lo_lo_6 = {dataInMem_hi_575, dataInMem_lo_447, dataInMem_hi_574, dataInMem_lo_446};
  wire [111:0]      dataInMem_lo_hi_hi_hi_lo_hi_6 = {dataInMem_hi_577, dataInMem_lo_449, dataInMem_hi_576, dataInMem_lo_448};
  wire [223:0]      dataInMem_lo_hi_hi_hi_lo_6 = {dataInMem_lo_hi_hi_hi_lo_hi_6, dataInMem_lo_hi_hi_hi_lo_lo_6};
  wire [111:0]      dataInMem_lo_hi_hi_hi_hi_lo_6 = {dataInMem_hi_579, dataInMem_lo_451, dataInMem_hi_578, dataInMem_lo_450};
  wire [111:0]      dataInMem_lo_hi_hi_hi_hi_hi_6 = {dataInMem_hi_581, dataInMem_lo_453, dataInMem_hi_580, dataInMem_lo_452};
  wire [223:0]      dataInMem_lo_hi_hi_hi_hi_6 = {dataInMem_lo_hi_hi_hi_hi_hi_6, dataInMem_lo_hi_hi_hi_hi_lo_6};
  wire [447:0]      dataInMem_lo_hi_hi_hi_6 = {dataInMem_lo_hi_hi_hi_hi_6, dataInMem_lo_hi_hi_hi_lo_6};
  wire [895:0]      dataInMem_lo_hi_hi_6 = {dataInMem_lo_hi_hi_hi_6, dataInMem_lo_hi_hi_lo_6};
  wire [1791:0]     dataInMem_lo_hi_262 = {dataInMem_lo_hi_hi_6, dataInMem_lo_hi_lo_6};
  wire [3583:0]     dataInMem_lo_518 = {dataInMem_lo_hi_262, dataInMem_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_lo_lo_lo_lo_6 = {dataInMem_hi_583, dataInMem_lo_455, dataInMem_hi_582, dataInMem_lo_454};
  wire [111:0]      dataInMem_hi_lo_lo_lo_lo_hi_6 = {dataInMem_hi_585, dataInMem_lo_457, dataInMem_hi_584, dataInMem_lo_456};
  wire [223:0]      dataInMem_hi_lo_lo_lo_lo_6 = {dataInMem_hi_lo_lo_lo_lo_hi_6, dataInMem_hi_lo_lo_lo_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_lo_lo_hi_lo_6 = {dataInMem_hi_587, dataInMem_lo_459, dataInMem_hi_586, dataInMem_lo_458};
  wire [111:0]      dataInMem_hi_lo_lo_lo_hi_hi_6 = {dataInMem_hi_589, dataInMem_lo_461, dataInMem_hi_588, dataInMem_lo_460};
  wire [223:0]      dataInMem_hi_lo_lo_lo_hi_6 = {dataInMem_hi_lo_lo_lo_hi_hi_6, dataInMem_hi_lo_lo_lo_hi_lo_6};
  wire [447:0]      dataInMem_hi_lo_lo_lo_6 = {dataInMem_hi_lo_lo_lo_hi_6, dataInMem_hi_lo_lo_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_lo_hi_lo_lo_6 = {dataInMem_hi_591, dataInMem_lo_463, dataInMem_hi_590, dataInMem_lo_462};
  wire [111:0]      dataInMem_hi_lo_lo_hi_lo_hi_6 = {dataInMem_hi_593, dataInMem_lo_465, dataInMem_hi_592, dataInMem_lo_464};
  wire [223:0]      dataInMem_hi_lo_lo_hi_lo_6 = {dataInMem_hi_lo_lo_hi_lo_hi_6, dataInMem_hi_lo_lo_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_lo_hi_hi_lo_6 = {dataInMem_hi_595, dataInMem_lo_467, dataInMem_hi_594, dataInMem_lo_466};
  wire [111:0]      dataInMem_hi_lo_lo_hi_hi_hi_6 = {dataInMem_hi_597, dataInMem_lo_469, dataInMem_hi_596, dataInMem_lo_468};
  wire [223:0]      dataInMem_hi_lo_lo_hi_hi_6 = {dataInMem_hi_lo_lo_hi_hi_hi_6, dataInMem_hi_lo_lo_hi_hi_lo_6};
  wire [447:0]      dataInMem_hi_lo_lo_hi_6 = {dataInMem_hi_lo_lo_hi_hi_6, dataInMem_hi_lo_lo_hi_lo_6};
  wire [895:0]      dataInMem_hi_lo_lo_6 = {dataInMem_hi_lo_lo_hi_6, dataInMem_hi_lo_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_hi_lo_lo_lo_6 = {dataInMem_hi_599, dataInMem_lo_471, dataInMem_hi_598, dataInMem_lo_470};
  wire [111:0]      dataInMem_hi_lo_hi_lo_lo_hi_6 = {dataInMem_hi_601, dataInMem_lo_473, dataInMem_hi_600, dataInMem_lo_472};
  wire [223:0]      dataInMem_hi_lo_hi_lo_lo_6 = {dataInMem_hi_lo_hi_lo_lo_hi_6, dataInMem_hi_lo_hi_lo_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_hi_lo_hi_lo_6 = {dataInMem_hi_603, dataInMem_lo_475, dataInMem_hi_602, dataInMem_lo_474};
  wire [111:0]      dataInMem_hi_lo_hi_lo_hi_hi_6 = {dataInMem_hi_605, dataInMem_lo_477, dataInMem_hi_604, dataInMem_lo_476};
  wire [223:0]      dataInMem_hi_lo_hi_lo_hi_6 = {dataInMem_hi_lo_hi_lo_hi_hi_6, dataInMem_hi_lo_hi_lo_hi_lo_6};
  wire [447:0]      dataInMem_hi_lo_hi_lo_6 = {dataInMem_hi_lo_hi_lo_hi_6, dataInMem_hi_lo_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_hi_hi_lo_lo_6 = {dataInMem_hi_607, dataInMem_lo_479, dataInMem_hi_606, dataInMem_lo_478};
  wire [111:0]      dataInMem_hi_lo_hi_hi_lo_hi_6 = {dataInMem_hi_609, dataInMem_lo_481, dataInMem_hi_608, dataInMem_lo_480};
  wire [223:0]      dataInMem_hi_lo_hi_hi_lo_6 = {dataInMem_hi_lo_hi_hi_lo_hi_6, dataInMem_hi_lo_hi_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_lo_hi_hi_hi_lo_6 = {dataInMem_hi_611, dataInMem_lo_483, dataInMem_hi_610, dataInMem_lo_482};
  wire [111:0]      dataInMem_hi_lo_hi_hi_hi_hi_6 = {dataInMem_hi_613, dataInMem_lo_485, dataInMem_hi_612, dataInMem_lo_484};
  wire [223:0]      dataInMem_hi_lo_hi_hi_hi_6 = {dataInMem_hi_lo_hi_hi_hi_hi_6, dataInMem_hi_lo_hi_hi_hi_lo_6};
  wire [447:0]      dataInMem_hi_lo_hi_hi_6 = {dataInMem_hi_lo_hi_hi_hi_6, dataInMem_hi_lo_hi_hi_lo_6};
  wire [895:0]      dataInMem_hi_lo_hi_6 = {dataInMem_hi_lo_hi_hi_6, dataInMem_hi_lo_hi_lo_6};
  wire [1791:0]     dataInMem_hi_lo_134 = {dataInMem_hi_lo_hi_6, dataInMem_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_lo_lo_lo_lo_6 = {dataInMem_hi_615, dataInMem_lo_487, dataInMem_hi_614, dataInMem_lo_486};
  wire [111:0]      dataInMem_hi_hi_lo_lo_lo_hi_6 = {dataInMem_hi_617, dataInMem_lo_489, dataInMem_hi_616, dataInMem_lo_488};
  wire [223:0]      dataInMem_hi_hi_lo_lo_lo_6 = {dataInMem_hi_hi_lo_lo_lo_hi_6, dataInMem_hi_hi_lo_lo_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_lo_lo_hi_lo_6 = {dataInMem_hi_619, dataInMem_lo_491, dataInMem_hi_618, dataInMem_lo_490};
  wire [111:0]      dataInMem_hi_hi_lo_lo_hi_hi_6 = {dataInMem_hi_621, dataInMem_lo_493, dataInMem_hi_620, dataInMem_lo_492};
  wire [223:0]      dataInMem_hi_hi_lo_lo_hi_6 = {dataInMem_hi_hi_lo_lo_hi_hi_6, dataInMem_hi_hi_lo_lo_hi_lo_6};
  wire [447:0]      dataInMem_hi_hi_lo_lo_6 = {dataInMem_hi_hi_lo_lo_hi_6, dataInMem_hi_hi_lo_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_lo_hi_lo_lo_6 = {dataInMem_hi_623, dataInMem_lo_495, dataInMem_hi_622, dataInMem_lo_494};
  wire [111:0]      dataInMem_hi_hi_lo_hi_lo_hi_6 = {dataInMem_hi_625, dataInMem_lo_497, dataInMem_hi_624, dataInMem_lo_496};
  wire [223:0]      dataInMem_hi_hi_lo_hi_lo_6 = {dataInMem_hi_hi_lo_hi_lo_hi_6, dataInMem_hi_hi_lo_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_lo_hi_hi_lo_6 = {dataInMem_hi_627, dataInMem_lo_499, dataInMem_hi_626, dataInMem_lo_498};
  wire [111:0]      dataInMem_hi_hi_lo_hi_hi_hi_6 = {dataInMem_hi_629, dataInMem_lo_501, dataInMem_hi_628, dataInMem_lo_500};
  wire [223:0]      dataInMem_hi_hi_lo_hi_hi_6 = {dataInMem_hi_hi_lo_hi_hi_hi_6, dataInMem_hi_hi_lo_hi_hi_lo_6};
  wire [447:0]      dataInMem_hi_hi_lo_hi_6 = {dataInMem_hi_hi_lo_hi_hi_6, dataInMem_hi_hi_lo_hi_lo_6};
  wire [895:0]      dataInMem_hi_hi_lo_6 = {dataInMem_hi_hi_lo_hi_6, dataInMem_hi_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_hi_lo_lo_lo_6 = {dataInMem_hi_631, dataInMem_lo_503, dataInMem_hi_630, dataInMem_lo_502};
  wire [111:0]      dataInMem_hi_hi_hi_lo_lo_hi_6 = {dataInMem_hi_633, dataInMem_lo_505, dataInMem_hi_632, dataInMem_lo_504};
  wire [223:0]      dataInMem_hi_hi_hi_lo_lo_6 = {dataInMem_hi_hi_hi_lo_lo_hi_6, dataInMem_hi_hi_hi_lo_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_hi_lo_hi_lo_6 = {dataInMem_hi_635, dataInMem_lo_507, dataInMem_hi_634, dataInMem_lo_506};
  wire [111:0]      dataInMem_hi_hi_hi_lo_hi_hi_6 = {dataInMem_hi_637, dataInMem_lo_509, dataInMem_hi_636, dataInMem_lo_508};
  wire [223:0]      dataInMem_hi_hi_hi_lo_hi_6 = {dataInMem_hi_hi_hi_lo_hi_hi_6, dataInMem_hi_hi_hi_lo_hi_lo_6};
  wire [447:0]      dataInMem_hi_hi_hi_lo_6 = {dataInMem_hi_hi_hi_lo_hi_6, dataInMem_hi_hi_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_hi_hi_lo_lo_6 = {dataInMem_hi_639, dataInMem_lo_511, dataInMem_hi_638, dataInMem_lo_510};
  wire [111:0]      dataInMem_hi_hi_hi_hi_lo_hi_6 = {dataInMem_hi_641, dataInMem_lo_513, dataInMem_hi_640, dataInMem_lo_512};
  wire [223:0]      dataInMem_hi_hi_hi_hi_lo_6 = {dataInMem_hi_hi_hi_hi_lo_hi_6, dataInMem_hi_hi_hi_hi_lo_lo_6};
  wire [111:0]      dataInMem_hi_hi_hi_hi_hi_lo_6 = {dataInMem_hi_643, dataInMem_lo_515, dataInMem_hi_642, dataInMem_lo_514};
  wire [111:0]      dataInMem_hi_hi_hi_hi_hi_hi_6 = {dataInMem_hi_645, dataInMem_lo_517, dataInMem_hi_644, dataInMem_lo_516};
  wire [223:0]      dataInMem_hi_hi_hi_hi_hi_6 = {dataInMem_hi_hi_hi_hi_hi_hi_6, dataInMem_hi_hi_hi_hi_hi_lo_6};
  wire [447:0]      dataInMem_hi_hi_hi_hi_6 = {dataInMem_hi_hi_hi_hi_hi_6, dataInMem_hi_hi_hi_hi_lo_6};
  wire [895:0]      dataInMem_hi_hi_hi_6 = {dataInMem_hi_hi_hi_hi_6, dataInMem_hi_hi_hi_lo_6};
  wire [1791:0]     dataInMem_hi_hi_390 = {dataInMem_hi_hi_hi_6, dataInMem_hi_hi_lo_6};
  wire [3583:0]     dataInMem_hi_646 = {dataInMem_hi_hi_390, dataInMem_hi_lo_134};
  wire [7167:0]     dataInMem_6 = {dataInMem_hi_646, dataInMem_lo_518};
  wire [1023:0]     regroupCacheLine_6_0 = dataInMem_6[1023:0];
  wire [1023:0]     regroupCacheLine_6_1 = dataInMem_6[2047:1024];
  wire [1023:0]     regroupCacheLine_6_2 = dataInMem_6[3071:2048];
  wire [1023:0]     regroupCacheLine_6_3 = dataInMem_6[4095:3072];
  wire [1023:0]     regroupCacheLine_6_4 = dataInMem_6[5119:4096];
  wire [1023:0]     regroupCacheLine_6_5 = dataInMem_6[6143:5120];
  wire [1023:0]     regroupCacheLine_6_6 = dataInMem_6[7167:6144];
  wire [1023:0]     res_48 = regroupCacheLine_6_0;
  wire [1023:0]     res_49 = regroupCacheLine_6_1;
  wire [1023:0]     res_50 = regroupCacheLine_6_2;
  wire [1023:0]     res_51 = regroupCacheLine_6_3;
  wire [1023:0]     res_52 = regroupCacheLine_6_4;
  wire [1023:0]     res_53 = regroupCacheLine_6_5;
  wire [1023:0]     res_54 = regroupCacheLine_6_6;
  wire [2047:0]     lo_lo_6 = {res_49, res_48};
  wire [2047:0]     lo_hi_6 = {res_51, res_50};
  wire [4095:0]     lo_6 = {lo_hi_6, lo_lo_6};
  wire [2047:0]     hi_lo_6 = {res_53, res_52};
  wire [2047:0]     hi_hi_6 = {1024'h0, res_54};
  wire [4095:0]     hi_6 = {hi_hi_6, hi_lo_6};
  wire [8191:0]     regroupLoadData_0_6 = {hi_6, lo_6};
  wire [31:0]       dataInMem_lo_519 = {dataInMem_lo_hi_263, dataInMem_lo_lo_7};
  wire [15:0]       dataInMem_hi_hi_391 = {dataRegroupBySew_7_0, dataRegroupBySew_6_0};
  wire [31:0]       dataInMem_hi_647 = {dataInMem_hi_hi_391, dataInMem_hi_lo_135};
  wire [31:0]       dataInMem_lo_520 = {dataInMem_lo_hi_264, dataInMem_lo_lo_8};
  wire [15:0]       dataInMem_hi_hi_392 = {dataRegroupBySew_7_1, dataRegroupBySew_6_1};
  wire [31:0]       dataInMem_hi_648 = {dataInMem_hi_hi_392, dataInMem_hi_lo_136};
  wire [31:0]       dataInMem_lo_521 = {dataInMem_lo_hi_265, dataInMem_lo_lo_9};
  wire [15:0]       dataInMem_hi_hi_393 = {dataRegroupBySew_7_2, dataRegroupBySew_6_2};
  wire [31:0]       dataInMem_hi_649 = {dataInMem_hi_hi_393, dataInMem_hi_lo_137};
  wire [31:0]       dataInMem_lo_522 = {dataInMem_lo_hi_266, dataInMem_lo_lo_10};
  wire [15:0]       dataInMem_hi_hi_394 = {dataRegroupBySew_7_3, dataRegroupBySew_6_3};
  wire [31:0]       dataInMem_hi_650 = {dataInMem_hi_hi_394, dataInMem_hi_lo_138};
  wire [31:0]       dataInMem_lo_523 = {dataInMem_lo_hi_267, dataInMem_lo_lo_11};
  wire [15:0]       dataInMem_hi_hi_395 = {dataRegroupBySew_7_4, dataRegroupBySew_6_4};
  wire [31:0]       dataInMem_hi_651 = {dataInMem_hi_hi_395, dataInMem_hi_lo_139};
  wire [31:0]       dataInMem_lo_524 = {dataInMem_lo_hi_268, dataInMem_lo_lo_12};
  wire [15:0]       dataInMem_hi_hi_396 = {dataRegroupBySew_7_5, dataRegroupBySew_6_5};
  wire [31:0]       dataInMem_hi_652 = {dataInMem_hi_hi_396, dataInMem_hi_lo_140};
  wire [31:0]       dataInMem_lo_525 = {dataInMem_lo_hi_269, dataInMem_lo_lo_13};
  wire [15:0]       dataInMem_hi_hi_397 = {dataRegroupBySew_7_6, dataRegroupBySew_6_6};
  wire [31:0]       dataInMem_hi_653 = {dataInMem_hi_hi_397, dataInMem_hi_lo_141};
  wire [31:0]       dataInMem_lo_526 = {dataInMem_lo_hi_270, dataInMem_lo_lo_14};
  wire [15:0]       dataInMem_hi_hi_398 = {dataRegroupBySew_7_7, dataRegroupBySew_6_7};
  wire [31:0]       dataInMem_hi_654 = {dataInMem_hi_hi_398, dataInMem_hi_lo_142};
  wire [31:0]       dataInMem_lo_527 = {dataInMem_lo_hi_271, dataInMem_lo_lo_15};
  wire [15:0]       dataInMem_hi_hi_399 = {dataRegroupBySew_7_8, dataRegroupBySew_6_8};
  wire [31:0]       dataInMem_hi_655 = {dataInMem_hi_hi_399, dataInMem_hi_lo_143};
  wire [31:0]       dataInMem_lo_528 = {dataInMem_lo_hi_272, dataInMem_lo_lo_16};
  wire [15:0]       dataInMem_hi_hi_400 = {dataRegroupBySew_7_9, dataRegroupBySew_6_9};
  wire [31:0]       dataInMem_hi_656 = {dataInMem_hi_hi_400, dataInMem_hi_lo_144};
  wire [31:0]       dataInMem_lo_529 = {dataInMem_lo_hi_273, dataInMem_lo_lo_17};
  wire [15:0]       dataInMem_hi_hi_401 = {dataRegroupBySew_7_10, dataRegroupBySew_6_10};
  wire [31:0]       dataInMem_hi_657 = {dataInMem_hi_hi_401, dataInMem_hi_lo_145};
  wire [31:0]       dataInMem_lo_530 = {dataInMem_lo_hi_274, dataInMem_lo_lo_18};
  wire [15:0]       dataInMem_hi_hi_402 = {dataRegroupBySew_7_11, dataRegroupBySew_6_11};
  wire [31:0]       dataInMem_hi_658 = {dataInMem_hi_hi_402, dataInMem_hi_lo_146};
  wire [31:0]       dataInMem_lo_531 = {dataInMem_lo_hi_275, dataInMem_lo_lo_19};
  wire [15:0]       dataInMem_hi_hi_403 = {dataRegroupBySew_7_12, dataRegroupBySew_6_12};
  wire [31:0]       dataInMem_hi_659 = {dataInMem_hi_hi_403, dataInMem_hi_lo_147};
  wire [31:0]       dataInMem_lo_532 = {dataInMem_lo_hi_276, dataInMem_lo_lo_20};
  wire [15:0]       dataInMem_hi_hi_404 = {dataRegroupBySew_7_13, dataRegroupBySew_6_13};
  wire [31:0]       dataInMem_hi_660 = {dataInMem_hi_hi_404, dataInMem_hi_lo_148};
  wire [31:0]       dataInMem_lo_533 = {dataInMem_lo_hi_277, dataInMem_lo_lo_21};
  wire [15:0]       dataInMem_hi_hi_405 = {dataRegroupBySew_7_14, dataRegroupBySew_6_14};
  wire [31:0]       dataInMem_hi_661 = {dataInMem_hi_hi_405, dataInMem_hi_lo_149};
  wire [31:0]       dataInMem_lo_534 = {dataInMem_lo_hi_278, dataInMem_lo_lo_22};
  wire [15:0]       dataInMem_hi_hi_406 = {dataRegroupBySew_7_15, dataRegroupBySew_6_15};
  wire [31:0]       dataInMem_hi_662 = {dataInMem_hi_hi_406, dataInMem_hi_lo_150};
  wire [31:0]       dataInMem_lo_535 = {dataInMem_lo_hi_279, dataInMem_lo_lo_23};
  wire [15:0]       dataInMem_hi_hi_407 = {dataRegroupBySew_7_16, dataRegroupBySew_6_16};
  wire [31:0]       dataInMem_hi_663 = {dataInMem_hi_hi_407, dataInMem_hi_lo_151};
  wire [31:0]       dataInMem_lo_536 = {dataInMem_lo_hi_280, dataInMem_lo_lo_24};
  wire [15:0]       dataInMem_hi_hi_408 = {dataRegroupBySew_7_17, dataRegroupBySew_6_17};
  wire [31:0]       dataInMem_hi_664 = {dataInMem_hi_hi_408, dataInMem_hi_lo_152};
  wire [31:0]       dataInMem_lo_537 = {dataInMem_lo_hi_281, dataInMem_lo_lo_25};
  wire [15:0]       dataInMem_hi_hi_409 = {dataRegroupBySew_7_18, dataRegroupBySew_6_18};
  wire [31:0]       dataInMem_hi_665 = {dataInMem_hi_hi_409, dataInMem_hi_lo_153};
  wire [31:0]       dataInMem_lo_538 = {dataInMem_lo_hi_282, dataInMem_lo_lo_26};
  wire [15:0]       dataInMem_hi_hi_410 = {dataRegroupBySew_7_19, dataRegroupBySew_6_19};
  wire [31:0]       dataInMem_hi_666 = {dataInMem_hi_hi_410, dataInMem_hi_lo_154};
  wire [31:0]       dataInMem_lo_539 = {dataInMem_lo_hi_283, dataInMem_lo_lo_27};
  wire [15:0]       dataInMem_hi_hi_411 = {dataRegroupBySew_7_20, dataRegroupBySew_6_20};
  wire [31:0]       dataInMem_hi_667 = {dataInMem_hi_hi_411, dataInMem_hi_lo_155};
  wire [31:0]       dataInMem_lo_540 = {dataInMem_lo_hi_284, dataInMem_lo_lo_28};
  wire [15:0]       dataInMem_hi_hi_412 = {dataRegroupBySew_7_21, dataRegroupBySew_6_21};
  wire [31:0]       dataInMem_hi_668 = {dataInMem_hi_hi_412, dataInMem_hi_lo_156};
  wire [31:0]       dataInMem_lo_541 = {dataInMem_lo_hi_285, dataInMem_lo_lo_29};
  wire [15:0]       dataInMem_hi_hi_413 = {dataRegroupBySew_7_22, dataRegroupBySew_6_22};
  wire [31:0]       dataInMem_hi_669 = {dataInMem_hi_hi_413, dataInMem_hi_lo_157};
  wire [31:0]       dataInMem_lo_542 = {dataInMem_lo_hi_286, dataInMem_lo_lo_30};
  wire [15:0]       dataInMem_hi_hi_414 = {dataRegroupBySew_7_23, dataRegroupBySew_6_23};
  wire [31:0]       dataInMem_hi_670 = {dataInMem_hi_hi_414, dataInMem_hi_lo_158};
  wire [31:0]       dataInMem_lo_543 = {dataInMem_lo_hi_287, dataInMem_lo_lo_31};
  wire [15:0]       dataInMem_hi_hi_415 = {dataRegroupBySew_7_24, dataRegroupBySew_6_24};
  wire [31:0]       dataInMem_hi_671 = {dataInMem_hi_hi_415, dataInMem_hi_lo_159};
  wire [31:0]       dataInMem_lo_544 = {dataInMem_lo_hi_288, dataInMem_lo_lo_32};
  wire [15:0]       dataInMem_hi_hi_416 = {dataRegroupBySew_7_25, dataRegroupBySew_6_25};
  wire [31:0]       dataInMem_hi_672 = {dataInMem_hi_hi_416, dataInMem_hi_lo_160};
  wire [31:0]       dataInMem_lo_545 = {dataInMem_lo_hi_289, dataInMem_lo_lo_33};
  wire [15:0]       dataInMem_hi_hi_417 = {dataRegroupBySew_7_26, dataRegroupBySew_6_26};
  wire [31:0]       dataInMem_hi_673 = {dataInMem_hi_hi_417, dataInMem_hi_lo_161};
  wire [31:0]       dataInMem_lo_546 = {dataInMem_lo_hi_290, dataInMem_lo_lo_34};
  wire [15:0]       dataInMem_hi_hi_418 = {dataRegroupBySew_7_27, dataRegroupBySew_6_27};
  wire [31:0]       dataInMem_hi_674 = {dataInMem_hi_hi_418, dataInMem_hi_lo_162};
  wire [31:0]       dataInMem_lo_547 = {dataInMem_lo_hi_291, dataInMem_lo_lo_35};
  wire [15:0]       dataInMem_hi_hi_419 = {dataRegroupBySew_7_28, dataRegroupBySew_6_28};
  wire [31:0]       dataInMem_hi_675 = {dataInMem_hi_hi_419, dataInMem_hi_lo_163};
  wire [31:0]       dataInMem_lo_548 = {dataInMem_lo_hi_292, dataInMem_lo_lo_36};
  wire [15:0]       dataInMem_hi_hi_420 = {dataRegroupBySew_7_29, dataRegroupBySew_6_29};
  wire [31:0]       dataInMem_hi_676 = {dataInMem_hi_hi_420, dataInMem_hi_lo_164};
  wire [31:0]       dataInMem_lo_549 = {dataInMem_lo_hi_293, dataInMem_lo_lo_37};
  wire [15:0]       dataInMem_hi_hi_421 = {dataRegroupBySew_7_30, dataRegroupBySew_6_30};
  wire [31:0]       dataInMem_hi_677 = {dataInMem_hi_hi_421, dataInMem_hi_lo_165};
  wire [31:0]       dataInMem_lo_550 = {dataInMem_lo_hi_294, dataInMem_lo_lo_38};
  wire [15:0]       dataInMem_hi_hi_422 = {dataRegroupBySew_7_31, dataRegroupBySew_6_31};
  wire [31:0]       dataInMem_hi_678 = {dataInMem_hi_hi_422, dataInMem_hi_lo_166};
  wire [31:0]       dataInMem_lo_551 = {dataInMem_lo_hi_295, dataInMem_lo_lo_39};
  wire [15:0]       dataInMem_hi_hi_423 = {dataRegroupBySew_7_32, dataRegroupBySew_6_32};
  wire [31:0]       dataInMem_hi_679 = {dataInMem_hi_hi_423, dataInMem_hi_lo_167};
  wire [31:0]       dataInMem_lo_552 = {dataInMem_lo_hi_296, dataInMem_lo_lo_40};
  wire [15:0]       dataInMem_hi_hi_424 = {dataRegroupBySew_7_33, dataRegroupBySew_6_33};
  wire [31:0]       dataInMem_hi_680 = {dataInMem_hi_hi_424, dataInMem_hi_lo_168};
  wire [31:0]       dataInMem_lo_553 = {dataInMem_lo_hi_297, dataInMem_lo_lo_41};
  wire [15:0]       dataInMem_hi_hi_425 = {dataRegroupBySew_7_34, dataRegroupBySew_6_34};
  wire [31:0]       dataInMem_hi_681 = {dataInMem_hi_hi_425, dataInMem_hi_lo_169};
  wire [31:0]       dataInMem_lo_554 = {dataInMem_lo_hi_298, dataInMem_lo_lo_42};
  wire [15:0]       dataInMem_hi_hi_426 = {dataRegroupBySew_7_35, dataRegroupBySew_6_35};
  wire [31:0]       dataInMem_hi_682 = {dataInMem_hi_hi_426, dataInMem_hi_lo_170};
  wire [31:0]       dataInMem_lo_555 = {dataInMem_lo_hi_299, dataInMem_lo_lo_43};
  wire [15:0]       dataInMem_hi_hi_427 = {dataRegroupBySew_7_36, dataRegroupBySew_6_36};
  wire [31:0]       dataInMem_hi_683 = {dataInMem_hi_hi_427, dataInMem_hi_lo_171};
  wire [31:0]       dataInMem_lo_556 = {dataInMem_lo_hi_300, dataInMem_lo_lo_44};
  wire [15:0]       dataInMem_hi_hi_428 = {dataRegroupBySew_7_37, dataRegroupBySew_6_37};
  wire [31:0]       dataInMem_hi_684 = {dataInMem_hi_hi_428, dataInMem_hi_lo_172};
  wire [31:0]       dataInMem_lo_557 = {dataInMem_lo_hi_301, dataInMem_lo_lo_45};
  wire [15:0]       dataInMem_hi_hi_429 = {dataRegroupBySew_7_38, dataRegroupBySew_6_38};
  wire [31:0]       dataInMem_hi_685 = {dataInMem_hi_hi_429, dataInMem_hi_lo_173};
  wire [31:0]       dataInMem_lo_558 = {dataInMem_lo_hi_302, dataInMem_lo_lo_46};
  wire [15:0]       dataInMem_hi_hi_430 = {dataRegroupBySew_7_39, dataRegroupBySew_6_39};
  wire [31:0]       dataInMem_hi_686 = {dataInMem_hi_hi_430, dataInMem_hi_lo_174};
  wire [31:0]       dataInMem_lo_559 = {dataInMem_lo_hi_303, dataInMem_lo_lo_47};
  wire [15:0]       dataInMem_hi_hi_431 = {dataRegroupBySew_7_40, dataRegroupBySew_6_40};
  wire [31:0]       dataInMem_hi_687 = {dataInMem_hi_hi_431, dataInMem_hi_lo_175};
  wire [31:0]       dataInMem_lo_560 = {dataInMem_lo_hi_304, dataInMem_lo_lo_48};
  wire [15:0]       dataInMem_hi_hi_432 = {dataRegroupBySew_7_41, dataRegroupBySew_6_41};
  wire [31:0]       dataInMem_hi_688 = {dataInMem_hi_hi_432, dataInMem_hi_lo_176};
  wire [31:0]       dataInMem_lo_561 = {dataInMem_lo_hi_305, dataInMem_lo_lo_49};
  wire [15:0]       dataInMem_hi_hi_433 = {dataRegroupBySew_7_42, dataRegroupBySew_6_42};
  wire [31:0]       dataInMem_hi_689 = {dataInMem_hi_hi_433, dataInMem_hi_lo_177};
  wire [31:0]       dataInMem_lo_562 = {dataInMem_lo_hi_306, dataInMem_lo_lo_50};
  wire [15:0]       dataInMem_hi_hi_434 = {dataRegroupBySew_7_43, dataRegroupBySew_6_43};
  wire [31:0]       dataInMem_hi_690 = {dataInMem_hi_hi_434, dataInMem_hi_lo_178};
  wire [31:0]       dataInMem_lo_563 = {dataInMem_lo_hi_307, dataInMem_lo_lo_51};
  wire [15:0]       dataInMem_hi_hi_435 = {dataRegroupBySew_7_44, dataRegroupBySew_6_44};
  wire [31:0]       dataInMem_hi_691 = {dataInMem_hi_hi_435, dataInMem_hi_lo_179};
  wire [31:0]       dataInMem_lo_564 = {dataInMem_lo_hi_308, dataInMem_lo_lo_52};
  wire [15:0]       dataInMem_hi_hi_436 = {dataRegroupBySew_7_45, dataRegroupBySew_6_45};
  wire [31:0]       dataInMem_hi_692 = {dataInMem_hi_hi_436, dataInMem_hi_lo_180};
  wire [31:0]       dataInMem_lo_565 = {dataInMem_lo_hi_309, dataInMem_lo_lo_53};
  wire [15:0]       dataInMem_hi_hi_437 = {dataRegroupBySew_7_46, dataRegroupBySew_6_46};
  wire [31:0]       dataInMem_hi_693 = {dataInMem_hi_hi_437, dataInMem_hi_lo_181};
  wire [31:0]       dataInMem_lo_566 = {dataInMem_lo_hi_310, dataInMem_lo_lo_54};
  wire [15:0]       dataInMem_hi_hi_438 = {dataRegroupBySew_7_47, dataRegroupBySew_6_47};
  wire [31:0]       dataInMem_hi_694 = {dataInMem_hi_hi_438, dataInMem_hi_lo_182};
  wire [31:0]       dataInMem_lo_567 = {dataInMem_lo_hi_311, dataInMem_lo_lo_55};
  wire [15:0]       dataInMem_hi_hi_439 = {dataRegroupBySew_7_48, dataRegroupBySew_6_48};
  wire [31:0]       dataInMem_hi_695 = {dataInMem_hi_hi_439, dataInMem_hi_lo_183};
  wire [31:0]       dataInMem_lo_568 = {dataInMem_lo_hi_312, dataInMem_lo_lo_56};
  wire [15:0]       dataInMem_hi_hi_440 = {dataRegroupBySew_7_49, dataRegroupBySew_6_49};
  wire [31:0]       dataInMem_hi_696 = {dataInMem_hi_hi_440, dataInMem_hi_lo_184};
  wire [31:0]       dataInMem_lo_569 = {dataInMem_lo_hi_313, dataInMem_lo_lo_57};
  wire [15:0]       dataInMem_hi_hi_441 = {dataRegroupBySew_7_50, dataRegroupBySew_6_50};
  wire [31:0]       dataInMem_hi_697 = {dataInMem_hi_hi_441, dataInMem_hi_lo_185};
  wire [31:0]       dataInMem_lo_570 = {dataInMem_lo_hi_314, dataInMem_lo_lo_58};
  wire [15:0]       dataInMem_hi_hi_442 = {dataRegroupBySew_7_51, dataRegroupBySew_6_51};
  wire [31:0]       dataInMem_hi_698 = {dataInMem_hi_hi_442, dataInMem_hi_lo_186};
  wire [31:0]       dataInMem_lo_571 = {dataInMem_lo_hi_315, dataInMem_lo_lo_59};
  wire [15:0]       dataInMem_hi_hi_443 = {dataRegroupBySew_7_52, dataRegroupBySew_6_52};
  wire [31:0]       dataInMem_hi_699 = {dataInMem_hi_hi_443, dataInMem_hi_lo_187};
  wire [31:0]       dataInMem_lo_572 = {dataInMem_lo_hi_316, dataInMem_lo_lo_60};
  wire [15:0]       dataInMem_hi_hi_444 = {dataRegroupBySew_7_53, dataRegroupBySew_6_53};
  wire [31:0]       dataInMem_hi_700 = {dataInMem_hi_hi_444, dataInMem_hi_lo_188};
  wire [31:0]       dataInMem_lo_573 = {dataInMem_lo_hi_317, dataInMem_lo_lo_61};
  wire [15:0]       dataInMem_hi_hi_445 = {dataRegroupBySew_7_54, dataRegroupBySew_6_54};
  wire [31:0]       dataInMem_hi_701 = {dataInMem_hi_hi_445, dataInMem_hi_lo_189};
  wire [31:0]       dataInMem_lo_574 = {dataInMem_lo_hi_318, dataInMem_lo_lo_62};
  wire [15:0]       dataInMem_hi_hi_446 = {dataRegroupBySew_7_55, dataRegroupBySew_6_55};
  wire [31:0]       dataInMem_hi_702 = {dataInMem_hi_hi_446, dataInMem_hi_lo_190};
  wire [31:0]       dataInMem_lo_575 = {dataInMem_lo_hi_319, dataInMem_lo_lo_63};
  wire [15:0]       dataInMem_hi_hi_447 = {dataRegroupBySew_7_56, dataRegroupBySew_6_56};
  wire [31:0]       dataInMem_hi_703 = {dataInMem_hi_hi_447, dataInMem_hi_lo_191};
  wire [31:0]       dataInMem_lo_576 = {dataInMem_lo_hi_320, dataInMem_lo_lo_64};
  wire [15:0]       dataInMem_hi_hi_448 = {dataRegroupBySew_7_57, dataRegroupBySew_6_57};
  wire [31:0]       dataInMem_hi_704 = {dataInMem_hi_hi_448, dataInMem_hi_lo_192};
  wire [31:0]       dataInMem_lo_577 = {dataInMem_lo_hi_321, dataInMem_lo_lo_65};
  wire [15:0]       dataInMem_hi_hi_449 = {dataRegroupBySew_7_58, dataRegroupBySew_6_58};
  wire [31:0]       dataInMem_hi_705 = {dataInMem_hi_hi_449, dataInMem_hi_lo_193};
  wire [31:0]       dataInMem_lo_578 = {dataInMem_lo_hi_322, dataInMem_lo_lo_66};
  wire [15:0]       dataInMem_hi_hi_450 = {dataRegroupBySew_7_59, dataRegroupBySew_6_59};
  wire [31:0]       dataInMem_hi_706 = {dataInMem_hi_hi_450, dataInMem_hi_lo_194};
  wire [31:0]       dataInMem_lo_579 = {dataInMem_lo_hi_323, dataInMem_lo_lo_67};
  wire [15:0]       dataInMem_hi_hi_451 = {dataRegroupBySew_7_60, dataRegroupBySew_6_60};
  wire [31:0]       dataInMem_hi_707 = {dataInMem_hi_hi_451, dataInMem_hi_lo_195};
  wire [31:0]       dataInMem_lo_580 = {dataInMem_lo_hi_324, dataInMem_lo_lo_68};
  wire [15:0]       dataInMem_hi_hi_452 = {dataRegroupBySew_7_61, dataRegroupBySew_6_61};
  wire [31:0]       dataInMem_hi_708 = {dataInMem_hi_hi_452, dataInMem_hi_lo_196};
  wire [31:0]       dataInMem_lo_581 = {dataInMem_lo_hi_325, dataInMem_lo_lo_69};
  wire [15:0]       dataInMem_hi_hi_453 = {dataRegroupBySew_7_62, dataRegroupBySew_6_62};
  wire [31:0]       dataInMem_hi_709 = {dataInMem_hi_hi_453, dataInMem_hi_lo_197};
  wire [31:0]       dataInMem_lo_582 = {dataInMem_lo_hi_326, dataInMem_lo_lo_70};
  wire [15:0]       dataInMem_hi_hi_454 = {dataRegroupBySew_7_63, dataRegroupBySew_6_63};
  wire [31:0]       dataInMem_hi_710 = {dataInMem_hi_hi_454, dataInMem_hi_lo_198};
  wire [31:0]       dataInMem_lo_583 = {dataInMem_lo_hi_327, dataInMem_lo_lo_71};
  wire [15:0]       dataInMem_hi_hi_455 = {dataRegroupBySew_7_64, dataRegroupBySew_6_64};
  wire [31:0]       dataInMem_hi_711 = {dataInMem_hi_hi_455, dataInMem_hi_lo_199};
  wire [31:0]       dataInMem_lo_584 = {dataInMem_lo_hi_328, dataInMem_lo_lo_72};
  wire [15:0]       dataInMem_hi_hi_456 = {dataRegroupBySew_7_65, dataRegroupBySew_6_65};
  wire [31:0]       dataInMem_hi_712 = {dataInMem_hi_hi_456, dataInMem_hi_lo_200};
  wire [31:0]       dataInMem_lo_585 = {dataInMem_lo_hi_329, dataInMem_lo_lo_73};
  wire [15:0]       dataInMem_hi_hi_457 = {dataRegroupBySew_7_66, dataRegroupBySew_6_66};
  wire [31:0]       dataInMem_hi_713 = {dataInMem_hi_hi_457, dataInMem_hi_lo_201};
  wire [31:0]       dataInMem_lo_586 = {dataInMem_lo_hi_330, dataInMem_lo_lo_74};
  wire [15:0]       dataInMem_hi_hi_458 = {dataRegroupBySew_7_67, dataRegroupBySew_6_67};
  wire [31:0]       dataInMem_hi_714 = {dataInMem_hi_hi_458, dataInMem_hi_lo_202};
  wire [31:0]       dataInMem_lo_587 = {dataInMem_lo_hi_331, dataInMem_lo_lo_75};
  wire [15:0]       dataInMem_hi_hi_459 = {dataRegroupBySew_7_68, dataRegroupBySew_6_68};
  wire [31:0]       dataInMem_hi_715 = {dataInMem_hi_hi_459, dataInMem_hi_lo_203};
  wire [31:0]       dataInMem_lo_588 = {dataInMem_lo_hi_332, dataInMem_lo_lo_76};
  wire [15:0]       dataInMem_hi_hi_460 = {dataRegroupBySew_7_69, dataRegroupBySew_6_69};
  wire [31:0]       dataInMem_hi_716 = {dataInMem_hi_hi_460, dataInMem_hi_lo_204};
  wire [31:0]       dataInMem_lo_589 = {dataInMem_lo_hi_333, dataInMem_lo_lo_77};
  wire [15:0]       dataInMem_hi_hi_461 = {dataRegroupBySew_7_70, dataRegroupBySew_6_70};
  wire [31:0]       dataInMem_hi_717 = {dataInMem_hi_hi_461, dataInMem_hi_lo_205};
  wire [31:0]       dataInMem_lo_590 = {dataInMem_lo_hi_334, dataInMem_lo_lo_78};
  wire [15:0]       dataInMem_hi_hi_462 = {dataRegroupBySew_7_71, dataRegroupBySew_6_71};
  wire [31:0]       dataInMem_hi_718 = {dataInMem_hi_hi_462, dataInMem_hi_lo_206};
  wire [31:0]       dataInMem_lo_591 = {dataInMem_lo_hi_335, dataInMem_lo_lo_79};
  wire [15:0]       dataInMem_hi_hi_463 = {dataRegroupBySew_7_72, dataRegroupBySew_6_72};
  wire [31:0]       dataInMem_hi_719 = {dataInMem_hi_hi_463, dataInMem_hi_lo_207};
  wire [31:0]       dataInMem_lo_592 = {dataInMem_lo_hi_336, dataInMem_lo_lo_80};
  wire [15:0]       dataInMem_hi_hi_464 = {dataRegroupBySew_7_73, dataRegroupBySew_6_73};
  wire [31:0]       dataInMem_hi_720 = {dataInMem_hi_hi_464, dataInMem_hi_lo_208};
  wire [31:0]       dataInMem_lo_593 = {dataInMem_lo_hi_337, dataInMem_lo_lo_81};
  wire [15:0]       dataInMem_hi_hi_465 = {dataRegroupBySew_7_74, dataRegroupBySew_6_74};
  wire [31:0]       dataInMem_hi_721 = {dataInMem_hi_hi_465, dataInMem_hi_lo_209};
  wire [31:0]       dataInMem_lo_594 = {dataInMem_lo_hi_338, dataInMem_lo_lo_82};
  wire [15:0]       dataInMem_hi_hi_466 = {dataRegroupBySew_7_75, dataRegroupBySew_6_75};
  wire [31:0]       dataInMem_hi_722 = {dataInMem_hi_hi_466, dataInMem_hi_lo_210};
  wire [31:0]       dataInMem_lo_595 = {dataInMem_lo_hi_339, dataInMem_lo_lo_83};
  wire [15:0]       dataInMem_hi_hi_467 = {dataRegroupBySew_7_76, dataRegroupBySew_6_76};
  wire [31:0]       dataInMem_hi_723 = {dataInMem_hi_hi_467, dataInMem_hi_lo_211};
  wire [31:0]       dataInMem_lo_596 = {dataInMem_lo_hi_340, dataInMem_lo_lo_84};
  wire [15:0]       dataInMem_hi_hi_468 = {dataRegroupBySew_7_77, dataRegroupBySew_6_77};
  wire [31:0]       dataInMem_hi_724 = {dataInMem_hi_hi_468, dataInMem_hi_lo_212};
  wire [31:0]       dataInMem_lo_597 = {dataInMem_lo_hi_341, dataInMem_lo_lo_85};
  wire [15:0]       dataInMem_hi_hi_469 = {dataRegroupBySew_7_78, dataRegroupBySew_6_78};
  wire [31:0]       dataInMem_hi_725 = {dataInMem_hi_hi_469, dataInMem_hi_lo_213};
  wire [31:0]       dataInMem_lo_598 = {dataInMem_lo_hi_342, dataInMem_lo_lo_86};
  wire [15:0]       dataInMem_hi_hi_470 = {dataRegroupBySew_7_79, dataRegroupBySew_6_79};
  wire [31:0]       dataInMem_hi_726 = {dataInMem_hi_hi_470, dataInMem_hi_lo_214};
  wire [31:0]       dataInMem_lo_599 = {dataInMem_lo_hi_343, dataInMem_lo_lo_87};
  wire [15:0]       dataInMem_hi_hi_471 = {dataRegroupBySew_7_80, dataRegroupBySew_6_80};
  wire [31:0]       dataInMem_hi_727 = {dataInMem_hi_hi_471, dataInMem_hi_lo_215};
  wire [31:0]       dataInMem_lo_600 = {dataInMem_lo_hi_344, dataInMem_lo_lo_88};
  wire [15:0]       dataInMem_hi_hi_472 = {dataRegroupBySew_7_81, dataRegroupBySew_6_81};
  wire [31:0]       dataInMem_hi_728 = {dataInMem_hi_hi_472, dataInMem_hi_lo_216};
  wire [31:0]       dataInMem_lo_601 = {dataInMem_lo_hi_345, dataInMem_lo_lo_89};
  wire [15:0]       dataInMem_hi_hi_473 = {dataRegroupBySew_7_82, dataRegroupBySew_6_82};
  wire [31:0]       dataInMem_hi_729 = {dataInMem_hi_hi_473, dataInMem_hi_lo_217};
  wire [31:0]       dataInMem_lo_602 = {dataInMem_lo_hi_346, dataInMem_lo_lo_90};
  wire [15:0]       dataInMem_hi_hi_474 = {dataRegroupBySew_7_83, dataRegroupBySew_6_83};
  wire [31:0]       dataInMem_hi_730 = {dataInMem_hi_hi_474, dataInMem_hi_lo_218};
  wire [31:0]       dataInMem_lo_603 = {dataInMem_lo_hi_347, dataInMem_lo_lo_91};
  wire [15:0]       dataInMem_hi_hi_475 = {dataRegroupBySew_7_84, dataRegroupBySew_6_84};
  wire [31:0]       dataInMem_hi_731 = {dataInMem_hi_hi_475, dataInMem_hi_lo_219};
  wire [31:0]       dataInMem_lo_604 = {dataInMem_lo_hi_348, dataInMem_lo_lo_92};
  wire [15:0]       dataInMem_hi_hi_476 = {dataRegroupBySew_7_85, dataRegroupBySew_6_85};
  wire [31:0]       dataInMem_hi_732 = {dataInMem_hi_hi_476, dataInMem_hi_lo_220};
  wire [31:0]       dataInMem_lo_605 = {dataInMem_lo_hi_349, dataInMem_lo_lo_93};
  wire [15:0]       dataInMem_hi_hi_477 = {dataRegroupBySew_7_86, dataRegroupBySew_6_86};
  wire [31:0]       dataInMem_hi_733 = {dataInMem_hi_hi_477, dataInMem_hi_lo_221};
  wire [31:0]       dataInMem_lo_606 = {dataInMem_lo_hi_350, dataInMem_lo_lo_94};
  wire [15:0]       dataInMem_hi_hi_478 = {dataRegroupBySew_7_87, dataRegroupBySew_6_87};
  wire [31:0]       dataInMem_hi_734 = {dataInMem_hi_hi_478, dataInMem_hi_lo_222};
  wire [31:0]       dataInMem_lo_607 = {dataInMem_lo_hi_351, dataInMem_lo_lo_95};
  wire [15:0]       dataInMem_hi_hi_479 = {dataRegroupBySew_7_88, dataRegroupBySew_6_88};
  wire [31:0]       dataInMem_hi_735 = {dataInMem_hi_hi_479, dataInMem_hi_lo_223};
  wire [31:0]       dataInMem_lo_608 = {dataInMem_lo_hi_352, dataInMem_lo_lo_96};
  wire [15:0]       dataInMem_hi_hi_480 = {dataRegroupBySew_7_89, dataRegroupBySew_6_89};
  wire [31:0]       dataInMem_hi_736 = {dataInMem_hi_hi_480, dataInMem_hi_lo_224};
  wire [31:0]       dataInMem_lo_609 = {dataInMem_lo_hi_353, dataInMem_lo_lo_97};
  wire [15:0]       dataInMem_hi_hi_481 = {dataRegroupBySew_7_90, dataRegroupBySew_6_90};
  wire [31:0]       dataInMem_hi_737 = {dataInMem_hi_hi_481, dataInMem_hi_lo_225};
  wire [31:0]       dataInMem_lo_610 = {dataInMem_lo_hi_354, dataInMem_lo_lo_98};
  wire [15:0]       dataInMem_hi_hi_482 = {dataRegroupBySew_7_91, dataRegroupBySew_6_91};
  wire [31:0]       dataInMem_hi_738 = {dataInMem_hi_hi_482, dataInMem_hi_lo_226};
  wire [31:0]       dataInMem_lo_611 = {dataInMem_lo_hi_355, dataInMem_lo_lo_99};
  wire [15:0]       dataInMem_hi_hi_483 = {dataRegroupBySew_7_92, dataRegroupBySew_6_92};
  wire [31:0]       dataInMem_hi_739 = {dataInMem_hi_hi_483, dataInMem_hi_lo_227};
  wire [31:0]       dataInMem_lo_612 = {dataInMem_lo_hi_356, dataInMem_lo_lo_100};
  wire [15:0]       dataInMem_hi_hi_484 = {dataRegroupBySew_7_93, dataRegroupBySew_6_93};
  wire [31:0]       dataInMem_hi_740 = {dataInMem_hi_hi_484, dataInMem_hi_lo_228};
  wire [31:0]       dataInMem_lo_613 = {dataInMem_lo_hi_357, dataInMem_lo_lo_101};
  wire [15:0]       dataInMem_hi_hi_485 = {dataRegroupBySew_7_94, dataRegroupBySew_6_94};
  wire [31:0]       dataInMem_hi_741 = {dataInMem_hi_hi_485, dataInMem_hi_lo_229};
  wire [31:0]       dataInMem_lo_614 = {dataInMem_lo_hi_358, dataInMem_lo_lo_102};
  wire [15:0]       dataInMem_hi_hi_486 = {dataRegroupBySew_7_95, dataRegroupBySew_6_95};
  wire [31:0]       dataInMem_hi_742 = {dataInMem_hi_hi_486, dataInMem_hi_lo_230};
  wire [31:0]       dataInMem_lo_615 = {dataInMem_lo_hi_359, dataInMem_lo_lo_103};
  wire [15:0]       dataInMem_hi_hi_487 = {dataRegroupBySew_7_96, dataRegroupBySew_6_96};
  wire [31:0]       dataInMem_hi_743 = {dataInMem_hi_hi_487, dataInMem_hi_lo_231};
  wire [31:0]       dataInMem_lo_616 = {dataInMem_lo_hi_360, dataInMem_lo_lo_104};
  wire [15:0]       dataInMem_hi_hi_488 = {dataRegroupBySew_7_97, dataRegroupBySew_6_97};
  wire [31:0]       dataInMem_hi_744 = {dataInMem_hi_hi_488, dataInMem_hi_lo_232};
  wire [31:0]       dataInMem_lo_617 = {dataInMem_lo_hi_361, dataInMem_lo_lo_105};
  wire [15:0]       dataInMem_hi_hi_489 = {dataRegroupBySew_7_98, dataRegroupBySew_6_98};
  wire [31:0]       dataInMem_hi_745 = {dataInMem_hi_hi_489, dataInMem_hi_lo_233};
  wire [31:0]       dataInMem_lo_618 = {dataInMem_lo_hi_362, dataInMem_lo_lo_106};
  wire [15:0]       dataInMem_hi_hi_490 = {dataRegroupBySew_7_99, dataRegroupBySew_6_99};
  wire [31:0]       dataInMem_hi_746 = {dataInMem_hi_hi_490, dataInMem_hi_lo_234};
  wire [31:0]       dataInMem_lo_619 = {dataInMem_lo_hi_363, dataInMem_lo_lo_107};
  wire [15:0]       dataInMem_hi_hi_491 = {dataRegroupBySew_7_100, dataRegroupBySew_6_100};
  wire [31:0]       dataInMem_hi_747 = {dataInMem_hi_hi_491, dataInMem_hi_lo_235};
  wire [31:0]       dataInMem_lo_620 = {dataInMem_lo_hi_364, dataInMem_lo_lo_108};
  wire [15:0]       dataInMem_hi_hi_492 = {dataRegroupBySew_7_101, dataRegroupBySew_6_101};
  wire [31:0]       dataInMem_hi_748 = {dataInMem_hi_hi_492, dataInMem_hi_lo_236};
  wire [31:0]       dataInMem_lo_621 = {dataInMem_lo_hi_365, dataInMem_lo_lo_109};
  wire [15:0]       dataInMem_hi_hi_493 = {dataRegroupBySew_7_102, dataRegroupBySew_6_102};
  wire [31:0]       dataInMem_hi_749 = {dataInMem_hi_hi_493, dataInMem_hi_lo_237};
  wire [31:0]       dataInMem_lo_622 = {dataInMem_lo_hi_366, dataInMem_lo_lo_110};
  wire [15:0]       dataInMem_hi_hi_494 = {dataRegroupBySew_7_103, dataRegroupBySew_6_103};
  wire [31:0]       dataInMem_hi_750 = {dataInMem_hi_hi_494, dataInMem_hi_lo_238};
  wire [31:0]       dataInMem_lo_623 = {dataInMem_lo_hi_367, dataInMem_lo_lo_111};
  wire [15:0]       dataInMem_hi_hi_495 = {dataRegroupBySew_7_104, dataRegroupBySew_6_104};
  wire [31:0]       dataInMem_hi_751 = {dataInMem_hi_hi_495, dataInMem_hi_lo_239};
  wire [31:0]       dataInMem_lo_624 = {dataInMem_lo_hi_368, dataInMem_lo_lo_112};
  wire [15:0]       dataInMem_hi_hi_496 = {dataRegroupBySew_7_105, dataRegroupBySew_6_105};
  wire [31:0]       dataInMem_hi_752 = {dataInMem_hi_hi_496, dataInMem_hi_lo_240};
  wire [31:0]       dataInMem_lo_625 = {dataInMem_lo_hi_369, dataInMem_lo_lo_113};
  wire [15:0]       dataInMem_hi_hi_497 = {dataRegroupBySew_7_106, dataRegroupBySew_6_106};
  wire [31:0]       dataInMem_hi_753 = {dataInMem_hi_hi_497, dataInMem_hi_lo_241};
  wire [31:0]       dataInMem_lo_626 = {dataInMem_lo_hi_370, dataInMem_lo_lo_114};
  wire [15:0]       dataInMem_hi_hi_498 = {dataRegroupBySew_7_107, dataRegroupBySew_6_107};
  wire [31:0]       dataInMem_hi_754 = {dataInMem_hi_hi_498, dataInMem_hi_lo_242};
  wire [31:0]       dataInMem_lo_627 = {dataInMem_lo_hi_371, dataInMem_lo_lo_115};
  wire [15:0]       dataInMem_hi_hi_499 = {dataRegroupBySew_7_108, dataRegroupBySew_6_108};
  wire [31:0]       dataInMem_hi_755 = {dataInMem_hi_hi_499, dataInMem_hi_lo_243};
  wire [31:0]       dataInMem_lo_628 = {dataInMem_lo_hi_372, dataInMem_lo_lo_116};
  wire [15:0]       dataInMem_hi_hi_500 = {dataRegroupBySew_7_109, dataRegroupBySew_6_109};
  wire [31:0]       dataInMem_hi_756 = {dataInMem_hi_hi_500, dataInMem_hi_lo_244};
  wire [31:0]       dataInMem_lo_629 = {dataInMem_lo_hi_373, dataInMem_lo_lo_117};
  wire [15:0]       dataInMem_hi_hi_501 = {dataRegroupBySew_7_110, dataRegroupBySew_6_110};
  wire [31:0]       dataInMem_hi_757 = {dataInMem_hi_hi_501, dataInMem_hi_lo_245};
  wire [31:0]       dataInMem_lo_630 = {dataInMem_lo_hi_374, dataInMem_lo_lo_118};
  wire [15:0]       dataInMem_hi_hi_502 = {dataRegroupBySew_7_111, dataRegroupBySew_6_111};
  wire [31:0]       dataInMem_hi_758 = {dataInMem_hi_hi_502, dataInMem_hi_lo_246};
  wire [31:0]       dataInMem_lo_631 = {dataInMem_lo_hi_375, dataInMem_lo_lo_119};
  wire [15:0]       dataInMem_hi_hi_503 = {dataRegroupBySew_7_112, dataRegroupBySew_6_112};
  wire [31:0]       dataInMem_hi_759 = {dataInMem_hi_hi_503, dataInMem_hi_lo_247};
  wire [31:0]       dataInMem_lo_632 = {dataInMem_lo_hi_376, dataInMem_lo_lo_120};
  wire [15:0]       dataInMem_hi_hi_504 = {dataRegroupBySew_7_113, dataRegroupBySew_6_113};
  wire [31:0]       dataInMem_hi_760 = {dataInMem_hi_hi_504, dataInMem_hi_lo_248};
  wire [31:0]       dataInMem_lo_633 = {dataInMem_lo_hi_377, dataInMem_lo_lo_121};
  wire [15:0]       dataInMem_hi_hi_505 = {dataRegroupBySew_7_114, dataRegroupBySew_6_114};
  wire [31:0]       dataInMem_hi_761 = {dataInMem_hi_hi_505, dataInMem_hi_lo_249};
  wire [31:0]       dataInMem_lo_634 = {dataInMem_lo_hi_378, dataInMem_lo_lo_122};
  wire [15:0]       dataInMem_hi_hi_506 = {dataRegroupBySew_7_115, dataRegroupBySew_6_115};
  wire [31:0]       dataInMem_hi_762 = {dataInMem_hi_hi_506, dataInMem_hi_lo_250};
  wire [31:0]       dataInMem_lo_635 = {dataInMem_lo_hi_379, dataInMem_lo_lo_123};
  wire [15:0]       dataInMem_hi_hi_507 = {dataRegroupBySew_7_116, dataRegroupBySew_6_116};
  wire [31:0]       dataInMem_hi_763 = {dataInMem_hi_hi_507, dataInMem_hi_lo_251};
  wire [31:0]       dataInMem_lo_636 = {dataInMem_lo_hi_380, dataInMem_lo_lo_124};
  wire [15:0]       dataInMem_hi_hi_508 = {dataRegroupBySew_7_117, dataRegroupBySew_6_117};
  wire [31:0]       dataInMem_hi_764 = {dataInMem_hi_hi_508, dataInMem_hi_lo_252};
  wire [31:0]       dataInMem_lo_637 = {dataInMem_lo_hi_381, dataInMem_lo_lo_125};
  wire [15:0]       dataInMem_hi_hi_509 = {dataRegroupBySew_7_118, dataRegroupBySew_6_118};
  wire [31:0]       dataInMem_hi_765 = {dataInMem_hi_hi_509, dataInMem_hi_lo_253};
  wire [31:0]       dataInMem_lo_638 = {dataInMem_lo_hi_382, dataInMem_lo_lo_126};
  wire [15:0]       dataInMem_hi_hi_510 = {dataRegroupBySew_7_119, dataRegroupBySew_6_119};
  wire [31:0]       dataInMem_hi_766 = {dataInMem_hi_hi_510, dataInMem_hi_lo_254};
  wire [31:0]       dataInMem_lo_639 = {dataInMem_lo_hi_383, dataInMem_lo_lo_127};
  wire [15:0]       dataInMem_hi_hi_511 = {dataRegroupBySew_7_120, dataRegroupBySew_6_120};
  wire [31:0]       dataInMem_hi_767 = {dataInMem_hi_hi_511, dataInMem_hi_lo_255};
  wire [31:0]       dataInMem_lo_640 = {dataInMem_lo_hi_384, dataInMem_lo_lo_128};
  wire [15:0]       dataInMem_hi_hi_512 = {dataRegroupBySew_7_121, dataRegroupBySew_6_121};
  wire [31:0]       dataInMem_hi_768 = {dataInMem_hi_hi_512, dataInMem_hi_lo_256};
  wire [31:0]       dataInMem_lo_641 = {dataInMem_lo_hi_385, dataInMem_lo_lo_129};
  wire [15:0]       dataInMem_hi_hi_513 = {dataRegroupBySew_7_122, dataRegroupBySew_6_122};
  wire [31:0]       dataInMem_hi_769 = {dataInMem_hi_hi_513, dataInMem_hi_lo_257};
  wire [31:0]       dataInMem_lo_642 = {dataInMem_lo_hi_386, dataInMem_lo_lo_130};
  wire [15:0]       dataInMem_hi_hi_514 = {dataRegroupBySew_7_123, dataRegroupBySew_6_123};
  wire [31:0]       dataInMem_hi_770 = {dataInMem_hi_hi_514, dataInMem_hi_lo_258};
  wire [31:0]       dataInMem_lo_643 = {dataInMem_lo_hi_387, dataInMem_lo_lo_131};
  wire [15:0]       dataInMem_hi_hi_515 = {dataRegroupBySew_7_124, dataRegroupBySew_6_124};
  wire [31:0]       dataInMem_hi_771 = {dataInMem_hi_hi_515, dataInMem_hi_lo_259};
  wire [31:0]       dataInMem_lo_644 = {dataInMem_lo_hi_388, dataInMem_lo_lo_132};
  wire [15:0]       dataInMem_hi_hi_516 = {dataRegroupBySew_7_125, dataRegroupBySew_6_125};
  wire [31:0]       dataInMem_hi_772 = {dataInMem_hi_hi_516, dataInMem_hi_lo_260};
  wire [31:0]       dataInMem_lo_645 = {dataInMem_lo_hi_389, dataInMem_lo_lo_133};
  wire [15:0]       dataInMem_hi_hi_517 = {dataRegroupBySew_7_126, dataRegroupBySew_6_126};
  wire [31:0]       dataInMem_hi_773 = {dataInMem_hi_hi_517, dataInMem_hi_lo_261};
  wire [31:0]       dataInMem_lo_646 = {dataInMem_lo_hi_390, dataInMem_lo_lo_134};
  wire [15:0]       dataInMem_hi_hi_518 = {dataRegroupBySew_7_127, dataRegroupBySew_6_127};
  wire [31:0]       dataInMem_hi_774 = {dataInMem_hi_hi_518, dataInMem_hi_lo_262};
  wire [127:0]      dataInMem_lo_lo_lo_lo_lo_lo_7 = {dataInMem_hi_648, dataInMem_lo_520, dataInMem_hi_647, dataInMem_lo_519};
  wire [127:0]      dataInMem_lo_lo_lo_lo_lo_hi_7 = {dataInMem_hi_650, dataInMem_lo_522, dataInMem_hi_649, dataInMem_lo_521};
  wire [255:0]      dataInMem_lo_lo_lo_lo_lo_7 = {dataInMem_lo_lo_lo_lo_lo_hi_7, dataInMem_lo_lo_lo_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_lo_lo_lo_hi_lo_7 = {dataInMem_hi_652, dataInMem_lo_524, dataInMem_hi_651, dataInMem_lo_523};
  wire [127:0]      dataInMem_lo_lo_lo_lo_hi_hi_7 = {dataInMem_hi_654, dataInMem_lo_526, dataInMem_hi_653, dataInMem_lo_525};
  wire [255:0]      dataInMem_lo_lo_lo_lo_hi_7 = {dataInMem_lo_lo_lo_lo_hi_hi_7, dataInMem_lo_lo_lo_lo_hi_lo_7};
  wire [511:0]      dataInMem_lo_lo_lo_lo_7 = {dataInMem_lo_lo_lo_lo_hi_7, dataInMem_lo_lo_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_lo_lo_hi_lo_lo_7 = {dataInMem_hi_656, dataInMem_lo_528, dataInMem_hi_655, dataInMem_lo_527};
  wire [127:0]      dataInMem_lo_lo_lo_hi_lo_hi_7 = {dataInMem_hi_658, dataInMem_lo_530, dataInMem_hi_657, dataInMem_lo_529};
  wire [255:0]      dataInMem_lo_lo_lo_hi_lo_7 = {dataInMem_lo_lo_lo_hi_lo_hi_7, dataInMem_lo_lo_lo_hi_lo_lo_7};
  wire [127:0]      dataInMem_lo_lo_lo_hi_hi_lo_7 = {dataInMem_hi_660, dataInMem_lo_532, dataInMem_hi_659, dataInMem_lo_531};
  wire [127:0]      dataInMem_lo_lo_lo_hi_hi_hi_7 = {dataInMem_hi_662, dataInMem_lo_534, dataInMem_hi_661, dataInMem_lo_533};
  wire [255:0]      dataInMem_lo_lo_lo_hi_hi_7 = {dataInMem_lo_lo_lo_hi_hi_hi_7, dataInMem_lo_lo_lo_hi_hi_lo_7};
  wire [511:0]      dataInMem_lo_lo_lo_hi_7 = {dataInMem_lo_lo_lo_hi_hi_7, dataInMem_lo_lo_lo_hi_lo_7};
  wire [1023:0]     dataInMem_lo_lo_lo_7 = {dataInMem_lo_lo_lo_hi_7, dataInMem_lo_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_lo_hi_lo_lo_lo_7 = {dataInMem_hi_664, dataInMem_lo_536, dataInMem_hi_663, dataInMem_lo_535};
  wire [127:0]      dataInMem_lo_lo_hi_lo_lo_hi_7 = {dataInMem_hi_666, dataInMem_lo_538, dataInMem_hi_665, dataInMem_lo_537};
  wire [255:0]      dataInMem_lo_lo_hi_lo_lo_7 = {dataInMem_lo_lo_hi_lo_lo_hi_7, dataInMem_lo_lo_hi_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_lo_hi_lo_hi_lo_7 = {dataInMem_hi_668, dataInMem_lo_540, dataInMem_hi_667, dataInMem_lo_539};
  wire [127:0]      dataInMem_lo_lo_hi_lo_hi_hi_7 = {dataInMem_hi_670, dataInMem_lo_542, dataInMem_hi_669, dataInMem_lo_541};
  wire [255:0]      dataInMem_lo_lo_hi_lo_hi_7 = {dataInMem_lo_lo_hi_lo_hi_hi_7, dataInMem_lo_lo_hi_lo_hi_lo_7};
  wire [511:0]      dataInMem_lo_lo_hi_lo_7 = {dataInMem_lo_lo_hi_lo_hi_7, dataInMem_lo_lo_hi_lo_lo_7};
  wire [127:0]      dataInMem_lo_lo_hi_hi_lo_lo_7 = {dataInMem_hi_672, dataInMem_lo_544, dataInMem_hi_671, dataInMem_lo_543};
  wire [127:0]      dataInMem_lo_lo_hi_hi_lo_hi_7 = {dataInMem_hi_674, dataInMem_lo_546, dataInMem_hi_673, dataInMem_lo_545};
  wire [255:0]      dataInMem_lo_lo_hi_hi_lo_7 = {dataInMem_lo_lo_hi_hi_lo_hi_7, dataInMem_lo_lo_hi_hi_lo_lo_7};
  wire [127:0]      dataInMem_lo_lo_hi_hi_hi_lo_7 = {dataInMem_hi_676, dataInMem_lo_548, dataInMem_hi_675, dataInMem_lo_547};
  wire [127:0]      dataInMem_lo_lo_hi_hi_hi_hi_7 = {dataInMem_hi_678, dataInMem_lo_550, dataInMem_hi_677, dataInMem_lo_549};
  wire [255:0]      dataInMem_lo_lo_hi_hi_hi_7 = {dataInMem_lo_lo_hi_hi_hi_hi_7, dataInMem_lo_lo_hi_hi_hi_lo_7};
  wire [511:0]      dataInMem_lo_lo_hi_hi_7 = {dataInMem_lo_lo_hi_hi_hi_7, dataInMem_lo_lo_hi_hi_lo_7};
  wire [1023:0]     dataInMem_lo_lo_hi_7 = {dataInMem_lo_lo_hi_hi_7, dataInMem_lo_lo_hi_lo_7};
  wire [2047:0]     dataInMem_lo_lo_135 = {dataInMem_lo_lo_hi_7, dataInMem_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_lo_lo_lo_lo_7 = {dataInMem_hi_680, dataInMem_lo_552, dataInMem_hi_679, dataInMem_lo_551};
  wire [127:0]      dataInMem_lo_hi_lo_lo_lo_hi_7 = {dataInMem_hi_682, dataInMem_lo_554, dataInMem_hi_681, dataInMem_lo_553};
  wire [255:0]      dataInMem_lo_hi_lo_lo_lo_7 = {dataInMem_lo_hi_lo_lo_lo_hi_7, dataInMem_lo_hi_lo_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_lo_lo_hi_lo_7 = {dataInMem_hi_684, dataInMem_lo_556, dataInMem_hi_683, dataInMem_lo_555};
  wire [127:0]      dataInMem_lo_hi_lo_lo_hi_hi_7 = {dataInMem_hi_686, dataInMem_lo_558, dataInMem_hi_685, dataInMem_lo_557};
  wire [255:0]      dataInMem_lo_hi_lo_lo_hi_7 = {dataInMem_lo_hi_lo_lo_hi_hi_7, dataInMem_lo_hi_lo_lo_hi_lo_7};
  wire [511:0]      dataInMem_lo_hi_lo_lo_7 = {dataInMem_lo_hi_lo_lo_hi_7, dataInMem_lo_hi_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_lo_hi_lo_lo_7 = {dataInMem_hi_688, dataInMem_lo_560, dataInMem_hi_687, dataInMem_lo_559};
  wire [127:0]      dataInMem_lo_hi_lo_hi_lo_hi_7 = {dataInMem_hi_690, dataInMem_lo_562, dataInMem_hi_689, dataInMem_lo_561};
  wire [255:0]      dataInMem_lo_hi_lo_hi_lo_7 = {dataInMem_lo_hi_lo_hi_lo_hi_7, dataInMem_lo_hi_lo_hi_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_lo_hi_hi_lo_7 = {dataInMem_hi_692, dataInMem_lo_564, dataInMem_hi_691, dataInMem_lo_563};
  wire [127:0]      dataInMem_lo_hi_lo_hi_hi_hi_7 = {dataInMem_hi_694, dataInMem_lo_566, dataInMem_hi_693, dataInMem_lo_565};
  wire [255:0]      dataInMem_lo_hi_lo_hi_hi_7 = {dataInMem_lo_hi_lo_hi_hi_hi_7, dataInMem_lo_hi_lo_hi_hi_lo_7};
  wire [511:0]      dataInMem_lo_hi_lo_hi_7 = {dataInMem_lo_hi_lo_hi_hi_7, dataInMem_lo_hi_lo_hi_lo_7};
  wire [1023:0]     dataInMem_lo_hi_lo_7 = {dataInMem_lo_hi_lo_hi_7, dataInMem_lo_hi_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_hi_lo_lo_lo_7 = {dataInMem_hi_696, dataInMem_lo_568, dataInMem_hi_695, dataInMem_lo_567};
  wire [127:0]      dataInMem_lo_hi_hi_lo_lo_hi_7 = {dataInMem_hi_698, dataInMem_lo_570, dataInMem_hi_697, dataInMem_lo_569};
  wire [255:0]      dataInMem_lo_hi_hi_lo_lo_7 = {dataInMem_lo_hi_hi_lo_lo_hi_7, dataInMem_lo_hi_hi_lo_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_hi_lo_hi_lo_7 = {dataInMem_hi_700, dataInMem_lo_572, dataInMem_hi_699, dataInMem_lo_571};
  wire [127:0]      dataInMem_lo_hi_hi_lo_hi_hi_7 = {dataInMem_hi_702, dataInMem_lo_574, dataInMem_hi_701, dataInMem_lo_573};
  wire [255:0]      dataInMem_lo_hi_hi_lo_hi_7 = {dataInMem_lo_hi_hi_lo_hi_hi_7, dataInMem_lo_hi_hi_lo_hi_lo_7};
  wire [511:0]      dataInMem_lo_hi_hi_lo_7 = {dataInMem_lo_hi_hi_lo_hi_7, dataInMem_lo_hi_hi_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_hi_hi_lo_lo_7 = {dataInMem_hi_704, dataInMem_lo_576, dataInMem_hi_703, dataInMem_lo_575};
  wire [127:0]      dataInMem_lo_hi_hi_hi_lo_hi_7 = {dataInMem_hi_706, dataInMem_lo_578, dataInMem_hi_705, dataInMem_lo_577};
  wire [255:0]      dataInMem_lo_hi_hi_hi_lo_7 = {dataInMem_lo_hi_hi_hi_lo_hi_7, dataInMem_lo_hi_hi_hi_lo_lo_7};
  wire [127:0]      dataInMem_lo_hi_hi_hi_hi_lo_7 = {dataInMem_hi_708, dataInMem_lo_580, dataInMem_hi_707, dataInMem_lo_579};
  wire [127:0]      dataInMem_lo_hi_hi_hi_hi_hi_7 = {dataInMem_hi_710, dataInMem_lo_582, dataInMem_hi_709, dataInMem_lo_581};
  wire [255:0]      dataInMem_lo_hi_hi_hi_hi_7 = {dataInMem_lo_hi_hi_hi_hi_hi_7, dataInMem_lo_hi_hi_hi_hi_lo_7};
  wire [511:0]      dataInMem_lo_hi_hi_hi_7 = {dataInMem_lo_hi_hi_hi_hi_7, dataInMem_lo_hi_hi_hi_lo_7};
  wire [1023:0]     dataInMem_lo_hi_hi_7 = {dataInMem_lo_hi_hi_hi_7, dataInMem_lo_hi_hi_lo_7};
  wire [2047:0]     dataInMem_lo_hi_391 = {dataInMem_lo_hi_hi_7, dataInMem_lo_hi_lo_7};
  wire [4095:0]     dataInMem_lo_647 = {dataInMem_lo_hi_391, dataInMem_lo_lo_135};
  wire [127:0]      dataInMem_hi_lo_lo_lo_lo_lo_7 = {dataInMem_hi_712, dataInMem_lo_584, dataInMem_hi_711, dataInMem_lo_583};
  wire [127:0]      dataInMem_hi_lo_lo_lo_lo_hi_7 = {dataInMem_hi_714, dataInMem_lo_586, dataInMem_hi_713, dataInMem_lo_585};
  wire [255:0]      dataInMem_hi_lo_lo_lo_lo_7 = {dataInMem_hi_lo_lo_lo_lo_hi_7, dataInMem_hi_lo_lo_lo_lo_lo_7};
  wire [127:0]      dataInMem_hi_lo_lo_lo_hi_lo_7 = {dataInMem_hi_716, dataInMem_lo_588, dataInMem_hi_715, dataInMem_lo_587};
  wire [127:0]      dataInMem_hi_lo_lo_lo_hi_hi_7 = {dataInMem_hi_718, dataInMem_lo_590, dataInMem_hi_717, dataInMem_lo_589};
  wire [255:0]      dataInMem_hi_lo_lo_lo_hi_7 = {dataInMem_hi_lo_lo_lo_hi_hi_7, dataInMem_hi_lo_lo_lo_hi_lo_7};
  wire [511:0]      dataInMem_hi_lo_lo_lo_7 = {dataInMem_hi_lo_lo_lo_hi_7, dataInMem_hi_lo_lo_lo_lo_7};
  wire [127:0]      dataInMem_hi_lo_lo_hi_lo_lo_7 = {dataInMem_hi_720, dataInMem_lo_592, dataInMem_hi_719, dataInMem_lo_591};
  wire [127:0]      dataInMem_hi_lo_lo_hi_lo_hi_7 = {dataInMem_hi_722, dataInMem_lo_594, dataInMem_hi_721, dataInMem_lo_593};
  wire [255:0]      dataInMem_hi_lo_lo_hi_lo_7 = {dataInMem_hi_lo_lo_hi_lo_hi_7, dataInMem_hi_lo_lo_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_lo_lo_hi_hi_lo_7 = {dataInMem_hi_724, dataInMem_lo_596, dataInMem_hi_723, dataInMem_lo_595};
  wire [127:0]      dataInMem_hi_lo_lo_hi_hi_hi_7 = {dataInMem_hi_726, dataInMem_lo_598, dataInMem_hi_725, dataInMem_lo_597};
  wire [255:0]      dataInMem_hi_lo_lo_hi_hi_7 = {dataInMem_hi_lo_lo_hi_hi_hi_7, dataInMem_hi_lo_lo_hi_hi_lo_7};
  wire [511:0]      dataInMem_hi_lo_lo_hi_7 = {dataInMem_hi_lo_lo_hi_hi_7, dataInMem_hi_lo_lo_hi_lo_7};
  wire [1023:0]     dataInMem_hi_lo_lo_7 = {dataInMem_hi_lo_lo_hi_7, dataInMem_hi_lo_lo_lo_7};
  wire [127:0]      dataInMem_hi_lo_hi_lo_lo_lo_7 = {dataInMem_hi_728, dataInMem_lo_600, dataInMem_hi_727, dataInMem_lo_599};
  wire [127:0]      dataInMem_hi_lo_hi_lo_lo_hi_7 = {dataInMem_hi_730, dataInMem_lo_602, dataInMem_hi_729, dataInMem_lo_601};
  wire [255:0]      dataInMem_hi_lo_hi_lo_lo_7 = {dataInMem_hi_lo_hi_lo_lo_hi_7, dataInMem_hi_lo_hi_lo_lo_lo_7};
  wire [127:0]      dataInMem_hi_lo_hi_lo_hi_lo_7 = {dataInMem_hi_732, dataInMem_lo_604, dataInMem_hi_731, dataInMem_lo_603};
  wire [127:0]      dataInMem_hi_lo_hi_lo_hi_hi_7 = {dataInMem_hi_734, dataInMem_lo_606, dataInMem_hi_733, dataInMem_lo_605};
  wire [255:0]      dataInMem_hi_lo_hi_lo_hi_7 = {dataInMem_hi_lo_hi_lo_hi_hi_7, dataInMem_hi_lo_hi_lo_hi_lo_7};
  wire [511:0]      dataInMem_hi_lo_hi_lo_7 = {dataInMem_hi_lo_hi_lo_hi_7, dataInMem_hi_lo_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_lo_hi_hi_lo_lo_7 = {dataInMem_hi_736, dataInMem_lo_608, dataInMem_hi_735, dataInMem_lo_607};
  wire [127:0]      dataInMem_hi_lo_hi_hi_lo_hi_7 = {dataInMem_hi_738, dataInMem_lo_610, dataInMem_hi_737, dataInMem_lo_609};
  wire [255:0]      dataInMem_hi_lo_hi_hi_lo_7 = {dataInMem_hi_lo_hi_hi_lo_hi_7, dataInMem_hi_lo_hi_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_lo_hi_hi_hi_lo_7 = {dataInMem_hi_740, dataInMem_lo_612, dataInMem_hi_739, dataInMem_lo_611};
  wire [127:0]      dataInMem_hi_lo_hi_hi_hi_hi_7 = {dataInMem_hi_742, dataInMem_lo_614, dataInMem_hi_741, dataInMem_lo_613};
  wire [255:0]      dataInMem_hi_lo_hi_hi_hi_7 = {dataInMem_hi_lo_hi_hi_hi_hi_7, dataInMem_hi_lo_hi_hi_hi_lo_7};
  wire [511:0]      dataInMem_hi_lo_hi_hi_7 = {dataInMem_hi_lo_hi_hi_hi_7, dataInMem_hi_lo_hi_hi_lo_7};
  wire [1023:0]     dataInMem_hi_lo_hi_7 = {dataInMem_hi_lo_hi_hi_7, dataInMem_hi_lo_hi_lo_7};
  wire [2047:0]     dataInMem_hi_lo_263 = {dataInMem_hi_lo_hi_7, dataInMem_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_lo_lo_lo_lo_7 = {dataInMem_hi_744, dataInMem_lo_616, dataInMem_hi_743, dataInMem_lo_615};
  wire [127:0]      dataInMem_hi_hi_lo_lo_lo_hi_7 = {dataInMem_hi_746, dataInMem_lo_618, dataInMem_hi_745, dataInMem_lo_617};
  wire [255:0]      dataInMem_hi_hi_lo_lo_lo_7 = {dataInMem_hi_hi_lo_lo_lo_hi_7, dataInMem_hi_hi_lo_lo_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_lo_lo_hi_lo_7 = {dataInMem_hi_748, dataInMem_lo_620, dataInMem_hi_747, dataInMem_lo_619};
  wire [127:0]      dataInMem_hi_hi_lo_lo_hi_hi_7 = {dataInMem_hi_750, dataInMem_lo_622, dataInMem_hi_749, dataInMem_lo_621};
  wire [255:0]      dataInMem_hi_hi_lo_lo_hi_7 = {dataInMem_hi_hi_lo_lo_hi_hi_7, dataInMem_hi_hi_lo_lo_hi_lo_7};
  wire [511:0]      dataInMem_hi_hi_lo_lo_7 = {dataInMem_hi_hi_lo_lo_hi_7, dataInMem_hi_hi_lo_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_lo_hi_lo_lo_7 = {dataInMem_hi_752, dataInMem_lo_624, dataInMem_hi_751, dataInMem_lo_623};
  wire [127:0]      dataInMem_hi_hi_lo_hi_lo_hi_7 = {dataInMem_hi_754, dataInMem_lo_626, dataInMem_hi_753, dataInMem_lo_625};
  wire [255:0]      dataInMem_hi_hi_lo_hi_lo_7 = {dataInMem_hi_hi_lo_hi_lo_hi_7, dataInMem_hi_hi_lo_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_lo_hi_hi_lo_7 = {dataInMem_hi_756, dataInMem_lo_628, dataInMem_hi_755, dataInMem_lo_627};
  wire [127:0]      dataInMem_hi_hi_lo_hi_hi_hi_7 = {dataInMem_hi_758, dataInMem_lo_630, dataInMem_hi_757, dataInMem_lo_629};
  wire [255:0]      dataInMem_hi_hi_lo_hi_hi_7 = {dataInMem_hi_hi_lo_hi_hi_hi_7, dataInMem_hi_hi_lo_hi_hi_lo_7};
  wire [511:0]      dataInMem_hi_hi_lo_hi_7 = {dataInMem_hi_hi_lo_hi_hi_7, dataInMem_hi_hi_lo_hi_lo_7};
  wire [1023:0]     dataInMem_hi_hi_lo_7 = {dataInMem_hi_hi_lo_hi_7, dataInMem_hi_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_hi_lo_lo_lo_7 = {dataInMem_hi_760, dataInMem_lo_632, dataInMem_hi_759, dataInMem_lo_631};
  wire [127:0]      dataInMem_hi_hi_hi_lo_lo_hi_7 = {dataInMem_hi_762, dataInMem_lo_634, dataInMem_hi_761, dataInMem_lo_633};
  wire [255:0]      dataInMem_hi_hi_hi_lo_lo_7 = {dataInMem_hi_hi_hi_lo_lo_hi_7, dataInMem_hi_hi_hi_lo_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_hi_lo_hi_lo_7 = {dataInMem_hi_764, dataInMem_lo_636, dataInMem_hi_763, dataInMem_lo_635};
  wire [127:0]      dataInMem_hi_hi_hi_lo_hi_hi_7 = {dataInMem_hi_766, dataInMem_lo_638, dataInMem_hi_765, dataInMem_lo_637};
  wire [255:0]      dataInMem_hi_hi_hi_lo_hi_7 = {dataInMem_hi_hi_hi_lo_hi_hi_7, dataInMem_hi_hi_hi_lo_hi_lo_7};
  wire [511:0]      dataInMem_hi_hi_hi_lo_7 = {dataInMem_hi_hi_hi_lo_hi_7, dataInMem_hi_hi_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_hi_hi_lo_lo_7 = {dataInMem_hi_768, dataInMem_lo_640, dataInMem_hi_767, dataInMem_lo_639};
  wire [127:0]      dataInMem_hi_hi_hi_hi_lo_hi_7 = {dataInMem_hi_770, dataInMem_lo_642, dataInMem_hi_769, dataInMem_lo_641};
  wire [255:0]      dataInMem_hi_hi_hi_hi_lo_7 = {dataInMem_hi_hi_hi_hi_lo_hi_7, dataInMem_hi_hi_hi_hi_lo_lo_7};
  wire [127:0]      dataInMem_hi_hi_hi_hi_hi_lo_7 = {dataInMem_hi_772, dataInMem_lo_644, dataInMem_hi_771, dataInMem_lo_643};
  wire [127:0]      dataInMem_hi_hi_hi_hi_hi_hi_7 = {dataInMem_hi_774, dataInMem_lo_646, dataInMem_hi_773, dataInMem_lo_645};
  wire [255:0]      dataInMem_hi_hi_hi_hi_hi_7 = {dataInMem_hi_hi_hi_hi_hi_hi_7, dataInMem_hi_hi_hi_hi_hi_lo_7};
  wire [511:0]      dataInMem_hi_hi_hi_hi_7 = {dataInMem_hi_hi_hi_hi_hi_7, dataInMem_hi_hi_hi_hi_lo_7};
  wire [1023:0]     dataInMem_hi_hi_hi_7 = {dataInMem_hi_hi_hi_hi_7, dataInMem_hi_hi_hi_lo_7};
  wire [2047:0]     dataInMem_hi_hi_519 = {dataInMem_hi_hi_hi_7, dataInMem_hi_hi_lo_7};
  wire [4095:0]     dataInMem_hi_775 = {dataInMem_hi_hi_519, dataInMem_hi_lo_263};
  wire [8191:0]     dataInMem_7 = {dataInMem_hi_775, dataInMem_lo_647};
  wire [1023:0]     regroupCacheLine_7_0 = dataInMem_7[1023:0];
  wire [1023:0]     regroupCacheLine_7_1 = dataInMem_7[2047:1024];
  wire [1023:0]     regroupCacheLine_7_2 = dataInMem_7[3071:2048];
  wire [1023:0]     regroupCacheLine_7_3 = dataInMem_7[4095:3072];
  wire [1023:0]     regroupCacheLine_7_4 = dataInMem_7[5119:4096];
  wire [1023:0]     regroupCacheLine_7_5 = dataInMem_7[6143:5120];
  wire [1023:0]     regroupCacheLine_7_6 = dataInMem_7[7167:6144];
  wire [1023:0]     regroupCacheLine_7_7 = dataInMem_7[8191:7168];
  wire [1023:0]     res_56 = regroupCacheLine_7_0;
  wire [1023:0]     res_57 = regroupCacheLine_7_1;
  wire [1023:0]     res_58 = regroupCacheLine_7_2;
  wire [1023:0]     res_59 = regroupCacheLine_7_3;
  wire [1023:0]     res_60 = regroupCacheLine_7_4;
  wire [1023:0]     res_61 = regroupCacheLine_7_5;
  wire [1023:0]     res_62 = regroupCacheLine_7_6;
  wire [1023:0]     res_63 = regroupCacheLine_7_7;
  wire [2047:0]     lo_lo_7 = {res_57, res_56};
  wire [2047:0]     lo_hi_7 = {res_59, res_58};
  wire [4095:0]     lo_7 = {lo_hi_7, lo_lo_7};
  wire [2047:0]     hi_lo_7 = {res_61, res_60};
  wire [2047:0]     hi_hi_7 = {res_63, res_62};
  wire [4095:0]     hi_7 = {hi_hi_7, hi_lo_7};
  wire [8191:0]     regroupLoadData_0_7 = {hi_7, lo_7};
  wire [15:0]       dataRegroupBySew_0_1_0 = bufferStageEnqueueData_0[15:0];
  wire [15:0]       dataRegroupBySew_0_1_1 = bufferStageEnqueueData_0[31:16];
  wire [15:0]       dataRegroupBySew_0_1_2 = bufferStageEnqueueData_0[47:32];
  wire [15:0]       dataRegroupBySew_0_1_3 = bufferStageEnqueueData_0[63:48];
  wire [15:0]       dataRegroupBySew_0_1_4 = bufferStageEnqueueData_0[79:64];
  wire [15:0]       dataRegroupBySew_0_1_5 = bufferStageEnqueueData_0[95:80];
  wire [15:0]       dataRegroupBySew_0_1_6 = bufferStageEnqueueData_0[111:96];
  wire [15:0]       dataRegroupBySew_0_1_7 = bufferStageEnqueueData_0[127:112];
  wire [15:0]       dataRegroupBySew_0_1_8 = bufferStageEnqueueData_0[143:128];
  wire [15:0]       dataRegroupBySew_0_1_9 = bufferStageEnqueueData_0[159:144];
  wire [15:0]       dataRegroupBySew_0_1_10 = bufferStageEnqueueData_0[175:160];
  wire [15:0]       dataRegroupBySew_0_1_11 = bufferStageEnqueueData_0[191:176];
  wire [15:0]       dataRegroupBySew_0_1_12 = bufferStageEnqueueData_0[207:192];
  wire [15:0]       dataRegroupBySew_0_1_13 = bufferStageEnqueueData_0[223:208];
  wire [15:0]       dataRegroupBySew_0_1_14 = bufferStageEnqueueData_0[239:224];
  wire [15:0]       dataRegroupBySew_0_1_15 = bufferStageEnqueueData_0[255:240];
  wire [15:0]       dataRegroupBySew_0_1_16 = bufferStageEnqueueData_0[271:256];
  wire [15:0]       dataRegroupBySew_0_1_17 = bufferStageEnqueueData_0[287:272];
  wire [15:0]       dataRegroupBySew_0_1_18 = bufferStageEnqueueData_0[303:288];
  wire [15:0]       dataRegroupBySew_0_1_19 = bufferStageEnqueueData_0[319:304];
  wire [15:0]       dataRegroupBySew_0_1_20 = bufferStageEnqueueData_0[335:320];
  wire [15:0]       dataRegroupBySew_0_1_21 = bufferStageEnqueueData_0[351:336];
  wire [15:0]       dataRegroupBySew_0_1_22 = bufferStageEnqueueData_0[367:352];
  wire [15:0]       dataRegroupBySew_0_1_23 = bufferStageEnqueueData_0[383:368];
  wire [15:0]       dataRegroupBySew_0_1_24 = bufferStageEnqueueData_0[399:384];
  wire [15:0]       dataRegroupBySew_0_1_25 = bufferStageEnqueueData_0[415:400];
  wire [15:0]       dataRegroupBySew_0_1_26 = bufferStageEnqueueData_0[431:416];
  wire [15:0]       dataRegroupBySew_0_1_27 = bufferStageEnqueueData_0[447:432];
  wire [15:0]       dataRegroupBySew_0_1_28 = bufferStageEnqueueData_0[463:448];
  wire [15:0]       dataRegroupBySew_0_1_29 = bufferStageEnqueueData_0[479:464];
  wire [15:0]       dataRegroupBySew_0_1_30 = bufferStageEnqueueData_0[495:480];
  wire [15:0]       dataRegroupBySew_0_1_31 = bufferStageEnqueueData_0[511:496];
  wire [15:0]       dataRegroupBySew_0_1_32 = bufferStageEnqueueData_0[527:512];
  wire [15:0]       dataRegroupBySew_0_1_33 = bufferStageEnqueueData_0[543:528];
  wire [15:0]       dataRegroupBySew_0_1_34 = bufferStageEnqueueData_0[559:544];
  wire [15:0]       dataRegroupBySew_0_1_35 = bufferStageEnqueueData_0[575:560];
  wire [15:0]       dataRegroupBySew_0_1_36 = bufferStageEnqueueData_0[591:576];
  wire [15:0]       dataRegroupBySew_0_1_37 = bufferStageEnqueueData_0[607:592];
  wire [15:0]       dataRegroupBySew_0_1_38 = bufferStageEnqueueData_0[623:608];
  wire [15:0]       dataRegroupBySew_0_1_39 = bufferStageEnqueueData_0[639:624];
  wire [15:0]       dataRegroupBySew_0_1_40 = bufferStageEnqueueData_0[655:640];
  wire [15:0]       dataRegroupBySew_0_1_41 = bufferStageEnqueueData_0[671:656];
  wire [15:0]       dataRegroupBySew_0_1_42 = bufferStageEnqueueData_0[687:672];
  wire [15:0]       dataRegroupBySew_0_1_43 = bufferStageEnqueueData_0[703:688];
  wire [15:0]       dataRegroupBySew_0_1_44 = bufferStageEnqueueData_0[719:704];
  wire [15:0]       dataRegroupBySew_0_1_45 = bufferStageEnqueueData_0[735:720];
  wire [15:0]       dataRegroupBySew_0_1_46 = bufferStageEnqueueData_0[751:736];
  wire [15:0]       dataRegroupBySew_0_1_47 = bufferStageEnqueueData_0[767:752];
  wire [15:0]       dataRegroupBySew_0_1_48 = bufferStageEnqueueData_0[783:768];
  wire [15:0]       dataRegroupBySew_0_1_49 = bufferStageEnqueueData_0[799:784];
  wire [15:0]       dataRegroupBySew_0_1_50 = bufferStageEnqueueData_0[815:800];
  wire [15:0]       dataRegroupBySew_0_1_51 = bufferStageEnqueueData_0[831:816];
  wire [15:0]       dataRegroupBySew_0_1_52 = bufferStageEnqueueData_0[847:832];
  wire [15:0]       dataRegroupBySew_0_1_53 = bufferStageEnqueueData_0[863:848];
  wire [15:0]       dataRegroupBySew_0_1_54 = bufferStageEnqueueData_0[879:864];
  wire [15:0]       dataRegroupBySew_0_1_55 = bufferStageEnqueueData_0[895:880];
  wire [15:0]       dataRegroupBySew_0_1_56 = bufferStageEnqueueData_0[911:896];
  wire [15:0]       dataRegroupBySew_0_1_57 = bufferStageEnqueueData_0[927:912];
  wire [15:0]       dataRegroupBySew_0_1_58 = bufferStageEnqueueData_0[943:928];
  wire [15:0]       dataRegroupBySew_0_1_59 = bufferStageEnqueueData_0[959:944];
  wire [15:0]       dataRegroupBySew_0_1_60 = bufferStageEnqueueData_0[975:960];
  wire [15:0]       dataRegroupBySew_0_1_61 = bufferStageEnqueueData_0[991:976];
  wire [15:0]       dataRegroupBySew_0_1_62 = bufferStageEnqueueData_0[1007:992];
  wire [15:0]       dataRegroupBySew_0_1_63 = bufferStageEnqueueData_0[1023:1008];
  wire [15:0]       dataRegroupBySew_1_1_0 = bufferStageEnqueueData_1[15:0];
  wire [15:0]       dataRegroupBySew_1_1_1 = bufferStageEnqueueData_1[31:16];
  wire [15:0]       dataRegroupBySew_1_1_2 = bufferStageEnqueueData_1[47:32];
  wire [15:0]       dataRegroupBySew_1_1_3 = bufferStageEnqueueData_1[63:48];
  wire [15:0]       dataRegroupBySew_1_1_4 = bufferStageEnqueueData_1[79:64];
  wire [15:0]       dataRegroupBySew_1_1_5 = bufferStageEnqueueData_1[95:80];
  wire [15:0]       dataRegroupBySew_1_1_6 = bufferStageEnqueueData_1[111:96];
  wire [15:0]       dataRegroupBySew_1_1_7 = bufferStageEnqueueData_1[127:112];
  wire [15:0]       dataRegroupBySew_1_1_8 = bufferStageEnqueueData_1[143:128];
  wire [15:0]       dataRegroupBySew_1_1_9 = bufferStageEnqueueData_1[159:144];
  wire [15:0]       dataRegroupBySew_1_1_10 = bufferStageEnqueueData_1[175:160];
  wire [15:0]       dataRegroupBySew_1_1_11 = bufferStageEnqueueData_1[191:176];
  wire [15:0]       dataRegroupBySew_1_1_12 = bufferStageEnqueueData_1[207:192];
  wire [15:0]       dataRegroupBySew_1_1_13 = bufferStageEnqueueData_1[223:208];
  wire [15:0]       dataRegroupBySew_1_1_14 = bufferStageEnqueueData_1[239:224];
  wire [15:0]       dataRegroupBySew_1_1_15 = bufferStageEnqueueData_1[255:240];
  wire [15:0]       dataRegroupBySew_1_1_16 = bufferStageEnqueueData_1[271:256];
  wire [15:0]       dataRegroupBySew_1_1_17 = bufferStageEnqueueData_1[287:272];
  wire [15:0]       dataRegroupBySew_1_1_18 = bufferStageEnqueueData_1[303:288];
  wire [15:0]       dataRegroupBySew_1_1_19 = bufferStageEnqueueData_1[319:304];
  wire [15:0]       dataRegroupBySew_1_1_20 = bufferStageEnqueueData_1[335:320];
  wire [15:0]       dataRegroupBySew_1_1_21 = bufferStageEnqueueData_1[351:336];
  wire [15:0]       dataRegroupBySew_1_1_22 = bufferStageEnqueueData_1[367:352];
  wire [15:0]       dataRegroupBySew_1_1_23 = bufferStageEnqueueData_1[383:368];
  wire [15:0]       dataRegroupBySew_1_1_24 = bufferStageEnqueueData_1[399:384];
  wire [15:0]       dataRegroupBySew_1_1_25 = bufferStageEnqueueData_1[415:400];
  wire [15:0]       dataRegroupBySew_1_1_26 = bufferStageEnqueueData_1[431:416];
  wire [15:0]       dataRegroupBySew_1_1_27 = bufferStageEnqueueData_1[447:432];
  wire [15:0]       dataRegroupBySew_1_1_28 = bufferStageEnqueueData_1[463:448];
  wire [15:0]       dataRegroupBySew_1_1_29 = bufferStageEnqueueData_1[479:464];
  wire [15:0]       dataRegroupBySew_1_1_30 = bufferStageEnqueueData_1[495:480];
  wire [15:0]       dataRegroupBySew_1_1_31 = bufferStageEnqueueData_1[511:496];
  wire [15:0]       dataRegroupBySew_1_1_32 = bufferStageEnqueueData_1[527:512];
  wire [15:0]       dataRegroupBySew_1_1_33 = bufferStageEnqueueData_1[543:528];
  wire [15:0]       dataRegroupBySew_1_1_34 = bufferStageEnqueueData_1[559:544];
  wire [15:0]       dataRegroupBySew_1_1_35 = bufferStageEnqueueData_1[575:560];
  wire [15:0]       dataRegroupBySew_1_1_36 = bufferStageEnqueueData_1[591:576];
  wire [15:0]       dataRegroupBySew_1_1_37 = bufferStageEnqueueData_1[607:592];
  wire [15:0]       dataRegroupBySew_1_1_38 = bufferStageEnqueueData_1[623:608];
  wire [15:0]       dataRegroupBySew_1_1_39 = bufferStageEnqueueData_1[639:624];
  wire [15:0]       dataRegroupBySew_1_1_40 = bufferStageEnqueueData_1[655:640];
  wire [15:0]       dataRegroupBySew_1_1_41 = bufferStageEnqueueData_1[671:656];
  wire [15:0]       dataRegroupBySew_1_1_42 = bufferStageEnqueueData_1[687:672];
  wire [15:0]       dataRegroupBySew_1_1_43 = bufferStageEnqueueData_1[703:688];
  wire [15:0]       dataRegroupBySew_1_1_44 = bufferStageEnqueueData_1[719:704];
  wire [15:0]       dataRegroupBySew_1_1_45 = bufferStageEnqueueData_1[735:720];
  wire [15:0]       dataRegroupBySew_1_1_46 = bufferStageEnqueueData_1[751:736];
  wire [15:0]       dataRegroupBySew_1_1_47 = bufferStageEnqueueData_1[767:752];
  wire [15:0]       dataRegroupBySew_1_1_48 = bufferStageEnqueueData_1[783:768];
  wire [15:0]       dataRegroupBySew_1_1_49 = bufferStageEnqueueData_1[799:784];
  wire [15:0]       dataRegroupBySew_1_1_50 = bufferStageEnqueueData_1[815:800];
  wire [15:0]       dataRegroupBySew_1_1_51 = bufferStageEnqueueData_1[831:816];
  wire [15:0]       dataRegroupBySew_1_1_52 = bufferStageEnqueueData_1[847:832];
  wire [15:0]       dataRegroupBySew_1_1_53 = bufferStageEnqueueData_1[863:848];
  wire [15:0]       dataRegroupBySew_1_1_54 = bufferStageEnqueueData_1[879:864];
  wire [15:0]       dataRegroupBySew_1_1_55 = bufferStageEnqueueData_1[895:880];
  wire [15:0]       dataRegroupBySew_1_1_56 = bufferStageEnqueueData_1[911:896];
  wire [15:0]       dataRegroupBySew_1_1_57 = bufferStageEnqueueData_1[927:912];
  wire [15:0]       dataRegroupBySew_1_1_58 = bufferStageEnqueueData_1[943:928];
  wire [15:0]       dataRegroupBySew_1_1_59 = bufferStageEnqueueData_1[959:944];
  wire [15:0]       dataRegroupBySew_1_1_60 = bufferStageEnqueueData_1[975:960];
  wire [15:0]       dataRegroupBySew_1_1_61 = bufferStageEnqueueData_1[991:976];
  wire [15:0]       dataRegroupBySew_1_1_62 = bufferStageEnqueueData_1[1007:992];
  wire [15:0]       dataRegroupBySew_1_1_63 = bufferStageEnqueueData_1[1023:1008];
  wire [15:0]       dataRegroupBySew_2_1_0 = bufferStageEnqueueData_2[15:0];
  wire [15:0]       dataRegroupBySew_2_1_1 = bufferStageEnqueueData_2[31:16];
  wire [15:0]       dataRegroupBySew_2_1_2 = bufferStageEnqueueData_2[47:32];
  wire [15:0]       dataRegroupBySew_2_1_3 = bufferStageEnqueueData_2[63:48];
  wire [15:0]       dataRegroupBySew_2_1_4 = bufferStageEnqueueData_2[79:64];
  wire [15:0]       dataRegroupBySew_2_1_5 = bufferStageEnqueueData_2[95:80];
  wire [15:0]       dataRegroupBySew_2_1_6 = bufferStageEnqueueData_2[111:96];
  wire [15:0]       dataRegroupBySew_2_1_7 = bufferStageEnqueueData_2[127:112];
  wire [15:0]       dataRegroupBySew_2_1_8 = bufferStageEnqueueData_2[143:128];
  wire [15:0]       dataRegroupBySew_2_1_9 = bufferStageEnqueueData_2[159:144];
  wire [15:0]       dataRegroupBySew_2_1_10 = bufferStageEnqueueData_2[175:160];
  wire [15:0]       dataRegroupBySew_2_1_11 = bufferStageEnqueueData_2[191:176];
  wire [15:0]       dataRegroupBySew_2_1_12 = bufferStageEnqueueData_2[207:192];
  wire [15:0]       dataRegroupBySew_2_1_13 = bufferStageEnqueueData_2[223:208];
  wire [15:0]       dataRegroupBySew_2_1_14 = bufferStageEnqueueData_2[239:224];
  wire [15:0]       dataRegroupBySew_2_1_15 = bufferStageEnqueueData_2[255:240];
  wire [15:0]       dataRegroupBySew_2_1_16 = bufferStageEnqueueData_2[271:256];
  wire [15:0]       dataRegroupBySew_2_1_17 = bufferStageEnqueueData_2[287:272];
  wire [15:0]       dataRegroupBySew_2_1_18 = bufferStageEnqueueData_2[303:288];
  wire [15:0]       dataRegroupBySew_2_1_19 = bufferStageEnqueueData_2[319:304];
  wire [15:0]       dataRegroupBySew_2_1_20 = bufferStageEnqueueData_2[335:320];
  wire [15:0]       dataRegroupBySew_2_1_21 = bufferStageEnqueueData_2[351:336];
  wire [15:0]       dataRegroupBySew_2_1_22 = bufferStageEnqueueData_2[367:352];
  wire [15:0]       dataRegroupBySew_2_1_23 = bufferStageEnqueueData_2[383:368];
  wire [15:0]       dataRegroupBySew_2_1_24 = bufferStageEnqueueData_2[399:384];
  wire [15:0]       dataRegroupBySew_2_1_25 = bufferStageEnqueueData_2[415:400];
  wire [15:0]       dataRegroupBySew_2_1_26 = bufferStageEnqueueData_2[431:416];
  wire [15:0]       dataRegroupBySew_2_1_27 = bufferStageEnqueueData_2[447:432];
  wire [15:0]       dataRegroupBySew_2_1_28 = bufferStageEnqueueData_2[463:448];
  wire [15:0]       dataRegroupBySew_2_1_29 = bufferStageEnqueueData_2[479:464];
  wire [15:0]       dataRegroupBySew_2_1_30 = bufferStageEnqueueData_2[495:480];
  wire [15:0]       dataRegroupBySew_2_1_31 = bufferStageEnqueueData_2[511:496];
  wire [15:0]       dataRegroupBySew_2_1_32 = bufferStageEnqueueData_2[527:512];
  wire [15:0]       dataRegroupBySew_2_1_33 = bufferStageEnqueueData_2[543:528];
  wire [15:0]       dataRegroupBySew_2_1_34 = bufferStageEnqueueData_2[559:544];
  wire [15:0]       dataRegroupBySew_2_1_35 = bufferStageEnqueueData_2[575:560];
  wire [15:0]       dataRegroupBySew_2_1_36 = bufferStageEnqueueData_2[591:576];
  wire [15:0]       dataRegroupBySew_2_1_37 = bufferStageEnqueueData_2[607:592];
  wire [15:0]       dataRegroupBySew_2_1_38 = bufferStageEnqueueData_2[623:608];
  wire [15:0]       dataRegroupBySew_2_1_39 = bufferStageEnqueueData_2[639:624];
  wire [15:0]       dataRegroupBySew_2_1_40 = bufferStageEnqueueData_2[655:640];
  wire [15:0]       dataRegroupBySew_2_1_41 = bufferStageEnqueueData_2[671:656];
  wire [15:0]       dataRegroupBySew_2_1_42 = bufferStageEnqueueData_2[687:672];
  wire [15:0]       dataRegroupBySew_2_1_43 = bufferStageEnqueueData_2[703:688];
  wire [15:0]       dataRegroupBySew_2_1_44 = bufferStageEnqueueData_2[719:704];
  wire [15:0]       dataRegroupBySew_2_1_45 = bufferStageEnqueueData_2[735:720];
  wire [15:0]       dataRegroupBySew_2_1_46 = bufferStageEnqueueData_2[751:736];
  wire [15:0]       dataRegroupBySew_2_1_47 = bufferStageEnqueueData_2[767:752];
  wire [15:0]       dataRegroupBySew_2_1_48 = bufferStageEnqueueData_2[783:768];
  wire [15:0]       dataRegroupBySew_2_1_49 = bufferStageEnqueueData_2[799:784];
  wire [15:0]       dataRegroupBySew_2_1_50 = bufferStageEnqueueData_2[815:800];
  wire [15:0]       dataRegroupBySew_2_1_51 = bufferStageEnqueueData_2[831:816];
  wire [15:0]       dataRegroupBySew_2_1_52 = bufferStageEnqueueData_2[847:832];
  wire [15:0]       dataRegroupBySew_2_1_53 = bufferStageEnqueueData_2[863:848];
  wire [15:0]       dataRegroupBySew_2_1_54 = bufferStageEnqueueData_2[879:864];
  wire [15:0]       dataRegroupBySew_2_1_55 = bufferStageEnqueueData_2[895:880];
  wire [15:0]       dataRegroupBySew_2_1_56 = bufferStageEnqueueData_2[911:896];
  wire [15:0]       dataRegroupBySew_2_1_57 = bufferStageEnqueueData_2[927:912];
  wire [15:0]       dataRegroupBySew_2_1_58 = bufferStageEnqueueData_2[943:928];
  wire [15:0]       dataRegroupBySew_2_1_59 = bufferStageEnqueueData_2[959:944];
  wire [15:0]       dataRegroupBySew_2_1_60 = bufferStageEnqueueData_2[975:960];
  wire [15:0]       dataRegroupBySew_2_1_61 = bufferStageEnqueueData_2[991:976];
  wire [15:0]       dataRegroupBySew_2_1_62 = bufferStageEnqueueData_2[1007:992];
  wire [15:0]       dataRegroupBySew_2_1_63 = bufferStageEnqueueData_2[1023:1008];
  wire [15:0]       dataRegroupBySew_3_1_0 = bufferStageEnqueueData_3[15:0];
  wire [15:0]       dataRegroupBySew_3_1_1 = bufferStageEnqueueData_3[31:16];
  wire [15:0]       dataRegroupBySew_3_1_2 = bufferStageEnqueueData_3[47:32];
  wire [15:0]       dataRegroupBySew_3_1_3 = bufferStageEnqueueData_3[63:48];
  wire [15:0]       dataRegroupBySew_3_1_4 = bufferStageEnqueueData_3[79:64];
  wire [15:0]       dataRegroupBySew_3_1_5 = bufferStageEnqueueData_3[95:80];
  wire [15:0]       dataRegroupBySew_3_1_6 = bufferStageEnqueueData_3[111:96];
  wire [15:0]       dataRegroupBySew_3_1_7 = bufferStageEnqueueData_3[127:112];
  wire [15:0]       dataRegroupBySew_3_1_8 = bufferStageEnqueueData_3[143:128];
  wire [15:0]       dataRegroupBySew_3_1_9 = bufferStageEnqueueData_3[159:144];
  wire [15:0]       dataRegroupBySew_3_1_10 = bufferStageEnqueueData_3[175:160];
  wire [15:0]       dataRegroupBySew_3_1_11 = bufferStageEnqueueData_3[191:176];
  wire [15:0]       dataRegroupBySew_3_1_12 = bufferStageEnqueueData_3[207:192];
  wire [15:0]       dataRegroupBySew_3_1_13 = bufferStageEnqueueData_3[223:208];
  wire [15:0]       dataRegroupBySew_3_1_14 = bufferStageEnqueueData_3[239:224];
  wire [15:0]       dataRegroupBySew_3_1_15 = bufferStageEnqueueData_3[255:240];
  wire [15:0]       dataRegroupBySew_3_1_16 = bufferStageEnqueueData_3[271:256];
  wire [15:0]       dataRegroupBySew_3_1_17 = bufferStageEnqueueData_3[287:272];
  wire [15:0]       dataRegroupBySew_3_1_18 = bufferStageEnqueueData_3[303:288];
  wire [15:0]       dataRegroupBySew_3_1_19 = bufferStageEnqueueData_3[319:304];
  wire [15:0]       dataRegroupBySew_3_1_20 = bufferStageEnqueueData_3[335:320];
  wire [15:0]       dataRegroupBySew_3_1_21 = bufferStageEnqueueData_3[351:336];
  wire [15:0]       dataRegroupBySew_3_1_22 = bufferStageEnqueueData_3[367:352];
  wire [15:0]       dataRegroupBySew_3_1_23 = bufferStageEnqueueData_3[383:368];
  wire [15:0]       dataRegroupBySew_3_1_24 = bufferStageEnqueueData_3[399:384];
  wire [15:0]       dataRegroupBySew_3_1_25 = bufferStageEnqueueData_3[415:400];
  wire [15:0]       dataRegroupBySew_3_1_26 = bufferStageEnqueueData_3[431:416];
  wire [15:0]       dataRegroupBySew_3_1_27 = bufferStageEnqueueData_3[447:432];
  wire [15:0]       dataRegroupBySew_3_1_28 = bufferStageEnqueueData_3[463:448];
  wire [15:0]       dataRegroupBySew_3_1_29 = bufferStageEnqueueData_3[479:464];
  wire [15:0]       dataRegroupBySew_3_1_30 = bufferStageEnqueueData_3[495:480];
  wire [15:0]       dataRegroupBySew_3_1_31 = bufferStageEnqueueData_3[511:496];
  wire [15:0]       dataRegroupBySew_3_1_32 = bufferStageEnqueueData_3[527:512];
  wire [15:0]       dataRegroupBySew_3_1_33 = bufferStageEnqueueData_3[543:528];
  wire [15:0]       dataRegroupBySew_3_1_34 = bufferStageEnqueueData_3[559:544];
  wire [15:0]       dataRegroupBySew_3_1_35 = bufferStageEnqueueData_3[575:560];
  wire [15:0]       dataRegroupBySew_3_1_36 = bufferStageEnqueueData_3[591:576];
  wire [15:0]       dataRegroupBySew_3_1_37 = bufferStageEnqueueData_3[607:592];
  wire [15:0]       dataRegroupBySew_3_1_38 = bufferStageEnqueueData_3[623:608];
  wire [15:0]       dataRegroupBySew_3_1_39 = bufferStageEnqueueData_3[639:624];
  wire [15:0]       dataRegroupBySew_3_1_40 = bufferStageEnqueueData_3[655:640];
  wire [15:0]       dataRegroupBySew_3_1_41 = bufferStageEnqueueData_3[671:656];
  wire [15:0]       dataRegroupBySew_3_1_42 = bufferStageEnqueueData_3[687:672];
  wire [15:0]       dataRegroupBySew_3_1_43 = bufferStageEnqueueData_3[703:688];
  wire [15:0]       dataRegroupBySew_3_1_44 = bufferStageEnqueueData_3[719:704];
  wire [15:0]       dataRegroupBySew_3_1_45 = bufferStageEnqueueData_3[735:720];
  wire [15:0]       dataRegroupBySew_3_1_46 = bufferStageEnqueueData_3[751:736];
  wire [15:0]       dataRegroupBySew_3_1_47 = bufferStageEnqueueData_3[767:752];
  wire [15:0]       dataRegroupBySew_3_1_48 = bufferStageEnqueueData_3[783:768];
  wire [15:0]       dataRegroupBySew_3_1_49 = bufferStageEnqueueData_3[799:784];
  wire [15:0]       dataRegroupBySew_3_1_50 = bufferStageEnqueueData_3[815:800];
  wire [15:0]       dataRegroupBySew_3_1_51 = bufferStageEnqueueData_3[831:816];
  wire [15:0]       dataRegroupBySew_3_1_52 = bufferStageEnqueueData_3[847:832];
  wire [15:0]       dataRegroupBySew_3_1_53 = bufferStageEnqueueData_3[863:848];
  wire [15:0]       dataRegroupBySew_3_1_54 = bufferStageEnqueueData_3[879:864];
  wire [15:0]       dataRegroupBySew_3_1_55 = bufferStageEnqueueData_3[895:880];
  wire [15:0]       dataRegroupBySew_3_1_56 = bufferStageEnqueueData_3[911:896];
  wire [15:0]       dataRegroupBySew_3_1_57 = bufferStageEnqueueData_3[927:912];
  wire [15:0]       dataRegroupBySew_3_1_58 = bufferStageEnqueueData_3[943:928];
  wire [15:0]       dataRegroupBySew_3_1_59 = bufferStageEnqueueData_3[959:944];
  wire [15:0]       dataRegroupBySew_3_1_60 = bufferStageEnqueueData_3[975:960];
  wire [15:0]       dataRegroupBySew_3_1_61 = bufferStageEnqueueData_3[991:976];
  wire [15:0]       dataRegroupBySew_3_1_62 = bufferStageEnqueueData_3[1007:992];
  wire [15:0]       dataRegroupBySew_3_1_63 = bufferStageEnqueueData_3[1023:1008];
  wire [15:0]       dataRegroupBySew_4_1_0 = bufferStageEnqueueData_4[15:0];
  wire [15:0]       dataRegroupBySew_4_1_1 = bufferStageEnqueueData_4[31:16];
  wire [15:0]       dataRegroupBySew_4_1_2 = bufferStageEnqueueData_4[47:32];
  wire [15:0]       dataRegroupBySew_4_1_3 = bufferStageEnqueueData_4[63:48];
  wire [15:0]       dataRegroupBySew_4_1_4 = bufferStageEnqueueData_4[79:64];
  wire [15:0]       dataRegroupBySew_4_1_5 = bufferStageEnqueueData_4[95:80];
  wire [15:0]       dataRegroupBySew_4_1_6 = bufferStageEnqueueData_4[111:96];
  wire [15:0]       dataRegroupBySew_4_1_7 = bufferStageEnqueueData_4[127:112];
  wire [15:0]       dataRegroupBySew_4_1_8 = bufferStageEnqueueData_4[143:128];
  wire [15:0]       dataRegroupBySew_4_1_9 = bufferStageEnqueueData_4[159:144];
  wire [15:0]       dataRegroupBySew_4_1_10 = bufferStageEnqueueData_4[175:160];
  wire [15:0]       dataRegroupBySew_4_1_11 = bufferStageEnqueueData_4[191:176];
  wire [15:0]       dataRegroupBySew_4_1_12 = bufferStageEnqueueData_4[207:192];
  wire [15:0]       dataRegroupBySew_4_1_13 = bufferStageEnqueueData_4[223:208];
  wire [15:0]       dataRegroupBySew_4_1_14 = bufferStageEnqueueData_4[239:224];
  wire [15:0]       dataRegroupBySew_4_1_15 = bufferStageEnqueueData_4[255:240];
  wire [15:0]       dataRegroupBySew_4_1_16 = bufferStageEnqueueData_4[271:256];
  wire [15:0]       dataRegroupBySew_4_1_17 = bufferStageEnqueueData_4[287:272];
  wire [15:0]       dataRegroupBySew_4_1_18 = bufferStageEnqueueData_4[303:288];
  wire [15:0]       dataRegroupBySew_4_1_19 = bufferStageEnqueueData_4[319:304];
  wire [15:0]       dataRegroupBySew_4_1_20 = bufferStageEnqueueData_4[335:320];
  wire [15:0]       dataRegroupBySew_4_1_21 = bufferStageEnqueueData_4[351:336];
  wire [15:0]       dataRegroupBySew_4_1_22 = bufferStageEnqueueData_4[367:352];
  wire [15:0]       dataRegroupBySew_4_1_23 = bufferStageEnqueueData_4[383:368];
  wire [15:0]       dataRegroupBySew_4_1_24 = bufferStageEnqueueData_4[399:384];
  wire [15:0]       dataRegroupBySew_4_1_25 = bufferStageEnqueueData_4[415:400];
  wire [15:0]       dataRegroupBySew_4_1_26 = bufferStageEnqueueData_4[431:416];
  wire [15:0]       dataRegroupBySew_4_1_27 = bufferStageEnqueueData_4[447:432];
  wire [15:0]       dataRegroupBySew_4_1_28 = bufferStageEnqueueData_4[463:448];
  wire [15:0]       dataRegroupBySew_4_1_29 = bufferStageEnqueueData_4[479:464];
  wire [15:0]       dataRegroupBySew_4_1_30 = bufferStageEnqueueData_4[495:480];
  wire [15:0]       dataRegroupBySew_4_1_31 = bufferStageEnqueueData_4[511:496];
  wire [15:0]       dataRegroupBySew_4_1_32 = bufferStageEnqueueData_4[527:512];
  wire [15:0]       dataRegroupBySew_4_1_33 = bufferStageEnqueueData_4[543:528];
  wire [15:0]       dataRegroupBySew_4_1_34 = bufferStageEnqueueData_4[559:544];
  wire [15:0]       dataRegroupBySew_4_1_35 = bufferStageEnqueueData_4[575:560];
  wire [15:0]       dataRegroupBySew_4_1_36 = bufferStageEnqueueData_4[591:576];
  wire [15:0]       dataRegroupBySew_4_1_37 = bufferStageEnqueueData_4[607:592];
  wire [15:0]       dataRegroupBySew_4_1_38 = bufferStageEnqueueData_4[623:608];
  wire [15:0]       dataRegroupBySew_4_1_39 = bufferStageEnqueueData_4[639:624];
  wire [15:0]       dataRegroupBySew_4_1_40 = bufferStageEnqueueData_4[655:640];
  wire [15:0]       dataRegroupBySew_4_1_41 = bufferStageEnqueueData_4[671:656];
  wire [15:0]       dataRegroupBySew_4_1_42 = bufferStageEnqueueData_4[687:672];
  wire [15:0]       dataRegroupBySew_4_1_43 = bufferStageEnqueueData_4[703:688];
  wire [15:0]       dataRegroupBySew_4_1_44 = bufferStageEnqueueData_4[719:704];
  wire [15:0]       dataRegroupBySew_4_1_45 = bufferStageEnqueueData_4[735:720];
  wire [15:0]       dataRegroupBySew_4_1_46 = bufferStageEnqueueData_4[751:736];
  wire [15:0]       dataRegroupBySew_4_1_47 = bufferStageEnqueueData_4[767:752];
  wire [15:0]       dataRegroupBySew_4_1_48 = bufferStageEnqueueData_4[783:768];
  wire [15:0]       dataRegroupBySew_4_1_49 = bufferStageEnqueueData_4[799:784];
  wire [15:0]       dataRegroupBySew_4_1_50 = bufferStageEnqueueData_4[815:800];
  wire [15:0]       dataRegroupBySew_4_1_51 = bufferStageEnqueueData_4[831:816];
  wire [15:0]       dataRegroupBySew_4_1_52 = bufferStageEnqueueData_4[847:832];
  wire [15:0]       dataRegroupBySew_4_1_53 = bufferStageEnqueueData_4[863:848];
  wire [15:0]       dataRegroupBySew_4_1_54 = bufferStageEnqueueData_4[879:864];
  wire [15:0]       dataRegroupBySew_4_1_55 = bufferStageEnqueueData_4[895:880];
  wire [15:0]       dataRegroupBySew_4_1_56 = bufferStageEnqueueData_4[911:896];
  wire [15:0]       dataRegroupBySew_4_1_57 = bufferStageEnqueueData_4[927:912];
  wire [15:0]       dataRegroupBySew_4_1_58 = bufferStageEnqueueData_4[943:928];
  wire [15:0]       dataRegroupBySew_4_1_59 = bufferStageEnqueueData_4[959:944];
  wire [15:0]       dataRegroupBySew_4_1_60 = bufferStageEnqueueData_4[975:960];
  wire [15:0]       dataRegroupBySew_4_1_61 = bufferStageEnqueueData_4[991:976];
  wire [15:0]       dataRegroupBySew_4_1_62 = bufferStageEnqueueData_4[1007:992];
  wire [15:0]       dataRegroupBySew_4_1_63 = bufferStageEnqueueData_4[1023:1008];
  wire [15:0]       dataRegroupBySew_5_1_0 = bufferStageEnqueueData_5[15:0];
  wire [15:0]       dataRegroupBySew_5_1_1 = bufferStageEnqueueData_5[31:16];
  wire [15:0]       dataRegroupBySew_5_1_2 = bufferStageEnqueueData_5[47:32];
  wire [15:0]       dataRegroupBySew_5_1_3 = bufferStageEnqueueData_5[63:48];
  wire [15:0]       dataRegroupBySew_5_1_4 = bufferStageEnqueueData_5[79:64];
  wire [15:0]       dataRegroupBySew_5_1_5 = bufferStageEnqueueData_5[95:80];
  wire [15:0]       dataRegroupBySew_5_1_6 = bufferStageEnqueueData_5[111:96];
  wire [15:0]       dataRegroupBySew_5_1_7 = bufferStageEnqueueData_5[127:112];
  wire [15:0]       dataRegroupBySew_5_1_8 = bufferStageEnqueueData_5[143:128];
  wire [15:0]       dataRegroupBySew_5_1_9 = bufferStageEnqueueData_5[159:144];
  wire [15:0]       dataRegroupBySew_5_1_10 = bufferStageEnqueueData_5[175:160];
  wire [15:0]       dataRegroupBySew_5_1_11 = bufferStageEnqueueData_5[191:176];
  wire [15:0]       dataRegroupBySew_5_1_12 = bufferStageEnqueueData_5[207:192];
  wire [15:0]       dataRegroupBySew_5_1_13 = bufferStageEnqueueData_5[223:208];
  wire [15:0]       dataRegroupBySew_5_1_14 = bufferStageEnqueueData_5[239:224];
  wire [15:0]       dataRegroupBySew_5_1_15 = bufferStageEnqueueData_5[255:240];
  wire [15:0]       dataRegroupBySew_5_1_16 = bufferStageEnqueueData_5[271:256];
  wire [15:0]       dataRegroupBySew_5_1_17 = bufferStageEnqueueData_5[287:272];
  wire [15:0]       dataRegroupBySew_5_1_18 = bufferStageEnqueueData_5[303:288];
  wire [15:0]       dataRegroupBySew_5_1_19 = bufferStageEnqueueData_5[319:304];
  wire [15:0]       dataRegroupBySew_5_1_20 = bufferStageEnqueueData_5[335:320];
  wire [15:0]       dataRegroupBySew_5_1_21 = bufferStageEnqueueData_5[351:336];
  wire [15:0]       dataRegroupBySew_5_1_22 = bufferStageEnqueueData_5[367:352];
  wire [15:0]       dataRegroupBySew_5_1_23 = bufferStageEnqueueData_5[383:368];
  wire [15:0]       dataRegroupBySew_5_1_24 = bufferStageEnqueueData_5[399:384];
  wire [15:0]       dataRegroupBySew_5_1_25 = bufferStageEnqueueData_5[415:400];
  wire [15:0]       dataRegroupBySew_5_1_26 = bufferStageEnqueueData_5[431:416];
  wire [15:0]       dataRegroupBySew_5_1_27 = bufferStageEnqueueData_5[447:432];
  wire [15:0]       dataRegroupBySew_5_1_28 = bufferStageEnqueueData_5[463:448];
  wire [15:0]       dataRegroupBySew_5_1_29 = bufferStageEnqueueData_5[479:464];
  wire [15:0]       dataRegroupBySew_5_1_30 = bufferStageEnqueueData_5[495:480];
  wire [15:0]       dataRegroupBySew_5_1_31 = bufferStageEnqueueData_5[511:496];
  wire [15:0]       dataRegroupBySew_5_1_32 = bufferStageEnqueueData_5[527:512];
  wire [15:0]       dataRegroupBySew_5_1_33 = bufferStageEnqueueData_5[543:528];
  wire [15:0]       dataRegroupBySew_5_1_34 = bufferStageEnqueueData_5[559:544];
  wire [15:0]       dataRegroupBySew_5_1_35 = bufferStageEnqueueData_5[575:560];
  wire [15:0]       dataRegroupBySew_5_1_36 = bufferStageEnqueueData_5[591:576];
  wire [15:0]       dataRegroupBySew_5_1_37 = bufferStageEnqueueData_5[607:592];
  wire [15:0]       dataRegroupBySew_5_1_38 = bufferStageEnqueueData_5[623:608];
  wire [15:0]       dataRegroupBySew_5_1_39 = bufferStageEnqueueData_5[639:624];
  wire [15:0]       dataRegroupBySew_5_1_40 = bufferStageEnqueueData_5[655:640];
  wire [15:0]       dataRegroupBySew_5_1_41 = bufferStageEnqueueData_5[671:656];
  wire [15:0]       dataRegroupBySew_5_1_42 = bufferStageEnqueueData_5[687:672];
  wire [15:0]       dataRegroupBySew_5_1_43 = bufferStageEnqueueData_5[703:688];
  wire [15:0]       dataRegroupBySew_5_1_44 = bufferStageEnqueueData_5[719:704];
  wire [15:0]       dataRegroupBySew_5_1_45 = bufferStageEnqueueData_5[735:720];
  wire [15:0]       dataRegroupBySew_5_1_46 = bufferStageEnqueueData_5[751:736];
  wire [15:0]       dataRegroupBySew_5_1_47 = bufferStageEnqueueData_5[767:752];
  wire [15:0]       dataRegroupBySew_5_1_48 = bufferStageEnqueueData_5[783:768];
  wire [15:0]       dataRegroupBySew_5_1_49 = bufferStageEnqueueData_5[799:784];
  wire [15:0]       dataRegroupBySew_5_1_50 = bufferStageEnqueueData_5[815:800];
  wire [15:0]       dataRegroupBySew_5_1_51 = bufferStageEnqueueData_5[831:816];
  wire [15:0]       dataRegroupBySew_5_1_52 = bufferStageEnqueueData_5[847:832];
  wire [15:0]       dataRegroupBySew_5_1_53 = bufferStageEnqueueData_5[863:848];
  wire [15:0]       dataRegroupBySew_5_1_54 = bufferStageEnqueueData_5[879:864];
  wire [15:0]       dataRegroupBySew_5_1_55 = bufferStageEnqueueData_5[895:880];
  wire [15:0]       dataRegroupBySew_5_1_56 = bufferStageEnqueueData_5[911:896];
  wire [15:0]       dataRegroupBySew_5_1_57 = bufferStageEnqueueData_5[927:912];
  wire [15:0]       dataRegroupBySew_5_1_58 = bufferStageEnqueueData_5[943:928];
  wire [15:0]       dataRegroupBySew_5_1_59 = bufferStageEnqueueData_5[959:944];
  wire [15:0]       dataRegroupBySew_5_1_60 = bufferStageEnqueueData_5[975:960];
  wire [15:0]       dataRegroupBySew_5_1_61 = bufferStageEnqueueData_5[991:976];
  wire [15:0]       dataRegroupBySew_5_1_62 = bufferStageEnqueueData_5[1007:992];
  wire [15:0]       dataRegroupBySew_5_1_63 = bufferStageEnqueueData_5[1023:1008];
  wire [15:0]       dataRegroupBySew_6_1_0 = bufferStageEnqueueData_6[15:0];
  wire [15:0]       dataRegroupBySew_6_1_1 = bufferStageEnqueueData_6[31:16];
  wire [15:0]       dataRegroupBySew_6_1_2 = bufferStageEnqueueData_6[47:32];
  wire [15:0]       dataRegroupBySew_6_1_3 = bufferStageEnqueueData_6[63:48];
  wire [15:0]       dataRegroupBySew_6_1_4 = bufferStageEnqueueData_6[79:64];
  wire [15:0]       dataRegroupBySew_6_1_5 = bufferStageEnqueueData_6[95:80];
  wire [15:0]       dataRegroupBySew_6_1_6 = bufferStageEnqueueData_6[111:96];
  wire [15:0]       dataRegroupBySew_6_1_7 = bufferStageEnqueueData_6[127:112];
  wire [15:0]       dataRegroupBySew_6_1_8 = bufferStageEnqueueData_6[143:128];
  wire [15:0]       dataRegroupBySew_6_1_9 = bufferStageEnqueueData_6[159:144];
  wire [15:0]       dataRegroupBySew_6_1_10 = bufferStageEnqueueData_6[175:160];
  wire [15:0]       dataRegroupBySew_6_1_11 = bufferStageEnqueueData_6[191:176];
  wire [15:0]       dataRegroupBySew_6_1_12 = bufferStageEnqueueData_6[207:192];
  wire [15:0]       dataRegroupBySew_6_1_13 = bufferStageEnqueueData_6[223:208];
  wire [15:0]       dataRegroupBySew_6_1_14 = bufferStageEnqueueData_6[239:224];
  wire [15:0]       dataRegroupBySew_6_1_15 = bufferStageEnqueueData_6[255:240];
  wire [15:0]       dataRegroupBySew_6_1_16 = bufferStageEnqueueData_6[271:256];
  wire [15:0]       dataRegroupBySew_6_1_17 = bufferStageEnqueueData_6[287:272];
  wire [15:0]       dataRegroupBySew_6_1_18 = bufferStageEnqueueData_6[303:288];
  wire [15:0]       dataRegroupBySew_6_1_19 = bufferStageEnqueueData_6[319:304];
  wire [15:0]       dataRegroupBySew_6_1_20 = bufferStageEnqueueData_6[335:320];
  wire [15:0]       dataRegroupBySew_6_1_21 = bufferStageEnqueueData_6[351:336];
  wire [15:0]       dataRegroupBySew_6_1_22 = bufferStageEnqueueData_6[367:352];
  wire [15:0]       dataRegroupBySew_6_1_23 = bufferStageEnqueueData_6[383:368];
  wire [15:0]       dataRegroupBySew_6_1_24 = bufferStageEnqueueData_6[399:384];
  wire [15:0]       dataRegroupBySew_6_1_25 = bufferStageEnqueueData_6[415:400];
  wire [15:0]       dataRegroupBySew_6_1_26 = bufferStageEnqueueData_6[431:416];
  wire [15:0]       dataRegroupBySew_6_1_27 = bufferStageEnqueueData_6[447:432];
  wire [15:0]       dataRegroupBySew_6_1_28 = bufferStageEnqueueData_6[463:448];
  wire [15:0]       dataRegroupBySew_6_1_29 = bufferStageEnqueueData_6[479:464];
  wire [15:0]       dataRegroupBySew_6_1_30 = bufferStageEnqueueData_6[495:480];
  wire [15:0]       dataRegroupBySew_6_1_31 = bufferStageEnqueueData_6[511:496];
  wire [15:0]       dataRegroupBySew_6_1_32 = bufferStageEnqueueData_6[527:512];
  wire [15:0]       dataRegroupBySew_6_1_33 = bufferStageEnqueueData_6[543:528];
  wire [15:0]       dataRegroupBySew_6_1_34 = bufferStageEnqueueData_6[559:544];
  wire [15:0]       dataRegroupBySew_6_1_35 = bufferStageEnqueueData_6[575:560];
  wire [15:0]       dataRegroupBySew_6_1_36 = bufferStageEnqueueData_6[591:576];
  wire [15:0]       dataRegroupBySew_6_1_37 = bufferStageEnqueueData_6[607:592];
  wire [15:0]       dataRegroupBySew_6_1_38 = bufferStageEnqueueData_6[623:608];
  wire [15:0]       dataRegroupBySew_6_1_39 = bufferStageEnqueueData_6[639:624];
  wire [15:0]       dataRegroupBySew_6_1_40 = bufferStageEnqueueData_6[655:640];
  wire [15:0]       dataRegroupBySew_6_1_41 = bufferStageEnqueueData_6[671:656];
  wire [15:0]       dataRegroupBySew_6_1_42 = bufferStageEnqueueData_6[687:672];
  wire [15:0]       dataRegroupBySew_6_1_43 = bufferStageEnqueueData_6[703:688];
  wire [15:0]       dataRegroupBySew_6_1_44 = bufferStageEnqueueData_6[719:704];
  wire [15:0]       dataRegroupBySew_6_1_45 = bufferStageEnqueueData_6[735:720];
  wire [15:0]       dataRegroupBySew_6_1_46 = bufferStageEnqueueData_6[751:736];
  wire [15:0]       dataRegroupBySew_6_1_47 = bufferStageEnqueueData_6[767:752];
  wire [15:0]       dataRegroupBySew_6_1_48 = bufferStageEnqueueData_6[783:768];
  wire [15:0]       dataRegroupBySew_6_1_49 = bufferStageEnqueueData_6[799:784];
  wire [15:0]       dataRegroupBySew_6_1_50 = bufferStageEnqueueData_6[815:800];
  wire [15:0]       dataRegroupBySew_6_1_51 = bufferStageEnqueueData_6[831:816];
  wire [15:0]       dataRegroupBySew_6_1_52 = bufferStageEnqueueData_6[847:832];
  wire [15:0]       dataRegroupBySew_6_1_53 = bufferStageEnqueueData_6[863:848];
  wire [15:0]       dataRegroupBySew_6_1_54 = bufferStageEnqueueData_6[879:864];
  wire [15:0]       dataRegroupBySew_6_1_55 = bufferStageEnqueueData_6[895:880];
  wire [15:0]       dataRegroupBySew_6_1_56 = bufferStageEnqueueData_6[911:896];
  wire [15:0]       dataRegroupBySew_6_1_57 = bufferStageEnqueueData_6[927:912];
  wire [15:0]       dataRegroupBySew_6_1_58 = bufferStageEnqueueData_6[943:928];
  wire [15:0]       dataRegroupBySew_6_1_59 = bufferStageEnqueueData_6[959:944];
  wire [15:0]       dataRegroupBySew_6_1_60 = bufferStageEnqueueData_6[975:960];
  wire [15:0]       dataRegroupBySew_6_1_61 = bufferStageEnqueueData_6[991:976];
  wire [15:0]       dataRegroupBySew_6_1_62 = bufferStageEnqueueData_6[1007:992];
  wire [15:0]       dataRegroupBySew_6_1_63 = bufferStageEnqueueData_6[1023:1008];
  wire [15:0]       dataRegroupBySew_7_1_0 = bufferStageEnqueueData_7[15:0];
  wire [15:0]       dataRegroupBySew_7_1_1 = bufferStageEnqueueData_7[31:16];
  wire [15:0]       dataRegroupBySew_7_1_2 = bufferStageEnqueueData_7[47:32];
  wire [15:0]       dataRegroupBySew_7_1_3 = bufferStageEnqueueData_7[63:48];
  wire [15:0]       dataRegroupBySew_7_1_4 = bufferStageEnqueueData_7[79:64];
  wire [15:0]       dataRegroupBySew_7_1_5 = bufferStageEnqueueData_7[95:80];
  wire [15:0]       dataRegroupBySew_7_1_6 = bufferStageEnqueueData_7[111:96];
  wire [15:0]       dataRegroupBySew_7_1_7 = bufferStageEnqueueData_7[127:112];
  wire [15:0]       dataRegroupBySew_7_1_8 = bufferStageEnqueueData_7[143:128];
  wire [15:0]       dataRegroupBySew_7_1_9 = bufferStageEnqueueData_7[159:144];
  wire [15:0]       dataRegroupBySew_7_1_10 = bufferStageEnqueueData_7[175:160];
  wire [15:0]       dataRegroupBySew_7_1_11 = bufferStageEnqueueData_7[191:176];
  wire [15:0]       dataRegroupBySew_7_1_12 = bufferStageEnqueueData_7[207:192];
  wire [15:0]       dataRegroupBySew_7_1_13 = bufferStageEnqueueData_7[223:208];
  wire [15:0]       dataRegroupBySew_7_1_14 = bufferStageEnqueueData_7[239:224];
  wire [15:0]       dataRegroupBySew_7_1_15 = bufferStageEnqueueData_7[255:240];
  wire [15:0]       dataRegroupBySew_7_1_16 = bufferStageEnqueueData_7[271:256];
  wire [15:0]       dataRegroupBySew_7_1_17 = bufferStageEnqueueData_7[287:272];
  wire [15:0]       dataRegroupBySew_7_1_18 = bufferStageEnqueueData_7[303:288];
  wire [15:0]       dataRegroupBySew_7_1_19 = bufferStageEnqueueData_7[319:304];
  wire [15:0]       dataRegroupBySew_7_1_20 = bufferStageEnqueueData_7[335:320];
  wire [15:0]       dataRegroupBySew_7_1_21 = bufferStageEnqueueData_7[351:336];
  wire [15:0]       dataRegroupBySew_7_1_22 = bufferStageEnqueueData_7[367:352];
  wire [15:0]       dataRegroupBySew_7_1_23 = bufferStageEnqueueData_7[383:368];
  wire [15:0]       dataRegroupBySew_7_1_24 = bufferStageEnqueueData_7[399:384];
  wire [15:0]       dataRegroupBySew_7_1_25 = bufferStageEnqueueData_7[415:400];
  wire [15:0]       dataRegroupBySew_7_1_26 = bufferStageEnqueueData_7[431:416];
  wire [15:0]       dataRegroupBySew_7_1_27 = bufferStageEnqueueData_7[447:432];
  wire [15:0]       dataRegroupBySew_7_1_28 = bufferStageEnqueueData_7[463:448];
  wire [15:0]       dataRegroupBySew_7_1_29 = bufferStageEnqueueData_7[479:464];
  wire [15:0]       dataRegroupBySew_7_1_30 = bufferStageEnqueueData_7[495:480];
  wire [15:0]       dataRegroupBySew_7_1_31 = bufferStageEnqueueData_7[511:496];
  wire [15:0]       dataRegroupBySew_7_1_32 = bufferStageEnqueueData_7[527:512];
  wire [15:0]       dataRegroupBySew_7_1_33 = bufferStageEnqueueData_7[543:528];
  wire [15:0]       dataRegroupBySew_7_1_34 = bufferStageEnqueueData_7[559:544];
  wire [15:0]       dataRegroupBySew_7_1_35 = bufferStageEnqueueData_7[575:560];
  wire [15:0]       dataRegroupBySew_7_1_36 = bufferStageEnqueueData_7[591:576];
  wire [15:0]       dataRegroupBySew_7_1_37 = bufferStageEnqueueData_7[607:592];
  wire [15:0]       dataRegroupBySew_7_1_38 = bufferStageEnqueueData_7[623:608];
  wire [15:0]       dataRegroupBySew_7_1_39 = bufferStageEnqueueData_7[639:624];
  wire [15:0]       dataRegroupBySew_7_1_40 = bufferStageEnqueueData_7[655:640];
  wire [15:0]       dataRegroupBySew_7_1_41 = bufferStageEnqueueData_7[671:656];
  wire [15:0]       dataRegroupBySew_7_1_42 = bufferStageEnqueueData_7[687:672];
  wire [15:0]       dataRegroupBySew_7_1_43 = bufferStageEnqueueData_7[703:688];
  wire [15:0]       dataRegroupBySew_7_1_44 = bufferStageEnqueueData_7[719:704];
  wire [15:0]       dataRegroupBySew_7_1_45 = bufferStageEnqueueData_7[735:720];
  wire [15:0]       dataRegroupBySew_7_1_46 = bufferStageEnqueueData_7[751:736];
  wire [15:0]       dataRegroupBySew_7_1_47 = bufferStageEnqueueData_7[767:752];
  wire [15:0]       dataRegroupBySew_7_1_48 = bufferStageEnqueueData_7[783:768];
  wire [15:0]       dataRegroupBySew_7_1_49 = bufferStageEnqueueData_7[799:784];
  wire [15:0]       dataRegroupBySew_7_1_50 = bufferStageEnqueueData_7[815:800];
  wire [15:0]       dataRegroupBySew_7_1_51 = bufferStageEnqueueData_7[831:816];
  wire [15:0]       dataRegroupBySew_7_1_52 = bufferStageEnqueueData_7[847:832];
  wire [15:0]       dataRegroupBySew_7_1_53 = bufferStageEnqueueData_7[863:848];
  wire [15:0]       dataRegroupBySew_7_1_54 = bufferStageEnqueueData_7[879:864];
  wire [15:0]       dataRegroupBySew_7_1_55 = bufferStageEnqueueData_7[895:880];
  wire [15:0]       dataRegroupBySew_7_1_56 = bufferStageEnqueueData_7[911:896];
  wire [15:0]       dataRegroupBySew_7_1_57 = bufferStageEnqueueData_7[927:912];
  wire [15:0]       dataRegroupBySew_7_1_58 = bufferStageEnqueueData_7[943:928];
  wire [15:0]       dataRegroupBySew_7_1_59 = bufferStageEnqueueData_7[959:944];
  wire [15:0]       dataRegroupBySew_7_1_60 = bufferStageEnqueueData_7[975:960];
  wire [15:0]       dataRegroupBySew_7_1_61 = bufferStageEnqueueData_7[991:976];
  wire [15:0]       dataRegroupBySew_7_1_62 = bufferStageEnqueueData_7[1007:992];
  wire [15:0]       dataRegroupBySew_7_1_63 = bufferStageEnqueueData_7[1023:1008];
  wire [31:0]       dataInMem_lo_lo_lo_lo_lo_8 = {dataRegroupBySew_0_1_1, dataRegroupBySew_0_1_0};
  wire [31:0]       dataInMem_lo_lo_lo_lo_hi_8 = {dataRegroupBySew_0_1_3, dataRegroupBySew_0_1_2};
  wire [63:0]       dataInMem_lo_lo_lo_lo_8 = {dataInMem_lo_lo_lo_lo_hi_8, dataInMem_lo_lo_lo_lo_lo_8};
  wire [31:0]       dataInMem_lo_lo_lo_hi_lo_8 = {dataRegroupBySew_0_1_5, dataRegroupBySew_0_1_4};
  wire [31:0]       dataInMem_lo_lo_lo_hi_hi_8 = {dataRegroupBySew_0_1_7, dataRegroupBySew_0_1_6};
  wire [63:0]       dataInMem_lo_lo_lo_hi_8 = {dataInMem_lo_lo_lo_hi_hi_8, dataInMem_lo_lo_lo_hi_lo_8};
  wire [127:0]      dataInMem_lo_lo_lo_8 = {dataInMem_lo_lo_lo_hi_8, dataInMem_lo_lo_lo_lo_8};
  wire [31:0]       dataInMem_lo_lo_hi_lo_lo_8 = {dataRegroupBySew_0_1_9, dataRegroupBySew_0_1_8};
  wire [31:0]       dataInMem_lo_lo_hi_lo_hi_8 = {dataRegroupBySew_0_1_11, dataRegroupBySew_0_1_10};
  wire [63:0]       dataInMem_lo_lo_hi_lo_8 = {dataInMem_lo_lo_hi_lo_hi_8, dataInMem_lo_lo_hi_lo_lo_8};
  wire [31:0]       dataInMem_lo_lo_hi_hi_lo_8 = {dataRegroupBySew_0_1_13, dataRegroupBySew_0_1_12};
  wire [31:0]       dataInMem_lo_lo_hi_hi_hi_8 = {dataRegroupBySew_0_1_15, dataRegroupBySew_0_1_14};
  wire [63:0]       dataInMem_lo_lo_hi_hi_8 = {dataInMem_lo_lo_hi_hi_hi_8, dataInMem_lo_lo_hi_hi_lo_8};
  wire [127:0]      dataInMem_lo_lo_hi_8 = {dataInMem_lo_lo_hi_hi_8, dataInMem_lo_lo_hi_lo_8};
  wire [255:0]      dataInMem_lo_lo_136 = {dataInMem_lo_lo_hi_8, dataInMem_lo_lo_lo_8};
  wire [31:0]       dataInMem_lo_hi_lo_lo_lo_8 = {dataRegroupBySew_0_1_17, dataRegroupBySew_0_1_16};
  wire [31:0]       dataInMem_lo_hi_lo_lo_hi_8 = {dataRegroupBySew_0_1_19, dataRegroupBySew_0_1_18};
  wire [63:0]       dataInMem_lo_hi_lo_lo_8 = {dataInMem_lo_hi_lo_lo_hi_8, dataInMem_lo_hi_lo_lo_lo_8};
  wire [31:0]       dataInMem_lo_hi_lo_hi_lo_8 = {dataRegroupBySew_0_1_21, dataRegroupBySew_0_1_20};
  wire [31:0]       dataInMem_lo_hi_lo_hi_hi_8 = {dataRegroupBySew_0_1_23, dataRegroupBySew_0_1_22};
  wire [63:0]       dataInMem_lo_hi_lo_hi_8 = {dataInMem_lo_hi_lo_hi_hi_8, dataInMem_lo_hi_lo_hi_lo_8};
  wire [127:0]      dataInMem_lo_hi_lo_8 = {dataInMem_lo_hi_lo_hi_8, dataInMem_lo_hi_lo_lo_8};
  wire [31:0]       dataInMem_lo_hi_hi_lo_lo_8 = {dataRegroupBySew_0_1_25, dataRegroupBySew_0_1_24};
  wire [31:0]       dataInMem_lo_hi_hi_lo_hi_8 = {dataRegroupBySew_0_1_27, dataRegroupBySew_0_1_26};
  wire [63:0]       dataInMem_lo_hi_hi_lo_8 = {dataInMem_lo_hi_hi_lo_hi_8, dataInMem_lo_hi_hi_lo_lo_8};
  wire [31:0]       dataInMem_lo_hi_hi_hi_lo_8 = {dataRegroupBySew_0_1_29, dataRegroupBySew_0_1_28};
  wire [31:0]       dataInMem_lo_hi_hi_hi_hi_8 = {dataRegroupBySew_0_1_31, dataRegroupBySew_0_1_30};
  wire [63:0]       dataInMem_lo_hi_hi_hi_8 = {dataInMem_lo_hi_hi_hi_hi_8, dataInMem_lo_hi_hi_hi_lo_8};
  wire [127:0]      dataInMem_lo_hi_hi_8 = {dataInMem_lo_hi_hi_hi_8, dataInMem_lo_hi_hi_lo_8};
  wire [255:0]      dataInMem_lo_hi_392 = {dataInMem_lo_hi_hi_8, dataInMem_lo_hi_lo_8};
  wire [511:0]      dataInMem_lo_648 = {dataInMem_lo_hi_392, dataInMem_lo_lo_136};
  wire [31:0]       dataInMem_hi_lo_lo_lo_lo_8 = {dataRegroupBySew_0_1_33, dataRegroupBySew_0_1_32};
  wire [31:0]       dataInMem_hi_lo_lo_lo_hi_8 = {dataRegroupBySew_0_1_35, dataRegroupBySew_0_1_34};
  wire [63:0]       dataInMem_hi_lo_lo_lo_8 = {dataInMem_hi_lo_lo_lo_hi_8, dataInMem_hi_lo_lo_lo_lo_8};
  wire [31:0]       dataInMem_hi_lo_lo_hi_lo_8 = {dataRegroupBySew_0_1_37, dataRegroupBySew_0_1_36};
  wire [31:0]       dataInMem_hi_lo_lo_hi_hi_8 = {dataRegroupBySew_0_1_39, dataRegroupBySew_0_1_38};
  wire [63:0]       dataInMem_hi_lo_lo_hi_8 = {dataInMem_hi_lo_lo_hi_hi_8, dataInMem_hi_lo_lo_hi_lo_8};
  wire [127:0]      dataInMem_hi_lo_lo_8 = {dataInMem_hi_lo_lo_hi_8, dataInMem_hi_lo_lo_lo_8};
  wire [31:0]       dataInMem_hi_lo_hi_lo_lo_8 = {dataRegroupBySew_0_1_41, dataRegroupBySew_0_1_40};
  wire [31:0]       dataInMem_hi_lo_hi_lo_hi_8 = {dataRegroupBySew_0_1_43, dataRegroupBySew_0_1_42};
  wire [63:0]       dataInMem_hi_lo_hi_lo_8 = {dataInMem_hi_lo_hi_lo_hi_8, dataInMem_hi_lo_hi_lo_lo_8};
  wire [31:0]       dataInMem_hi_lo_hi_hi_lo_8 = {dataRegroupBySew_0_1_45, dataRegroupBySew_0_1_44};
  wire [31:0]       dataInMem_hi_lo_hi_hi_hi_8 = {dataRegroupBySew_0_1_47, dataRegroupBySew_0_1_46};
  wire [63:0]       dataInMem_hi_lo_hi_hi_8 = {dataInMem_hi_lo_hi_hi_hi_8, dataInMem_hi_lo_hi_hi_lo_8};
  wire [127:0]      dataInMem_hi_lo_hi_8 = {dataInMem_hi_lo_hi_hi_8, dataInMem_hi_lo_hi_lo_8};
  wire [255:0]      dataInMem_hi_lo_264 = {dataInMem_hi_lo_hi_8, dataInMem_hi_lo_lo_8};
  wire [31:0]       dataInMem_hi_hi_lo_lo_lo_8 = {dataRegroupBySew_0_1_49, dataRegroupBySew_0_1_48};
  wire [31:0]       dataInMem_hi_hi_lo_lo_hi_8 = {dataRegroupBySew_0_1_51, dataRegroupBySew_0_1_50};
  wire [63:0]       dataInMem_hi_hi_lo_lo_8 = {dataInMem_hi_hi_lo_lo_hi_8, dataInMem_hi_hi_lo_lo_lo_8};
  wire [31:0]       dataInMem_hi_hi_lo_hi_lo_8 = {dataRegroupBySew_0_1_53, dataRegroupBySew_0_1_52};
  wire [31:0]       dataInMem_hi_hi_lo_hi_hi_8 = {dataRegroupBySew_0_1_55, dataRegroupBySew_0_1_54};
  wire [63:0]       dataInMem_hi_hi_lo_hi_8 = {dataInMem_hi_hi_lo_hi_hi_8, dataInMem_hi_hi_lo_hi_lo_8};
  wire [127:0]      dataInMem_hi_hi_lo_8 = {dataInMem_hi_hi_lo_hi_8, dataInMem_hi_hi_lo_lo_8};
  wire [31:0]       dataInMem_hi_hi_hi_lo_lo_8 = {dataRegroupBySew_0_1_57, dataRegroupBySew_0_1_56};
  wire [31:0]       dataInMem_hi_hi_hi_lo_hi_8 = {dataRegroupBySew_0_1_59, dataRegroupBySew_0_1_58};
  wire [63:0]       dataInMem_hi_hi_hi_lo_8 = {dataInMem_hi_hi_hi_lo_hi_8, dataInMem_hi_hi_hi_lo_lo_8};
  wire [31:0]       dataInMem_hi_hi_hi_hi_lo_8 = {dataRegroupBySew_0_1_61, dataRegroupBySew_0_1_60};
  wire [31:0]       dataInMem_hi_hi_hi_hi_hi_8 = {dataRegroupBySew_0_1_63, dataRegroupBySew_0_1_62};
  wire [63:0]       dataInMem_hi_hi_hi_hi_8 = {dataInMem_hi_hi_hi_hi_hi_8, dataInMem_hi_hi_hi_hi_lo_8};
  wire [127:0]      dataInMem_hi_hi_hi_8 = {dataInMem_hi_hi_hi_hi_8, dataInMem_hi_hi_hi_lo_8};
  wire [255:0]      dataInMem_hi_hi_520 = {dataInMem_hi_hi_hi_8, dataInMem_hi_hi_lo_8};
  wire [511:0]      dataInMem_hi_776 = {dataInMem_hi_hi_520, dataInMem_hi_lo_264};
  wire [1023:0]     dataInMem_8 = {dataInMem_hi_776, dataInMem_lo_648};
  wire [1023:0]     regroupCacheLine_8_0 = dataInMem_8;
  wire [1023:0]     res_64 = regroupCacheLine_8_0;
  wire [2047:0]     lo_lo_8 = {1024'h0, res_64};
  wire [4095:0]     lo_8 = {2048'h0, lo_lo_8};
  wire [8191:0]     regroupLoadData_1_0 = {4096'h0, lo_8};
  wire [63:0]       dataInMem_lo_lo_lo_lo_lo_9 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1, dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [63:0]       dataInMem_lo_lo_lo_lo_hi_9 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3, dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [127:0]      dataInMem_lo_lo_lo_lo_9 = {dataInMem_lo_lo_lo_lo_hi_9, dataInMem_lo_lo_lo_lo_lo_9};
  wire [63:0]       dataInMem_lo_lo_lo_hi_lo_9 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5, dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [63:0]       dataInMem_lo_lo_lo_hi_hi_9 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7, dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [127:0]      dataInMem_lo_lo_lo_hi_9 = {dataInMem_lo_lo_lo_hi_hi_9, dataInMem_lo_lo_lo_hi_lo_9};
  wire [255:0]      dataInMem_lo_lo_lo_9 = {dataInMem_lo_lo_lo_hi_9, dataInMem_lo_lo_lo_lo_9};
  wire [63:0]       dataInMem_lo_lo_hi_lo_lo_9 = {dataRegroupBySew_1_1_9, dataRegroupBySew_0_1_9, dataRegroupBySew_1_1_8, dataRegroupBySew_0_1_8};
  wire [63:0]       dataInMem_lo_lo_hi_lo_hi_9 = {dataRegroupBySew_1_1_11, dataRegroupBySew_0_1_11, dataRegroupBySew_1_1_10, dataRegroupBySew_0_1_10};
  wire [127:0]      dataInMem_lo_lo_hi_lo_9 = {dataInMem_lo_lo_hi_lo_hi_9, dataInMem_lo_lo_hi_lo_lo_9};
  wire [63:0]       dataInMem_lo_lo_hi_hi_lo_9 = {dataRegroupBySew_1_1_13, dataRegroupBySew_0_1_13, dataRegroupBySew_1_1_12, dataRegroupBySew_0_1_12};
  wire [63:0]       dataInMem_lo_lo_hi_hi_hi_9 = {dataRegroupBySew_1_1_15, dataRegroupBySew_0_1_15, dataRegroupBySew_1_1_14, dataRegroupBySew_0_1_14};
  wire [127:0]      dataInMem_lo_lo_hi_hi_9 = {dataInMem_lo_lo_hi_hi_hi_9, dataInMem_lo_lo_hi_hi_lo_9};
  wire [255:0]      dataInMem_lo_lo_hi_9 = {dataInMem_lo_lo_hi_hi_9, dataInMem_lo_lo_hi_lo_9};
  wire [511:0]      dataInMem_lo_lo_137 = {dataInMem_lo_lo_hi_9, dataInMem_lo_lo_lo_9};
  wire [63:0]       dataInMem_lo_hi_lo_lo_lo_9 = {dataRegroupBySew_1_1_17, dataRegroupBySew_0_1_17, dataRegroupBySew_1_1_16, dataRegroupBySew_0_1_16};
  wire [63:0]       dataInMem_lo_hi_lo_lo_hi_9 = {dataRegroupBySew_1_1_19, dataRegroupBySew_0_1_19, dataRegroupBySew_1_1_18, dataRegroupBySew_0_1_18};
  wire [127:0]      dataInMem_lo_hi_lo_lo_9 = {dataInMem_lo_hi_lo_lo_hi_9, dataInMem_lo_hi_lo_lo_lo_9};
  wire [63:0]       dataInMem_lo_hi_lo_hi_lo_9 = {dataRegroupBySew_1_1_21, dataRegroupBySew_0_1_21, dataRegroupBySew_1_1_20, dataRegroupBySew_0_1_20};
  wire [63:0]       dataInMem_lo_hi_lo_hi_hi_9 = {dataRegroupBySew_1_1_23, dataRegroupBySew_0_1_23, dataRegroupBySew_1_1_22, dataRegroupBySew_0_1_22};
  wire [127:0]      dataInMem_lo_hi_lo_hi_9 = {dataInMem_lo_hi_lo_hi_hi_9, dataInMem_lo_hi_lo_hi_lo_9};
  wire [255:0]      dataInMem_lo_hi_lo_9 = {dataInMem_lo_hi_lo_hi_9, dataInMem_lo_hi_lo_lo_9};
  wire [63:0]       dataInMem_lo_hi_hi_lo_lo_9 = {dataRegroupBySew_1_1_25, dataRegroupBySew_0_1_25, dataRegroupBySew_1_1_24, dataRegroupBySew_0_1_24};
  wire [63:0]       dataInMem_lo_hi_hi_lo_hi_9 = {dataRegroupBySew_1_1_27, dataRegroupBySew_0_1_27, dataRegroupBySew_1_1_26, dataRegroupBySew_0_1_26};
  wire [127:0]      dataInMem_lo_hi_hi_lo_9 = {dataInMem_lo_hi_hi_lo_hi_9, dataInMem_lo_hi_hi_lo_lo_9};
  wire [63:0]       dataInMem_lo_hi_hi_hi_lo_9 = {dataRegroupBySew_1_1_29, dataRegroupBySew_0_1_29, dataRegroupBySew_1_1_28, dataRegroupBySew_0_1_28};
  wire [63:0]       dataInMem_lo_hi_hi_hi_hi_9 = {dataRegroupBySew_1_1_31, dataRegroupBySew_0_1_31, dataRegroupBySew_1_1_30, dataRegroupBySew_0_1_30};
  wire [127:0]      dataInMem_lo_hi_hi_hi_9 = {dataInMem_lo_hi_hi_hi_hi_9, dataInMem_lo_hi_hi_hi_lo_9};
  wire [255:0]      dataInMem_lo_hi_hi_9 = {dataInMem_lo_hi_hi_hi_9, dataInMem_lo_hi_hi_lo_9};
  wire [511:0]      dataInMem_lo_hi_393 = {dataInMem_lo_hi_hi_9, dataInMem_lo_hi_lo_9};
  wire [1023:0]     dataInMem_lo_649 = {dataInMem_lo_hi_393, dataInMem_lo_lo_137};
  wire [63:0]       dataInMem_hi_lo_lo_lo_lo_9 = {dataRegroupBySew_1_1_33, dataRegroupBySew_0_1_33, dataRegroupBySew_1_1_32, dataRegroupBySew_0_1_32};
  wire [63:0]       dataInMem_hi_lo_lo_lo_hi_9 = {dataRegroupBySew_1_1_35, dataRegroupBySew_0_1_35, dataRegroupBySew_1_1_34, dataRegroupBySew_0_1_34};
  wire [127:0]      dataInMem_hi_lo_lo_lo_9 = {dataInMem_hi_lo_lo_lo_hi_9, dataInMem_hi_lo_lo_lo_lo_9};
  wire [63:0]       dataInMem_hi_lo_lo_hi_lo_9 = {dataRegroupBySew_1_1_37, dataRegroupBySew_0_1_37, dataRegroupBySew_1_1_36, dataRegroupBySew_0_1_36};
  wire [63:0]       dataInMem_hi_lo_lo_hi_hi_9 = {dataRegroupBySew_1_1_39, dataRegroupBySew_0_1_39, dataRegroupBySew_1_1_38, dataRegroupBySew_0_1_38};
  wire [127:0]      dataInMem_hi_lo_lo_hi_9 = {dataInMem_hi_lo_lo_hi_hi_9, dataInMem_hi_lo_lo_hi_lo_9};
  wire [255:0]      dataInMem_hi_lo_lo_9 = {dataInMem_hi_lo_lo_hi_9, dataInMem_hi_lo_lo_lo_9};
  wire [63:0]       dataInMem_hi_lo_hi_lo_lo_9 = {dataRegroupBySew_1_1_41, dataRegroupBySew_0_1_41, dataRegroupBySew_1_1_40, dataRegroupBySew_0_1_40};
  wire [63:0]       dataInMem_hi_lo_hi_lo_hi_9 = {dataRegroupBySew_1_1_43, dataRegroupBySew_0_1_43, dataRegroupBySew_1_1_42, dataRegroupBySew_0_1_42};
  wire [127:0]      dataInMem_hi_lo_hi_lo_9 = {dataInMem_hi_lo_hi_lo_hi_9, dataInMem_hi_lo_hi_lo_lo_9};
  wire [63:0]       dataInMem_hi_lo_hi_hi_lo_9 = {dataRegroupBySew_1_1_45, dataRegroupBySew_0_1_45, dataRegroupBySew_1_1_44, dataRegroupBySew_0_1_44};
  wire [63:0]       dataInMem_hi_lo_hi_hi_hi_9 = {dataRegroupBySew_1_1_47, dataRegroupBySew_0_1_47, dataRegroupBySew_1_1_46, dataRegroupBySew_0_1_46};
  wire [127:0]      dataInMem_hi_lo_hi_hi_9 = {dataInMem_hi_lo_hi_hi_hi_9, dataInMem_hi_lo_hi_hi_lo_9};
  wire [255:0]      dataInMem_hi_lo_hi_9 = {dataInMem_hi_lo_hi_hi_9, dataInMem_hi_lo_hi_lo_9};
  wire [511:0]      dataInMem_hi_lo_265 = {dataInMem_hi_lo_hi_9, dataInMem_hi_lo_lo_9};
  wire [63:0]       dataInMem_hi_hi_lo_lo_lo_9 = {dataRegroupBySew_1_1_49, dataRegroupBySew_0_1_49, dataRegroupBySew_1_1_48, dataRegroupBySew_0_1_48};
  wire [63:0]       dataInMem_hi_hi_lo_lo_hi_9 = {dataRegroupBySew_1_1_51, dataRegroupBySew_0_1_51, dataRegroupBySew_1_1_50, dataRegroupBySew_0_1_50};
  wire [127:0]      dataInMem_hi_hi_lo_lo_9 = {dataInMem_hi_hi_lo_lo_hi_9, dataInMem_hi_hi_lo_lo_lo_9};
  wire [63:0]       dataInMem_hi_hi_lo_hi_lo_9 = {dataRegroupBySew_1_1_53, dataRegroupBySew_0_1_53, dataRegroupBySew_1_1_52, dataRegroupBySew_0_1_52};
  wire [63:0]       dataInMem_hi_hi_lo_hi_hi_9 = {dataRegroupBySew_1_1_55, dataRegroupBySew_0_1_55, dataRegroupBySew_1_1_54, dataRegroupBySew_0_1_54};
  wire [127:0]      dataInMem_hi_hi_lo_hi_9 = {dataInMem_hi_hi_lo_hi_hi_9, dataInMem_hi_hi_lo_hi_lo_9};
  wire [255:0]      dataInMem_hi_hi_lo_9 = {dataInMem_hi_hi_lo_hi_9, dataInMem_hi_hi_lo_lo_9};
  wire [63:0]       dataInMem_hi_hi_hi_lo_lo_9 = {dataRegroupBySew_1_1_57, dataRegroupBySew_0_1_57, dataRegroupBySew_1_1_56, dataRegroupBySew_0_1_56};
  wire [63:0]       dataInMem_hi_hi_hi_lo_hi_9 = {dataRegroupBySew_1_1_59, dataRegroupBySew_0_1_59, dataRegroupBySew_1_1_58, dataRegroupBySew_0_1_58};
  wire [127:0]      dataInMem_hi_hi_hi_lo_9 = {dataInMem_hi_hi_hi_lo_hi_9, dataInMem_hi_hi_hi_lo_lo_9};
  wire [63:0]       dataInMem_hi_hi_hi_hi_lo_9 = {dataRegroupBySew_1_1_61, dataRegroupBySew_0_1_61, dataRegroupBySew_1_1_60, dataRegroupBySew_0_1_60};
  wire [63:0]       dataInMem_hi_hi_hi_hi_hi_9 = {dataRegroupBySew_1_1_63, dataRegroupBySew_0_1_63, dataRegroupBySew_1_1_62, dataRegroupBySew_0_1_62};
  wire [127:0]      dataInMem_hi_hi_hi_hi_9 = {dataInMem_hi_hi_hi_hi_hi_9, dataInMem_hi_hi_hi_hi_lo_9};
  wire [255:0]      dataInMem_hi_hi_hi_9 = {dataInMem_hi_hi_hi_hi_9, dataInMem_hi_hi_hi_lo_9};
  wire [511:0]      dataInMem_hi_hi_521 = {dataInMem_hi_hi_hi_9, dataInMem_hi_hi_lo_9};
  wire [1023:0]     dataInMem_hi_777 = {dataInMem_hi_hi_521, dataInMem_hi_lo_265};
  wire [2047:0]     dataInMem_9 = {dataInMem_hi_777, dataInMem_lo_649};
  wire [1023:0]     regroupCacheLine_9_0 = dataInMem_9[1023:0];
  wire [1023:0]     regroupCacheLine_9_1 = dataInMem_9[2047:1024];
  wire [1023:0]     res_72 = regroupCacheLine_9_0;
  wire [1023:0]     res_73 = regroupCacheLine_9_1;
  wire [2047:0]     lo_lo_9 = {res_73, res_72};
  wire [4095:0]     lo_9 = {2048'h0, lo_lo_9};
  wire [8191:0]     regroupLoadData_1_1 = {4096'h0, lo_9};
  wire [31:0]       _GEN_646 = {dataRegroupBySew_2_1_0, dataRegroupBySew_1_1_0};
  wire [31:0]       dataInMem_hi_778;
  assign dataInMem_hi_778 = _GEN_646;
  wire [31:0]       dataInMem_lo_hi_397;
  assign dataInMem_lo_hi_397 = _GEN_646;
  wire [31:0]       dataInMem_lo_hi_462;
  assign dataInMem_lo_hi_462 = _GEN_646;
  wire [31:0]       _GEN_647 = {dataRegroupBySew_2_1_1, dataRegroupBySew_1_1_1};
  wire [31:0]       dataInMem_hi_779;
  assign dataInMem_hi_779 = _GEN_647;
  wire [31:0]       dataInMem_lo_hi_398;
  assign dataInMem_lo_hi_398 = _GEN_647;
  wire [31:0]       dataInMem_lo_hi_463;
  assign dataInMem_lo_hi_463 = _GEN_647;
  wire [31:0]       _GEN_648 = {dataRegroupBySew_2_1_2, dataRegroupBySew_1_1_2};
  wire [31:0]       dataInMem_hi_780;
  assign dataInMem_hi_780 = _GEN_648;
  wire [31:0]       dataInMem_lo_hi_399;
  assign dataInMem_lo_hi_399 = _GEN_648;
  wire [31:0]       dataInMem_lo_hi_464;
  assign dataInMem_lo_hi_464 = _GEN_648;
  wire [31:0]       _GEN_649 = {dataRegroupBySew_2_1_3, dataRegroupBySew_1_1_3};
  wire [31:0]       dataInMem_hi_781;
  assign dataInMem_hi_781 = _GEN_649;
  wire [31:0]       dataInMem_lo_hi_400;
  assign dataInMem_lo_hi_400 = _GEN_649;
  wire [31:0]       dataInMem_lo_hi_465;
  assign dataInMem_lo_hi_465 = _GEN_649;
  wire [31:0]       _GEN_650 = {dataRegroupBySew_2_1_4, dataRegroupBySew_1_1_4};
  wire [31:0]       dataInMem_hi_782;
  assign dataInMem_hi_782 = _GEN_650;
  wire [31:0]       dataInMem_lo_hi_401;
  assign dataInMem_lo_hi_401 = _GEN_650;
  wire [31:0]       dataInMem_lo_hi_466;
  assign dataInMem_lo_hi_466 = _GEN_650;
  wire [31:0]       _GEN_651 = {dataRegroupBySew_2_1_5, dataRegroupBySew_1_1_5};
  wire [31:0]       dataInMem_hi_783;
  assign dataInMem_hi_783 = _GEN_651;
  wire [31:0]       dataInMem_lo_hi_402;
  assign dataInMem_lo_hi_402 = _GEN_651;
  wire [31:0]       dataInMem_lo_hi_467;
  assign dataInMem_lo_hi_467 = _GEN_651;
  wire [31:0]       _GEN_652 = {dataRegroupBySew_2_1_6, dataRegroupBySew_1_1_6};
  wire [31:0]       dataInMem_hi_784;
  assign dataInMem_hi_784 = _GEN_652;
  wire [31:0]       dataInMem_lo_hi_403;
  assign dataInMem_lo_hi_403 = _GEN_652;
  wire [31:0]       dataInMem_lo_hi_468;
  assign dataInMem_lo_hi_468 = _GEN_652;
  wire [31:0]       _GEN_653 = {dataRegroupBySew_2_1_7, dataRegroupBySew_1_1_7};
  wire [31:0]       dataInMem_hi_785;
  assign dataInMem_hi_785 = _GEN_653;
  wire [31:0]       dataInMem_lo_hi_404;
  assign dataInMem_lo_hi_404 = _GEN_653;
  wire [31:0]       dataInMem_lo_hi_469;
  assign dataInMem_lo_hi_469 = _GEN_653;
  wire [31:0]       _GEN_654 = {dataRegroupBySew_2_1_8, dataRegroupBySew_1_1_8};
  wire [31:0]       dataInMem_hi_786;
  assign dataInMem_hi_786 = _GEN_654;
  wire [31:0]       dataInMem_lo_hi_405;
  assign dataInMem_lo_hi_405 = _GEN_654;
  wire [31:0]       dataInMem_lo_hi_470;
  assign dataInMem_lo_hi_470 = _GEN_654;
  wire [31:0]       _GEN_655 = {dataRegroupBySew_2_1_9, dataRegroupBySew_1_1_9};
  wire [31:0]       dataInMem_hi_787;
  assign dataInMem_hi_787 = _GEN_655;
  wire [31:0]       dataInMem_lo_hi_406;
  assign dataInMem_lo_hi_406 = _GEN_655;
  wire [31:0]       dataInMem_lo_hi_471;
  assign dataInMem_lo_hi_471 = _GEN_655;
  wire [31:0]       _GEN_656 = {dataRegroupBySew_2_1_10, dataRegroupBySew_1_1_10};
  wire [31:0]       dataInMem_hi_788;
  assign dataInMem_hi_788 = _GEN_656;
  wire [31:0]       dataInMem_lo_hi_407;
  assign dataInMem_lo_hi_407 = _GEN_656;
  wire [31:0]       dataInMem_lo_hi_472;
  assign dataInMem_lo_hi_472 = _GEN_656;
  wire [31:0]       _GEN_657 = {dataRegroupBySew_2_1_11, dataRegroupBySew_1_1_11};
  wire [31:0]       dataInMem_hi_789;
  assign dataInMem_hi_789 = _GEN_657;
  wire [31:0]       dataInMem_lo_hi_408;
  assign dataInMem_lo_hi_408 = _GEN_657;
  wire [31:0]       dataInMem_lo_hi_473;
  assign dataInMem_lo_hi_473 = _GEN_657;
  wire [31:0]       _GEN_658 = {dataRegroupBySew_2_1_12, dataRegroupBySew_1_1_12};
  wire [31:0]       dataInMem_hi_790;
  assign dataInMem_hi_790 = _GEN_658;
  wire [31:0]       dataInMem_lo_hi_409;
  assign dataInMem_lo_hi_409 = _GEN_658;
  wire [31:0]       dataInMem_lo_hi_474;
  assign dataInMem_lo_hi_474 = _GEN_658;
  wire [31:0]       _GEN_659 = {dataRegroupBySew_2_1_13, dataRegroupBySew_1_1_13};
  wire [31:0]       dataInMem_hi_791;
  assign dataInMem_hi_791 = _GEN_659;
  wire [31:0]       dataInMem_lo_hi_410;
  assign dataInMem_lo_hi_410 = _GEN_659;
  wire [31:0]       dataInMem_lo_hi_475;
  assign dataInMem_lo_hi_475 = _GEN_659;
  wire [31:0]       _GEN_660 = {dataRegroupBySew_2_1_14, dataRegroupBySew_1_1_14};
  wire [31:0]       dataInMem_hi_792;
  assign dataInMem_hi_792 = _GEN_660;
  wire [31:0]       dataInMem_lo_hi_411;
  assign dataInMem_lo_hi_411 = _GEN_660;
  wire [31:0]       dataInMem_lo_hi_476;
  assign dataInMem_lo_hi_476 = _GEN_660;
  wire [31:0]       _GEN_661 = {dataRegroupBySew_2_1_15, dataRegroupBySew_1_1_15};
  wire [31:0]       dataInMem_hi_793;
  assign dataInMem_hi_793 = _GEN_661;
  wire [31:0]       dataInMem_lo_hi_412;
  assign dataInMem_lo_hi_412 = _GEN_661;
  wire [31:0]       dataInMem_lo_hi_477;
  assign dataInMem_lo_hi_477 = _GEN_661;
  wire [31:0]       _GEN_662 = {dataRegroupBySew_2_1_16, dataRegroupBySew_1_1_16};
  wire [31:0]       dataInMem_hi_794;
  assign dataInMem_hi_794 = _GEN_662;
  wire [31:0]       dataInMem_lo_hi_413;
  assign dataInMem_lo_hi_413 = _GEN_662;
  wire [31:0]       dataInMem_lo_hi_478;
  assign dataInMem_lo_hi_478 = _GEN_662;
  wire [31:0]       _GEN_663 = {dataRegroupBySew_2_1_17, dataRegroupBySew_1_1_17};
  wire [31:0]       dataInMem_hi_795;
  assign dataInMem_hi_795 = _GEN_663;
  wire [31:0]       dataInMem_lo_hi_414;
  assign dataInMem_lo_hi_414 = _GEN_663;
  wire [31:0]       dataInMem_lo_hi_479;
  assign dataInMem_lo_hi_479 = _GEN_663;
  wire [31:0]       _GEN_664 = {dataRegroupBySew_2_1_18, dataRegroupBySew_1_1_18};
  wire [31:0]       dataInMem_hi_796;
  assign dataInMem_hi_796 = _GEN_664;
  wire [31:0]       dataInMem_lo_hi_415;
  assign dataInMem_lo_hi_415 = _GEN_664;
  wire [31:0]       dataInMem_lo_hi_480;
  assign dataInMem_lo_hi_480 = _GEN_664;
  wire [31:0]       _GEN_665 = {dataRegroupBySew_2_1_19, dataRegroupBySew_1_1_19};
  wire [31:0]       dataInMem_hi_797;
  assign dataInMem_hi_797 = _GEN_665;
  wire [31:0]       dataInMem_lo_hi_416;
  assign dataInMem_lo_hi_416 = _GEN_665;
  wire [31:0]       dataInMem_lo_hi_481;
  assign dataInMem_lo_hi_481 = _GEN_665;
  wire [31:0]       _GEN_666 = {dataRegroupBySew_2_1_20, dataRegroupBySew_1_1_20};
  wire [31:0]       dataInMem_hi_798;
  assign dataInMem_hi_798 = _GEN_666;
  wire [31:0]       dataInMem_lo_hi_417;
  assign dataInMem_lo_hi_417 = _GEN_666;
  wire [31:0]       dataInMem_lo_hi_482;
  assign dataInMem_lo_hi_482 = _GEN_666;
  wire [31:0]       _GEN_667 = {dataRegroupBySew_2_1_21, dataRegroupBySew_1_1_21};
  wire [31:0]       dataInMem_hi_799;
  assign dataInMem_hi_799 = _GEN_667;
  wire [31:0]       dataInMem_lo_hi_418;
  assign dataInMem_lo_hi_418 = _GEN_667;
  wire [31:0]       dataInMem_lo_hi_483;
  assign dataInMem_lo_hi_483 = _GEN_667;
  wire [31:0]       _GEN_668 = {dataRegroupBySew_2_1_22, dataRegroupBySew_1_1_22};
  wire [31:0]       dataInMem_hi_800;
  assign dataInMem_hi_800 = _GEN_668;
  wire [31:0]       dataInMem_lo_hi_419;
  assign dataInMem_lo_hi_419 = _GEN_668;
  wire [31:0]       dataInMem_lo_hi_484;
  assign dataInMem_lo_hi_484 = _GEN_668;
  wire [31:0]       _GEN_669 = {dataRegroupBySew_2_1_23, dataRegroupBySew_1_1_23};
  wire [31:0]       dataInMem_hi_801;
  assign dataInMem_hi_801 = _GEN_669;
  wire [31:0]       dataInMem_lo_hi_420;
  assign dataInMem_lo_hi_420 = _GEN_669;
  wire [31:0]       dataInMem_lo_hi_485;
  assign dataInMem_lo_hi_485 = _GEN_669;
  wire [31:0]       _GEN_670 = {dataRegroupBySew_2_1_24, dataRegroupBySew_1_1_24};
  wire [31:0]       dataInMem_hi_802;
  assign dataInMem_hi_802 = _GEN_670;
  wire [31:0]       dataInMem_lo_hi_421;
  assign dataInMem_lo_hi_421 = _GEN_670;
  wire [31:0]       dataInMem_lo_hi_486;
  assign dataInMem_lo_hi_486 = _GEN_670;
  wire [31:0]       _GEN_671 = {dataRegroupBySew_2_1_25, dataRegroupBySew_1_1_25};
  wire [31:0]       dataInMem_hi_803;
  assign dataInMem_hi_803 = _GEN_671;
  wire [31:0]       dataInMem_lo_hi_422;
  assign dataInMem_lo_hi_422 = _GEN_671;
  wire [31:0]       dataInMem_lo_hi_487;
  assign dataInMem_lo_hi_487 = _GEN_671;
  wire [31:0]       _GEN_672 = {dataRegroupBySew_2_1_26, dataRegroupBySew_1_1_26};
  wire [31:0]       dataInMem_hi_804;
  assign dataInMem_hi_804 = _GEN_672;
  wire [31:0]       dataInMem_lo_hi_423;
  assign dataInMem_lo_hi_423 = _GEN_672;
  wire [31:0]       dataInMem_lo_hi_488;
  assign dataInMem_lo_hi_488 = _GEN_672;
  wire [31:0]       _GEN_673 = {dataRegroupBySew_2_1_27, dataRegroupBySew_1_1_27};
  wire [31:0]       dataInMem_hi_805;
  assign dataInMem_hi_805 = _GEN_673;
  wire [31:0]       dataInMem_lo_hi_424;
  assign dataInMem_lo_hi_424 = _GEN_673;
  wire [31:0]       dataInMem_lo_hi_489;
  assign dataInMem_lo_hi_489 = _GEN_673;
  wire [31:0]       _GEN_674 = {dataRegroupBySew_2_1_28, dataRegroupBySew_1_1_28};
  wire [31:0]       dataInMem_hi_806;
  assign dataInMem_hi_806 = _GEN_674;
  wire [31:0]       dataInMem_lo_hi_425;
  assign dataInMem_lo_hi_425 = _GEN_674;
  wire [31:0]       dataInMem_lo_hi_490;
  assign dataInMem_lo_hi_490 = _GEN_674;
  wire [31:0]       _GEN_675 = {dataRegroupBySew_2_1_29, dataRegroupBySew_1_1_29};
  wire [31:0]       dataInMem_hi_807;
  assign dataInMem_hi_807 = _GEN_675;
  wire [31:0]       dataInMem_lo_hi_426;
  assign dataInMem_lo_hi_426 = _GEN_675;
  wire [31:0]       dataInMem_lo_hi_491;
  assign dataInMem_lo_hi_491 = _GEN_675;
  wire [31:0]       _GEN_676 = {dataRegroupBySew_2_1_30, dataRegroupBySew_1_1_30};
  wire [31:0]       dataInMem_hi_808;
  assign dataInMem_hi_808 = _GEN_676;
  wire [31:0]       dataInMem_lo_hi_427;
  assign dataInMem_lo_hi_427 = _GEN_676;
  wire [31:0]       dataInMem_lo_hi_492;
  assign dataInMem_lo_hi_492 = _GEN_676;
  wire [31:0]       _GEN_677 = {dataRegroupBySew_2_1_31, dataRegroupBySew_1_1_31};
  wire [31:0]       dataInMem_hi_809;
  assign dataInMem_hi_809 = _GEN_677;
  wire [31:0]       dataInMem_lo_hi_428;
  assign dataInMem_lo_hi_428 = _GEN_677;
  wire [31:0]       dataInMem_lo_hi_493;
  assign dataInMem_lo_hi_493 = _GEN_677;
  wire [31:0]       _GEN_678 = {dataRegroupBySew_2_1_32, dataRegroupBySew_1_1_32};
  wire [31:0]       dataInMem_hi_810;
  assign dataInMem_hi_810 = _GEN_678;
  wire [31:0]       dataInMem_lo_hi_429;
  assign dataInMem_lo_hi_429 = _GEN_678;
  wire [31:0]       dataInMem_lo_hi_494;
  assign dataInMem_lo_hi_494 = _GEN_678;
  wire [31:0]       _GEN_679 = {dataRegroupBySew_2_1_33, dataRegroupBySew_1_1_33};
  wire [31:0]       dataInMem_hi_811;
  assign dataInMem_hi_811 = _GEN_679;
  wire [31:0]       dataInMem_lo_hi_430;
  assign dataInMem_lo_hi_430 = _GEN_679;
  wire [31:0]       dataInMem_lo_hi_495;
  assign dataInMem_lo_hi_495 = _GEN_679;
  wire [31:0]       _GEN_680 = {dataRegroupBySew_2_1_34, dataRegroupBySew_1_1_34};
  wire [31:0]       dataInMem_hi_812;
  assign dataInMem_hi_812 = _GEN_680;
  wire [31:0]       dataInMem_lo_hi_431;
  assign dataInMem_lo_hi_431 = _GEN_680;
  wire [31:0]       dataInMem_lo_hi_496;
  assign dataInMem_lo_hi_496 = _GEN_680;
  wire [31:0]       _GEN_681 = {dataRegroupBySew_2_1_35, dataRegroupBySew_1_1_35};
  wire [31:0]       dataInMem_hi_813;
  assign dataInMem_hi_813 = _GEN_681;
  wire [31:0]       dataInMem_lo_hi_432;
  assign dataInMem_lo_hi_432 = _GEN_681;
  wire [31:0]       dataInMem_lo_hi_497;
  assign dataInMem_lo_hi_497 = _GEN_681;
  wire [31:0]       _GEN_682 = {dataRegroupBySew_2_1_36, dataRegroupBySew_1_1_36};
  wire [31:0]       dataInMem_hi_814;
  assign dataInMem_hi_814 = _GEN_682;
  wire [31:0]       dataInMem_lo_hi_433;
  assign dataInMem_lo_hi_433 = _GEN_682;
  wire [31:0]       dataInMem_lo_hi_498;
  assign dataInMem_lo_hi_498 = _GEN_682;
  wire [31:0]       _GEN_683 = {dataRegroupBySew_2_1_37, dataRegroupBySew_1_1_37};
  wire [31:0]       dataInMem_hi_815;
  assign dataInMem_hi_815 = _GEN_683;
  wire [31:0]       dataInMem_lo_hi_434;
  assign dataInMem_lo_hi_434 = _GEN_683;
  wire [31:0]       dataInMem_lo_hi_499;
  assign dataInMem_lo_hi_499 = _GEN_683;
  wire [31:0]       _GEN_684 = {dataRegroupBySew_2_1_38, dataRegroupBySew_1_1_38};
  wire [31:0]       dataInMem_hi_816;
  assign dataInMem_hi_816 = _GEN_684;
  wire [31:0]       dataInMem_lo_hi_435;
  assign dataInMem_lo_hi_435 = _GEN_684;
  wire [31:0]       dataInMem_lo_hi_500;
  assign dataInMem_lo_hi_500 = _GEN_684;
  wire [31:0]       _GEN_685 = {dataRegroupBySew_2_1_39, dataRegroupBySew_1_1_39};
  wire [31:0]       dataInMem_hi_817;
  assign dataInMem_hi_817 = _GEN_685;
  wire [31:0]       dataInMem_lo_hi_436;
  assign dataInMem_lo_hi_436 = _GEN_685;
  wire [31:0]       dataInMem_lo_hi_501;
  assign dataInMem_lo_hi_501 = _GEN_685;
  wire [31:0]       _GEN_686 = {dataRegroupBySew_2_1_40, dataRegroupBySew_1_1_40};
  wire [31:0]       dataInMem_hi_818;
  assign dataInMem_hi_818 = _GEN_686;
  wire [31:0]       dataInMem_lo_hi_437;
  assign dataInMem_lo_hi_437 = _GEN_686;
  wire [31:0]       dataInMem_lo_hi_502;
  assign dataInMem_lo_hi_502 = _GEN_686;
  wire [31:0]       _GEN_687 = {dataRegroupBySew_2_1_41, dataRegroupBySew_1_1_41};
  wire [31:0]       dataInMem_hi_819;
  assign dataInMem_hi_819 = _GEN_687;
  wire [31:0]       dataInMem_lo_hi_438;
  assign dataInMem_lo_hi_438 = _GEN_687;
  wire [31:0]       dataInMem_lo_hi_503;
  assign dataInMem_lo_hi_503 = _GEN_687;
  wire [31:0]       _GEN_688 = {dataRegroupBySew_2_1_42, dataRegroupBySew_1_1_42};
  wire [31:0]       dataInMem_hi_820;
  assign dataInMem_hi_820 = _GEN_688;
  wire [31:0]       dataInMem_lo_hi_439;
  assign dataInMem_lo_hi_439 = _GEN_688;
  wire [31:0]       dataInMem_lo_hi_504;
  assign dataInMem_lo_hi_504 = _GEN_688;
  wire [31:0]       _GEN_689 = {dataRegroupBySew_2_1_43, dataRegroupBySew_1_1_43};
  wire [31:0]       dataInMem_hi_821;
  assign dataInMem_hi_821 = _GEN_689;
  wire [31:0]       dataInMem_lo_hi_440;
  assign dataInMem_lo_hi_440 = _GEN_689;
  wire [31:0]       dataInMem_lo_hi_505;
  assign dataInMem_lo_hi_505 = _GEN_689;
  wire [31:0]       _GEN_690 = {dataRegroupBySew_2_1_44, dataRegroupBySew_1_1_44};
  wire [31:0]       dataInMem_hi_822;
  assign dataInMem_hi_822 = _GEN_690;
  wire [31:0]       dataInMem_lo_hi_441;
  assign dataInMem_lo_hi_441 = _GEN_690;
  wire [31:0]       dataInMem_lo_hi_506;
  assign dataInMem_lo_hi_506 = _GEN_690;
  wire [31:0]       _GEN_691 = {dataRegroupBySew_2_1_45, dataRegroupBySew_1_1_45};
  wire [31:0]       dataInMem_hi_823;
  assign dataInMem_hi_823 = _GEN_691;
  wire [31:0]       dataInMem_lo_hi_442;
  assign dataInMem_lo_hi_442 = _GEN_691;
  wire [31:0]       dataInMem_lo_hi_507;
  assign dataInMem_lo_hi_507 = _GEN_691;
  wire [31:0]       _GEN_692 = {dataRegroupBySew_2_1_46, dataRegroupBySew_1_1_46};
  wire [31:0]       dataInMem_hi_824;
  assign dataInMem_hi_824 = _GEN_692;
  wire [31:0]       dataInMem_lo_hi_443;
  assign dataInMem_lo_hi_443 = _GEN_692;
  wire [31:0]       dataInMem_lo_hi_508;
  assign dataInMem_lo_hi_508 = _GEN_692;
  wire [31:0]       _GEN_693 = {dataRegroupBySew_2_1_47, dataRegroupBySew_1_1_47};
  wire [31:0]       dataInMem_hi_825;
  assign dataInMem_hi_825 = _GEN_693;
  wire [31:0]       dataInMem_lo_hi_444;
  assign dataInMem_lo_hi_444 = _GEN_693;
  wire [31:0]       dataInMem_lo_hi_509;
  assign dataInMem_lo_hi_509 = _GEN_693;
  wire [31:0]       _GEN_694 = {dataRegroupBySew_2_1_48, dataRegroupBySew_1_1_48};
  wire [31:0]       dataInMem_hi_826;
  assign dataInMem_hi_826 = _GEN_694;
  wire [31:0]       dataInMem_lo_hi_445;
  assign dataInMem_lo_hi_445 = _GEN_694;
  wire [31:0]       dataInMem_lo_hi_510;
  assign dataInMem_lo_hi_510 = _GEN_694;
  wire [31:0]       _GEN_695 = {dataRegroupBySew_2_1_49, dataRegroupBySew_1_1_49};
  wire [31:0]       dataInMem_hi_827;
  assign dataInMem_hi_827 = _GEN_695;
  wire [31:0]       dataInMem_lo_hi_446;
  assign dataInMem_lo_hi_446 = _GEN_695;
  wire [31:0]       dataInMem_lo_hi_511;
  assign dataInMem_lo_hi_511 = _GEN_695;
  wire [31:0]       _GEN_696 = {dataRegroupBySew_2_1_50, dataRegroupBySew_1_1_50};
  wire [31:0]       dataInMem_hi_828;
  assign dataInMem_hi_828 = _GEN_696;
  wire [31:0]       dataInMem_lo_hi_447;
  assign dataInMem_lo_hi_447 = _GEN_696;
  wire [31:0]       dataInMem_lo_hi_512;
  assign dataInMem_lo_hi_512 = _GEN_696;
  wire [31:0]       _GEN_697 = {dataRegroupBySew_2_1_51, dataRegroupBySew_1_1_51};
  wire [31:0]       dataInMem_hi_829;
  assign dataInMem_hi_829 = _GEN_697;
  wire [31:0]       dataInMem_lo_hi_448;
  assign dataInMem_lo_hi_448 = _GEN_697;
  wire [31:0]       dataInMem_lo_hi_513;
  assign dataInMem_lo_hi_513 = _GEN_697;
  wire [31:0]       _GEN_698 = {dataRegroupBySew_2_1_52, dataRegroupBySew_1_1_52};
  wire [31:0]       dataInMem_hi_830;
  assign dataInMem_hi_830 = _GEN_698;
  wire [31:0]       dataInMem_lo_hi_449;
  assign dataInMem_lo_hi_449 = _GEN_698;
  wire [31:0]       dataInMem_lo_hi_514;
  assign dataInMem_lo_hi_514 = _GEN_698;
  wire [31:0]       _GEN_699 = {dataRegroupBySew_2_1_53, dataRegroupBySew_1_1_53};
  wire [31:0]       dataInMem_hi_831;
  assign dataInMem_hi_831 = _GEN_699;
  wire [31:0]       dataInMem_lo_hi_450;
  assign dataInMem_lo_hi_450 = _GEN_699;
  wire [31:0]       dataInMem_lo_hi_515;
  assign dataInMem_lo_hi_515 = _GEN_699;
  wire [31:0]       _GEN_700 = {dataRegroupBySew_2_1_54, dataRegroupBySew_1_1_54};
  wire [31:0]       dataInMem_hi_832;
  assign dataInMem_hi_832 = _GEN_700;
  wire [31:0]       dataInMem_lo_hi_451;
  assign dataInMem_lo_hi_451 = _GEN_700;
  wire [31:0]       dataInMem_lo_hi_516;
  assign dataInMem_lo_hi_516 = _GEN_700;
  wire [31:0]       _GEN_701 = {dataRegroupBySew_2_1_55, dataRegroupBySew_1_1_55};
  wire [31:0]       dataInMem_hi_833;
  assign dataInMem_hi_833 = _GEN_701;
  wire [31:0]       dataInMem_lo_hi_452;
  assign dataInMem_lo_hi_452 = _GEN_701;
  wire [31:0]       dataInMem_lo_hi_517;
  assign dataInMem_lo_hi_517 = _GEN_701;
  wire [31:0]       _GEN_702 = {dataRegroupBySew_2_1_56, dataRegroupBySew_1_1_56};
  wire [31:0]       dataInMem_hi_834;
  assign dataInMem_hi_834 = _GEN_702;
  wire [31:0]       dataInMem_lo_hi_453;
  assign dataInMem_lo_hi_453 = _GEN_702;
  wire [31:0]       dataInMem_lo_hi_518;
  assign dataInMem_lo_hi_518 = _GEN_702;
  wire [31:0]       _GEN_703 = {dataRegroupBySew_2_1_57, dataRegroupBySew_1_1_57};
  wire [31:0]       dataInMem_hi_835;
  assign dataInMem_hi_835 = _GEN_703;
  wire [31:0]       dataInMem_lo_hi_454;
  assign dataInMem_lo_hi_454 = _GEN_703;
  wire [31:0]       dataInMem_lo_hi_519;
  assign dataInMem_lo_hi_519 = _GEN_703;
  wire [31:0]       _GEN_704 = {dataRegroupBySew_2_1_58, dataRegroupBySew_1_1_58};
  wire [31:0]       dataInMem_hi_836;
  assign dataInMem_hi_836 = _GEN_704;
  wire [31:0]       dataInMem_lo_hi_455;
  assign dataInMem_lo_hi_455 = _GEN_704;
  wire [31:0]       dataInMem_lo_hi_520;
  assign dataInMem_lo_hi_520 = _GEN_704;
  wire [31:0]       _GEN_705 = {dataRegroupBySew_2_1_59, dataRegroupBySew_1_1_59};
  wire [31:0]       dataInMem_hi_837;
  assign dataInMem_hi_837 = _GEN_705;
  wire [31:0]       dataInMem_lo_hi_456;
  assign dataInMem_lo_hi_456 = _GEN_705;
  wire [31:0]       dataInMem_lo_hi_521;
  assign dataInMem_lo_hi_521 = _GEN_705;
  wire [31:0]       _GEN_706 = {dataRegroupBySew_2_1_60, dataRegroupBySew_1_1_60};
  wire [31:0]       dataInMem_hi_838;
  assign dataInMem_hi_838 = _GEN_706;
  wire [31:0]       dataInMem_lo_hi_457;
  assign dataInMem_lo_hi_457 = _GEN_706;
  wire [31:0]       dataInMem_lo_hi_522;
  assign dataInMem_lo_hi_522 = _GEN_706;
  wire [31:0]       _GEN_707 = {dataRegroupBySew_2_1_61, dataRegroupBySew_1_1_61};
  wire [31:0]       dataInMem_hi_839;
  assign dataInMem_hi_839 = _GEN_707;
  wire [31:0]       dataInMem_lo_hi_458;
  assign dataInMem_lo_hi_458 = _GEN_707;
  wire [31:0]       dataInMem_lo_hi_523;
  assign dataInMem_lo_hi_523 = _GEN_707;
  wire [31:0]       _GEN_708 = {dataRegroupBySew_2_1_62, dataRegroupBySew_1_1_62};
  wire [31:0]       dataInMem_hi_840;
  assign dataInMem_hi_840 = _GEN_708;
  wire [31:0]       dataInMem_lo_hi_459;
  assign dataInMem_lo_hi_459 = _GEN_708;
  wire [31:0]       dataInMem_lo_hi_524;
  assign dataInMem_lo_hi_524 = _GEN_708;
  wire [31:0]       _GEN_709 = {dataRegroupBySew_2_1_63, dataRegroupBySew_1_1_63};
  wire [31:0]       dataInMem_hi_841;
  assign dataInMem_hi_841 = _GEN_709;
  wire [31:0]       dataInMem_lo_hi_460;
  assign dataInMem_lo_hi_460 = _GEN_709;
  wire [31:0]       dataInMem_lo_hi_525;
  assign dataInMem_lo_hi_525 = _GEN_709;
  wire [95:0]       dataInMem_lo_lo_lo_lo_lo_10 = {dataInMem_hi_779, dataRegroupBySew_0_1_1, dataInMem_hi_778, dataRegroupBySew_0_1_0};
  wire [95:0]       dataInMem_lo_lo_lo_lo_hi_10 = {dataInMem_hi_781, dataRegroupBySew_0_1_3, dataInMem_hi_780, dataRegroupBySew_0_1_2};
  wire [191:0]      dataInMem_lo_lo_lo_lo_10 = {dataInMem_lo_lo_lo_lo_hi_10, dataInMem_lo_lo_lo_lo_lo_10};
  wire [95:0]       dataInMem_lo_lo_lo_hi_lo_10 = {dataInMem_hi_783, dataRegroupBySew_0_1_5, dataInMem_hi_782, dataRegroupBySew_0_1_4};
  wire [95:0]       dataInMem_lo_lo_lo_hi_hi_10 = {dataInMem_hi_785, dataRegroupBySew_0_1_7, dataInMem_hi_784, dataRegroupBySew_0_1_6};
  wire [191:0]      dataInMem_lo_lo_lo_hi_10 = {dataInMem_lo_lo_lo_hi_hi_10, dataInMem_lo_lo_lo_hi_lo_10};
  wire [383:0]      dataInMem_lo_lo_lo_10 = {dataInMem_lo_lo_lo_hi_10, dataInMem_lo_lo_lo_lo_10};
  wire [95:0]       dataInMem_lo_lo_hi_lo_lo_10 = {dataInMem_hi_787, dataRegroupBySew_0_1_9, dataInMem_hi_786, dataRegroupBySew_0_1_8};
  wire [95:0]       dataInMem_lo_lo_hi_lo_hi_10 = {dataInMem_hi_789, dataRegroupBySew_0_1_11, dataInMem_hi_788, dataRegroupBySew_0_1_10};
  wire [191:0]      dataInMem_lo_lo_hi_lo_10 = {dataInMem_lo_lo_hi_lo_hi_10, dataInMem_lo_lo_hi_lo_lo_10};
  wire [95:0]       dataInMem_lo_lo_hi_hi_lo_10 = {dataInMem_hi_791, dataRegroupBySew_0_1_13, dataInMem_hi_790, dataRegroupBySew_0_1_12};
  wire [95:0]       dataInMem_lo_lo_hi_hi_hi_10 = {dataInMem_hi_793, dataRegroupBySew_0_1_15, dataInMem_hi_792, dataRegroupBySew_0_1_14};
  wire [191:0]      dataInMem_lo_lo_hi_hi_10 = {dataInMem_lo_lo_hi_hi_hi_10, dataInMem_lo_lo_hi_hi_lo_10};
  wire [383:0]      dataInMem_lo_lo_hi_10 = {dataInMem_lo_lo_hi_hi_10, dataInMem_lo_lo_hi_lo_10};
  wire [767:0]      dataInMem_lo_lo_138 = {dataInMem_lo_lo_hi_10, dataInMem_lo_lo_lo_10};
  wire [95:0]       dataInMem_lo_hi_lo_lo_lo_10 = {dataInMem_hi_795, dataRegroupBySew_0_1_17, dataInMem_hi_794, dataRegroupBySew_0_1_16};
  wire [95:0]       dataInMem_lo_hi_lo_lo_hi_10 = {dataInMem_hi_797, dataRegroupBySew_0_1_19, dataInMem_hi_796, dataRegroupBySew_0_1_18};
  wire [191:0]      dataInMem_lo_hi_lo_lo_10 = {dataInMem_lo_hi_lo_lo_hi_10, dataInMem_lo_hi_lo_lo_lo_10};
  wire [95:0]       dataInMem_lo_hi_lo_hi_lo_10 = {dataInMem_hi_799, dataRegroupBySew_0_1_21, dataInMem_hi_798, dataRegroupBySew_0_1_20};
  wire [95:0]       dataInMem_lo_hi_lo_hi_hi_10 = {dataInMem_hi_801, dataRegroupBySew_0_1_23, dataInMem_hi_800, dataRegroupBySew_0_1_22};
  wire [191:0]      dataInMem_lo_hi_lo_hi_10 = {dataInMem_lo_hi_lo_hi_hi_10, dataInMem_lo_hi_lo_hi_lo_10};
  wire [383:0]      dataInMem_lo_hi_lo_10 = {dataInMem_lo_hi_lo_hi_10, dataInMem_lo_hi_lo_lo_10};
  wire [95:0]       dataInMem_lo_hi_hi_lo_lo_10 = {dataInMem_hi_803, dataRegroupBySew_0_1_25, dataInMem_hi_802, dataRegroupBySew_0_1_24};
  wire [95:0]       dataInMem_lo_hi_hi_lo_hi_10 = {dataInMem_hi_805, dataRegroupBySew_0_1_27, dataInMem_hi_804, dataRegroupBySew_0_1_26};
  wire [191:0]      dataInMem_lo_hi_hi_lo_10 = {dataInMem_lo_hi_hi_lo_hi_10, dataInMem_lo_hi_hi_lo_lo_10};
  wire [95:0]       dataInMem_lo_hi_hi_hi_lo_10 = {dataInMem_hi_807, dataRegroupBySew_0_1_29, dataInMem_hi_806, dataRegroupBySew_0_1_28};
  wire [95:0]       dataInMem_lo_hi_hi_hi_hi_10 = {dataInMem_hi_809, dataRegroupBySew_0_1_31, dataInMem_hi_808, dataRegroupBySew_0_1_30};
  wire [191:0]      dataInMem_lo_hi_hi_hi_10 = {dataInMem_lo_hi_hi_hi_hi_10, dataInMem_lo_hi_hi_hi_lo_10};
  wire [383:0]      dataInMem_lo_hi_hi_10 = {dataInMem_lo_hi_hi_hi_10, dataInMem_lo_hi_hi_lo_10};
  wire [767:0]      dataInMem_lo_hi_394 = {dataInMem_lo_hi_hi_10, dataInMem_lo_hi_lo_10};
  wire [1535:0]     dataInMem_lo_650 = {dataInMem_lo_hi_394, dataInMem_lo_lo_138};
  wire [95:0]       dataInMem_hi_lo_lo_lo_lo_10 = {dataInMem_hi_811, dataRegroupBySew_0_1_33, dataInMem_hi_810, dataRegroupBySew_0_1_32};
  wire [95:0]       dataInMem_hi_lo_lo_lo_hi_10 = {dataInMem_hi_813, dataRegroupBySew_0_1_35, dataInMem_hi_812, dataRegroupBySew_0_1_34};
  wire [191:0]      dataInMem_hi_lo_lo_lo_10 = {dataInMem_hi_lo_lo_lo_hi_10, dataInMem_hi_lo_lo_lo_lo_10};
  wire [95:0]       dataInMem_hi_lo_lo_hi_lo_10 = {dataInMem_hi_815, dataRegroupBySew_0_1_37, dataInMem_hi_814, dataRegroupBySew_0_1_36};
  wire [95:0]       dataInMem_hi_lo_lo_hi_hi_10 = {dataInMem_hi_817, dataRegroupBySew_0_1_39, dataInMem_hi_816, dataRegroupBySew_0_1_38};
  wire [191:0]      dataInMem_hi_lo_lo_hi_10 = {dataInMem_hi_lo_lo_hi_hi_10, dataInMem_hi_lo_lo_hi_lo_10};
  wire [383:0]      dataInMem_hi_lo_lo_10 = {dataInMem_hi_lo_lo_hi_10, dataInMem_hi_lo_lo_lo_10};
  wire [95:0]       dataInMem_hi_lo_hi_lo_lo_10 = {dataInMem_hi_819, dataRegroupBySew_0_1_41, dataInMem_hi_818, dataRegroupBySew_0_1_40};
  wire [95:0]       dataInMem_hi_lo_hi_lo_hi_10 = {dataInMem_hi_821, dataRegroupBySew_0_1_43, dataInMem_hi_820, dataRegroupBySew_0_1_42};
  wire [191:0]      dataInMem_hi_lo_hi_lo_10 = {dataInMem_hi_lo_hi_lo_hi_10, dataInMem_hi_lo_hi_lo_lo_10};
  wire [95:0]       dataInMem_hi_lo_hi_hi_lo_10 = {dataInMem_hi_823, dataRegroupBySew_0_1_45, dataInMem_hi_822, dataRegroupBySew_0_1_44};
  wire [95:0]       dataInMem_hi_lo_hi_hi_hi_10 = {dataInMem_hi_825, dataRegroupBySew_0_1_47, dataInMem_hi_824, dataRegroupBySew_0_1_46};
  wire [191:0]      dataInMem_hi_lo_hi_hi_10 = {dataInMem_hi_lo_hi_hi_hi_10, dataInMem_hi_lo_hi_hi_lo_10};
  wire [383:0]      dataInMem_hi_lo_hi_10 = {dataInMem_hi_lo_hi_hi_10, dataInMem_hi_lo_hi_lo_10};
  wire [767:0]      dataInMem_hi_lo_266 = {dataInMem_hi_lo_hi_10, dataInMem_hi_lo_lo_10};
  wire [95:0]       dataInMem_hi_hi_lo_lo_lo_10 = {dataInMem_hi_827, dataRegroupBySew_0_1_49, dataInMem_hi_826, dataRegroupBySew_0_1_48};
  wire [95:0]       dataInMem_hi_hi_lo_lo_hi_10 = {dataInMem_hi_829, dataRegroupBySew_0_1_51, dataInMem_hi_828, dataRegroupBySew_0_1_50};
  wire [191:0]      dataInMem_hi_hi_lo_lo_10 = {dataInMem_hi_hi_lo_lo_hi_10, dataInMem_hi_hi_lo_lo_lo_10};
  wire [95:0]       dataInMem_hi_hi_lo_hi_lo_10 = {dataInMem_hi_831, dataRegroupBySew_0_1_53, dataInMem_hi_830, dataRegroupBySew_0_1_52};
  wire [95:0]       dataInMem_hi_hi_lo_hi_hi_10 = {dataInMem_hi_833, dataRegroupBySew_0_1_55, dataInMem_hi_832, dataRegroupBySew_0_1_54};
  wire [191:0]      dataInMem_hi_hi_lo_hi_10 = {dataInMem_hi_hi_lo_hi_hi_10, dataInMem_hi_hi_lo_hi_lo_10};
  wire [383:0]      dataInMem_hi_hi_lo_10 = {dataInMem_hi_hi_lo_hi_10, dataInMem_hi_hi_lo_lo_10};
  wire [95:0]       dataInMem_hi_hi_hi_lo_lo_10 = {dataInMem_hi_835, dataRegroupBySew_0_1_57, dataInMem_hi_834, dataRegroupBySew_0_1_56};
  wire [95:0]       dataInMem_hi_hi_hi_lo_hi_10 = {dataInMem_hi_837, dataRegroupBySew_0_1_59, dataInMem_hi_836, dataRegroupBySew_0_1_58};
  wire [191:0]      dataInMem_hi_hi_hi_lo_10 = {dataInMem_hi_hi_hi_lo_hi_10, dataInMem_hi_hi_hi_lo_lo_10};
  wire [95:0]       dataInMem_hi_hi_hi_hi_lo_10 = {dataInMem_hi_839, dataRegroupBySew_0_1_61, dataInMem_hi_838, dataRegroupBySew_0_1_60};
  wire [95:0]       dataInMem_hi_hi_hi_hi_hi_10 = {dataInMem_hi_841, dataRegroupBySew_0_1_63, dataInMem_hi_840, dataRegroupBySew_0_1_62};
  wire [191:0]      dataInMem_hi_hi_hi_hi_10 = {dataInMem_hi_hi_hi_hi_hi_10, dataInMem_hi_hi_hi_hi_lo_10};
  wire [383:0]      dataInMem_hi_hi_hi_10 = {dataInMem_hi_hi_hi_hi_10, dataInMem_hi_hi_hi_lo_10};
  wire [767:0]      dataInMem_hi_hi_522 = {dataInMem_hi_hi_hi_10, dataInMem_hi_hi_lo_10};
  wire [1535:0]     dataInMem_hi_842 = {dataInMem_hi_hi_522, dataInMem_hi_lo_266};
  wire [3071:0]     dataInMem_10 = {dataInMem_hi_842, dataInMem_lo_650};
  wire [1023:0]     regroupCacheLine_10_0 = dataInMem_10[1023:0];
  wire [1023:0]     regroupCacheLine_10_1 = dataInMem_10[2047:1024];
  wire [1023:0]     regroupCacheLine_10_2 = dataInMem_10[3071:2048];
  wire [1023:0]     res_80 = regroupCacheLine_10_0;
  wire [1023:0]     res_81 = regroupCacheLine_10_1;
  wire [1023:0]     res_82 = regroupCacheLine_10_2;
  wire [2047:0]     lo_lo_10 = {res_81, res_80};
  wire [2047:0]     lo_hi_10 = {1024'h0, res_82};
  wire [4095:0]     lo_10 = {lo_hi_10, lo_lo_10};
  wire [8191:0]     regroupLoadData_1_2 = {4096'h0, lo_10};
  wire [31:0]       _GEN_710 = {dataRegroupBySew_1_1_0, dataRegroupBySew_0_1_0};
  wire [31:0]       dataInMem_lo_651;
  assign dataInMem_lo_651 = _GEN_710;
  wire [31:0]       dataInMem_lo_716;
  assign dataInMem_lo_716 = _GEN_710;
  wire [31:0]       dataInMem_lo_lo_143;
  assign dataInMem_lo_lo_143 = _GEN_710;
  wire [31:0]       _GEN_711 = {dataRegroupBySew_3_1_0, dataRegroupBySew_2_1_0};
  wire [31:0]       dataInMem_hi_843;
  assign dataInMem_hi_843 = _GEN_711;
  wire [31:0]       dataInMem_lo_hi_527;
  assign dataInMem_lo_hi_527 = _GEN_711;
  wire [31:0]       _GEN_712 = {dataRegroupBySew_1_1_1, dataRegroupBySew_0_1_1};
  wire [31:0]       dataInMem_lo_652;
  assign dataInMem_lo_652 = _GEN_712;
  wire [31:0]       dataInMem_lo_717;
  assign dataInMem_lo_717 = _GEN_712;
  wire [31:0]       dataInMem_lo_lo_144;
  assign dataInMem_lo_lo_144 = _GEN_712;
  wire [31:0]       _GEN_713 = {dataRegroupBySew_3_1_1, dataRegroupBySew_2_1_1};
  wire [31:0]       dataInMem_hi_844;
  assign dataInMem_hi_844 = _GEN_713;
  wire [31:0]       dataInMem_lo_hi_528;
  assign dataInMem_lo_hi_528 = _GEN_713;
  wire [31:0]       _GEN_714 = {dataRegroupBySew_1_1_2, dataRegroupBySew_0_1_2};
  wire [31:0]       dataInMem_lo_653;
  assign dataInMem_lo_653 = _GEN_714;
  wire [31:0]       dataInMem_lo_718;
  assign dataInMem_lo_718 = _GEN_714;
  wire [31:0]       dataInMem_lo_lo_145;
  assign dataInMem_lo_lo_145 = _GEN_714;
  wire [31:0]       _GEN_715 = {dataRegroupBySew_3_1_2, dataRegroupBySew_2_1_2};
  wire [31:0]       dataInMem_hi_845;
  assign dataInMem_hi_845 = _GEN_715;
  wire [31:0]       dataInMem_lo_hi_529;
  assign dataInMem_lo_hi_529 = _GEN_715;
  wire [31:0]       _GEN_716 = {dataRegroupBySew_1_1_3, dataRegroupBySew_0_1_3};
  wire [31:0]       dataInMem_lo_654;
  assign dataInMem_lo_654 = _GEN_716;
  wire [31:0]       dataInMem_lo_719;
  assign dataInMem_lo_719 = _GEN_716;
  wire [31:0]       dataInMem_lo_lo_146;
  assign dataInMem_lo_lo_146 = _GEN_716;
  wire [31:0]       _GEN_717 = {dataRegroupBySew_3_1_3, dataRegroupBySew_2_1_3};
  wire [31:0]       dataInMem_hi_846;
  assign dataInMem_hi_846 = _GEN_717;
  wire [31:0]       dataInMem_lo_hi_530;
  assign dataInMem_lo_hi_530 = _GEN_717;
  wire [31:0]       _GEN_718 = {dataRegroupBySew_1_1_4, dataRegroupBySew_0_1_4};
  wire [31:0]       dataInMem_lo_655;
  assign dataInMem_lo_655 = _GEN_718;
  wire [31:0]       dataInMem_lo_720;
  assign dataInMem_lo_720 = _GEN_718;
  wire [31:0]       dataInMem_lo_lo_147;
  assign dataInMem_lo_lo_147 = _GEN_718;
  wire [31:0]       _GEN_719 = {dataRegroupBySew_3_1_4, dataRegroupBySew_2_1_4};
  wire [31:0]       dataInMem_hi_847;
  assign dataInMem_hi_847 = _GEN_719;
  wire [31:0]       dataInMem_lo_hi_531;
  assign dataInMem_lo_hi_531 = _GEN_719;
  wire [31:0]       _GEN_720 = {dataRegroupBySew_1_1_5, dataRegroupBySew_0_1_5};
  wire [31:0]       dataInMem_lo_656;
  assign dataInMem_lo_656 = _GEN_720;
  wire [31:0]       dataInMem_lo_721;
  assign dataInMem_lo_721 = _GEN_720;
  wire [31:0]       dataInMem_lo_lo_148;
  assign dataInMem_lo_lo_148 = _GEN_720;
  wire [31:0]       _GEN_721 = {dataRegroupBySew_3_1_5, dataRegroupBySew_2_1_5};
  wire [31:0]       dataInMem_hi_848;
  assign dataInMem_hi_848 = _GEN_721;
  wire [31:0]       dataInMem_lo_hi_532;
  assign dataInMem_lo_hi_532 = _GEN_721;
  wire [31:0]       _GEN_722 = {dataRegroupBySew_1_1_6, dataRegroupBySew_0_1_6};
  wire [31:0]       dataInMem_lo_657;
  assign dataInMem_lo_657 = _GEN_722;
  wire [31:0]       dataInMem_lo_722;
  assign dataInMem_lo_722 = _GEN_722;
  wire [31:0]       dataInMem_lo_lo_149;
  assign dataInMem_lo_lo_149 = _GEN_722;
  wire [31:0]       _GEN_723 = {dataRegroupBySew_3_1_6, dataRegroupBySew_2_1_6};
  wire [31:0]       dataInMem_hi_849;
  assign dataInMem_hi_849 = _GEN_723;
  wire [31:0]       dataInMem_lo_hi_533;
  assign dataInMem_lo_hi_533 = _GEN_723;
  wire [31:0]       _GEN_724 = {dataRegroupBySew_1_1_7, dataRegroupBySew_0_1_7};
  wire [31:0]       dataInMem_lo_658;
  assign dataInMem_lo_658 = _GEN_724;
  wire [31:0]       dataInMem_lo_723;
  assign dataInMem_lo_723 = _GEN_724;
  wire [31:0]       dataInMem_lo_lo_150;
  assign dataInMem_lo_lo_150 = _GEN_724;
  wire [31:0]       _GEN_725 = {dataRegroupBySew_3_1_7, dataRegroupBySew_2_1_7};
  wire [31:0]       dataInMem_hi_850;
  assign dataInMem_hi_850 = _GEN_725;
  wire [31:0]       dataInMem_lo_hi_534;
  assign dataInMem_lo_hi_534 = _GEN_725;
  wire [31:0]       _GEN_726 = {dataRegroupBySew_1_1_8, dataRegroupBySew_0_1_8};
  wire [31:0]       dataInMem_lo_659;
  assign dataInMem_lo_659 = _GEN_726;
  wire [31:0]       dataInMem_lo_724;
  assign dataInMem_lo_724 = _GEN_726;
  wire [31:0]       dataInMem_lo_lo_151;
  assign dataInMem_lo_lo_151 = _GEN_726;
  wire [31:0]       _GEN_727 = {dataRegroupBySew_3_1_8, dataRegroupBySew_2_1_8};
  wire [31:0]       dataInMem_hi_851;
  assign dataInMem_hi_851 = _GEN_727;
  wire [31:0]       dataInMem_lo_hi_535;
  assign dataInMem_lo_hi_535 = _GEN_727;
  wire [31:0]       _GEN_728 = {dataRegroupBySew_1_1_9, dataRegroupBySew_0_1_9};
  wire [31:0]       dataInMem_lo_660;
  assign dataInMem_lo_660 = _GEN_728;
  wire [31:0]       dataInMem_lo_725;
  assign dataInMem_lo_725 = _GEN_728;
  wire [31:0]       dataInMem_lo_lo_152;
  assign dataInMem_lo_lo_152 = _GEN_728;
  wire [31:0]       _GEN_729 = {dataRegroupBySew_3_1_9, dataRegroupBySew_2_1_9};
  wire [31:0]       dataInMem_hi_852;
  assign dataInMem_hi_852 = _GEN_729;
  wire [31:0]       dataInMem_lo_hi_536;
  assign dataInMem_lo_hi_536 = _GEN_729;
  wire [31:0]       _GEN_730 = {dataRegroupBySew_1_1_10, dataRegroupBySew_0_1_10};
  wire [31:0]       dataInMem_lo_661;
  assign dataInMem_lo_661 = _GEN_730;
  wire [31:0]       dataInMem_lo_726;
  assign dataInMem_lo_726 = _GEN_730;
  wire [31:0]       dataInMem_lo_lo_153;
  assign dataInMem_lo_lo_153 = _GEN_730;
  wire [31:0]       _GEN_731 = {dataRegroupBySew_3_1_10, dataRegroupBySew_2_1_10};
  wire [31:0]       dataInMem_hi_853;
  assign dataInMem_hi_853 = _GEN_731;
  wire [31:0]       dataInMem_lo_hi_537;
  assign dataInMem_lo_hi_537 = _GEN_731;
  wire [31:0]       _GEN_732 = {dataRegroupBySew_1_1_11, dataRegroupBySew_0_1_11};
  wire [31:0]       dataInMem_lo_662;
  assign dataInMem_lo_662 = _GEN_732;
  wire [31:0]       dataInMem_lo_727;
  assign dataInMem_lo_727 = _GEN_732;
  wire [31:0]       dataInMem_lo_lo_154;
  assign dataInMem_lo_lo_154 = _GEN_732;
  wire [31:0]       _GEN_733 = {dataRegroupBySew_3_1_11, dataRegroupBySew_2_1_11};
  wire [31:0]       dataInMem_hi_854;
  assign dataInMem_hi_854 = _GEN_733;
  wire [31:0]       dataInMem_lo_hi_538;
  assign dataInMem_lo_hi_538 = _GEN_733;
  wire [31:0]       _GEN_734 = {dataRegroupBySew_1_1_12, dataRegroupBySew_0_1_12};
  wire [31:0]       dataInMem_lo_663;
  assign dataInMem_lo_663 = _GEN_734;
  wire [31:0]       dataInMem_lo_728;
  assign dataInMem_lo_728 = _GEN_734;
  wire [31:0]       dataInMem_lo_lo_155;
  assign dataInMem_lo_lo_155 = _GEN_734;
  wire [31:0]       _GEN_735 = {dataRegroupBySew_3_1_12, dataRegroupBySew_2_1_12};
  wire [31:0]       dataInMem_hi_855;
  assign dataInMem_hi_855 = _GEN_735;
  wire [31:0]       dataInMem_lo_hi_539;
  assign dataInMem_lo_hi_539 = _GEN_735;
  wire [31:0]       _GEN_736 = {dataRegroupBySew_1_1_13, dataRegroupBySew_0_1_13};
  wire [31:0]       dataInMem_lo_664;
  assign dataInMem_lo_664 = _GEN_736;
  wire [31:0]       dataInMem_lo_729;
  assign dataInMem_lo_729 = _GEN_736;
  wire [31:0]       dataInMem_lo_lo_156;
  assign dataInMem_lo_lo_156 = _GEN_736;
  wire [31:0]       _GEN_737 = {dataRegroupBySew_3_1_13, dataRegroupBySew_2_1_13};
  wire [31:0]       dataInMem_hi_856;
  assign dataInMem_hi_856 = _GEN_737;
  wire [31:0]       dataInMem_lo_hi_540;
  assign dataInMem_lo_hi_540 = _GEN_737;
  wire [31:0]       _GEN_738 = {dataRegroupBySew_1_1_14, dataRegroupBySew_0_1_14};
  wire [31:0]       dataInMem_lo_665;
  assign dataInMem_lo_665 = _GEN_738;
  wire [31:0]       dataInMem_lo_730;
  assign dataInMem_lo_730 = _GEN_738;
  wire [31:0]       dataInMem_lo_lo_157;
  assign dataInMem_lo_lo_157 = _GEN_738;
  wire [31:0]       _GEN_739 = {dataRegroupBySew_3_1_14, dataRegroupBySew_2_1_14};
  wire [31:0]       dataInMem_hi_857;
  assign dataInMem_hi_857 = _GEN_739;
  wire [31:0]       dataInMem_lo_hi_541;
  assign dataInMem_lo_hi_541 = _GEN_739;
  wire [31:0]       _GEN_740 = {dataRegroupBySew_1_1_15, dataRegroupBySew_0_1_15};
  wire [31:0]       dataInMem_lo_666;
  assign dataInMem_lo_666 = _GEN_740;
  wire [31:0]       dataInMem_lo_731;
  assign dataInMem_lo_731 = _GEN_740;
  wire [31:0]       dataInMem_lo_lo_158;
  assign dataInMem_lo_lo_158 = _GEN_740;
  wire [31:0]       _GEN_741 = {dataRegroupBySew_3_1_15, dataRegroupBySew_2_1_15};
  wire [31:0]       dataInMem_hi_858;
  assign dataInMem_hi_858 = _GEN_741;
  wire [31:0]       dataInMem_lo_hi_542;
  assign dataInMem_lo_hi_542 = _GEN_741;
  wire [31:0]       _GEN_742 = {dataRegroupBySew_1_1_16, dataRegroupBySew_0_1_16};
  wire [31:0]       dataInMem_lo_667;
  assign dataInMem_lo_667 = _GEN_742;
  wire [31:0]       dataInMem_lo_732;
  assign dataInMem_lo_732 = _GEN_742;
  wire [31:0]       dataInMem_lo_lo_159;
  assign dataInMem_lo_lo_159 = _GEN_742;
  wire [31:0]       _GEN_743 = {dataRegroupBySew_3_1_16, dataRegroupBySew_2_1_16};
  wire [31:0]       dataInMem_hi_859;
  assign dataInMem_hi_859 = _GEN_743;
  wire [31:0]       dataInMem_lo_hi_543;
  assign dataInMem_lo_hi_543 = _GEN_743;
  wire [31:0]       _GEN_744 = {dataRegroupBySew_1_1_17, dataRegroupBySew_0_1_17};
  wire [31:0]       dataInMem_lo_668;
  assign dataInMem_lo_668 = _GEN_744;
  wire [31:0]       dataInMem_lo_733;
  assign dataInMem_lo_733 = _GEN_744;
  wire [31:0]       dataInMem_lo_lo_160;
  assign dataInMem_lo_lo_160 = _GEN_744;
  wire [31:0]       _GEN_745 = {dataRegroupBySew_3_1_17, dataRegroupBySew_2_1_17};
  wire [31:0]       dataInMem_hi_860;
  assign dataInMem_hi_860 = _GEN_745;
  wire [31:0]       dataInMem_lo_hi_544;
  assign dataInMem_lo_hi_544 = _GEN_745;
  wire [31:0]       _GEN_746 = {dataRegroupBySew_1_1_18, dataRegroupBySew_0_1_18};
  wire [31:0]       dataInMem_lo_669;
  assign dataInMem_lo_669 = _GEN_746;
  wire [31:0]       dataInMem_lo_734;
  assign dataInMem_lo_734 = _GEN_746;
  wire [31:0]       dataInMem_lo_lo_161;
  assign dataInMem_lo_lo_161 = _GEN_746;
  wire [31:0]       _GEN_747 = {dataRegroupBySew_3_1_18, dataRegroupBySew_2_1_18};
  wire [31:0]       dataInMem_hi_861;
  assign dataInMem_hi_861 = _GEN_747;
  wire [31:0]       dataInMem_lo_hi_545;
  assign dataInMem_lo_hi_545 = _GEN_747;
  wire [31:0]       _GEN_748 = {dataRegroupBySew_1_1_19, dataRegroupBySew_0_1_19};
  wire [31:0]       dataInMem_lo_670;
  assign dataInMem_lo_670 = _GEN_748;
  wire [31:0]       dataInMem_lo_735;
  assign dataInMem_lo_735 = _GEN_748;
  wire [31:0]       dataInMem_lo_lo_162;
  assign dataInMem_lo_lo_162 = _GEN_748;
  wire [31:0]       _GEN_749 = {dataRegroupBySew_3_1_19, dataRegroupBySew_2_1_19};
  wire [31:0]       dataInMem_hi_862;
  assign dataInMem_hi_862 = _GEN_749;
  wire [31:0]       dataInMem_lo_hi_546;
  assign dataInMem_lo_hi_546 = _GEN_749;
  wire [31:0]       _GEN_750 = {dataRegroupBySew_1_1_20, dataRegroupBySew_0_1_20};
  wire [31:0]       dataInMem_lo_671;
  assign dataInMem_lo_671 = _GEN_750;
  wire [31:0]       dataInMem_lo_736;
  assign dataInMem_lo_736 = _GEN_750;
  wire [31:0]       dataInMem_lo_lo_163;
  assign dataInMem_lo_lo_163 = _GEN_750;
  wire [31:0]       _GEN_751 = {dataRegroupBySew_3_1_20, dataRegroupBySew_2_1_20};
  wire [31:0]       dataInMem_hi_863;
  assign dataInMem_hi_863 = _GEN_751;
  wire [31:0]       dataInMem_lo_hi_547;
  assign dataInMem_lo_hi_547 = _GEN_751;
  wire [31:0]       _GEN_752 = {dataRegroupBySew_1_1_21, dataRegroupBySew_0_1_21};
  wire [31:0]       dataInMem_lo_672;
  assign dataInMem_lo_672 = _GEN_752;
  wire [31:0]       dataInMem_lo_737;
  assign dataInMem_lo_737 = _GEN_752;
  wire [31:0]       dataInMem_lo_lo_164;
  assign dataInMem_lo_lo_164 = _GEN_752;
  wire [31:0]       _GEN_753 = {dataRegroupBySew_3_1_21, dataRegroupBySew_2_1_21};
  wire [31:0]       dataInMem_hi_864;
  assign dataInMem_hi_864 = _GEN_753;
  wire [31:0]       dataInMem_lo_hi_548;
  assign dataInMem_lo_hi_548 = _GEN_753;
  wire [31:0]       _GEN_754 = {dataRegroupBySew_1_1_22, dataRegroupBySew_0_1_22};
  wire [31:0]       dataInMem_lo_673;
  assign dataInMem_lo_673 = _GEN_754;
  wire [31:0]       dataInMem_lo_738;
  assign dataInMem_lo_738 = _GEN_754;
  wire [31:0]       dataInMem_lo_lo_165;
  assign dataInMem_lo_lo_165 = _GEN_754;
  wire [31:0]       _GEN_755 = {dataRegroupBySew_3_1_22, dataRegroupBySew_2_1_22};
  wire [31:0]       dataInMem_hi_865;
  assign dataInMem_hi_865 = _GEN_755;
  wire [31:0]       dataInMem_lo_hi_549;
  assign dataInMem_lo_hi_549 = _GEN_755;
  wire [31:0]       _GEN_756 = {dataRegroupBySew_1_1_23, dataRegroupBySew_0_1_23};
  wire [31:0]       dataInMem_lo_674;
  assign dataInMem_lo_674 = _GEN_756;
  wire [31:0]       dataInMem_lo_739;
  assign dataInMem_lo_739 = _GEN_756;
  wire [31:0]       dataInMem_lo_lo_166;
  assign dataInMem_lo_lo_166 = _GEN_756;
  wire [31:0]       _GEN_757 = {dataRegroupBySew_3_1_23, dataRegroupBySew_2_1_23};
  wire [31:0]       dataInMem_hi_866;
  assign dataInMem_hi_866 = _GEN_757;
  wire [31:0]       dataInMem_lo_hi_550;
  assign dataInMem_lo_hi_550 = _GEN_757;
  wire [31:0]       _GEN_758 = {dataRegroupBySew_1_1_24, dataRegroupBySew_0_1_24};
  wire [31:0]       dataInMem_lo_675;
  assign dataInMem_lo_675 = _GEN_758;
  wire [31:0]       dataInMem_lo_740;
  assign dataInMem_lo_740 = _GEN_758;
  wire [31:0]       dataInMem_lo_lo_167;
  assign dataInMem_lo_lo_167 = _GEN_758;
  wire [31:0]       _GEN_759 = {dataRegroupBySew_3_1_24, dataRegroupBySew_2_1_24};
  wire [31:0]       dataInMem_hi_867;
  assign dataInMem_hi_867 = _GEN_759;
  wire [31:0]       dataInMem_lo_hi_551;
  assign dataInMem_lo_hi_551 = _GEN_759;
  wire [31:0]       _GEN_760 = {dataRegroupBySew_1_1_25, dataRegroupBySew_0_1_25};
  wire [31:0]       dataInMem_lo_676;
  assign dataInMem_lo_676 = _GEN_760;
  wire [31:0]       dataInMem_lo_741;
  assign dataInMem_lo_741 = _GEN_760;
  wire [31:0]       dataInMem_lo_lo_168;
  assign dataInMem_lo_lo_168 = _GEN_760;
  wire [31:0]       _GEN_761 = {dataRegroupBySew_3_1_25, dataRegroupBySew_2_1_25};
  wire [31:0]       dataInMem_hi_868;
  assign dataInMem_hi_868 = _GEN_761;
  wire [31:0]       dataInMem_lo_hi_552;
  assign dataInMem_lo_hi_552 = _GEN_761;
  wire [31:0]       _GEN_762 = {dataRegroupBySew_1_1_26, dataRegroupBySew_0_1_26};
  wire [31:0]       dataInMem_lo_677;
  assign dataInMem_lo_677 = _GEN_762;
  wire [31:0]       dataInMem_lo_742;
  assign dataInMem_lo_742 = _GEN_762;
  wire [31:0]       dataInMem_lo_lo_169;
  assign dataInMem_lo_lo_169 = _GEN_762;
  wire [31:0]       _GEN_763 = {dataRegroupBySew_3_1_26, dataRegroupBySew_2_1_26};
  wire [31:0]       dataInMem_hi_869;
  assign dataInMem_hi_869 = _GEN_763;
  wire [31:0]       dataInMem_lo_hi_553;
  assign dataInMem_lo_hi_553 = _GEN_763;
  wire [31:0]       _GEN_764 = {dataRegroupBySew_1_1_27, dataRegroupBySew_0_1_27};
  wire [31:0]       dataInMem_lo_678;
  assign dataInMem_lo_678 = _GEN_764;
  wire [31:0]       dataInMem_lo_743;
  assign dataInMem_lo_743 = _GEN_764;
  wire [31:0]       dataInMem_lo_lo_170;
  assign dataInMem_lo_lo_170 = _GEN_764;
  wire [31:0]       _GEN_765 = {dataRegroupBySew_3_1_27, dataRegroupBySew_2_1_27};
  wire [31:0]       dataInMem_hi_870;
  assign dataInMem_hi_870 = _GEN_765;
  wire [31:0]       dataInMem_lo_hi_554;
  assign dataInMem_lo_hi_554 = _GEN_765;
  wire [31:0]       _GEN_766 = {dataRegroupBySew_1_1_28, dataRegroupBySew_0_1_28};
  wire [31:0]       dataInMem_lo_679;
  assign dataInMem_lo_679 = _GEN_766;
  wire [31:0]       dataInMem_lo_744;
  assign dataInMem_lo_744 = _GEN_766;
  wire [31:0]       dataInMem_lo_lo_171;
  assign dataInMem_lo_lo_171 = _GEN_766;
  wire [31:0]       _GEN_767 = {dataRegroupBySew_3_1_28, dataRegroupBySew_2_1_28};
  wire [31:0]       dataInMem_hi_871;
  assign dataInMem_hi_871 = _GEN_767;
  wire [31:0]       dataInMem_lo_hi_555;
  assign dataInMem_lo_hi_555 = _GEN_767;
  wire [31:0]       _GEN_768 = {dataRegroupBySew_1_1_29, dataRegroupBySew_0_1_29};
  wire [31:0]       dataInMem_lo_680;
  assign dataInMem_lo_680 = _GEN_768;
  wire [31:0]       dataInMem_lo_745;
  assign dataInMem_lo_745 = _GEN_768;
  wire [31:0]       dataInMem_lo_lo_172;
  assign dataInMem_lo_lo_172 = _GEN_768;
  wire [31:0]       _GEN_769 = {dataRegroupBySew_3_1_29, dataRegroupBySew_2_1_29};
  wire [31:0]       dataInMem_hi_872;
  assign dataInMem_hi_872 = _GEN_769;
  wire [31:0]       dataInMem_lo_hi_556;
  assign dataInMem_lo_hi_556 = _GEN_769;
  wire [31:0]       _GEN_770 = {dataRegroupBySew_1_1_30, dataRegroupBySew_0_1_30};
  wire [31:0]       dataInMem_lo_681;
  assign dataInMem_lo_681 = _GEN_770;
  wire [31:0]       dataInMem_lo_746;
  assign dataInMem_lo_746 = _GEN_770;
  wire [31:0]       dataInMem_lo_lo_173;
  assign dataInMem_lo_lo_173 = _GEN_770;
  wire [31:0]       _GEN_771 = {dataRegroupBySew_3_1_30, dataRegroupBySew_2_1_30};
  wire [31:0]       dataInMem_hi_873;
  assign dataInMem_hi_873 = _GEN_771;
  wire [31:0]       dataInMem_lo_hi_557;
  assign dataInMem_lo_hi_557 = _GEN_771;
  wire [31:0]       _GEN_772 = {dataRegroupBySew_1_1_31, dataRegroupBySew_0_1_31};
  wire [31:0]       dataInMem_lo_682;
  assign dataInMem_lo_682 = _GEN_772;
  wire [31:0]       dataInMem_lo_747;
  assign dataInMem_lo_747 = _GEN_772;
  wire [31:0]       dataInMem_lo_lo_174;
  assign dataInMem_lo_lo_174 = _GEN_772;
  wire [31:0]       _GEN_773 = {dataRegroupBySew_3_1_31, dataRegroupBySew_2_1_31};
  wire [31:0]       dataInMem_hi_874;
  assign dataInMem_hi_874 = _GEN_773;
  wire [31:0]       dataInMem_lo_hi_558;
  assign dataInMem_lo_hi_558 = _GEN_773;
  wire [31:0]       _GEN_774 = {dataRegroupBySew_1_1_32, dataRegroupBySew_0_1_32};
  wire [31:0]       dataInMem_lo_683;
  assign dataInMem_lo_683 = _GEN_774;
  wire [31:0]       dataInMem_lo_748;
  assign dataInMem_lo_748 = _GEN_774;
  wire [31:0]       dataInMem_lo_lo_175;
  assign dataInMem_lo_lo_175 = _GEN_774;
  wire [31:0]       _GEN_775 = {dataRegroupBySew_3_1_32, dataRegroupBySew_2_1_32};
  wire [31:0]       dataInMem_hi_875;
  assign dataInMem_hi_875 = _GEN_775;
  wire [31:0]       dataInMem_lo_hi_559;
  assign dataInMem_lo_hi_559 = _GEN_775;
  wire [31:0]       _GEN_776 = {dataRegroupBySew_1_1_33, dataRegroupBySew_0_1_33};
  wire [31:0]       dataInMem_lo_684;
  assign dataInMem_lo_684 = _GEN_776;
  wire [31:0]       dataInMem_lo_749;
  assign dataInMem_lo_749 = _GEN_776;
  wire [31:0]       dataInMem_lo_lo_176;
  assign dataInMem_lo_lo_176 = _GEN_776;
  wire [31:0]       _GEN_777 = {dataRegroupBySew_3_1_33, dataRegroupBySew_2_1_33};
  wire [31:0]       dataInMem_hi_876;
  assign dataInMem_hi_876 = _GEN_777;
  wire [31:0]       dataInMem_lo_hi_560;
  assign dataInMem_lo_hi_560 = _GEN_777;
  wire [31:0]       _GEN_778 = {dataRegroupBySew_1_1_34, dataRegroupBySew_0_1_34};
  wire [31:0]       dataInMem_lo_685;
  assign dataInMem_lo_685 = _GEN_778;
  wire [31:0]       dataInMem_lo_750;
  assign dataInMem_lo_750 = _GEN_778;
  wire [31:0]       dataInMem_lo_lo_177;
  assign dataInMem_lo_lo_177 = _GEN_778;
  wire [31:0]       _GEN_779 = {dataRegroupBySew_3_1_34, dataRegroupBySew_2_1_34};
  wire [31:0]       dataInMem_hi_877;
  assign dataInMem_hi_877 = _GEN_779;
  wire [31:0]       dataInMem_lo_hi_561;
  assign dataInMem_lo_hi_561 = _GEN_779;
  wire [31:0]       _GEN_780 = {dataRegroupBySew_1_1_35, dataRegroupBySew_0_1_35};
  wire [31:0]       dataInMem_lo_686;
  assign dataInMem_lo_686 = _GEN_780;
  wire [31:0]       dataInMem_lo_751;
  assign dataInMem_lo_751 = _GEN_780;
  wire [31:0]       dataInMem_lo_lo_178;
  assign dataInMem_lo_lo_178 = _GEN_780;
  wire [31:0]       _GEN_781 = {dataRegroupBySew_3_1_35, dataRegroupBySew_2_1_35};
  wire [31:0]       dataInMem_hi_878;
  assign dataInMem_hi_878 = _GEN_781;
  wire [31:0]       dataInMem_lo_hi_562;
  assign dataInMem_lo_hi_562 = _GEN_781;
  wire [31:0]       _GEN_782 = {dataRegroupBySew_1_1_36, dataRegroupBySew_0_1_36};
  wire [31:0]       dataInMem_lo_687;
  assign dataInMem_lo_687 = _GEN_782;
  wire [31:0]       dataInMem_lo_752;
  assign dataInMem_lo_752 = _GEN_782;
  wire [31:0]       dataInMem_lo_lo_179;
  assign dataInMem_lo_lo_179 = _GEN_782;
  wire [31:0]       _GEN_783 = {dataRegroupBySew_3_1_36, dataRegroupBySew_2_1_36};
  wire [31:0]       dataInMem_hi_879;
  assign dataInMem_hi_879 = _GEN_783;
  wire [31:0]       dataInMem_lo_hi_563;
  assign dataInMem_lo_hi_563 = _GEN_783;
  wire [31:0]       _GEN_784 = {dataRegroupBySew_1_1_37, dataRegroupBySew_0_1_37};
  wire [31:0]       dataInMem_lo_688;
  assign dataInMem_lo_688 = _GEN_784;
  wire [31:0]       dataInMem_lo_753;
  assign dataInMem_lo_753 = _GEN_784;
  wire [31:0]       dataInMem_lo_lo_180;
  assign dataInMem_lo_lo_180 = _GEN_784;
  wire [31:0]       _GEN_785 = {dataRegroupBySew_3_1_37, dataRegroupBySew_2_1_37};
  wire [31:0]       dataInMem_hi_880;
  assign dataInMem_hi_880 = _GEN_785;
  wire [31:0]       dataInMem_lo_hi_564;
  assign dataInMem_lo_hi_564 = _GEN_785;
  wire [31:0]       _GEN_786 = {dataRegroupBySew_1_1_38, dataRegroupBySew_0_1_38};
  wire [31:0]       dataInMem_lo_689;
  assign dataInMem_lo_689 = _GEN_786;
  wire [31:0]       dataInMem_lo_754;
  assign dataInMem_lo_754 = _GEN_786;
  wire [31:0]       dataInMem_lo_lo_181;
  assign dataInMem_lo_lo_181 = _GEN_786;
  wire [31:0]       _GEN_787 = {dataRegroupBySew_3_1_38, dataRegroupBySew_2_1_38};
  wire [31:0]       dataInMem_hi_881;
  assign dataInMem_hi_881 = _GEN_787;
  wire [31:0]       dataInMem_lo_hi_565;
  assign dataInMem_lo_hi_565 = _GEN_787;
  wire [31:0]       _GEN_788 = {dataRegroupBySew_1_1_39, dataRegroupBySew_0_1_39};
  wire [31:0]       dataInMem_lo_690;
  assign dataInMem_lo_690 = _GEN_788;
  wire [31:0]       dataInMem_lo_755;
  assign dataInMem_lo_755 = _GEN_788;
  wire [31:0]       dataInMem_lo_lo_182;
  assign dataInMem_lo_lo_182 = _GEN_788;
  wire [31:0]       _GEN_789 = {dataRegroupBySew_3_1_39, dataRegroupBySew_2_1_39};
  wire [31:0]       dataInMem_hi_882;
  assign dataInMem_hi_882 = _GEN_789;
  wire [31:0]       dataInMem_lo_hi_566;
  assign dataInMem_lo_hi_566 = _GEN_789;
  wire [31:0]       _GEN_790 = {dataRegroupBySew_1_1_40, dataRegroupBySew_0_1_40};
  wire [31:0]       dataInMem_lo_691;
  assign dataInMem_lo_691 = _GEN_790;
  wire [31:0]       dataInMem_lo_756;
  assign dataInMem_lo_756 = _GEN_790;
  wire [31:0]       dataInMem_lo_lo_183;
  assign dataInMem_lo_lo_183 = _GEN_790;
  wire [31:0]       _GEN_791 = {dataRegroupBySew_3_1_40, dataRegroupBySew_2_1_40};
  wire [31:0]       dataInMem_hi_883;
  assign dataInMem_hi_883 = _GEN_791;
  wire [31:0]       dataInMem_lo_hi_567;
  assign dataInMem_lo_hi_567 = _GEN_791;
  wire [31:0]       _GEN_792 = {dataRegroupBySew_1_1_41, dataRegroupBySew_0_1_41};
  wire [31:0]       dataInMem_lo_692;
  assign dataInMem_lo_692 = _GEN_792;
  wire [31:0]       dataInMem_lo_757;
  assign dataInMem_lo_757 = _GEN_792;
  wire [31:0]       dataInMem_lo_lo_184;
  assign dataInMem_lo_lo_184 = _GEN_792;
  wire [31:0]       _GEN_793 = {dataRegroupBySew_3_1_41, dataRegroupBySew_2_1_41};
  wire [31:0]       dataInMem_hi_884;
  assign dataInMem_hi_884 = _GEN_793;
  wire [31:0]       dataInMem_lo_hi_568;
  assign dataInMem_lo_hi_568 = _GEN_793;
  wire [31:0]       _GEN_794 = {dataRegroupBySew_1_1_42, dataRegroupBySew_0_1_42};
  wire [31:0]       dataInMem_lo_693;
  assign dataInMem_lo_693 = _GEN_794;
  wire [31:0]       dataInMem_lo_758;
  assign dataInMem_lo_758 = _GEN_794;
  wire [31:0]       dataInMem_lo_lo_185;
  assign dataInMem_lo_lo_185 = _GEN_794;
  wire [31:0]       _GEN_795 = {dataRegroupBySew_3_1_42, dataRegroupBySew_2_1_42};
  wire [31:0]       dataInMem_hi_885;
  assign dataInMem_hi_885 = _GEN_795;
  wire [31:0]       dataInMem_lo_hi_569;
  assign dataInMem_lo_hi_569 = _GEN_795;
  wire [31:0]       _GEN_796 = {dataRegroupBySew_1_1_43, dataRegroupBySew_0_1_43};
  wire [31:0]       dataInMem_lo_694;
  assign dataInMem_lo_694 = _GEN_796;
  wire [31:0]       dataInMem_lo_759;
  assign dataInMem_lo_759 = _GEN_796;
  wire [31:0]       dataInMem_lo_lo_186;
  assign dataInMem_lo_lo_186 = _GEN_796;
  wire [31:0]       _GEN_797 = {dataRegroupBySew_3_1_43, dataRegroupBySew_2_1_43};
  wire [31:0]       dataInMem_hi_886;
  assign dataInMem_hi_886 = _GEN_797;
  wire [31:0]       dataInMem_lo_hi_570;
  assign dataInMem_lo_hi_570 = _GEN_797;
  wire [31:0]       _GEN_798 = {dataRegroupBySew_1_1_44, dataRegroupBySew_0_1_44};
  wire [31:0]       dataInMem_lo_695;
  assign dataInMem_lo_695 = _GEN_798;
  wire [31:0]       dataInMem_lo_760;
  assign dataInMem_lo_760 = _GEN_798;
  wire [31:0]       dataInMem_lo_lo_187;
  assign dataInMem_lo_lo_187 = _GEN_798;
  wire [31:0]       _GEN_799 = {dataRegroupBySew_3_1_44, dataRegroupBySew_2_1_44};
  wire [31:0]       dataInMem_hi_887;
  assign dataInMem_hi_887 = _GEN_799;
  wire [31:0]       dataInMem_lo_hi_571;
  assign dataInMem_lo_hi_571 = _GEN_799;
  wire [31:0]       _GEN_800 = {dataRegroupBySew_1_1_45, dataRegroupBySew_0_1_45};
  wire [31:0]       dataInMem_lo_696;
  assign dataInMem_lo_696 = _GEN_800;
  wire [31:0]       dataInMem_lo_761;
  assign dataInMem_lo_761 = _GEN_800;
  wire [31:0]       dataInMem_lo_lo_188;
  assign dataInMem_lo_lo_188 = _GEN_800;
  wire [31:0]       _GEN_801 = {dataRegroupBySew_3_1_45, dataRegroupBySew_2_1_45};
  wire [31:0]       dataInMem_hi_888;
  assign dataInMem_hi_888 = _GEN_801;
  wire [31:0]       dataInMem_lo_hi_572;
  assign dataInMem_lo_hi_572 = _GEN_801;
  wire [31:0]       _GEN_802 = {dataRegroupBySew_1_1_46, dataRegroupBySew_0_1_46};
  wire [31:0]       dataInMem_lo_697;
  assign dataInMem_lo_697 = _GEN_802;
  wire [31:0]       dataInMem_lo_762;
  assign dataInMem_lo_762 = _GEN_802;
  wire [31:0]       dataInMem_lo_lo_189;
  assign dataInMem_lo_lo_189 = _GEN_802;
  wire [31:0]       _GEN_803 = {dataRegroupBySew_3_1_46, dataRegroupBySew_2_1_46};
  wire [31:0]       dataInMem_hi_889;
  assign dataInMem_hi_889 = _GEN_803;
  wire [31:0]       dataInMem_lo_hi_573;
  assign dataInMem_lo_hi_573 = _GEN_803;
  wire [31:0]       _GEN_804 = {dataRegroupBySew_1_1_47, dataRegroupBySew_0_1_47};
  wire [31:0]       dataInMem_lo_698;
  assign dataInMem_lo_698 = _GEN_804;
  wire [31:0]       dataInMem_lo_763;
  assign dataInMem_lo_763 = _GEN_804;
  wire [31:0]       dataInMem_lo_lo_190;
  assign dataInMem_lo_lo_190 = _GEN_804;
  wire [31:0]       _GEN_805 = {dataRegroupBySew_3_1_47, dataRegroupBySew_2_1_47};
  wire [31:0]       dataInMem_hi_890;
  assign dataInMem_hi_890 = _GEN_805;
  wire [31:0]       dataInMem_lo_hi_574;
  assign dataInMem_lo_hi_574 = _GEN_805;
  wire [31:0]       _GEN_806 = {dataRegroupBySew_1_1_48, dataRegroupBySew_0_1_48};
  wire [31:0]       dataInMem_lo_699;
  assign dataInMem_lo_699 = _GEN_806;
  wire [31:0]       dataInMem_lo_764;
  assign dataInMem_lo_764 = _GEN_806;
  wire [31:0]       dataInMem_lo_lo_191;
  assign dataInMem_lo_lo_191 = _GEN_806;
  wire [31:0]       _GEN_807 = {dataRegroupBySew_3_1_48, dataRegroupBySew_2_1_48};
  wire [31:0]       dataInMem_hi_891;
  assign dataInMem_hi_891 = _GEN_807;
  wire [31:0]       dataInMem_lo_hi_575;
  assign dataInMem_lo_hi_575 = _GEN_807;
  wire [31:0]       _GEN_808 = {dataRegroupBySew_1_1_49, dataRegroupBySew_0_1_49};
  wire [31:0]       dataInMem_lo_700;
  assign dataInMem_lo_700 = _GEN_808;
  wire [31:0]       dataInMem_lo_765;
  assign dataInMem_lo_765 = _GEN_808;
  wire [31:0]       dataInMem_lo_lo_192;
  assign dataInMem_lo_lo_192 = _GEN_808;
  wire [31:0]       _GEN_809 = {dataRegroupBySew_3_1_49, dataRegroupBySew_2_1_49};
  wire [31:0]       dataInMem_hi_892;
  assign dataInMem_hi_892 = _GEN_809;
  wire [31:0]       dataInMem_lo_hi_576;
  assign dataInMem_lo_hi_576 = _GEN_809;
  wire [31:0]       _GEN_810 = {dataRegroupBySew_1_1_50, dataRegroupBySew_0_1_50};
  wire [31:0]       dataInMem_lo_701;
  assign dataInMem_lo_701 = _GEN_810;
  wire [31:0]       dataInMem_lo_766;
  assign dataInMem_lo_766 = _GEN_810;
  wire [31:0]       dataInMem_lo_lo_193;
  assign dataInMem_lo_lo_193 = _GEN_810;
  wire [31:0]       _GEN_811 = {dataRegroupBySew_3_1_50, dataRegroupBySew_2_1_50};
  wire [31:0]       dataInMem_hi_893;
  assign dataInMem_hi_893 = _GEN_811;
  wire [31:0]       dataInMem_lo_hi_577;
  assign dataInMem_lo_hi_577 = _GEN_811;
  wire [31:0]       _GEN_812 = {dataRegroupBySew_1_1_51, dataRegroupBySew_0_1_51};
  wire [31:0]       dataInMem_lo_702;
  assign dataInMem_lo_702 = _GEN_812;
  wire [31:0]       dataInMem_lo_767;
  assign dataInMem_lo_767 = _GEN_812;
  wire [31:0]       dataInMem_lo_lo_194;
  assign dataInMem_lo_lo_194 = _GEN_812;
  wire [31:0]       _GEN_813 = {dataRegroupBySew_3_1_51, dataRegroupBySew_2_1_51};
  wire [31:0]       dataInMem_hi_894;
  assign dataInMem_hi_894 = _GEN_813;
  wire [31:0]       dataInMem_lo_hi_578;
  assign dataInMem_lo_hi_578 = _GEN_813;
  wire [31:0]       _GEN_814 = {dataRegroupBySew_1_1_52, dataRegroupBySew_0_1_52};
  wire [31:0]       dataInMem_lo_703;
  assign dataInMem_lo_703 = _GEN_814;
  wire [31:0]       dataInMem_lo_768;
  assign dataInMem_lo_768 = _GEN_814;
  wire [31:0]       dataInMem_lo_lo_195;
  assign dataInMem_lo_lo_195 = _GEN_814;
  wire [31:0]       _GEN_815 = {dataRegroupBySew_3_1_52, dataRegroupBySew_2_1_52};
  wire [31:0]       dataInMem_hi_895;
  assign dataInMem_hi_895 = _GEN_815;
  wire [31:0]       dataInMem_lo_hi_579;
  assign dataInMem_lo_hi_579 = _GEN_815;
  wire [31:0]       _GEN_816 = {dataRegroupBySew_1_1_53, dataRegroupBySew_0_1_53};
  wire [31:0]       dataInMem_lo_704;
  assign dataInMem_lo_704 = _GEN_816;
  wire [31:0]       dataInMem_lo_769;
  assign dataInMem_lo_769 = _GEN_816;
  wire [31:0]       dataInMem_lo_lo_196;
  assign dataInMem_lo_lo_196 = _GEN_816;
  wire [31:0]       _GEN_817 = {dataRegroupBySew_3_1_53, dataRegroupBySew_2_1_53};
  wire [31:0]       dataInMem_hi_896;
  assign dataInMem_hi_896 = _GEN_817;
  wire [31:0]       dataInMem_lo_hi_580;
  assign dataInMem_lo_hi_580 = _GEN_817;
  wire [31:0]       _GEN_818 = {dataRegroupBySew_1_1_54, dataRegroupBySew_0_1_54};
  wire [31:0]       dataInMem_lo_705;
  assign dataInMem_lo_705 = _GEN_818;
  wire [31:0]       dataInMem_lo_770;
  assign dataInMem_lo_770 = _GEN_818;
  wire [31:0]       dataInMem_lo_lo_197;
  assign dataInMem_lo_lo_197 = _GEN_818;
  wire [31:0]       _GEN_819 = {dataRegroupBySew_3_1_54, dataRegroupBySew_2_1_54};
  wire [31:0]       dataInMem_hi_897;
  assign dataInMem_hi_897 = _GEN_819;
  wire [31:0]       dataInMem_lo_hi_581;
  assign dataInMem_lo_hi_581 = _GEN_819;
  wire [31:0]       _GEN_820 = {dataRegroupBySew_1_1_55, dataRegroupBySew_0_1_55};
  wire [31:0]       dataInMem_lo_706;
  assign dataInMem_lo_706 = _GEN_820;
  wire [31:0]       dataInMem_lo_771;
  assign dataInMem_lo_771 = _GEN_820;
  wire [31:0]       dataInMem_lo_lo_198;
  assign dataInMem_lo_lo_198 = _GEN_820;
  wire [31:0]       _GEN_821 = {dataRegroupBySew_3_1_55, dataRegroupBySew_2_1_55};
  wire [31:0]       dataInMem_hi_898;
  assign dataInMem_hi_898 = _GEN_821;
  wire [31:0]       dataInMem_lo_hi_582;
  assign dataInMem_lo_hi_582 = _GEN_821;
  wire [31:0]       _GEN_822 = {dataRegroupBySew_1_1_56, dataRegroupBySew_0_1_56};
  wire [31:0]       dataInMem_lo_707;
  assign dataInMem_lo_707 = _GEN_822;
  wire [31:0]       dataInMem_lo_772;
  assign dataInMem_lo_772 = _GEN_822;
  wire [31:0]       dataInMem_lo_lo_199;
  assign dataInMem_lo_lo_199 = _GEN_822;
  wire [31:0]       _GEN_823 = {dataRegroupBySew_3_1_56, dataRegroupBySew_2_1_56};
  wire [31:0]       dataInMem_hi_899;
  assign dataInMem_hi_899 = _GEN_823;
  wire [31:0]       dataInMem_lo_hi_583;
  assign dataInMem_lo_hi_583 = _GEN_823;
  wire [31:0]       _GEN_824 = {dataRegroupBySew_1_1_57, dataRegroupBySew_0_1_57};
  wire [31:0]       dataInMem_lo_708;
  assign dataInMem_lo_708 = _GEN_824;
  wire [31:0]       dataInMem_lo_773;
  assign dataInMem_lo_773 = _GEN_824;
  wire [31:0]       dataInMem_lo_lo_200;
  assign dataInMem_lo_lo_200 = _GEN_824;
  wire [31:0]       _GEN_825 = {dataRegroupBySew_3_1_57, dataRegroupBySew_2_1_57};
  wire [31:0]       dataInMem_hi_900;
  assign dataInMem_hi_900 = _GEN_825;
  wire [31:0]       dataInMem_lo_hi_584;
  assign dataInMem_lo_hi_584 = _GEN_825;
  wire [31:0]       _GEN_826 = {dataRegroupBySew_1_1_58, dataRegroupBySew_0_1_58};
  wire [31:0]       dataInMem_lo_709;
  assign dataInMem_lo_709 = _GEN_826;
  wire [31:0]       dataInMem_lo_774;
  assign dataInMem_lo_774 = _GEN_826;
  wire [31:0]       dataInMem_lo_lo_201;
  assign dataInMem_lo_lo_201 = _GEN_826;
  wire [31:0]       _GEN_827 = {dataRegroupBySew_3_1_58, dataRegroupBySew_2_1_58};
  wire [31:0]       dataInMem_hi_901;
  assign dataInMem_hi_901 = _GEN_827;
  wire [31:0]       dataInMem_lo_hi_585;
  assign dataInMem_lo_hi_585 = _GEN_827;
  wire [31:0]       _GEN_828 = {dataRegroupBySew_1_1_59, dataRegroupBySew_0_1_59};
  wire [31:0]       dataInMem_lo_710;
  assign dataInMem_lo_710 = _GEN_828;
  wire [31:0]       dataInMem_lo_775;
  assign dataInMem_lo_775 = _GEN_828;
  wire [31:0]       dataInMem_lo_lo_202;
  assign dataInMem_lo_lo_202 = _GEN_828;
  wire [31:0]       _GEN_829 = {dataRegroupBySew_3_1_59, dataRegroupBySew_2_1_59};
  wire [31:0]       dataInMem_hi_902;
  assign dataInMem_hi_902 = _GEN_829;
  wire [31:0]       dataInMem_lo_hi_586;
  assign dataInMem_lo_hi_586 = _GEN_829;
  wire [31:0]       _GEN_830 = {dataRegroupBySew_1_1_60, dataRegroupBySew_0_1_60};
  wire [31:0]       dataInMem_lo_711;
  assign dataInMem_lo_711 = _GEN_830;
  wire [31:0]       dataInMem_lo_776;
  assign dataInMem_lo_776 = _GEN_830;
  wire [31:0]       dataInMem_lo_lo_203;
  assign dataInMem_lo_lo_203 = _GEN_830;
  wire [31:0]       _GEN_831 = {dataRegroupBySew_3_1_60, dataRegroupBySew_2_1_60};
  wire [31:0]       dataInMem_hi_903;
  assign dataInMem_hi_903 = _GEN_831;
  wire [31:0]       dataInMem_lo_hi_587;
  assign dataInMem_lo_hi_587 = _GEN_831;
  wire [31:0]       _GEN_832 = {dataRegroupBySew_1_1_61, dataRegroupBySew_0_1_61};
  wire [31:0]       dataInMem_lo_712;
  assign dataInMem_lo_712 = _GEN_832;
  wire [31:0]       dataInMem_lo_777;
  assign dataInMem_lo_777 = _GEN_832;
  wire [31:0]       dataInMem_lo_lo_204;
  assign dataInMem_lo_lo_204 = _GEN_832;
  wire [31:0]       _GEN_833 = {dataRegroupBySew_3_1_61, dataRegroupBySew_2_1_61};
  wire [31:0]       dataInMem_hi_904;
  assign dataInMem_hi_904 = _GEN_833;
  wire [31:0]       dataInMem_lo_hi_588;
  assign dataInMem_lo_hi_588 = _GEN_833;
  wire [31:0]       _GEN_834 = {dataRegroupBySew_1_1_62, dataRegroupBySew_0_1_62};
  wire [31:0]       dataInMem_lo_713;
  assign dataInMem_lo_713 = _GEN_834;
  wire [31:0]       dataInMem_lo_778;
  assign dataInMem_lo_778 = _GEN_834;
  wire [31:0]       dataInMem_lo_lo_205;
  assign dataInMem_lo_lo_205 = _GEN_834;
  wire [31:0]       _GEN_835 = {dataRegroupBySew_3_1_62, dataRegroupBySew_2_1_62};
  wire [31:0]       dataInMem_hi_905;
  assign dataInMem_hi_905 = _GEN_835;
  wire [31:0]       dataInMem_lo_hi_589;
  assign dataInMem_lo_hi_589 = _GEN_835;
  wire [31:0]       _GEN_836 = {dataRegroupBySew_1_1_63, dataRegroupBySew_0_1_63};
  wire [31:0]       dataInMem_lo_714;
  assign dataInMem_lo_714 = _GEN_836;
  wire [31:0]       dataInMem_lo_779;
  assign dataInMem_lo_779 = _GEN_836;
  wire [31:0]       dataInMem_lo_lo_206;
  assign dataInMem_lo_lo_206 = _GEN_836;
  wire [31:0]       _GEN_837 = {dataRegroupBySew_3_1_63, dataRegroupBySew_2_1_63};
  wire [31:0]       dataInMem_hi_906;
  assign dataInMem_hi_906 = _GEN_837;
  wire [31:0]       dataInMem_lo_hi_590;
  assign dataInMem_lo_hi_590 = _GEN_837;
  wire [127:0]      dataInMem_lo_lo_lo_lo_lo_11 = {dataInMem_hi_844, dataInMem_lo_652, dataInMem_hi_843, dataInMem_lo_651};
  wire [127:0]      dataInMem_lo_lo_lo_lo_hi_11 = {dataInMem_hi_846, dataInMem_lo_654, dataInMem_hi_845, dataInMem_lo_653};
  wire [255:0]      dataInMem_lo_lo_lo_lo_11 = {dataInMem_lo_lo_lo_lo_hi_11, dataInMem_lo_lo_lo_lo_lo_11};
  wire [127:0]      dataInMem_lo_lo_lo_hi_lo_11 = {dataInMem_hi_848, dataInMem_lo_656, dataInMem_hi_847, dataInMem_lo_655};
  wire [127:0]      dataInMem_lo_lo_lo_hi_hi_11 = {dataInMem_hi_850, dataInMem_lo_658, dataInMem_hi_849, dataInMem_lo_657};
  wire [255:0]      dataInMem_lo_lo_lo_hi_11 = {dataInMem_lo_lo_lo_hi_hi_11, dataInMem_lo_lo_lo_hi_lo_11};
  wire [511:0]      dataInMem_lo_lo_lo_11 = {dataInMem_lo_lo_lo_hi_11, dataInMem_lo_lo_lo_lo_11};
  wire [127:0]      dataInMem_lo_lo_hi_lo_lo_11 = {dataInMem_hi_852, dataInMem_lo_660, dataInMem_hi_851, dataInMem_lo_659};
  wire [127:0]      dataInMem_lo_lo_hi_lo_hi_11 = {dataInMem_hi_854, dataInMem_lo_662, dataInMem_hi_853, dataInMem_lo_661};
  wire [255:0]      dataInMem_lo_lo_hi_lo_11 = {dataInMem_lo_lo_hi_lo_hi_11, dataInMem_lo_lo_hi_lo_lo_11};
  wire [127:0]      dataInMem_lo_lo_hi_hi_lo_11 = {dataInMem_hi_856, dataInMem_lo_664, dataInMem_hi_855, dataInMem_lo_663};
  wire [127:0]      dataInMem_lo_lo_hi_hi_hi_11 = {dataInMem_hi_858, dataInMem_lo_666, dataInMem_hi_857, dataInMem_lo_665};
  wire [255:0]      dataInMem_lo_lo_hi_hi_11 = {dataInMem_lo_lo_hi_hi_hi_11, dataInMem_lo_lo_hi_hi_lo_11};
  wire [511:0]      dataInMem_lo_lo_hi_11 = {dataInMem_lo_lo_hi_hi_11, dataInMem_lo_lo_hi_lo_11};
  wire [1023:0]     dataInMem_lo_lo_139 = {dataInMem_lo_lo_hi_11, dataInMem_lo_lo_lo_11};
  wire [127:0]      dataInMem_lo_hi_lo_lo_lo_11 = {dataInMem_hi_860, dataInMem_lo_668, dataInMem_hi_859, dataInMem_lo_667};
  wire [127:0]      dataInMem_lo_hi_lo_lo_hi_11 = {dataInMem_hi_862, dataInMem_lo_670, dataInMem_hi_861, dataInMem_lo_669};
  wire [255:0]      dataInMem_lo_hi_lo_lo_11 = {dataInMem_lo_hi_lo_lo_hi_11, dataInMem_lo_hi_lo_lo_lo_11};
  wire [127:0]      dataInMem_lo_hi_lo_hi_lo_11 = {dataInMem_hi_864, dataInMem_lo_672, dataInMem_hi_863, dataInMem_lo_671};
  wire [127:0]      dataInMem_lo_hi_lo_hi_hi_11 = {dataInMem_hi_866, dataInMem_lo_674, dataInMem_hi_865, dataInMem_lo_673};
  wire [255:0]      dataInMem_lo_hi_lo_hi_11 = {dataInMem_lo_hi_lo_hi_hi_11, dataInMem_lo_hi_lo_hi_lo_11};
  wire [511:0]      dataInMem_lo_hi_lo_11 = {dataInMem_lo_hi_lo_hi_11, dataInMem_lo_hi_lo_lo_11};
  wire [127:0]      dataInMem_lo_hi_hi_lo_lo_11 = {dataInMem_hi_868, dataInMem_lo_676, dataInMem_hi_867, dataInMem_lo_675};
  wire [127:0]      dataInMem_lo_hi_hi_lo_hi_11 = {dataInMem_hi_870, dataInMem_lo_678, dataInMem_hi_869, dataInMem_lo_677};
  wire [255:0]      dataInMem_lo_hi_hi_lo_11 = {dataInMem_lo_hi_hi_lo_hi_11, dataInMem_lo_hi_hi_lo_lo_11};
  wire [127:0]      dataInMem_lo_hi_hi_hi_lo_11 = {dataInMem_hi_872, dataInMem_lo_680, dataInMem_hi_871, dataInMem_lo_679};
  wire [127:0]      dataInMem_lo_hi_hi_hi_hi_11 = {dataInMem_hi_874, dataInMem_lo_682, dataInMem_hi_873, dataInMem_lo_681};
  wire [255:0]      dataInMem_lo_hi_hi_hi_11 = {dataInMem_lo_hi_hi_hi_hi_11, dataInMem_lo_hi_hi_hi_lo_11};
  wire [511:0]      dataInMem_lo_hi_hi_11 = {dataInMem_lo_hi_hi_hi_11, dataInMem_lo_hi_hi_lo_11};
  wire [1023:0]     dataInMem_lo_hi_395 = {dataInMem_lo_hi_hi_11, dataInMem_lo_hi_lo_11};
  wire [2047:0]     dataInMem_lo_715 = {dataInMem_lo_hi_395, dataInMem_lo_lo_139};
  wire [127:0]      dataInMem_hi_lo_lo_lo_lo_11 = {dataInMem_hi_876, dataInMem_lo_684, dataInMem_hi_875, dataInMem_lo_683};
  wire [127:0]      dataInMem_hi_lo_lo_lo_hi_11 = {dataInMem_hi_878, dataInMem_lo_686, dataInMem_hi_877, dataInMem_lo_685};
  wire [255:0]      dataInMem_hi_lo_lo_lo_11 = {dataInMem_hi_lo_lo_lo_hi_11, dataInMem_hi_lo_lo_lo_lo_11};
  wire [127:0]      dataInMem_hi_lo_lo_hi_lo_11 = {dataInMem_hi_880, dataInMem_lo_688, dataInMem_hi_879, dataInMem_lo_687};
  wire [127:0]      dataInMem_hi_lo_lo_hi_hi_11 = {dataInMem_hi_882, dataInMem_lo_690, dataInMem_hi_881, dataInMem_lo_689};
  wire [255:0]      dataInMem_hi_lo_lo_hi_11 = {dataInMem_hi_lo_lo_hi_hi_11, dataInMem_hi_lo_lo_hi_lo_11};
  wire [511:0]      dataInMem_hi_lo_lo_11 = {dataInMem_hi_lo_lo_hi_11, dataInMem_hi_lo_lo_lo_11};
  wire [127:0]      dataInMem_hi_lo_hi_lo_lo_11 = {dataInMem_hi_884, dataInMem_lo_692, dataInMem_hi_883, dataInMem_lo_691};
  wire [127:0]      dataInMem_hi_lo_hi_lo_hi_11 = {dataInMem_hi_886, dataInMem_lo_694, dataInMem_hi_885, dataInMem_lo_693};
  wire [255:0]      dataInMem_hi_lo_hi_lo_11 = {dataInMem_hi_lo_hi_lo_hi_11, dataInMem_hi_lo_hi_lo_lo_11};
  wire [127:0]      dataInMem_hi_lo_hi_hi_lo_11 = {dataInMem_hi_888, dataInMem_lo_696, dataInMem_hi_887, dataInMem_lo_695};
  wire [127:0]      dataInMem_hi_lo_hi_hi_hi_11 = {dataInMem_hi_890, dataInMem_lo_698, dataInMem_hi_889, dataInMem_lo_697};
  wire [255:0]      dataInMem_hi_lo_hi_hi_11 = {dataInMem_hi_lo_hi_hi_hi_11, dataInMem_hi_lo_hi_hi_lo_11};
  wire [511:0]      dataInMem_hi_lo_hi_11 = {dataInMem_hi_lo_hi_hi_11, dataInMem_hi_lo_hi_lo_11};
  wire [1023:0]     dataInMem_hi_lo_267 = {dataInMem_hi_lo_hi_11, dataInMem_hi_lo_lo_11};
  wire [127:0]      dataInMem_hi_hi_lo_lo_lo_11 = {dataInMem_hi_892, dataInMem_lo_700, dataInMem_hi_891, dataInMem_lo_699};
  wire [127:0]      dataInMem_hi_hi_lo_lo_hi_11 = {dataInMem_hi_894, dataInMem_lo_702, dataInMem_hi_893, dataInMem_lo_701};
  wire [255:0]      dataInMem_hi_hi_lo_lo_11 = {dataInMem_hi_hi_lo_lo_hi_11, dataInMem_hi_hi_lo_lo_lo_11};
  wire [127:0]      dataInMem_hi_hi_lo_hi_lo_11 = {dataInMem_hi_896, dataInMem_lo_704, dataInMem_hi_895, dataInMem_lo_703};
  wire [127:0]      dataInMem_hi_hi_lo_hi_hi_11 = {dataInMem_hi_898, dataInMem_lo_706, dataInMem_hi_897, dataInMem_lo_705};
  wire [255:0]      dataInMem_hi_hi_lo_hi_11 = {dataInMem_hi_hi_lo_hi_hi_11, dataInMem_hi_hi_lo_hi_lo_11};
  wire [511:0]      dataInMem_hi_hi_lo_11 = {dataInMem_hi_hi_lo_hi_11, dataInMem_hi_hi_lo_lo_11};
  wire [127:0]      dataInMem_hi_hi_hi_lo_lo_11 = {dataInMem_hi_900, dataInMem_lo_708, dataInMem_hi_899, dataInMem_lo_707};
  wire [127:0]      dataInMem_hi_hi_hi_lo_hi_11 = {dataInMem_hi_902, dataInMem_lo_710, dataInMem_hi_901, dataInMem_lo_709};
  wire [255:0]      dataInMem_hi_hi_hi_lo_11 = {dataInMem_hi_hi_hi_lo_hi_11, dataInMem_hi_hi_hi_lo_lo_11};
  wire [127:0]      dataInMem_hi_hi_hi_hi_lo_11 = {dataInMem_hi_904, dataInMem_lo_712, dataInMem_hi_903, dataInMem_lo_711};
  wire [127:0]      dataInMem_hi_hi_hi_hi_hi_11 = {dataInMem_hi_906, dataInMem_lo_714, dataInMem_hi_905, dataInMem_lo_713};
  wire [255:0]      dataInMem_hi_hi_hi_hi_11 = {dataInMem_hi_hi_hi_hi_hi_11, dataInMem_hi_hi_hi_hi_lo_11};
  wire [511:0]      dataInMem_hi_hi_hi_11 = {dataInMem_hi_hi_hi_hi_11, dataInMem_hi_hi_hi_lo_11};
  wire [1023:0]     dataInMem_hi_hi_523 = {dataInMem_hi_hi_hi_11, dataInMem_hi_hi_lo_11};
  wire [2047:0]     dataInMem_hi_907 = {dataInMem_hi_hi_523, dataInMem_hi_lo_267};
  wire [4095:0]     dataInMem_11 = {dataInMem_hi_907, dataInMem_lo_715};
  wire [1023:0]     regroupCacheLine_11_0 = dataInMem_11[1023:0];
  wire [1023:0]     regroupCacheLine_11_1 = dataInMem_11[2047:1024];
  wire [1023:0]     regroupCacheLine_11_2 = dataInMem_11[3071:2048];
  wire [1023:0]     regroupCacheLine_11_3 = dataInMem_11[4095:3072];
  wire [1023:0]     res_88 = regroupCacheLine_11_0;
  wire [1023:0]     res_89 = regroupCacheLine_11_1;
  wire [1023:0]     res_90 = regroupCacheLine_11_2;
  wire [1023:0]     res_91 = regroupCacheLine_11_3;
  wire [2047:0]     lo_lo_11 = {res_89, res_88};
  wire [2047:0]     lo_hi_11 = {res_91, res_90};
  wire [4095:0]     lo_11 = {lo_hi_11, lo_lo_11};
  wire [8191:0]     regroupLoadData_1_3 = {4096'h0, lo_11};
  wire [31:0]       _GEN_838 = {dataRegroupBySew_4_1_0, dataRegroupBySew_3_1_0};
  wire [31:0]       dataInMem_hi_hi_524;
  assign dataInMem_hi_hi_524 = _GEN_838;
  wire [31:0]       dataInMem_hi_lo_270;
  assign dataInMem_hi_lo_270 = _GEN_838;
  wire [47:0]       dataInMem_hi_908 = {dataInMem_hi_hi_524, dataRegroupBySew_2_1_0};
  wire [31:0]       _GEN_839 = {dataRegroupBySew_4_1_1, dataRegroupBySew_3_1_1};
  wire [31:0]       dataInMem_hi_hi_525;
  assign dataInMem_hi_hi_525 = _GEN_839;
  wire [31:0]       dataInMem_hi_lo_271;
  assign dataInMem_hi_lo_271 = _GEN_839;
  wire [47:0]       dataInMem_hi_909 = {dataInMem_hi_hi_525, dataRegroupBySew_2_1_1};
  wire [31:0]       _GEN_840 = {dataRegroupBySew_4_1_2, dataRegroupBySew_3_1_2};
  wire [31:0]       dataInMem_hi_hi_526;
  assign dataInMem_hi_hi_526 = _GEN_840;
  wire [31:0]       dataInMem_hi_lo_272;
  assign dataInMem_hi_lo_272 = _GEN_840;
  wire [47:0]       dataInMem_hi_910 = {dataInMem_hi_hi_526, dataRegroupBySew_2_1_2};
  wire [31:0]       _GEN_841 = {dataRegroupBySew_4_1_3, dataRegroupBySew_3_1_3};
  wire [31:0]       dataInMem_hi_hi_527;
  assign dataInMem_hi_hi_527 = _GEN_841;
  wire [31:0]       dataInMem_hi_lo_273;
  assign dataInMem_hi_lo_273 = _GEN_841;
  wire [47:0]       dataInMem_hi_911 = {dataInMem_hi_hi_527, dataRegroupBySew_2_1_3};
  wire [31:0]       _GEN_842 = {dataRegroupBySew_4_1_4, dataRegroupBySew_3_1_4};
  wire [31:0]       dataInMem_hi_hi_528;
  assign dataInMem_hi_hi_528 = _GEN_842;
  wire [31:0]       dataInMem_hi_lo_274;
  assign dataInMem_hi_lo_274 = _GEN_842;
  wire [47:0]       dataInMem_hi_912 = {dataInMem_hi_hi_528, dataRegroupBySew_2_1_4};
  wire [31:0]       _GEN_843 = {dataRegroupBySew_4_1_5, dataRegroupBySew_3_1_5};
  wire [31:0]       dataInMem_hi_hi_529;
  assign dataInMem_hi_hi_529 = _GEN_843;
  wire [31:0]       dataInMem_hi_lo_275;
  assign dataInMem_hi_lo_275 = _GEN_843;
  wire [47:0]       dataInMem_hi_913 = {dataInMem_hi_hi_529, dataRegroupBySew_2_1_5};
  wire [31:0]       _GEN_844 = {dataRegroupBySew_4_1_6, dataRegroupBySew_3_1_6};
  wire [31:0]       dataInMem_hi_hi_530;
  assign dataInMem_hi_hi_530 = _GEN_844;
  wire [31:0]       dataInMem_hi_lo_276;
  assign dataInMem_hi_lo_276 = _GEN_844;
  wire [47:0]       dataInMem_hi_914 = {dataInMem_hi_hi_530, dataRegroupBySew_2_1_6};
  wire [31:0]       _GEN_845 = {dataRegroupBySew_4_1_7, dataRegroupBySew_3_1_7};
  wire [31:0]       dataInMem_hi_hi_531;
  assign dataInMem_hi_hi_531 = _GEN_845;
  wire [31:0]       dataInMem_hi_lo_277;
  assign dataInMem_hi_lo_277 = _GEN_845;
  wire [47:0]       dataInMem_hi_915 = {dataInMem_hi_hi_531, dataRegroupBySew_2_1_7};
  wire [31:0]       _GEN_846 = {dataRegroupBySew_4_1_8, dataRegroupBySew_3_1_8};
  wire [31:0]       dataInMem_hi_hi_532;
  assign dataInMem_hi_hi_532 = _GEN_846;
  wire [31:0]       dataInMem_hi_lo_278;
  assign dataInMem_hi_lo_278 = _GEN_846;
  wire [47:0]       dataInMem_hi_916 = {dataInMem_hi_hi_532, dataRegroupBySew_2_1_8};
  wire [31:0]       _GEN_847 = {dataRegroupBySew_4_1_9, dataRegroupBySew_3_1_9};
  wire [31:0]       dataInMem_hi_hi_533;
  assign dataInMem_hi_hi_533 = _GEN_847;
  wire [31:0]       dataInMem_hi_lo_279;
  assign dataInMem_hi_lo_279 = _GEN_847;
  wire [47:0]       dataInMem_hi_917 = {dataInMem_hi_hi_533, dataRegroupBySew_2_1_9};
  wire [31:0]       _GEN_848 = {dataRegroupBySew_4_1_10, dataRegroupBySew_3_1_10};
  wire [31:0]       dataInMem_hi_hi_534;
  assign dataInMem_hi_hi_534 = _GEN_848;
  wire [31:0]       dataInMem_hi_lo_280;
  assign dataInMem_hi_lo_280 = _GEN_848;
  wire [47:0]       dataInMem_hi_918 = {dataInMem_hi_hi_534, dataRegroupBySew_2_1_10};
  wire [31:0]       _GEN_849 = {dataRegroupBySew_4_1_11, dataRegroupBySew_3_1_11};
  wire [31:0]       dataInMem_hi_hi_535;
  assign dataInMem_hi_hi_535 = _GEN_849;
  wire [31:0]       dataInMem_hi_lo_281;
  assign dataInMem_hi_lo_281 = _GEN_849;
  wire [47:0]       dataInMem_hi_919 = {dataInMem_hi_hi_535, dataRegroupBySew_2_1_11};
  wire [31:0]       _GEN_850 = {dataRegroupBySew_4_1_12, dataRegroupBySew_3_1_12};
  wire [31:0]       dataInMem_hi_hi_536;
  assign dataInMem_hi_hi_536 = _GEN_850;
  wire [31:0]       dataInMem_hi_lo_282;
  assign dataInMem_hi_lo_282 = _GEN_850;
  wire [47:0]       dataInMem_hi_920 = {dataInMem_hi_hi_536, dataRegroupBySew_2_1_12};
  wire [31:0]       _GEN_851 = {dataRegroupBySew_4_1_13, dataRegroupBySew_3_1_13};
  wire [31:0]       dataInMem_hi_hi_537;
  assign dataInMem_hi_hi_537 = _GEN_851;
  wire [31:0]       dataInMem_hi_lo_283;
  assign dataInMem_hi_lo_283 = _GEN_851;
  wire [47:0]       dataInMem_hi_921 = {dataInMem_hi_hi_537, dataRegroupBySew_2_1_13};
  wire [31:0]       _GEN_852 = {dataRegroupBySew_4_1_14, dataRegroupBySew_3_1_14};
  wire [31:0]       dataInMem_hi_hi_538;
  assign dataInMem_hi_hi_538 = _GEN_852;
  wire [31:0]       dataInMem_hi_lo_284;
  assign dataInMem_hi_lo_284 = _GEN_852;
  wire [47:0]       dataInMem_hi_922 = {dataInMem_hi_hi_538, dataRegroupBySew_2_1_14};
  wire [31:0]       _GEN_853 = {dataRegroupBySew_4_1_15, dataRegroupBySew_3_1_15};
  wire [31:0]       dataInMem_hi_hi_539;
  assign dataInMem_hi_hi_539 = _GEN_853;
  wire [31:0]       dataInMem_hi_lo_285;
  assign dataInMem_hi_lo_285 = _GEN_853;
  wire [47:0]       dataInMem_hi_923 = {dataInMem_hi_hi_539, dataRegroupBySew_2_1_15};
  wire [31:0]       _GEN_854 = {dataRegroupBySew_4_1_16, dataRegroupBySew_3_1_16};
  wire [31:0]       dataInMem_hi_hi_540;
  assign dataInMem_hi_hi_540 = _GEN_854;
  wire [31:0]       dataInMem_hi_lo_286;
  assign dataInMem_hi_lo_286 = _GEN_854;
  wire [47:0]       dataInMem_hi_924 = {dataInMem_hi_hi_540, dataRegroupBySew_2_1_16};
  wire [31:0]       _GEN_855 = {dataRegroupBySew_4_1_17, dataRegroupBySew_3_1_17};
  wire [31:0]       dataInMem_hi_hi_541;
  assign dataInMem_hi_hi_541 = _GEN_855;
  wire [31:0]       dataInMem_hi_lo_287;
  assign dataInMem_hi_lo_287 = _GEN_855;
  wire [47:0]       dataInMem_hi_925 = {dataInMem_hi_hi_541, dataRegroupBySew_2_1_17};
  wire [31:0]       _GEN_856 = {dataRegroupBySew_4_1_18, dataRegroupBySew_3_1_18};
  wire [31:0]       dataInMem_hi_hi_542;
  assign dataInMem_hi_hi_542 = _GEN_856;
  wire [31:0]       dataInMem_hi_lo_288;
  assign dataInMem_hi_lo_288 = _GEN_856;
  wire [47:0]       dataInMem_hi_926 = {dataInMem_hi_hi_542, dataRegroupBySew_2_1_18};
  wire [31:0]       _GEN_857 = {dataRegroupBySew_4_1_19, dataRegroupBySew_3_1_19};
  wire [31:0]       dataInMem_hi_hi_543;
  assign dataInMem_hi_hi_543 = _GEN_857;
  wire [31:0]       dataInMem_hi_lo_289;
  assign dataInMem_hi_lo_289 = _GEN_857;
  wire [47:0]       dataInMem_hi_927 = {dataInMem_hi_hi_543, dataRegroupBySew_2_1_19};
  wire [31:0]       _GEN_858 = {dataRegroupBySew_4_1_20, dataRegroupBySew_3_1_20};
  wire [31:0]       dataInMem_hi_hi_544;
  assign dataInMem_hi_hi_544 = _GEN_858;
  wire [31:0]       dataInMem_hi_lo_290;
  assign dataInMem_hi_lo_290 = _GEN_858;
  wire [47:0]       dataInMem_hi_928 = {dataInMem_hi_hi_544, dataRegroupBySew_2_1_20};
  wire [31:0]       _GEN_859 = {dataRegroupBySew_4_1_21, dataRegroupBySew_3_1_21};
  wire [31:0]       dataInMem_hi_hi_545;
  assign dataInMem_hi_hi_545 = _GEN_859;
  wire [31:0]       dataInMem_hi_lo_291;
  assign dataInMem_hi_lo_291 = _GEN_859;
  wire [47:0]       dataInMem_hi_929 = {dataInMem_hi_hi_545, dataRegroupBySew_2_1_21};
  wire [31:0]       _GEN_860 = {dataRegroupBySew_4_1_22, dataRegroupBySew_3_1_22};
  wire [31:0]       dataInMem_hi_hi_546;
  assign dataInMem_hi_hi_546 = _GEN_860;
  wire [31:0]       dataInMem_hi_lo_292;
  assign dataInMem_hi_lo_292 = _GEN_860;
  wire [47:0]       dataInMem_hi_930 = {dataInMem_hi_hi_546, dataRegroupBySew_2_1_22};
  wire [31:0]       _GEN_861 = {dataRegroupBySew_4_1_23, dataRegroupBySew_3_1_23};
  wire [31:0]       dataInMem_hi_hi_547;
  assign dataInMem_hi_hi_547 = _GEN_861;
  wire [31:0]       dataInMem_hi_lo_293;
  assign dataInMem_hi_lo_293 = _GEN_861;
  wire [47:0]       dataInMem_hi_931 = {dataInMem_hi_hi_547, dataRegroupBySew_2_1_23};
  wire [31:0]       _GEN_862 = {dataRegroupBySew_4_1_24, dataRegroupBySew_3_1_24};
  wire [31:0]       dataInMem_hi_hi_548;
  assign dataInMem_hi_hi_548 = _GEN_862;
  wire [31:0]       dataInMem_hi_lo_294;
  assign dataInMem_hi_lo_294 = _GEN_862;
  wire [47:0]       dataInMem_hi_932 = {dataInMem_hi_hi_548, dataRegroupBySew_2_1_24};
  wire [31:0]       _GEN_863 = {dataRegroupBySew_4_1_25, dataRegroupBySew_3_1_25};
  wire [31:0]       dataInMem_hi_hi_549;
  assign dataInMem_hi_hi_549 = _GEN_863;
  wire [31:0]       dataInMem_hi_lo_295;
  assign dataInMem_hi_lo_295 = _GEN_863;
  wire [47:0]       dataInMem_hi_933 = {dataInMem_hi_hi_549, dataRegroupBySew_2_1_25};
  wire [31:0]       _GEN_864 = {dataRegroupBySew_4_1_26, dataRegroupBySew_3_1_26};
  wire [31:0]       dataInMem_hi_hi_550;
  assign dataInMem_hi_hi_550 = _GEN_864;
  wire [31:0]       dataInMem_hi_lo_296;
  assign dataInMem_hi_lo_296 = _GEN_864;
  wire [47:0]       dataInMem_hi_934 = {dataInMem_hi_hi_550, dataRegroupBySew_2_1_26};
  wire [31:0]       _GEN_865 = {dataRegroupBySew_4_1_27, dataRegroupBySew_3_1_27};
  wire [31:0]       dataInMem_hi_hi_551;
  assign dataInMem_hi_hi_551 = _GEN_865;
  wire [31:0]       dataInMem_hi_lo_297;
  assign dataInMem_hi_lo_297 = _GEN_865;
  wire [47:0]       dataInMem_hi_935 = {dataInMem_hi_hi_551, dataRegroupBySew_2_1_27};
  wire [31:0]       _GEN_866 = {dataRegroupBySew_4_1_28, dataRegroupBySew_3_1_28};
  wire [31:0]       dataInMem_hi_hi_552;
  assign dataInMem_hi_hi_552 = _GEN_866;
  wire [31:0]       dataInMem_hi_lo_298;
  assign dataInMem_hi_lo_298 = _GEN_866;
  wire [47:0]       dataInMem_hi_936 = {dataInMem_hi_hi_552, dataRegroupBySew_2_1_28};
  wire [31:0]       _GEN_867 = {dataRegroupBySew_4_1_29, dataRegroupBySew_3_1_29};
  wire [31:0]       dataInMem_hi_hi_553;
  assign dataInMem_hi_hi_553 = _GEN_867;
  wire [31:0]       dataInMem_hi_lo_299;
  assign dataInMem_hi_lo_299 = _GEN_867;
  wire [47:0]       dataInMem_hi_937 = {dataInMem_hi_hi_553, dataRegroupBySew_2_1_29};
  wire [31:0]       _GEN_868 = {dataRegroupBySew_4_1_30, dataRegroupBySew_3_1_30};
  wire [31:0]       dataInMem_hi_hi_554;
  assign dataInMem_hi_hi_554 = _GEN_868;
  wire [31:0]       dataInMem_hi_lo_300;
  assign dataInMem_hi_lo_300 = _GEN_868;
  wire [47:0]       dataInMem_hi_938 = {dataInMem_hi_hi_554, dataRegroupBySew_2_1_30};
  wire [31:0]       _GEN_869 = {dataRegroupBySew_4_1_31, dataRegroupBySew_3_1_31};
  wire [31:0]       dataInMem_hi_hi_555;
  assign dataInMem_hi_hi_555 = _GEN_869;
  wire [31:0]       dataInMem_hi_lo_301;
  assign dataInMem_hi_lo_301 = _GEN_869;
  wire [47:0]       dataInMem_hi_939 = {dataInMem_hi_hi_555, dataRegroupBySew_2_1_31};
  wire [31:0]       _GEN_870 = {dataRegroupBySew_4_1_32, dataRegroupBySew_3_1_32};
  wire [31:0]       dataInMem_hi_hi_556;
  assign dataInMem_hi_hi_556 = _GEN_870;
  wire [31:0]       dataInMem_hi_lo_302;
  assign dataInMem_hi_lo_302 = _GEN_870;
  wire [47:0]       dataInMem_hi_940 = {dataInMem_hi_hi_556, dataRegroupBySew_2_1_32};
  wire [31:0]       _GEN_871 = {dataRegroupBySew_4_1_33, dataRegroupBySew_3_1_33};
  wire [31:0]       dataInMem_hi_hi_557;
  assign dataInMem_hi_hi_557 = _GEN_871;
  wire [31:0]       dataInMem_hi_lo_303;
  assign dataInMem_hi_lo_303 = _GEN_871;
  wire [47:0]       dataInMem_hi_941 = {dataInMem_hi_hi_557, dataRegroupBySew_2_1_33};
  wire [31:0]       _GEN_872 = {dataRegroupBySew_4_1_34, dataRegroupBySew_3_1_34};
  wire [31:0]       dataInMem_hi_hi_558;
  assign dataInMem_hi_hi_558 = _GEN_872;
  wire [31:0]       dataInMem_hi_lo_304;
  assign dataInMem_hi_lo_304 = _GEN_872;
  wire [47:0]       dataInMem_hi_942 = {dataInMem_hi_hi_558, dataRegroupBySew_2_1_34};
  wire [31:0]       _GEN_873 = {dataRegroupBySew_4_1_35, dataRegroupBySew_3_1_35};
  wire [31:0]       dataInMem_hi_hi_559;
  assign dataInMem_hi_hi_559 = _GEN_873;
  wire [31:0]       dataInMem_hi_lo_305;
  assign dataInMem_hi_lo_305 = _GEN_873;
  wire [47:0]       dataInMem_hi_943 = {dataInMem_hi_hi_559, dataRegroupBySew_2_1_35};
  wire [31:0]       _GEN_874 = {dataRegroupBySew_4_1_36, dataRegroupBySew_3_1_36};
  wire [31:0]       dataInMem_hi_hi_560;
  assign dataInMem_hi_hi_560 = _GEN_874;
  wire [31:0]       dataInMem_hi_lo_306;
  assign dataInMem_hi_lo_306 = _GEN_874;
  wire [47:0]       dataInMem_hi_944 = {dataInMem_hi_hi_560, dataRegroupBySew_2_1_36};
  wire [31:0]       _GEN_875 = {dataRegroupBySew_4_1_37, dataRegroupBySew_3_1_37};
  wire [31:0]       dataInMem_hi_hi_561;
  assign dataInMem_hi_hi_561 = _GEN_875;
  wire [31:0]       dataInMem_hi_lo_307;
  assign dataInMem_hi_lo_307 = _GEN_875;
  wire [47:0]       dataInMem_hi_945 = {dataInMem_hi_hi_561, dataRegroupBySew_2_1_37};
  wire [31:0]       _GEN_876 = {dataRegroupBySew_4_1_38, dataRegroupBySew_3_1_38};
  wire [31:0]       dataInMem_hi_hi_562;
  assign dataInMem_hi_hi_562 = _GEN_876;
  wire [31:0]       dataInMem_hi_lo_308;
  assign dataInMem_hi_lo_308 = _GEN_876;
  wire [47:0]       dataInMem_hi_946 = {dataInMem_hi_hi_562, dataRegroupBySew_2_1_38};
  wire [31:0]       _GEN_877 = {dataRegroupBySew_4_1_39, dataRegroupBySew_3_1_39};
  wire [31:0]       dataInMem_hi_hi_563;
  assign dataInMem_hi_hi_563 = _GEN_877;
  wire [31:0]       dataInMem_hi_lo_309;
  assign dataInMem_hi_lo_309 = _GEN_877;
  wire [47:0]       dataInMem_hi_947 = {dataInMem_hi_hi_563, dataRegroupBySew_2_1_39};
  wire [31:0]       _GEN_878 = {dataRegroupBySew_4_1_40, dataRegroupBySew_3_1_40};
  wire [31:0]       dataInMem_hi_hi_564;
  assign dataInMem_hi_hi_564 = _GEN_878;
  wire [31:0]       dataInMem_hi_lo_310;
  assign dataInMem_hi_lo_310 = _GEN_878;
  wire [47:0]       dataInMem_hi_948 = {dataInMem_hi_hi_564, dataRegroupBySew_2_1_40};
  wire [31:0]       _GEN_879 = {dataRegroupBySew_4_1_41, dataRegroupBySew_3_1_41};
  wire [31:0]       dataInMem_hi_hi_565;
  assign dataInMem_hi_hi_565 = _GEN_879;
  wire [31:0]       dataInMem_hi_lo_311;
  assign dataInMem_hi_lo_311 = _GEN_879;
  wire [47:0]       dataInMem_hi_949 = {dataInMem_hi_hi_565, dataRegroupBySew_2_1_41};
  wire [31:0]       _GEN_880 = {dataRegroupBySew_4_1_42, dataRegroupBySew_3_1_42};
  wire [31:0]       dataInMem_hi_hi_566;
  assign dataInMem_hi_hi_566 = _GEN_880;
  wire [31:0]       dataInMem_hi_lo_312;
  assign dataInMem_hi_lo_312 = _GEN_880;
  wire [47:0]       dataInMem_hi_950 = {dataInMem_hi_hi_566, dataRegroupBySew_2_1_42};
  wire [31:0]       _GEN_881 = {dataRegroupBySew_4_1_43, dataRegroupBySew_3_1_43};
  wire [31:0]       dataInMem_hi_hi_567;
  assign dataInMem_hi_hi_567 = _GEN_881;
  wire [31:0]       dataInMem_hi_lo_313;
  assign dataInMem_hi_lo_313 = _GEN_881;
  wire [47:0]       dataInMem_hi_951 = {dataInMem_hi_hi_567, dataRegroupBySew_2_1_43};
  wire [31:0]       _GEN_882 = {dataRegroupBySew_4_1_44, dataRegroupBySew_3_1_44};
  wire [31:0]       dataInMem_hi_hi_568;
  assign dataInMem_hi_hi_568 = _GEN_882;
  wire [31:0]       dataInMem_hi_lo_314;
  assign dataInMem_hi_lo_314 = _GEN_882;
  wire [47:0]       dataInMem_hi_952 = {dataInMem_hi_hi_568, dataRegroupBySew_2_1_44};
  wire [31:0]       _GEN_883 = {dataRegroupBySew_4_1_45, dataRegroupBySew_3_1_45};
  wire [31:0]       dataInMem_hi_hi_569;
  assign dataInMem_hi_hi_569 = _GEN_883;
  wire [31:0]       dataInMem_hi_lo_315;
  assign dataInMem_hi_lo_315 = _GEN_883;
  wire [47:0]       dataInMem_hi_953 = {dataInMem_hi_hi_569, dataRegroupBySew_2_1_45};
  wire [31:0]       _GEN_884 = {dataRegroupBySew_4_1_46, dataRegroupBySew_3_1_46};
  wire [31:0]       dataInMem_hi_hi_570;
  assign dataInMem_hi_hi_570 = _GEN_884;
  wire [31:0]       dataInMem_hi_lo_316;
  assign dataInMem_hi_lo_316 = _GEN_884;
  wire [47:0]       dataInMem_hi_954 = {dataInMem_hi_hi_570, dataRegroupBySew_2_1_46};
  wire [31:0]       _GEN_885 = {dataRegroupBySew_4_1_47, dataRegroupBySew_3_1_47};
  wire [31:0]       dataInMem_hi_hi_571;
  assign dataInMem_hi_hi_571 = _GEN_885;
  wire [31:0]       dataInMem_hi_lo_317;
  assign dataInMem_hi_lo_317 = _GEN_885;
  wire [47:0]       dataInMem_hi_955 = {dataInMem_hi_hi_571, dataRegroupBySew_2_1_47};
  wire [31:0]       _GEN_886 = {dataRegroupBySew_4_1_48, dataRegroupBySew_3_1_48};
  wire [31:0]       dataInMem_hi_hi_572;
  assign dataInMem_hi_hi_572 = _GEN_886;
  wire [31:0]       dataInMem_hi_lo_318;
  assign dataInMem_hi_lo_318 = _GEN_886;
  wire [47:0]       dataInMem_hi_956 = {dataInMem_hi_hi_572, dataRegroupBySew_2_1_48};
  wire [31:0]       _GEN_887 = {dataRegroupBySew_4_1_49, dataRegroupBySew_3_1_49};
  wire [31:0]       dataInMem_hi_hi_573;
  assign dataInMem_hi_hi_573 = _GEN_887;
  wire [31:0]       dataInMem_hi_lo_319;
  assign dataInMem_hi_lo_319 = _GEN_887;
  wire [47:0]       dataInMem_hi_957 = {dataInMem_hi_hi_573, dataRegroupBySew_2_1_49};
  wire [31:0]       _GEN_888 = {dataRegroupBySew_4_1_50, dataRegroupBySew_3_1_50};
  wire [31:0]       dataInMem_hi_hi_574;
  assign dataInMem_hi_hi_574 = _GEN_888;
  wire [31:0]       dataInMem_hi_lo_320;
  assign dataInMem_hi_lo_320 = _GEN_888;
  wire [47:0]       dataInMem_hi_958 = {dataInMem_hi_hi_574, dataRegroupBySew_2_1_50};
  wire [31:0]       _GEN_889 = {dataRegroupBySew_4_1_51, dataRegroupBySew_3_1_51};
  wire [31:0]       dataInMem_hi_hi_575;
  assign dataInMem_hi_hi_575 = _GEN_889;
  wire [31:0]       dataInMem_hi_lo_321;
  assign dataInMem_hi_lo_321 = _GEN_889;
  wire [47:0]       dataInMem_hi_959 = {dataInMem_hi_hi_575, dataRegroupBySew_2_1_51};
  wire [31:0]       _GEN_890 = {dataRegroupBySew_4_1_52, dataRegroupBySew_3_1_52};
  wire [31:0]       dataInMem_hi_hi_576;
  assign dataInMem_hi_hi_576 = _GEN_890;
  wire [31:0]       dataInMem_hi_lo_322;
  assign dataInMem_hi_lo_322 = _GEN_890;
  wire [47:0]       dataInMem_hi_960 = {dataInMem_hi_hi_576, dataRegroupBySew_2_1_52};
  wire [31:0]       _GEN_891 = {dataRegroupBySew_4_1_53, dataRegroupBySew_3_1_53};
  wire [31:0]       dataInMem_hi_hi_577;
  assign dataInMem_hi_hi_577 = _GEN_891;
  wire [31:0]       dataInMem_hi_lo_323;
  assign dataInMem_hi_lo_323 = _GEN_891;
  wire [47:0]       dataInMem_hi_961 = {dataInMem_hi_hi_577, dataRegroupBySew_2_1_53};
  wire [31:0]       _GEN_892 = {dataRegroupBySew_4_1_54, dataRegroupBySew_3_1_54};
  wire [31:0]       dataInMem_hi_hi_578;
  assign dataInMem_hi_hi_578 = _GEN_892;
  wire [31:0]       dataInMem_hi_lo_324;
  assign dataInMem_hi_lo_324 = _GEN_892;
  wire [47:0]       dataInMem_hi_962 = {dataInMem_hi_hi_578, dataRegroupBySew_2_1_54};
  wire [31:0]       _GEN_893 = {dataRegroupBySew_4_1_55, dataRegroupBySew_3_1_55};
  wire [31:0]       dataInMem_hi_hi_579;
  assign dataInMem_hi_hi_579 = _GEN_893;
  wire [31:0]       dataInMem_hi_lo_325;
  assign dataInMem_hi_lo_325 = _GEN_893;
  wire [47:0]       dataInMem_hi_963 = {dataInMem_hi_hi_579, dataRegroupBySew_2_1_55};
  wire [31:0]       _GEN_894 = {dataRegroupBySew_4_1_56, dataRegroupBySew_3_1_56};
  wire [31:0]       dataInMem_hi_hi_580;
  assign dataInMem_hi_hi_580 = _GEN_894;
  wire [31:0]       dataInMem_hi_lo_326;
  assign dataInMem_hi_lo_326 = _GEN_894;
  wire [47:0]       dataInMem_hi_964 = {dataInMem_hi_hi_580, dataRegroupBySew_2_1_56};
  wire [31:0]       _GEN_895 = {dataRegroupBySew_4_1_57, dataRegroupBySew_3_1_57};
  wire [31:0]       dataInMem_hi_hi_581;
  assign dataInMem_hi_hi_581 = _GEN_895;
  wire [31:0]       dataInMem_hi_lo_327;
  assign dataInMem_hi_lo_327 = _GEN_895;
  wire [47:0]       dataInMem_hi_965 = {dataInMem_hi_hi_581, dataRegroupBySew_2_1_57};
  wire [31:0]       _GEN_896 = {dataRegroupBySew_4_1_58, dataRegroupBySew_3_1_58};
  wire [31:0]       dataInMem_hi_hi_582;
  assign dataInMem_hi_hi_582 = _GEN_896;
  wire [31:0]       dataInMem_hi_lo_328;
  assign dataInMem_hi_lo_328 = _GEN_896;
  wire [47:0]       dataInMem_hi_966 = {dataInMem_hi_hi_582, dataRegroupBySew_2_1_58};
  wire [31:0]       _GEN_897 = {dataRegroupBySew_4_1_59, dataRegroupBySew_3_1_59};
  wire [31:0]       dataInMem_hi_hi_583;
  assign dataInMem_hi_hi_583 = _GEN_897;
  wire [31:0]       dataInMem_hi_lo_329;
  assign dataInMem_hi_lo_329 = _GEN_897;
  wire [47:0]       dataInMem_hi_967 = {dataInMem_hi_hi_583, dataRegroupBySew_2_1_59};
  wire [31:0]       _GEN_898 = {dataRegroupBySew_4_1_60, dataRegroupBySew_3_1_60};
  wire [31:0]       dataInMem_hi_hi_584;
  assign dataInMem_hi_hi_584 = _GEN_898;
  wire [31:0]       dataInMem_hi_lo_330;
  assign dataInMem_hi_lo_330 = _GEN_898;
  wire [47:0]       dataInMem_hi_968 = {dataInMem_hi_hi_584, dataRegroupBySew_2_1_60};
  wire [31:0]       _GEN_899 = {dataRegroupBySew_4_1_61, dataRegroupBySew_3_1_61};
  wire [31:0]       dataInMem_hi_hi_585;
  assign dataInMem_hi_hi_585 = _GEN_899;
  wire [31:0]       dataInMem_hi_lo_331;
  assign dataInMem_hi_lo_331 = _GEN_899;
  wire [47:0]       dataInMem_hi_969 = {dataInMem_hi_hi_585, dataRegroupBySew_2_1_61};
  wire [31:0]       _GEN_900 = {dataRegroupBySew_4_1_62, dataRegroupBySew_3_1_62};
  wire [31:0]       dataInMem_hi_hi_586;
  assign dataInMem_hi_hi_586 = _GEN_900;
  wire [31:0]       dataInMem_hi_lo_332;
  assign dataInMem_hi_lo_332 = _GEN_900;
  wire [47:0]       dataInMem_hi_970 = {dataInMem_hi_hi_586, dataRegroupBySew_2_1_62};
  wire [31:0]       _GEN_901 = {dataRegroupBySew_4_1_63, dataRegroupBySew_3_1_63};
  wire [31:0]       dataInMem_hi_hi_587;
  assign dataInMem_hi_hi_587 = _GEN_901;
  wire [31:0]       dataInMem_hi_lo_333;
  assign dataInMem_hi_lo_333 = _GEN_901;
  wire [47:0]       dataInMem_hi_971 = {dataInMem_hi_hi_587, dataRegroupBySew_2_1_63};
  wire [159:0]      dataInMem_lo_lo_lo_lo_lo_12 = {dataInMem_hi_909, dataInMem_lo_717, dataInMem_hi_908, dataInMem_lo_716};
  wire [159:0]      dataInMem_lo_lo_lo_lo_hi_12 = {dataInMem_hi_911, dataInMem_lo_719, dataInMem_hi_910, dataInMem_lo_718};
  wire [319:0]      dataInMem_lo_lo_lo_lo_12 = {dataInMem_lo_lo_lo_lo_hi_12, dataInMem_lo_lo_lo_lo_lo_12};
  wire [159:0]      dataInMem_lo_lo_lo_hi_lo_12 = {dataInMem_hi_913, dataInMem_lo_721, dataInMem_hi_912, dataInMem_lo_720};
  wire [159:0]      dataInMem_lo_lo_lo_hi_hi_12 = {dataInMem_hi_915, dataInMem_lo_723, dataInMem_hi_914, dataInMem_lo_722};
  wire [319:0]      dataInMem_lo_lo_lo_hi_12 = {dataInMem_lo_lo_lo_hi_hi_12, dataInMem_lo_lo_lo_hi_lo_12};
  wire [639:0]      dataInMem_lo_lo_lo_12 = {dataInMem_lo_lo_lo_hi_12, dataInMem_lo_lo_lo_lo_12};
  wire [159:0]      dataInMem_lo_lo_hi_lo_lo_12 = {dataInMem_hi_917, dataInMem_lo_725, dataInMem_hi_916, dataInMem_lo_724};
  wire [159:0]      dataInMem_lo_lo_hi_lo_hi_12 = {dataInMem_hi_919, dataInMem_lo_727, dataInMem_hi_918, dataInMem_lo_726};
  wire [319:0]      dataInMem_lo_lo_hi_lo_12 = {dataInMem_lo_lo_hi_lo_hi_12, dataInMem_lo_lo_hi_lo_lo_12};
  wire [159:0]      dataInMem_lo_lo_hi_hi_lo_12 = {dataInMem_hi_921, dataInMem_lo_729, dataInMem_hi_920, dataInMem_lo_728};
  wire [159:0]      dataInMem_lo_lo_hi_hi_hi_12 = {dataInMem_hi_923, dataInMem_lo_731, dataInMem_hi_922, dataInMem_lo_730};
  wire [319:0]      dataInMem_lo_lo_hi_hi_12 = {dataInMem_lo_lo_hi_hi_hi_12, dataInMem_lo_lo_hi_hi_lo_12};
  wire [639:0]      dataInMem_lo_lo_hi_12 = {dataInMem_lo_lo_hi_hi_12, dataInMem_lo_lo_hi_lo_12};
  wire [1279:0]     dataInMem_lo_lo_140 = {dataInMem_lo_lo_hi_12, dataInMem_lo_lo_lo_12};
  wire [159:0]      dataInMem_lo_hi_lo_lo_lo_12 = {dataInMem_hi_925, dataInMem_lo_733, dataInMem_hi_924, dataInMem_lo_732};
  wire [159:0]      dataInMem_lo_hi_lo_lo_hi_12 = {dataInMem_hi_927, dataInMem_lo_735, dataInMem_hi_926, dataInMem_lo_734};
  wire [319:0]      dataInMem_lo_hi_lo_lo_12 = {dataInMem_lo_hi_lo_lo_hi_12, dataInMem_lo_hi_lo_lo_lo_12};
  wire [159:0]      dataInMem_lo_hi_lo_hi_lo_12 = {dataInMem_hi_929, dataInMem_lo_737, dataInMem_hi_928, dataInMem_lo_736};
  wire [159:0]      dataInMem_lo_hi_lo_hi_hi_12 = {dataInMem_hi_931, dataInMem_lo_739, dataInMem_hi_930, dataInMem_lo_738};
  wire [319:0]      dataInMem_lo_hi_lo_hi_12 = {dataInMem_lo_hi_lo_hi_hi_12, dataInMem_lo_hi_lo_hi_lo_12};
  wire [639:0]      dataInMem_lo_hi_lo_12 = {dataInMem_lo_hi_lo_hi_12, dataInMem_lo_hi_lo_lo_12};
  wire [159:0]      dataInMem_lo_hi_hi_lo_lo_12 = {dataInMem_hi_933, dataInMem_lo_741, dataInMem_hi_932, dataInMem_lo_740};
  wire [159:0]      dataInMem_lo_hi_hi_lo_hi_12 = {dataInMem_hi_935, dataInMem_lo_743, dataInMem_hi_934, dataInMem_lo_742};
  wire [319:0]      dataInMem_lo_hi_hi_lo_12 = {dataInMem_lo_hi_hi_lo_hi_12, dataInMem_lo_hi_hi_lo_lo_12};
  wire [159:0]      dataInMem_lo_hi_hi_hi_lo_12 = {dataInMem_hi_937, dataInMem_lo_745, dataInMem_hi_936, dataInMem_lo_744};
  wire [159:0]      dataInMem_lo_hi_hi_hi_hi_12 = {dataInMem_hi_939, dataInMem_lo_747, dataInMem_hi_938, dataInMem_lo_746};
  wire [319:0]      dataInMem_lo_hi_hi_hi_12 = {dataInMem_lo_hi_hi_hi_hi_12, dataInMem_lo_hi_hi_hi_lo_12};
  wire [639:0]      dataInMem_lo_hi_hi_12 = {dataInMem_lo_hi_hi_hi_12, dataInMem_lo_hi_hi_lo_12};
  wire [1279:0]     dataInMem_lo_hi_396 = {dataInMem_lo_hi_hi_12, dataInMem_lo_hi_lo_12};
  wire [2559:0]     dataInMem_lo_780 = {dataInMem_lo_hi_396, dataInMem_lo_lo_140};
  wire [159:0]      dataInMem_hi_lo_lo_lo_lo_12 = {dataInMem_hi_941, dataInMem_lo_749, dataInMem_hi_940, dataInMem_lo_748};
  wire [159:0]      dataInMem_hi_lo_lo_lo_hi_12 = {dataInMem_hi_943, dataInMem_lo_751, dataInMem_hi_942, dataInMem_lo_750};
  wire [319:0]      dataInMem_hi_lo_lo_lo_12 = {dataInMem_hi_lo_lo_lo_hi_12, dataInMem_hi_lo_lo_lo_lo_12};
  wire [159:0]      dataInMem_hi_lo_lo_hi_lo_12 = {dataInMem_hi_945, dataInMem_lo_753, dataInMem_hi_944, dataInMem_lo_752};
  wire [159:0]      dataInMem_hi_lo_lo_hi_hi_12 = {dataInMem_hi_947, dataInMem_lo_755, dataInMem_hi_946, dataInMem_lo_754};
  wire [319:0]      dataInMem_hi_lo_lo_hi_12 = {dataInMem_hi_lo_lo_hi_hi_12, dataInMem_hi_lo_lo_hi_lo_12};
  wire [639:0]      dataInMem_hi_lo_lo_12 = {dataInMem_hi_lo_lo_hi_12, dataInMem_hi_lo_lo_lo_12};
  wire [159:0]      dataInMem_hi_lo_hi_lo_lo_12 = {dataInMem_hi_949, dataInMem_lo_757, dataInMem_hi_948, dataInMem_lo_756};
  wire [159:0]      dataInMem_hi_lo_hi_lo_hi_12 = {dataInMem_hi_951, dataInMem_lo_759, dataInMem_hi_950, dataInMem_lo_758};
  wire [319:0]      dataInMem_hi_lo_hi_lo_12 = {dataInMem_hi_lo_hi_lo_hi_12, dataInMem_hi_lo_hi_lo_lo_12};
  wire [159:0]      dataInMem_hi_lo_hi_hi_lo_12 = {dataInMem_hi_953, dataInMem_lo_761, dataInMem_hi_952, dataInMem_lo_760};
  wire [159:0]      dataInMem_hi_lo_hi_hi_hi_12 = {dataInMem_hi_955, dataInMem_lo_763, dataInMem_hi_954, dataInMem_lo_762};
  wire [319:0]      dataInMem_hi_lo_hi_hi_12 = {dataInMem_hi_lo_hi_hi_hi_12, dataInMem_hi_lo_hi_hi_lo_12};
  wire [639:0]      dataInMem_hi_lo_hi_12 = {dataInMem_hi_lo_hi_hi_12, dataInMem_hi_lo_hi_lo_12};
  wire [1279:0]     dataInMem_hi_lo_268 = {dataInMem_hi_lo_hi_12, dataInMem_hi_lo_lo_12};
  wire [159:0]      dataInMem_hi_hi_lo_lo_lo_12 = {dataInMem_hi_957, dataInMem_lo_765, dataInMem_hi_956, dataInMem_lo_764};
  wire [159:0]      dataInMem_hi_hi_lo_lo_hi_12 = {dataInMem_hi_959, dataInMem_lo_767, dataInMem_hi_958, dataInMem_lo_766};
  wire [319:0]      dataInMem_hi_hi_lo_lo_12 = {dataInMem_hi_hi_lo_lo_hi_12, dataInMem_hi_hi_lo_lo_lo_12};
  wire [159:0]      dataInMem_hi_hi_lo_hi_lo_12 = {dataInMem_hi_961, dataInMem_lo_769, dataInMem_hi_960, dataInMem_lo_768};
  wire [159:0]      dataInMem_hi_hi_lo_hi_hi_12 = {dataInMem_hi_963, dataInMem_lo_771, dataInMem_hi_962, dataInMem_lo_770};
  wire [319:0]      dataInMem_hi_hi_lo_hi_12 = {dataInMem_hi_hi_lo_hi_hi_12, dataInMem_hi_hi_lo_hi_lo_12};
  wire [639:0]      dataInMem_hi_hi_lo_12 = {dataInMem_hi_hi_lo_hi_12, dataInMem_hi_hi_lo_lo_12};
  wire [159:0]      dataInMem_hi_hi_hi_lo_lo_12 = {dataInMem_hi_965, dataInMem_lo_773, dataInMem_hi_964, dataInMem_lo_772};
  wire [159:0]      dataInMem_hi_hi_hi_lo_hi_12 = {dataInMem_hi_967, dataInMem_lo_775, dataInMem_hi_966, dataInMem_lo_774};
  wire [319:0]      dataInMem_hi_hi_hi_lo_12 = {dataInMem_hi_hi_hi_lo_hi_12, dataInMem_hi_hi_hi_lo_lo_12};
  wire [159:0]      dataInMem_hi_hi_hi_hi_lo_12 = {dataInMem_hi_969, dataInMem_lo_777, dataInMem_hi_968, dataInMem_lo_776};
  wire [159:0]      dataInMem_hi_hi_hi_hi_hi_12 = {dataInMem_hi_971, dataInMem_lo_779, dataInMem_hi_970, dataInMem_lo_778};
  wire [319:0]      dataInMem_hi_hi_hi_hi_12 = {dataInMem_hi_hi_hi_hi_hi_12, dataInMem_hi_hi_hi_hi_lo_12};
  wire [639:0]      dataInMem_hi_hi_hi_12 = {dataInMem_hi_hi_hi_hi_12, dataInMem_hi_hi_hi_lo_12};
  wire [1279:0]     dataInMem_hi_hi_588 = {dataInMem_hi_hi_hi_12, dataInMem_hi_hi_lo_12};
  wire [2559:0]     dataInMem_hi_972 = {dataInMem_hi_hi_588, dataInMem_hi_lo_268};
  wire [5119:0]     dataInMem_12 = {dataInMem_hi_972, dataInMem_lo_780};
  wire [1023:0]     regroupCacheLine_12_0 = dataInMem_12[1023:0];
  wire [1023:0]     regroupCacheLine_12_1 = dataInMem_12[2047:1024];
  wire [1023:0]     regroupCacheLine_12_2 = dataInMem_12[3071:2048];
  wire [1023:0]     regroupCacheLine_12_3 = dataInMem_12[4095:3072];
  wire [1023:0]     regroupCacheLine_12_4 = dataInMem_12[5119:4096];
  wire [1023:0]     res_96 = regroupCacheLine_12_0;
  wire [1023:0]     res_97 = regroupCacheLine_12_1;
  wire [1023:0]     res_98 = regroupCacheLine_12_2;
  wire [1023:0]     res_99 = regroupCacheLine_12_3;
  wire [1023:0]     res_100 = regroupCacheLine_12_4;
  wire [2047:0]     lo_lo_12 = {res_97, res_96};
  wire [2047:0]     lo_hi_12 = {res_99, res_98};
  wire [4095:0]     lo_12 = {lo_hi_12, lo_lo_12};
  wire [2047:0]     hi_lo_12 = {1024'h0, res_100};
  wire [4095:0]     hi_12 = {2048'h0, hi_lo_12};
  wire [8191:0]     regroupLoadData_1_4 = {hi_12, lo_12};
  wire [47:0]       dataInMem_lo_781 = {dataInMem_lo_hi_397, dataRegroupBySew_0_1_0};
  wire [31:0]       _GEN_902 = {dataRegroupBySew_5_1_0, dataRegroupBySew_4_1_0};
  wire [31:0]       dataInMem_hi_hi_589;
  assign dataInMem_hi_hi_589 = _GEN_902;
  wire [31:0]       dataInMem_hi_lo_335;
  assign dataInMem_hi_lo_335 = _GEN_902;
  wire [47:0]       dataInMem_hi_973 = {dataInMem_hi_hi_589, dataRegroupBySew_3_1_0};
  wire [47:0]       dataInMem_lo_782 = {dataInMem_lo_hi_398, dataRegroupBySew_0_1_1};
  wire [31:0]       _GEN_903 = {dataRegroupBySew_5_1_1, dataRegroupBySew_4_1_1};
  wire [31:0]       dataInMem_hi_hi_590;
  assign dataInMem_hi_hi_590 = _GEN_903;
  wire [31:0]       dataInMem_hi_lo_336;
  assign dataInMem_hi_lo_336 = _GEN_903;
  wire [47:0]       dataInMem_hi_974 = {dataInMem_hi_hi_590, dataRegroupBySew_3_1_1};
  wire [47:0]       dataInMem_lo_783 = {dataInMem_lo_hi_399, dataRegroupBySew_0_1_2};
  wire [31:0]       _GEN_904 = {dataRegroupBySew_5_1_2, dataRegroupBySew_4_1_2};
  wire [31:0]       dataInMem_hi_hi_591;
  assign dataInMem_hi_hi_591 = _GEN_904;
  wire [31:0]       dataInMem_hi_lo_337;
  assign dataInMem_hi_lo_337 = _GEN_904;
  wire [47:0]       dataInMem_hi_975 = {dataInMem_hi_hi_591, dataRegroupBySew_3_1_2};
  wire [47:0]       dataInMem_lo_784 = {dataInMem_lo_hi_400, dataRegroupBySew_0_1_3};
  wire [31:0]       _GEN_905 = {dataRegroupBySew_5_1_3, dataRegroupBySew_4_1_3};
  wire [31:0]       dataInMem_hi_hi_592;
  assign dataInMem_hi_hi_592 = _GEN_905;
  wire [31:0]       dataInMem_hi_lo_338;
  assign dataInMem_hi_lo_338 = _GEN_905;
  wire [47:0]       dataInMem_hi_976 = {dataInMem_hi_hi_592, dataRegroupBySew_3_1_3};
  wire [47:0]       dataInMem_lo_785 = {dataInMem_lo_hi_401, dataRegroupBySew_0_1_4};
  wire [31:0]       _GEN_906 = {dataRegroupBySew_5_1_4, dataRegroupBySew_4_1_4};
  wire [31:0]       dataInMem_hi_hi_593;
  assign dataInMem_hi_hi_593 = _GEN_906;
  wire [31:0]       dataInMem_hi_lo_339;
  assign dataInMem_hi_lo_339 = _GEN_906;
  wire [47:0]       dataInMem_hi_977 = {dataInMem_hi_hi_593, dataRegroupBySew_3_1_4};
  wire [47:0]       dataInMem_lo_786 = {dataInMem_lo_hi_402, dataRegroupBySew_0_1_5};
  wire [31:0]       _GEN_907 = {dataRegroupBySew_5_1_5, dataRegroupBySew_4_1_5};
  wire [31:0]       dataInMem_hi_hi_594;
  assign dataInMem_hi_hi_594 = _GEN_907;
  wire [31:0]       dataInMem_hi_lo_340;
  assign dataInMem_hi_lo_340 = _GEN_907;
  wire [47:0]       dataInMem_hi_978 = {dataInMem_hi_hi_594, dataRegroupBySew_3_1_5};
  wire [47:0]       dataInMem_lo_787 = {dataInMem_lo_hi_403, dataRegroupBySew_0_1_6};
  wire [31:0]       _GEN_908 = {dataRegroupBySew_5_1_6, dataRegroupBySew_4_1_6};
  wire [31:0]       dataInMem_hi_hi_595;
  assign dataInMem_hi_hi_595 = _GEN_908;
  wire [31:0]       dataInMem_hi_lo_341;
  assign dataInMem_hi_lo_341 = _GEN_908;
  wire [47:0]       dataInMem_hi_979 = {dataInMem_hi_hi_595, dataRegroupBySew_3_1_6};
  wire [47:0]       dataInMem_lo_788 = {dataInMem_lo_hi_404, dataRegroupBySew_0_1_7};
  wire [31:0]       _GEN_909 = {dataRegroupBySew_5_1_7, dataRegroupBySew_4_1_7};
  wire [31:0]       dataInMem_hi_hi_596;
  assign dataInMem_hi_hi_596 = _GEN_909;
  wire [31:0]       dataInMem_hi_lo_342;
  assign dataInMem_hi_lo_342 = _GEN_909;
  wire [47:0]       dataInMem_hi_980 = {dataInMem_hi_hi_596, dataRegroupBySew_3_1_7};
  wire [47:0]       dataInMem_lo_789 = {dataInMem_lo_hi_405, dataRegroupBySew_0_1_8};
  wire [31:0]       _GEN_910 = {dataRegroupBySew_5_1_8, dataRegroupBySew_4_1_8};
  wire [31:0]       dataInMem_hi_hi_597;
  assign dataInMem_hi_hi_597 = _GEN_910;
  wire [31:0]       dataInMem_hi_lo_343;
  assign dataInMem_hi_lo_343 = _GEN_910;
  wire [47:0]       dataInMem_hi_981 = {dataInMem_hi_hi_597, dataRegroupBySew_3_1_8};
  wire [47:0]       dataInMem_lo_790 = {dataInMem_lo_hi_406, dataRegroupBySew_0_1_9};
  wire [31:0]       _GEN_911 = {dataRegroupBySew_5_1_9, dataRegroupBySew_4_1_9};
  wire [31:0]       dataInMem_hi_hi_598;
  assign dataInMem_hi_hi_598 = _GEN_911;
  wire [31:0]       dataInMem_hi_lo_344;
  assign dataInMem_hi_lo_344 = _GEN_911;
  wire [47:0]       dataInMem_hi_982 = {dataInMem_hi_hi_598, dataRegroupBySew_3_1_9};
  wire [47:0]       dataInMem_lo_791 = {dataInMem_lo_hi_407, dataRegroupBySew_0_1_10};
  wire [31:0]       _GEN_912 = {dataRegroupBySew_5_1_10, dataRegroupBySew_4_1_10};
  wire [31:0]       dataInMem_hi_hi_599;
  assign dataInMem_hi_hi_599 = _GEN_912;
  wire [31:0]       dataInMem_hi_lo_345;
  assign dataInMem_hi_lo_345 = _GEN_912;
  wire [47:0]       dataInMem_hi_983 = {dataInMem_hi_hi_599, dataRegroupBySew_3_1_10};
  wire [47:0]       dataInMem_lo_792 = {dataInMem_lo_hi_408, dataRegroupBySew_0_1_11};
  wire [31:0]       _GEN_913 = {dataRegroupBySew_5_1_11, dataRegroupBySew_4_1_11};
  wire [31:0]       dataInMem_hi_hi_600;
  assign dataInMem_hi_hi_600 = _GEN_913;
  wire [31:0]       dataInMem_hi_lo_346;
  assign dataInMem_hi_lo_346 = _GEN_913;
  wire [47:0]       dataInMem_hi_984 = {dataInMem_hi_hi_600, dataRegroupBySew_3_1_11};
  wire [47:0]       dataInMem_lo_793 = {dataInMem_lo_hi_409, dataRegroupBySew_0_1_12};
  wire [31:0]       _GEN_914 = {dataRegroupBySew_5_1_12, dataRegroupBySew_4_1_12};
  wire [31:0]       dataInMem_hi_hi_601;
  assign dataInMem_hi_hi_601 = _GEN_914;
  wire [31:0]       dataInMem_hi_lo_347;
  assign dataInMem_hi_lo_347 = _GEN_914;
  wire [47:0]       dataInMem_hi_985 = {dataInMem_hi_hi_601, dataRegroupBySew_3_1_12};
  wire [47:0]       dataInMem_lo_794 = {dataInMem_lo_hi_410, dataRegroupBySew_0_1_13};
  wire [31:0]       _GEN_915 = {dataRegroupBySew_5_1_13, dataRegroupBySew_4_1_13};
  wire [31:0]       dataInMem_hi_hi_602;
  assign dataInMem_hi_hi_602 = _GEN_915;
  wire [31:0]       dataInMem_hi_lo_348;
  assign dataInMem_hi_lo_348 = _GEN_915;
  wire [47:0]       dataInMem_hi_986 = {dataInMem_hi_hi_602, dataRegroupBySew_3_1_13};
  wire [47:0]       dataInMem_lo_795 = {dataInMem_lo_hi_411, dataRegroupBySew_0_1_14};
  wire [31:0]       _GEN_916 = {dataRegroupBySew_5_1_14, dataRegroupBySew_4_1_14};
  wire [31:0]       dataInMem_hi_hi_603;
  assign dataInMem_hi_hi_603 = _GEN_916;
  wire [31:0]       dataInMem_hi_lo_349;
  assign dataInMem_hi_lo_349 = _GEN_916;
  wire [47:0]       dataInMem_hi_987 = {dataInMem_hi_hi_603, dataRegroupBySew_3_1_14};
  wire [47:0]       dataInMem_lo_796 = {dataInMem_lo_hi_412, dataRegroupBySew_0_1_15};
  wire [31:0]       _GEN_917 = {dataRegroupBySew_5_1_15, dataRegroupBySew_4_1_15};
  wire [31:0]       dataInMem_hi_hi_604;
  assign dataInMem_hi_hi_604 = _GEN_917;
  wire [31:0]       dataInMem_hi_lo_350;
  assign dataInMem_hi_lo_350 = _GEN_917;
  wire [47:0]       dataInMem_hi_988 = {dataInMem_hi_hi_604, dataRegroupBySew_3_1_15};
  wire [47:0]       dataInMem_lo_797 = {dataInMem_lo_hi_413, dataRegroupBySew_0_1_16};
  wire [31:0]       _GEN_918 = {dataRegroupBySew_5_1_16, dataRegroupBySew_4_1_16};
  wire [31:0]       dataInMem_hi_hi_605;
  assign dataInMem_hi_hi_605 = _GEN_918;
  wire [31:0]       dataInMem_hi_lo_351;
  assign dataInMem_hi_lo_351 = _GEN_918;
  wire [47:0]       dataInMem_hi_989 = {dataInMem_hi_hi_605, dataRegroupBySew_3_1_16};
  wire [47:0]       dataInMem_lo_798 = {dataInMem_lo_hi_414, dataRegroupBySew_0_1_17};
  wire [31:0]       _GEN_919 = {dataRegroupBySew_5_1_17, dataRegroupBySew_4_1_17};
  wire [31:0]       dataInMem_hi_hi_606;
  assign dataInMem_hi_hi_606 = _GEN_919;
  wire [31:0]       dataInMem_hi_lo_352;
  assign dataInMem_hi_lo_352 = _GEN_919;
  wire [47:0]       dataInMem_hi_990 = {dataInMem_hi_hi_606, dataRegroupBySew_3_1_17};
  wire [47:0]       dataInMem_lo_799 = {dataInMem_lo_hi_415, dataRegroupBySew_0_1_18};
  wire [31:0]       _GEN_920 = {dataRegroupBySew_5_1_18, dataRegroupBySew_4_1_18};
  wire [31:0]       dataInMem_hi_hi_607;
  assign dataInMem_hi_hi_607 = _GEN_920;
  wire [31:0]       dataInMem_hi_lo_353;
  assign dataInMem_hi_lo_353 = _GEN_920;
  wire [47:0]       dataInMem_hi_991 = {dataInMem_hi_hi_607, dataRegroupBySew_3_1_18};
  wire [47:0]       dataInMem_lo_800 = {dataInMem_lo_hi_416, dataRegroupBySew_0_1_19};
  wire [31:0]       _GEN_921 = {dataRegroupBySew_5_1_19, dataRegroupBySew_4_1_19};
  wire [31:0]       dataInMem_hi_hi_608;
  assign dataInMem_hi_hi_608 = _GEN_921;
  wire [31:0]       dataInMem_hi_lo_354;
  assign dataInMem_hi_lo_354 = _GEN_921;
  wire [47:0]       dataInMem_hi_992 = {dataInMem_hi_hi_608, dataRegroupBySew_3_1_19};
  wire [47:0]       dataInMem_lo_801 = {dataInMem_lo_hi_417, dataRegroupBySew_0_1_20};
  wire [31:0]       _GEN_922 = {dataRegroupBySew_5_1_20, dataRegroupBySew_4_1_20};
  wire [31:0]       dataInMem_hi_hi_609;
  assign dataInMem_hi_hi_609 = _GEN_922;
  wire [31:0]       dataInMem_hi_lo_355;
  assign dataInMem_hi_lo_355 = _GEN_922;
  wire [47:0]       dataInMem_hi_993 = {dataInMem_hi_hi_609, dataRegroupBySew_3_1_20};
  wire [47:0]       dataInMem_lo_802 = {dataInMem_lo_hi_418, dataRegroupBySew_0_1_21};
  wire [31:0]       _GEN_923 = {dataRegroupBySew_5_1_21, dataRegroupBySew_4_1_21};
  wire [31:0]       dataInMem_hi_hi_610;
  assign dataInMem_hi_hi_610 = _GEN_923;
  wire [31:0]       dataInMem_hi_lo_356;
  assign dataInMem_hi_lo_356 = _GEN_923;
  wire [47:0]       dataInMem_hi_994 = {dataInMem_hi_hi_610, dataRegroupBySew_3_1_21};
  wire [47:0]       dataInMem_lo_803 = {dataInMem_lo_hi_419, dataRegroupBySew_0_1_22};
  wire [31:0]       _GEN_924 = {dataRegroupBySew_5_1_22, dataRegroupBySew_4_1_22};
  wire [31:0]       dataInMem_hi_hi_611;
  assign dataInMem_hi_hi_611 = _GEN_924;
  wire [31:0]       dataInMem_hi_lo_357;
  assign dataInMem_hi_lo_357 = _GEN_924;
  wire [47:0]       dataInMem_hi_995 = {dataInMem_hi_hi_611, dataRegroupBySew_3_1_22};
  wire [47:0]       dataInMem_lo_804 = {dataInMem_lo_hi_420, dataRegroupBySew_0_1_23};
  wire [31:0]       _GEN_925 = {dataRegroupBySew_5_1_23, dataRegroupBySew_4_1_23};
  wire [31:0]       dataInMem_hi_hi_612;
  assign dataInMem_hi_hi_612 = _GEN_925;
  wire [31:0]       dataInMem_hi_lo_358;
  assign dataInMem_hi_lo_358 = _GEN_925;
  wire [47:0]       dataInMem_hi_996 = {dataInMem_hi_hi_612, dataRegroupBySew_3_1_23};
  wire [47:0]       dataInMem_lo_805 = {dataInMem_lo_hi_421, dataRegroupBySew_0_1_24};
  wire [31:0]       _GEN_926 = {dataRegroupBySew_5_1_24, dataRegroupBySew_4_1_24};
  wire [31:0]       dataInMem_hi_hi_613;
  assign dataInMem_hi_hi_613 = _GEN_926;
  wire [31:0]       dataInMem_hi_lo_359;
  assign dataInMem_hi_lo_359 = _GEN_926;
  wire [47:0]       dataInMem_hi_997 = {dataInMem_hi_hi_613, dataRegroupBySew_3_1_24};
  wire [47:0]       dataInMem_lo_806 = {dataInMem_lo_hi_422, dataRegroupBySew_0_1_25};
  wire [31:0]       _GEN_927 = {dataRegroupBySew_5_1_25, dataRegroupBySew_4_1_25};
  wire [31:0]       dataInMem_hi_hi_614;
  assign dataInMem_hi_hi_614 = _GEN_927;
  wire [31:0]       dataInMem_hi_lo_360;
  assign dataInMem_hi_lo_360 = _GEN_927;
  wire [47:0]       dataInMem_hi_998 = {dataInMem_hi_hi_614, dataRegroupBySew_3_1_25};
  wire [47:0]       dataInMem_lo_807 = {dataInMem_lo_hi_423, dataRegroupBySew_0_1_26};
  wire [31:0]       _GEN_928 = {dataRegroupBySew_5_1_26, dataRegroupBySew_4_1_26};
  wire [31:0]       dataInMem_hi_hi_615;
  assign dataInMem_hi_hi_615 = _GEN_928;
  wire [31:0]       dataInMem_hi_lo_361;
  assign dataInMem_hi_lo_361 = _GEN_928;
  wire [47:0]       dataInMem_hi_999 = {dataInMem_hi_hi_615, dataRegroupBySew_3_1_26};
  wire [47:0]       dataInMem_lo_808 = {dataInMem_lo_hi_424, dataRegroupBySew_0_1_27};
  wire [31:0]       _GEN_929 = {dataRegroupBySew_5_1_27, dataRegroupBySew_4_1_27};
  wire [31:0]       dataInMem_hi_hi_616;
  assign dataInMem_hi_hi_616 = _GEN_929;
  wire [31:0]       dataInMem_hi_lo_362;
  assign dataInMem_hi_lo_362 = _GEN_929;
  wire [47:0]       dataInMem_hi_1000 = {dataInMem_hi_hi_616, dataRegroupBySew_3_1_27};
  wire [47:0]       dataInMem_lo_809 = {dataInMem_lo_hi_425, dataRegroupBySew_0_1_28};
  wire [31:0]       _GEN_930 = {dataRegroupBySew_5_1_28, dataRegroupBySew_4_1_28};
  wire [31:0]       dataInMem_hi_hi_617;
  assign dataInMem_hi_hi_617 = _GEN_930;
  wire [31:0]       dataInMem_hi_lo_363;
  assign dataInMem_hi_lo_363 = _GEN_930;
  wire [47:0]       dataInMem_hi_1001 = {dataInMem_hi_hi_617, dataRegroupBySew_3_1_28};
  wire [47:0]       dataInMem_lo_810 = {dataInMem_lo_hi_426, dataRegroupBySew_0_1_29};
  wire [31:0]       _GEN_931 = {dataRegroupBySew_5_1_29, dataRegroupBySew_4_1_29};
  wire [31:0]       dataInMem_hi_hi_618;
  assign dataInMem_hi_hi_618 = _GEN_931;
  wire [31:0]       dataInMem_hi_lo_364;
  assign dataInMem_hi_lo_364 = _GEN_931;
  wire [47:0]       dataInMem_hi_1002 = {dataInMem_hi_hi_618, dataRegroupBySew_3_1_29};
  wire [47:0]       dataInMem_lo_811 = {dataInMem_lo_hi_427, dataRegroupBySew_0_1_30};
  wire [31:0]       _GEN_932 = {dataRegroupBySew_5_1_30, dataRegroupBySew_4_1_30};
  wire [31:0]       dataInMem_hi_hi_619;
  assign dataInMem_hi_hi_619 = _GEN_932;
  wire [31:0]       dataInMem_hi_lo_365;
  assign dataInMem_hi_lo_365 = _GEN_932;
  wire [47:0]       dataInMem_hi_1003 = {dataInMem_hi_hi_619, dataRegroupBySew_3_1_30};
  wire [47:0]       dataInMem_lo_812 = {dataInMem_lo_hi_428, dataRegroupBySew_0_1_31};
  wire [31:0]       _GEN_933 = {dataRegroupBySew_5_1_31, dataRegroupBySew_4_1_31};
  wire [31:0]       dataInMem_hi_hi_620;
  assign dataInMem_hi_hi_620 = _GEN_933;
  wire [31:0]       dataInMem_hi_lo_366;
  assign dataInMem_hi_lo_366 = _GEN_933;
  wire [47:0]       dataInMem_hi_1004 = {dataInMem_hi_hi_620, dataRegroupBySew_3_1_31};
  wire [47:0]       dataInMem_lo_813 = {dataInMem_lo_hi_429, dataRegroupBySew_0_1_32};
  wire [31:0]       _GEN_934 = {dataRegroupBySew_5_1_32, dataRegroupBySew_4_1_32};
  wire [31:0]       dataInMem_hi_hi_621;
  assign dataInMem_hi_hi_621 = _GEN_934;
  wire [31:0]       dataInMem_hi_lo_367;
  assign dataInMem_hi_lo_367 = _GEN_934;
  wire [47:0]       dataInMem_hi_1005 = {dataInMem_hi_hi_621, dataRegroupBySew_3_1_32};
  wire [47:0]       dataInMem_lo_814 = {dataInMem_lo_hi_430, dataRegroupBySew_0_1_33};
  wire [31:0]       _GEN_935 = {dataRegroupBySew_5_1_33, dataRegroupBySew_4_1_33};
  wire [31:0]       dataInMem_hi_hi_622;
  assign dataInMem_hi_hi_622 = _GEN_935;
  wire [31:0]       dataInMem_hi_lo_368;
  assign dataInMem_hi_lo_368 = _GEN_935;
  wire [47:0]       dataInMem_hi_1006 = {dataInMem_hi_hi_622, dataRegroupBySew_3_1_33};
  wire [47:0]       dataInMem_lo_815 = {dataInMem_lo_hi_431, dataRegroupBySew_0_1_34};
  wire [31:0]       _GEN_936 = {dataRegroupBySew_5_1_34, dataRegroupBySew_4_1_34};
  wire [31:0]       dataInMem_hi_hi_623;
  assign dataInMem_hi_hi_623 = _GEN_936;
  wire [31:0]       dataInMem_hi_lo_369;
  assign dataInMem_hi_lo_369 = _GEN_936;
  wire [47:0]       dataInMem_hi_1007 = {dataInMem_hi_hi_623, dataRegroupBySew_3_1_34};
  wire [47:0]       dataInMem_lo_816 = {dataInMem_lo_hi_432, dataRegroupBySew_0_1_35};
  wire [31:0]       _GEN_937 = {dataRegroupBySew_5_1_35, dataRegroupBySew_4_1_35};
  wire [31:0]       dataInMem_hi_hi_624;
  assign dataInMem_hi_hi_624 = _GEN_937;
  wire [31:0]       dataInMem_hi_lo_370;
  assign dataInMem_hi_lo_370 = _GEN_937;
  wire [47:0]       dataInMem_hi_1008 = {dataInMem_hi_hi_624, dataRegroupBySew_3_1_35};
  wire [47:0]       dataInMem_lo_817 = {dataInMem_lo_hi_433, dataRegroupBySew_0_1_36};
  wire [31:0]       _GEN_938 = {dataRegroupBySew_5_1_36, dataRegroupBySew_4_1_36};
  wire [31:0]       dataInMem_hi_hi_625;
  assign dataInMem_hi_hi_625 = _GEN_938;
  wire [31:0]       dataInMem_hi_lo_371;
  assign dataInMem_hi_lo_371 = _GEN_938;
  wire [47:0]       dataInMem_hi_1009 = {dataInMem_hi_hi_625, dataRegroupBySew_3_1_36};
  wire [47:0]       dataInMem_lo_818 = {dataInMem_lo_hi_434, dataRegroupBySew_0_1_37};
  wire [31:0]       _GEN_939 = {dataRegroupBySew_5_1_37, dataRegroupBySew_4_1_37};
  wire [31:0]       dataInMem_hi_hi_626;
  assign dataInMem_hi_hi_626 = _GEN_939;
  wire [31:0]       dataInMem_hi_lo_372;
  assign dataInMem_hi_lo_372 = _GEN_939;
  wire [47:0]       dataInMem_hi_1010 = {dataInMem_hi_hi_626, dataRegroupBySew_3_1_37};
  wire [47:0]       dataInMem_lo_819 = {dataInMem_lo_hi_435, dataRegroupBySew_0_1_38};
  wire [31:0]       _GEN_940 = {dataRegroupBySew_5_1_38, dataRegroupBySew_4_1_38};
  wire [31:0]       dataInMem_hi_hi_627;
  assign dataInMem_hi_hi_627 = _GEN_940;
  wire [31:0]       dataInMem_hi_lo_373;
  assign dataInMem_hi_lo_373 = _GEN_940;
  wire [47:0]       dataInMem_hi_1011 = {dataInMem_hi_hi_627, dataRegroupBySew_3_1_38};
  wire [47:0]       dataInMem_lo_820 = {dataInMem_lo_hi_436, dataRegroupBySew_0_1_39};
  wire [31:0]       _GEN_941 = {dataRegroupBySew_5_1_39, dataRegroupBySew_4_1_39};
  wire [31:0]       dataInMem_hi_hi_628;
  assign dataInMem_hi_hi_628 = _GEN_941;
  wire [31:0]       dataInMem_hi_lo_374;
  assign dataInMem_hi_lo_374 = _GEN_941;
  wire [47:0]       dataInMem_hi_1012 = {dataInMem_hi_hi_628, dataRegroupBySew_3_1_39};
  wire [47:0]       dataInMem_lo_821 = {dataInMem_lo_hi_437, dataRegroupBySew_0_1_40};
  wire [31:0]       _GEN_942 = {dataRegroupBySew_5_1_40, dataRegroupBySew_4_1_40};
  wire [31:0]       dataInMem_hi_hi_629;
  assign dataInMem_hi_hi_629 = _GEN_942;
  wire [31:0]       dataInMem_hi_lo_375;
  assign dataInMem_hi_lo_375 = _GEN_942;
  wire [47:0]       dataInMem_hi_1013 = {dataInMem_hi_hi_629, dataRegroupBySew_3_1_40};
  wire [47:0]       dataInMem_lo_822 = {dataInMem_lo_hi_438, dataRegroupBySew_0_1_41};
  wire [31:0]       _GEN_943 = {dataRegroupBySew_5_1_41, dataRegroupBySew_4_1_41};
  wire [31:0]       dataInMem_hi_hi_630;
  assign dataInMem_hi_hi_630 = _GEN_943;
  wire [31:0]       dataInMem_hi_lo_376;
  assign dataInMem_hi_lo_376 = _GEN_943;
  wire [47:0]       dataInMem_hi_1014 = {dataInMem_hi_hi_630, dataRegroupBySew_3_1_41};
  wire [47:0]       dataInMem_lo_823 = {dataInMem_lo_hi_439, dataRegroupBySew_0_1_42};
  wire [31:0]       _GEN_944 = {dataRegroupBySew_5_1_42, dataRegroupBySew_4_1_42};
  wire [31:0]       dataInMem_hi_hi_631;
  assign dataInMem_hi_hi_631 = _GEN_944;
  wire [31:0]       dataInMem_hi_lo_377;
  assign dataInMem_hi_lo_377 = _GEN_944;
  wire [47:0]       dataInMem_hi_1015 = {dataInMem_hi_hi_631, dataRegroupBySew_3_1_42};
  wire [47:0]       dataInMem_lo_824 = {dataInMem_lo_hi_440, dataRegroupBySew_0_1_43};
  wire [31:0]       _GEN_945 = {dataRegroupBySew_5_1_43, dataRegroupBySew_4_1_43};
  wire [31:0]       dataInMem_hi_hi_632;
  assign dataInMem_hi_hi_632 = _GEN_945;
  wire [31:0]       dataInMem_hi_lo_378;
  assign dataInMem_hi_lo_378 = _GEN_945;
  wire [47:0]       dataInMem_hi_1016 = {dataInMem_hi_hi_632, dataRegroupBySew_3_1_43};
  wire [47:0]       dataInMem_lo_825 = {dataInMem_lo_hi_441, dataRegroupBySew_0_1_44};
  wire [31:0]       _GEN_946 = {dataRegroupBySew_5_1_44, dataRegroupBySew_4_1_44};
  wire [31:0]       dataInMem_hi_hi_633;
  assign dataInMem_hi_hi_633 = _GEN_946;
  wire [31:0]       dataInMem_hi_lo_379;
  assign dataInMem_hi_lo_379 = _GEN_946;
  wire [47:0]       dataInMem_hi_1017 = {dataInMem_hi_hi_633, dataRegroupBySew_3_1_44};
  wire [47:0]       dataInMem_lo_826 = {dataInMem_lo_hi_442, dataRegroupBySew_0_1_45};
  wire [31:0]       _GEN_947 = {dataRegroupBySew_5_1_45, dataRegroupBySew_4_1_45};
  wire [31:0]       dataInMem_hi_hi_634;
  assign dataInMem_hi_hi_634 = _GEN_947;
  wire [31:0]       dataInMem_hi_lo_380;
  assign dataInMem_hi_lo_380 = _GEN_947;
  wire [47:0]       dataInMem_hi_1018 = {dataInMem_hi_hi_634, dataRegroupBySew_3_1_45};
  wire [47:0]       dataInMem_lo_827 = {dataInMem_lo_hi_443, dataRegroupBySew_0_1_46};
  wire [31:0]       _GEN_948 = {dataRegroupBySew_5_1_46, dataRegroupBySew_4_1_46};
  wire [31:0]       dataInMem_hi_hi_635;
  assign dataInMem_hi_hi_635 = _GEN_948;
  wire [31:0]       dataInMem_hi_lo_381;
  assign dataInMem_hi_lo_381 = _GEN_948;
  wire [47:0]       dataInMem_hi_1019 = {dataInMem_hi_hi_635, dataRegroupBySew_3_1_46};
  wire [47:0]       dataInMem_lo_828 = {dataInMem_lo_hi_444, dataRegroupBySew_0_1_47};
  wire [31:0]       _GEN_949 = {dataRegroupBySew_5_1_47, dataRegroupBySew_4_1_47};
  wire [31:0]       dataInMem_hi_hi_636;
  assign dataInMem_hi_hi_636 = _GEN_949;
  wire [31:0]       dataInMem_hi_lo_382;
  assign dataInMem_hi_lo_382 = _GEN_949;
  wire [47:0]       dataInMem_hi_1020 = {dataInMem_hi_hi_636, dataRegroupBySew_3_1_47};
  wire [47:0]       dataInMem_lo_829 = {dataInMem_lo_hi_445, dataRegroupBySew_0_1_48};
  wire [31:0]       _GEN_950 = {dataRegroupBySew_5_1_48, dataRegroupBySew_4_1_48};
  wire [31:0]       dataInMem_hi_hi_637;
  assign dataInMem_hi_hi_637 = _GEN_950;
  wire [31:0]       dataInMem_hi_lo_383;
  assign dataInMem_hi_lo_383 = _GEN_950;
  wire [47:0]       dataInMem_hi_1021 = {dataInMem_hi_hi_637, dataRegroupBySew_3_1_48};
  wire [47:0]       dataInMem_lo_830 = {dataInMem_lo_hi_446, dataRegroupBySew_0_1_49};
  wire [31:0]       _GEN_951 = {dataRegroupBySew_5_1_49, dataRegroupBySew_4_1_49};
  wire [31:0]       dataInMem_hi_hi_638;
  assign dataInMem_hi_hi_638 = _GEN_951;
  wire [31:0]       dataInMem_hi_lo_384;
  assign dataInMem_hi_lo_384 = _GEN_951;
  wire [47:0]       dataInMem_hi_1022 = {dataInMem_hi_hi_638, dataRegroupBySew_3_1_49};
  wire [47:0]       dataInMem_lo_831 = {dataInMem_lo_hi_447, dataRegroupBySew_0_1_50};
  wire [31:0]       _GEN_952 = {dataRegroupBySew_5_1_50, dataRegroupBySew_4_1_50};
  wire [31:0]       dataInMem_hi_hi_639;
  assign dataInMem_hi_hi_639 = _GEN_952;
  wire [31:0]       dataInMem_hi_lo_385;
  assign dataInMem_hi_lo_385 = _GEN_952;
  wire [47:0]       dataInMem_hi_1023 = {dataInMem_hi_hi_639, dataRegroupBySew_3_1_50};
  wire [47:0]       dataInMem_lo_832 = {dataInMem_lo_hi_448, dataRegroupBySew_0_1_51};
  wire [31:0]       _GEN_953 = {dataRegroupBySew_5_1_51, dataRegroupBySew_4_1_51};
  wire [31:0]       dataInMem_hi_hi_640;
  assign dataInMem_hi_hi_640 = _GEN_953;
  wire [31:0]       dataInMem_hi_lo_386;
  assign dataInMem_hi_lo_386 = _GEN_953;
  wire [47:0]       dataInMem_hi_1024 = {dataInMem_hi_hi_640, dataRegroupBySew_3_1_51};
  wire [47:0]       dataInMem_lo_833 = {dataInMem_lo_hi_449, dataRegroupBySew_0_1_52};
  wire [31:0]       _GEN_954 = {dataRegroupBySew_5_1_52, dataRegroupBySew_4_1_52};
  wire [31:0]       dataInMem_hi_hi_641;
  assign dataInMem_hi_hi_641 = _GEN_954;
  wire [31:0]       dataInMem_hi_lo_387;
  assign dataInMem_hi_lo_387 = _GEN_954;
  wire [47:0]       dataInMem_hi_1025 = {dataInMem_hi_hi_641, dataRegroupBySew_3_1_52};
  wire [47:0]       dataInMem_lo_834 = {dataInMem_lo_hi_450, dataRegroupBySew_0_1_53};
  wire [31:0]       _GEN_955 = {dataRegroupBySew_5_1_53, dataRegroupBySew_4_1_53};
  wire [31:0]       dataInMem_hi_hi_642;
  assign dataInMem_hi_hi_642 = _GEN_955;
  wire [31:0]       dataInMem_hi_lo_388;
  assign dataInMem_hi_lo_388 = _GEN_955;
  wire [47:0]       dataInMem_hi_1026 = {dataInMem_hi_hi_642, dataRegroupBySew_3_1_53};
  wire [47:0]       dataInMem_lo_835 = {dataInMem_lo_hi_451, dataRegroupBySew_0_1_54};
  wire [31:0]       _GEN_956 = {dataRegroupBySew_5_1_54, dataRegroupBySew_4_1_54};
  wire [31:0]       dataInMem_hi_hi_643;
  assign dataInMem_hi_hi_643 = _GEN_956;
  wire [31:0]       dataInMem_hi_lo_389;
  assign dataInMem_hi_lo_389 = _GEN_956;
  wire [47:0]       dataInMem_hi_1027 = {dataInMem_hi_hi_643, dataRegroupBySew_3_1_54};
  wire [47:0]       dataInMem_lo_836 = {dataInMem_lo_hi_452, dataRegroupBySew_0_1_55};
  wire [31:0]       _GEN_957 = {dataRegroupBySew_5_1_55, dataRegroupBySew_4_1_55};
  wire [31:0]       dataInMem_hi_hi_644;
  assign dataInMem_hi_hi_644 = _GEN_957;
  wire [31:0]       dataInMem_hi_lo_390;
  assign dataInMem_hi_lo_390 = _GEN_957;
  wire [47:0]       dataInMem_hi_1028 = {dataInMem_hi_hi_644, dataRegroupBySew_3_1_55};
  wire [47:0]       dataInMem_lo_837 = {dataInMem_lo_hi_453, dataRegroupBySew_0_1_56};
  wire [31:0]       _GEN_958 = {dataRegroupBySew_5_1_56, dataRegroupBySew_4_1_56};
  wire [31:0]       dataInMem_hi_hi_645;
  assign dataInMem_hi_hi_645 = _GEN_958;
  wire [31:0]       dataInMem_hi_lo_391;
  assign dataInMem_hi_lo_391 = _GEN_958;
  wire [47:0]       dataInMem_hi_1029 = {dataInMem_hi_hi_645, dataRegroupBySew_3_1_56};
  wire [47:0]       dataInMem_lo_838 = {dataInMem_lo_hi_454, dataRegroupBySew_0_1_57};
  wire [31:0]       _GEN_959 = {dataRegroupBySew_5_1_57, dataRegroupBySew_4_1_57};
  wire [31:0]       dataInMem_hi_hi_646;
  assign dataInMem_hi_hi_646 = _GEN_959;
  wire [31:0]       dataInMem_hi_lo_392;
  assign dataInMem_hi_lo_392 = _GEN_959;
  wire [47:0]       dataInMem_hi_1030 = {dataInMem_hi_hi_646, dataRegroupBySew_3_1_57};
  wire [47:0]       dataInMem_lo_839 = {dataInMem_lo_hi_455, dataRegroupBySew_0_1_58};
  wire [31:0]       _GEN_960 = {dataRegroupBySew_5_1_58, dataRegroupBySew_4_1_58};
  wire [31:0]       dataInMem_hi_hi_647;
  assign dataInMem_hi_hi_647 = _GEN_960;
  wire [31:0]       dataInMem_hi_lo_393;
  assign dataInMem_hi_lo_393 = _GEN_960;
  wire [47:0]       dataInMem_hi_1031 = {dataInMem_hi_hi_647, dataRegroupBySew_3_1_58};
  wire [47:0]       dataInMem_lo_840 = {dataInMem_lo_hi_456, dataRegroupBySew_0_1_59};
  wire [31:0]       _GEN_961 = {dataRegroupBySew_5_1_59, dataRegroupBySew_4_1_59};
  wire [31:0]       dataInMem_hi_hi_648;
  assign dataInMem_hi_hi_648 = _GEN_961;
  wire [31:0]       dataInMem_hi_lo_394;
  assign dataInMem_hi_lo_394 = _GEN_961;
  wire [47:0]       dataInMem_hi_1032 = {dataInMem_hi_hi_648, dataRegroupBySew_3_1_59};
  wire [47:0]       dataInMem_lo_841 = {dataInMem_lo_hi_457, dataRegroupBySew_0_1_60};
  wire [31:0]       _GEN_962 = {dataRegroupBySew_5_1_60, dataRegroupBySew_4_1_60};
  wire [31:0]       dataInMem_hi_hi_649;
  assign dataInMem_hi_hi_649 = _GEN_962;
  wire [31:0]       dataInMem_hi_lo_395;
  assign dataInMem_hi_lo_395 = _GEN_962;
  wire [47:0]       dataInMem_hi_1033 = {dataInMem_hi_hi_649, dataRegroupBySew_3_1_60};
  wire [47:0]       dataInMem_lo_842 = {dataInMem_lo_hi_458, dataRegroupBySew_0_1_61};
  wire [31:0]       _GEN_963 = {dataRegroupBySew_5_1_61, dataRegroupBySew_4_1_61};
  wire [31:0]       dataInMem_hi_hi_650;
  assign dataInMem_hi_hi_650 = _GEN_963;
  wire [31:0]       dataInMem_hi_lo_396;
  assign dataInMem_hi_lo_396 = _GEN_963;
  wire [47:0]       dataInMem_hi_1034 = {dataInMem_hi_hi_650, dataRegroupBySew_3_1_61};
  wire [47:0]       dataInMem_lo_843 = {dataInMem_lo_hi_459, dataRegroupBySew_0_1_62};
  wire [31:0]       _GEN_964 = {dataRegroupBySew_5_1_62, dataRegroupBySew_4_1_62};
  wire [31:0]       dataInMem_hi_hi_651;
  assign dataInMem_hi_hi_651 = _GEN_964;
  wire [31:0]       dataInMem_hi_lo_397;
  assign dataInMem_hi_lo_397 = _GEN_964;
  wire [47:0]       dataInMem_hi_1035 = {dataInMem_hi_hi_651, dataRegroupBySew_3_1_62};
  wire [47:0]       dataInMem_lo_844 = {dataInMem_lo_hi_460, dataRegroupBySew_0_1_63};
  wire [31:0]       _GEN_965 = {dataRegroupBySew_5_1_63, dataRegroupBySew_4_1_63};
  wire [31:0]       dataInMem_hi_hi_652;
  assign dataInMem_hi_hi_652 = _GEN_965;
  wire [31:0]       dataInMem_hi_lo_398;
  assign dataInMem_hi_lo_398 = _GEN_965;
  wire [47:0]       dataInMem_hi_1036 = {dataInMem_hi_hi_652, dataRegroupBySew_3_1_63};
  wire [191:0]      dataInMem_lo_lo_lo_lo_lo_13 = {dataInMem_hi_974, dataInMem_lo_782, dataInMem_hi_973, dataInMem_lo_781};
  wire [191:0]      dataInMem_lo_lo_lo_lo_hi_13 = {dataInMem_hi_976, dataInMem_lo_784, dataInMem_hi_975, dataInMem_lo_783};
  wire [383:0]      dataInMem_lo_lo_lo_lo_13 = {dataInMem_lo_lo_lo_lo_hi_13, dataInMem_lo_lo_lo_lo_lo_13};
  wire [191:0]      dataInMem_lo_lo_lo_hi_lo_13 = {dataInMem_hi_978, dataInMem_lo_786, dataInMem_hi_977, dataInMem_lo_785};
  wire [191:0]      dataInMem_lo_lo_lo_hi_hi_13 = {dataInMem_hi_980, dataInMem_lo_788, dataInMem_hi_979, dataInMem_lo_787};
  wire [383:0]      dataInMem_lo_lo_lo_hi_13 = {dataInMem_lo_lo_lo_hi_hi_13, dataInMem_lo_lo_lo_hi_lo_13};
  wire [767:0]      dataInMem_lo_lo_lo_13 = {dataInMem_lo_lo_lo_hi_13, dataInMem_lo_lo_lo_lo_13};
  wire [191:0]      dataInMem_lo_lo_hi_lo_lo_13 = {dataInMem_hi_982, dataInMem_lo_790, dataInMem_hi_981, dataInMem_lo_789};
  wire [191:0]      dataInMem_lo_lo_hi_lo_hi_13 = {dataInMem_hi_984, dataInMem_lo_792, dataInMem_hi_983, dataInMem_lo_791};
  wire [383:0]      dataInMem_lo_lo_hi_lo_13 = {dataInMem_lo_lo_hi_lo_hi_13, dataInMem_lo_lo_hi_lo_lo_13};
  wire [191:0]      dataInMem_lo_lo_hi_hi_lo_13 = {dataInMem_hi_986, dataInMem_lo_794, dataInMem_hi_985, dataInMem_lo_793};
  wire [191:0]      dataInMem_lo_lo_hi_hi_hi_13 = {dataInMem_hi_988, dataInMem_lo_796, dataInMem_hi_987, dataInMem_lo_795};
  wire [383:0]      dataInMem_lo_lo_hi_hi_13 = {dataInMem_lo_lo_hi_hi_hi_13, dataInMem_lo_lo_hi_hi_lo_13};
  wire [767:0]      dataInMem_lo_lo_hi_13 = {dataInMem_lo_lo_hi_hi_13, dataInMem_lo_lo_hi_lo_13};
  wire [1535:0]     dataInMem_lo_lo_141 = {dataInMem_lo_lo_hi_13, dataInMem_lo_lo_lo_13};
  wire [191:0]      dataInMem_lo_hi_lo_lo_lo_13 = {dataInMem_hi_990, dataInMem_lo_798, dataInMem_hi_989, dataInMem_lo_797};
  wire [191:0]      dataInMem_lo_hi_lo_lo_hi_13 = {dataInMem_hi_992, dataInMem_lo_800, dataInMem_hi_991, dataInMem_lo_799};
  wire [383:0]      dataInMem_lo_hi_lo_lo_13 = {dataInMem_lo_hi_lo_lo_hi_13, dataInMem_lo_hi_lo_lo_lo_13};
  wire [191:0]      dataInMem_lo_hi_lo_hi_lo_13 = {dataInMem_hi_994, dataInMem_lo_802, dataInMem_hi_993, dataInMem_lo_801};
  wire [191:0]      dataInMem_lo_hi_lo_hi_hi_13 = {dataInMem_hi_996, dataInMem_lo_804, dataInMem_hi_995, dataInMem_lo_803};
  wire [383:0]      dataInMem_lo_hi_lo_hi_13 = {dataInMem_lo_hi_lo_hi_hi_13, dataInMem_lo_hi_lo_hi_lo_13};
  wire [767:0]      dataInMem_lo_hi_lo_13 = {dataInMem_lo_hi_lo_hi_13, dataInMem_lo_hi_lo_lo_13};
  wire [191:0]      dataInMem_lo_hi_hi_lo_lo_13 = {dataInMem_hi_998, dataInMem_lo_806, dataInMem_hi_997, dataInMem_lo_805};
  wire [191:0]      dataInMem_lo_hi_hi_lo_hi_13 = {dataInMem_hi_1000, dataInMem_lo_808, dataInMem_hi_999, dataInMem_lo_807};
  wire [383:0]      dataInMem_lo_hi_hi_lo_13 = {dataInMem_lo_hi_hi_lo_hi_13, dataInMem_lo_hi_hi_lo_lo_13};
  wire [191:0]      dataInMem_lo_hi_hi_hi_lo_13 = {dataInMem_hi_1002, dataInMem_lo_810, dataInMem_hi_1001, dataInMem_lo_809};
  wire [191:0]      dataInMem_lo_hi_hi_hi_hi_13 = {dataInMem_hi_1004, dataInMem_lo_812, dataInMem_hi_1003, dataInMem_lo_811};
  wire [383:0]      dataInMem_lo_hi_hi_hi_13 = {dataInMem_lo_hi_hi_hi_hi_13, dataInMem_lo_hi_hi_hi_lo_13};
  wire [767:0]      dataInMem_lo_hi_hi_13 = {dataInMem_lo_hi_hi_hi_13, dataInMem_lo_hi_hi_lo_13};
  wire [1535:0]     dataInMem_lo_hi_461 = {dataInMem_lo_hi_hi_13, dataInMem_lo_hi_lo_13};
  wire [3071:0]     dataInMem_lo_845 = {dataInMem_lo_hi_461, dataInMem_lo_lo_141};
  wire [191:0]      dataInMem_hi_lo_lo_lo_lo_13 = {dataInMem_hi_1006, dataInMem_lo_814, dataInMem_hi_1005, dataInMem_lo_813};
  wire [191:0]      dataInMem_hi_lo_lo_lo_hi_13 = {dataInMem_hi_1008, dataInMem_lo_816, dataInMem_hi_1007, dataInMem_lo_815};
  wire [383:0]      dataInMem_hi_lo_lo_lo_13 = {dataInMem_hi_lo_lo_lo_hi_13, dataInMem_hi_lo_lo_lo_lo_13};
  wire [191:0]      dataInMem_hi_lo_lo_hi_lo_13 = {dataInMem_hi_1010, dataInMem_lo_818, dataInMem_hi_1009, dataInMem_lo_817};
  wire [191:0]      dataInMem_hi_lo_lo_hi_hi_13 = {dataInMem_hi_1012, dataInMem_lo_820, dataInMem_hi_1011, dataInMem_lo_819};
  wire [383:0]      dataInMem_hi_lo_lo_hi_13 = {dataInMem_hi_lo_lo_hi_hi_13, dataInMem_hi_lo_lo_hi_lo_13};
  wire [767:0]      dataInMem_hi_lo_lo_13 = {dataInMem_hi_lo_lo_hi_13, dataInMem_hi_lo_lo_lo_13};
  wire [191:0]      dataInMem_hi_lo_hi_lo_lo_13 = {dataInMem_hi_1014, dataInMem_lo_822, dataInMem_hi_1013, dataInMem_lo_821};
  wire [191:0]      dataInMem_hi_lo_hi_lo_hi_13 = {dataInMem_hi_1016, dataInMem_lo_824, dataInMem_hi_1015, dataInMem_lo_823};
  wire [383:0]      dataInMem_hi_lo_hi_lo_13 = {dataInMem_hi_lo_hi_lo_hi_13, dataInMem_hi_lo_hi_lo_lo_13};
  wire [191:0]      dataInMem_hi_lo_hi_hi_lo_13 = {dataInMem_hi_1018, dataInMem_lo_826, dataInMem_hi_1017, dataInMem_lo_825};
  wire [191:0]      dataInMem_hi_lo_hi_hi_hi_13 = {dataInMem_hi_1020, dataInMem_lo_828, dataInMem_hi_1019, dataInMem_lo_827};
  wire [383:0]      dataInMem_hi_lo_hi_hi_13 = {dataInMem_hi_lo_hi_hi_hi_13, dataInMem_hi_lo_hi_hi_lo_13};
  wire [767:0]      dataInMem_hi_lo_hi_13 = {dataInMem_hi_lo_hi_hi_13, dataInMem_hi_lo_hi_lo_13};
  wire [1535:0]     dataInMem_hi_lo_269 = {dataInMem_hi_lo_hi_13, dataInMem_hi_lo_lo_13};
  wire [191:0]      dataInMem_hi_hi_lo_lo_lo_13 = {dataInMem_hi_1022, dataInMem_lo_830, dataInMem_hi_1021, dataInMem_lo_829};
  wire [191:0]      dataInMem_hi_hi_lo_lo_hi_13 = {dataInMem_hi_1024, dataInMem_lo_832, dataInMem_hi_1023, dataInMem_lo_831};
  wire [383:0]      dataInMem_hi_hi_lo_lo_13 = {dataInMem_hi_hi_lo_lo_hi_13, dataInMem_hi_hi_lo_lo_lo_13};
  wire [191:0]      dataInMem_hi_hi_lo_hi_lo_13 = {dataInMem_hi_1026, dataInMem_lo_834, dataInMem_hi_1025, dataInMem_lo_833};
  wire [191:0]      dataInMem_hi_hi_lo_hi_hi_13 = {dataInMem_hi_1028, dataInMem_lo_836, dataInMem_hi_1027, dataInMem_lo_835};
  wire [383:0]      dataInMem_hi_hi_lo_hi_13 = {dataInMem_hi_hi_lo_hi_hi_13, dataInMem_hi_hi_lo_hi_lo_13};
  wire [767:0]      dataInMem_hi_hi_lo_13 = {dataInMem_hi_hi_lo_hi_13, dataInMem_hi_hi_lo_lo_13};
  wire [191:0]      dataInMem_hi_hi_hi_lo_lo_13 = {dataInMem_hi_1030, dataInMem_lo_838, dataInMem_hi_1029, dataInMem_lo_837};
  wire [191:0]      dataInMem_hi_hi_hi_lo_hi_13 = {dataInMem_hi_1032, dataInMem_lo_840, dataInMem_hi_1031, dataInMem_lo_839};
  wire [383:0]      dataInMem_hi_hi_hi_lo_13 = {dataInMem_hi_hi_hi_lo_hi_13, dataInMem_hi_hi_hi_lo_lo_13};
  wire [191:0]      dataInMem_hi_hi_hi_hi_lo_13 = {dataInMem_hi_1034, dataInMem_lo_842, dataInMem_hi_1033, dataInMem_lo_841};
  wire [191:0]      dataInMem_hi_hi_hi_hi_hi_13 = {dataInMem_hi_1036, dataInMem_lo_844, dataInMem_hi_1035, dataInMem_lo_843};
  wire [383:0]      dataInMem_hi_hi_hi_hi_13 = {dataInMem_hi_hi_hi_hi_hi_13, dataInMem_hi_hi_hi_hi_lo_13};
  wire [767:0]      dataInMem_hi_hi_hi_13 = {dataInMem_hi_hi_hi_hi_13, dataInMem_hi_hi_hi_lo_13};
  wire [1535:0]     dataInMem_hi_hi_653 = {dataInMem_hi_hi_hi_13, dataInMem_hi_hi_lo_13};
  wire [3071:0]     dataInMem_hi_1037 = {dataInMem_hi_hi_653, dataInMem_hi_lo_269};
  wire [6143:0]     dataInMem_13 = {dataInMem_hi_1037, dataInMem_lo_845};
  wire [1023:0]     regroupCacheLine_13_0 = dataInMem_13[1023:0];
  wire [1023:0]     regroupCacheLine_13_1 = dataInMem_13[2047:1024];
  wire [1023:0]     regroupCacheLine_13_2 = dataInMem_13[3071:2048];
  wire [1023:0]     regroupCacheLine_13_3 = dataInMem_13[4095:3072];
  wire [1023:0]     regroupCacheLine_13_4 = dataInMem_13[5119:4096];
  wire [1023:0]     regroupCacheLine_13_5 = dataInMem_13[6143:5120];
  wire [1023:0]     res_104 = regroupCacheLine_13_0;
  wire [1023:0]     res_105 = regroupCacheLine_13_1;
  wire [1023:0]     res_106 = regroupCacheLine_13_2;
  wire [1023:0]     res_107 = regroupCacheLine_13_3;
  wire [1023:0]     res_108 = regroupCacheLine_13_4;
  wire [1023:0]     res_109 = regroupCacheLine_13_5;
  wire [2047:0]     lo_lo_13 = {res_105, res_104};
  wire [2047:0]     lo_hi_13 = {res_107, res_106};
  wire [4095:0]     lo_13 = {lo_hi_13, lo_lo_13};
  wire [2047:0]     hi_lo_13 = {res_109, res_108};
  wire [4095:0]     hi_13 = {2048'h0, hi_lo_13};
  wire [8191:0]     regroupLoadData_1_5 = {hi_13, lo_13};
  wire [47:0]       dataInMem_lo_846 = {dataInMem_lo_hi_462, dataRegroupBySew_0_1_0};
  wire [31:0]       dataInMem_hi_hi_654 = {dataRegroupBySew_6_1_0, dataRegroupBySew_5_1_0};
  wire [63:0]       dataInMem_hi_1038 = {dataInMem_hi_hi_654, dataInMem_hi_lo_270};
  wire [47:0]       dataInMem_lo_847 = {dataInMem_lo_hi_463, dataRegroupBySew_0_1_1};
  wire [31:0]       dataInMem_hi_hi_655 = {dataRegroupBySew_6_1_1, dataRegroupBySew_5_1_1};
  wire [63:0]       dataInMem_hi_1039 = {dataInMem_hi_hi_655, dataInMem_hi_lo_271};
  wire [47:0]       dataInMem_lo_848 = {dataInMem_lo_hi_464, dataRegroupBySew_0_1_2};
  wire [31:0]       dataInMem_hi_hi_656 = {dataRegroupBySew_6_1_2, dataRegroupBySew_5_1_2};
  wire [63:0]       dataInMem_hi_1040 = {dataInMem_hi_hi_656, dataInMem_hi_lo_272};
  wire [47:0]       dataInMem_lo_849 = {dataInMem_lo_hi_465, dataRegroupBySew_0_1_3};
  wire [31:0]       dataInMem_hi_hi_657 = {dataRegroupBySew_6_1_3, dataRegroupBySew_5_1_3};
  wire [63:0]       dataInMem_hi_1041 = {dataInMem_hi_hi_657, dataInMem_hi_lo_273};
  wire [47:0]       dataInMem_lo_850 = {dataInMem_lo_hi_466, dataRegroupBySew_0_1_4};
  wire [31:0]       dataInMem_hi_hi_658 = {dataRegroupBySew_6_1_4, dataRegroupBySew_5_1_4};
  wire [63:0]       dataInMem_hi_1042 = {dataInMem_hi_hi_658, dataInMem_hi_lo_274};
  wire [47:0]       dataInMem_lo_851 = {dataInMem_lo_hi_467, dataRegroupBySew_0_1_5};
  wire [31:0]       dataInMem_hi_hi_659 = {dataRegroupBySew_6_1_5, dataRegroupBySew_5_1_5};
  wire [63:0]       dataInMem_hi_1043 = {dataInMem_hi_hi_659, dataInMem_hi_lo_275};
  wire [47:0]       dataInMem_lo_852 = {dataInMem_lo_hi_468, dataRegroupBySew_0_1_6};
  wire [31:0]       dataInMem_hi_hi_660 = {dataRegroupBySew_6_1_6, dataRegroupBySew_5_1_6};
  wire [63:0]       dataInMem_hi_1044 = {dataInMem_hi_hi_660, dataInMem_hi_lo_276};
  wire [47:0]       dataInMem_lo_853 = {dataInMem_lo_hi_469, dataRegroupBySew_0_1_7};
  wire [31:0]       dataInMem_hi_hi_661 = {dataRegroupBySew_6_1_7, dataRegroupBySew_5_1_7};
  wire [63:0]       dataInMem_hi_1045 = {dataInMem_hi_hi_661, dataInMem_hi_lo_277};
  wire [47:0]       dataInMem_lo_854 = {dataInMem_lo_hi_470, dataRegroupBySew_0_1_8};
  wire [31:0]       dataInMem_hi_hi_662 = {dataRegroupBySew_6_1_8, dataRegroupBySew_5_1_8};
  wire [63:0]       dataInMem_hi_1046 = {dataInMem_hi_hi_662, dataInMem_hi_lo_278};
  wire [47:0]       dataInMem_lo_855 = {dataInMem_lo_hi_471, dataRegroupBySew_0_1_9};
  wire [31:0]       dataInMem_hi_hi_663 = {dataRegroupBySew_6_1_9, dataRegroupBySew_5_1_9};
  wire [63:0]       dataInMem_hi_1047 = {dataInMem_hi_hi_663, dataInMem_hi_lo_279};
  wire [47:0]       dataInMem_lo_856 = {dataInMem_lo_hi_472, dataRegroupBySew_0_1_10};
  wire [31:0]       dataInMem_hi_hi_664 = {dataRegroupBySew_6_1_10, dataRegroupBySew_5_1_10};
  wire [63:0]       dataInMem_hi_1048 = {dataInMem_hi_hi_664, dataInMem_hi_lo_280};
  wire [47:0]       dataInMem_lo_857 = {dataInMem_lo_hi_473, dataRegroupBySew_0_1_11};
  wire [31:0]       dataInMem_hi_hi_665 = {dataRegroupBySew_6_1_11, dataRegroupBySew_5_1_11};
  wire [63:0]       dataInMem_hi_1049 = {dataInMem_hi_hi_665, dataInMem_hi_lo_281};
  wire [47:0]       dataInMem_lo_858 = {dataInMem_lo_hi_474, dataRegroupBySew_0_1_12};
  wire [31:0]       dataInMem_hi_hi_666 = {dataRegroupBySew_6_1_12, dataRegroupBySew_5_1_12};
  wire [63:0]       dataInMem_hi_1050 = {dataInMem_hi_hi_666, dataInMem_hi_lo_282};
  wire [47:0]       dataInMem_lo_859 = {dataInMem_lo_hi_475, dataRegroupBySew_0_1_13};
  wire [31:0]       dataInMem_hi_hi_667 = {dataRegroupBySew_6_1_13, dataRegroupBySew_5_1_13};
  wire [63:0]       dataInMem_hi_1051 = {dataInMem_hi_hi_667, dataInMem_hi_lo_283};
  wire [47:0]       dataInMem_lo_860 = {dataInMem_lo_hi_476, dataRegroupBySew_0_1_14};
  wire [31:0]       dataInMem_hi_hi_668 = {dataRegroupBySew_6_1_14, dataRegroupBySew_5_1_14};
  wire [63:0]       dataInMem_hi_1052 = {dataInMem_hi_hi_668, dataInMem_hi_lo_284};
  wire [47:0]       dataInMem_lo_861 = {dataInMem_lo_hi_477, dataRegroupBySew_0_1_15};
  wire [31:0]       dataInMem_hi_hi_669 = {dataRegroupBySew_6_1_15, dataRegroupBySew_5_1_15};
  wire [63:0]       dataInMem_hi_1053 = {dataInMem_hi_hi_669, dataInMem_hi_lo_285};
  wire [47:0]       dataInMem_lo_862 = {dataInMem_lo_hi_478, dataRegroupBySew_0_1_16};
  wire [31:0]       dataInMem_hi_hi_670 = {dataRegroupBySew_6_1_16, dataRegroupBySew_5_1_16};
  wire [63:0]       dataInMem_hi_1054 = {dataInMem_hi_hi_670, dataInMem_hi_lo_286};
  wire [47:0]       dataInMem_lo_863 = {dataInMem_lo_hi_479, dataRegroupBySew_0_1_17};
  wire [31:0]       dataInMem_hi_hi_671 = {dataRegroupBySew_6_1_17, dataRegroupBySew_5_1_17};
  wire [63:0]       dataInMem_hi_1055 = {dataInMem_hi_hi_671, dataInMem_hi_lo_287};
  wire [47:0]       dataInMem_lo_864 = {dataInMem_lo_hi_480, dataRegroupBySew_0_1_18};
  wire [31:0]       dataInMem_hi_hi_672 = {dataRegroupBySew_6_1_18, dataRegroupBySew_5_1_18};
  wire [63:0]       dataInMem_hi_1056 = {dataInMem_hi_hi_672, dataInMem_hi_lo_288};
  wire [47:0]       dataInMem_lo_865 = {dataInMem_lo_hi_481, dataRegroupBySew_0_1_19};
  wire [31:0]       dataInMem_hi_hi_673 = {dataRegroupBySew_6_1_19, dataRegroupBySew_5_1_19};
  wire [63:0]       dataInMem_hi_1057 = {dataInMem_hi_hi_673, dataInMem_hi_lo_289};
  wire [47:0]       dataInMem_lo_866 = {dataInMem_lo_hi_482, dataRegroupBySew_0_1_20};
  wire [31:0]       dataInMem_hi_hi_674 = {dataRegroupBySew_6_1_20, dataRegroupBySew_5_1_20};
  wire [63:0]       dataInMem_hi_1058 = {dataInMem_hi_hi_674, dataInMem_hi_lo_290};
  wire [47:0]       dataInMem_lo_867 = {dataInMem_lo_hi_483, dataRegroupBySew_0_1_21};
  wire [31:0]       dataInMem_hi_hi_675 = {dataRegroupBySew_6_1_21, dataRegroupBySew_5_1_21};
  wire [63:0]       dataInMem_hi_1059 = {dataInMem_hi_hi_675, dataInMem_hi_lo_291};
  wire [47:0]       dataInMem_lo_868 = {dataInMem_lo_hi_484, dataRegroupBySew_0_1_22};
  wire [31:0]       dataInMem_hi_hi_676 = {dataRegroupBySew_6_1_22, dataRegroupBySew_5_1_22};
  wire [63:0]       dataInMem_hi_1060 = {dataInMem_hi_hi_676, dataInMem_hi_lo_292};
  wire [47:0]       dataInMem_lo_869 = {dataInMem_lo_hi_485, dataRegroupBySew_0_1_23};
  wire [31:0]       dataInMem_hi_hi_677 = {dataRegroupBySew_6_1_23, dataRegroupBySew_5_1_23};
  wire [63:0]       dataInMem_hi_1061 = {dataInMem_hi_hi_677, dataInMem_hi_lo_293};
  wire [47:0]       dataInMem_lo_870 = {dataInMem_lo_hi_486, dataRegroupBySew_0_1_24};
  wire [31:0]       dataInMem_hi_hi_678 = {dataRegroupBySew_6_1_24, dataRegroupBySew_5_1_24};
  wire [63:0]       dataInMem_hi_1062 = {dataInMem_hi_hi_678, dataInMem_hi_lo_294};
  wire [47:0]       dataInMem_lo_871 = {dataInMem_lo_hi_487, dataRegroupBySew_0_1_25};
  wire [31:0]       dataInMem_hi_hi_679 = {dataRegroupBySew_6_1_25, dataRegroupBySew_5_1_25};
  wire [63:0]       dataInMem_hi_1063 = {dataInMem_hi_hi_679, dataInMem_hi_lo_295};
  wire [47:0]       dataInMem_lo_872 = {dataInMem_lo_hi_488, dataRegroupBySew_0_1_26};
  wire [31:0]       dataInMem_hi_hi_680 = {dataRegroupBySew_6_1_26, dataRegroupBySew_5_1_26};
  wire [63:0]       dataInMem_hi_1064 = {dataInMem_hi_hi_680, dataInMem_hi_lo_296};
  wire [47:0]       dataInMem_lo_873 = {dataInMem_lo_hi_489, dataRegroupBySew_0_1_27};
  wire [31:0]       dataInMem_hi_hi_681 = {dataRegroupBySew_6_1_27, dataRegroupBySew_5_1_27};
  wire [63:0]       dataInMem_hi_1065 = {dataInMem_hi_hi_681, dataInMem_hi_lo_297};
  wire [47:0]       dataInMem_lo_874 = {dataInMem_lo_hi_490, dataRegroupBySew_0_1_28};
  wire [31:0]       dataInMem_hi_hi_682 = {dataRegroupBySew_6_1_28, dataRegroupBySew_5_1_28};
  wire [63:0]       dataInMem_hi_1066 = {dataInMem_hi_hi_682, dataInMem_hi_lo_298};
  wire [47:0]       dataInMem_lo_875 = {dataInMem_lo_hi_491, dataRegroupBySew_0_1_29};
  wire [31:0]       dataInMem_hi_hi_683 = {dataRegroupBySew_6_1_29, dataRegroupBySew_5_1_29};
  wire [63:0]       dataInMem_hi_1067 = {dataInMem_hi_hi_683, dataInMem_hi_lo_299};
  wire [47:0]       dataInMem_lo_876 = {dataInMem_lo_hi_492, dataRegroupBySew_0_1_30};
  wire [31:0]       dataInMem_hi_hi_684 = {dataRegroupBySew_6_1_30, dataRegroupBySew_5_1_30};
  wire [63:0]       dataInMem_hi_1068 = {dataInMem_hi_hi_684, dataInMem_hi_lo_300};
  wire [47:0]       dataInMem_lo_877 = {dataInMem_lo_hi_493, dataRegroupBySew_0_1_31};
  wire [31:0]       dataInMem_hi_hi_685 = {dataRegroupBySew_6_1_31, dataRegroupBySew_5_1_31};
  wire [63:0]       dataInMem_hi_1069 = {dataInMem_hi_hi_685, dataInMem_hi_lo_301};
  wire [47:0]       dataInMem_lo_878 = {dataInMem_lo_hi_494, dataRegroupBySew_0_1_32};
  wire [31:0]       dataInMem_hi_hi_686 = {dataRegroupBySew_6_1_32, dataRegroupBySew_5_1_32};
  wire [63:0]       dataInMem_hi_1070 = {dataInMem_hi_hi_686, dataInMem_hi_lo_302};
  wire [47:0]       dataInMem_lo_879 = {dataInMem_lo_hi_495, dataRegroupBySew_0_1_33};
  wire [31:0]       dataInMem_hi_hi_687 = {dataRegroupBySew_6_1_33, dataRegroupBySew_5_1_33};
  wire [63:0]       dataInMem_hi_1071 = {dataInMem_hi_hi_687, dataInMem_hi_lo_303};
  wire [47:0]       dataInMem_lo_880 = {dataInMem_lo_hi_496, dataRegroupBySew_0_1_34};
  wire [31:0]       dataInMem_hi_hi_688 = {dataRegroupBySew_6_1_34, dataRegroupBySew_5_1_34};
  wire [63:0]       dataInMem_hi_1072 = {dataInMem_hi_hi_688, dataInMem_hi_lo_304};
  wire [47:0]       dataInMem_lo_881 = {dataInMem_lo_hi_497, dataRegroupBySew_0_1_35};
  wire [31:0]       dataInMem_hi_hi_689 = {dataRegroupBySew_6_1_35, dataRegroupBySew_5_1_35};
  wire [63:0]       dataInMem_hi_1073 = {dataInMem_hi_hi_689, dataInMem_hi_lo_305};
  wire [47:0]       dataInMem_lo_882 = {dataInMem_lo_hi_498, dataRegroupBySew_0_1_36};
  wire [31:0]       dataInMem_hi_hi_690 = {dataRegroupBySew_6_1_36, dataRegroupBySew_5_1_36};
  wire [63:0]       dataInMem_hi_1074 = {dataInMem_hi_hi_690, dataInMem_hi_lo_306};
  wire [47:0]       dataInMem_lo_883 = {dataInMem_lo_hi_499, dataRegroupBySew_0_1_37};
  wire [31:0]       dataInMem_hi_hi_691 = {dataRegroupBySew_6_1_37, dataRegroupBySew_5_1_37};
  wire [63:0]       dataInMem_hi_1075 = {dataInMem_hi_hi_691, dataInMem_hi_lo_307};
  wire [47:0]       dataInMem_lo_884 = {dataInMem_lo_hi_500, dataRegroupBySew_0_1_38};
  wire [31:0]       dataInMem_hi_hi_692 = {dataRegroupBySew_6_1_38, dataRegroupBySew_5_1_38};
  wire [63:0]       dataInMem_hi_1076 = {dataInMem_hi_hi_692, dataInMem_hi_lo_308};
  wire [47:0]       dataInMem_lo_885 = {dataInMem_lo_hi_501, dataRegroupBySew_0_1_39};
  wire [31:0]       dataInMem_hi_hi_693 = {dataRegroupBySew_6_1_39, dataRegroupBySew_5_1_39};
  wire [63:0]       dataInMem_hi_1077 = {dataInMem_hi_hi_693, dataInMem_hi_lo_309};
  wire [47:0]       dataInMem_lo_886 = {dataInMem_lo_hi_502, dataRegroupBySew_0_1_40};
  wire [31:0]       dataInMem_hi_hi_694 = {dataRegroupBySew_6_1_40, dataRegroupBySew_5_1_40};
  wire [63:0]       dataInMem_hi_1078 = {dataInMem_hi_hi_694, dataInMem_hi_lo_310};
  wire [47:0]       dataInMem_lo_887 = {dataInMem_lo_hi_503, dataRegroupBySew_0_1_41};
  wire [31:0]       dataInMem_hi_hi_695 = {dataRegroupBySew_6_1_41, dataRegroupBySew_5_1_41};
  wire [63:0]       dataInMem_hi_1079 = {dataInMem_hi_hi_695, dataInMem_hi_lo_311};
  wire [47:0]       dataInMem_lo_888 = {dataInMem_lo_hi_504, dataRegroupBySew_0_1_42};
  wire [31:0]       dataInMem_hi_hi_696 = {dataRegroupBySew_6_1_42, dataRegroupBySew_5_1_42};
  wire [63:0]       dataInMem_hi_1080 = {dataInMem_hi_hi_696, dataInMem_hi_lo_312};
  wire [47:0]       dataInMem_lo_889 = {dataInMem_lo_hi_505, dataRegroupBySew_0_1_43};
  wire [31:0]       dataInMem_hi_hi_697 = {dataRegroupBySew_6_1_43, dataRegroupBySew_5_1_43};
  wire [63:0]       dataInMem_hi_1081 = {dataInMem_hi_hi_697, dataInMem_hi_lo_313};
  wire [47:0]       dataInMem_lo_890 = {dataInMem_lo_hi_506, dataRegroupBySew_0_1_44};
  wire [31:0]       dataInMem_hi_hi_698 = {dataRegroupBySew_6_1_44, dataRegroupBySew_5_1_44};
  wire [63:0]       dataInMem_hi_1082 = {dataInMem_hi_hi_698, dataInMem_hi_lo_314};
  wire [47:0]       dataInMem_lo_891 = {dataInMem_lo_hi_507, dataRegroupBySew_0_1_45};
  wire [31:0]       dataInMem_hi_hi_699 = {dataRegroupBySew_6_1_45, dataRegroupBySew_5_1_45};
  wire [63:0]       dataInMem_hi_1083 = {dataInMem_hi_hi_699, dataInMem_hi_lo_315};
  wire [47:0]       dataInMem_lo_892 = {dataInMem_lo_hi_508, dataRegroupBySew_0_1_46};
  wire [31:0]       dataInMem_hi_hi_700 = {dataRegroupBySew_6_1_46, dataRegroupBySew_5_1_46};
  wire [63:0]       dataInMem_hi_1084 = {dataInMem_hi_hi_700, dataInMem_hi_lo_316};
  wire [47:0]       dataInMem_lo_893 = {dataInMem_lo_hi_509, dataRegroupBySew_0_1_47};
  wire [31:0]       dataInMem_hi_hi_701 = {dataRegroupBySew_6_1_47, dataRegroupBySew_5_1_47};
  wire [63:0]       dataInMem_hi_1085 = {dataInMem_hi_hi_701, dataInMem_hi_lo_317};
  wire [47:0]       dataInMem_lo_894 = {dataInMem_lo_hi_510, dataRegroupBySew_0_1_48};
  wire [31:0]       dataInMem_hi_hi_702 = {dataRegroupBySew_6_1_48, dataRegroupBySew_5_1_48};
  wire [63:0]       dataInMem_hi_1086 = {dataInMem_hi_hi_702, dataInMem_hi_lo_318};
  wire [47:0]       dataInMem_lo_895 = {dataInMem_lo_hi_511, dataRegroupBySew_0_1_49};
  wire [31:0]       dataInMem_hi_hi_703 = {dataRegroupBySew_6_1_49, dataRegroupBySew_5_1_49};
  wire [63:0]       dataInMem_hi_1087 = {dataInMem_hi_hi_703, dataInMem_hi_lo_319};
  wire [47:0]       dataInMem_lo_896 = {dataInMem_lo_hi_512, dataRegroupBySew_0_1_50};
  wire [31:0]       dataInMem_hi_hi_704 = {dataRegroupBySew_6_1_50, dataRegroupBySew_5_1_50};
  wire [63:0]       dataInMem_hi_1088 = {dataInMem_hi_hi_704, dataInMem_hi_lo_320};
  wire [47:0]       dataInMem_lo_897 = {dataInMem_lo_hi_513, dataRegroupBySew_0_1_51};
  wire [31:0]       dataInMem_hi_hi_705 = {dataRegroupBySew_6_1_51, dataRegroupBySew_5_1_51};
  wire [63:0]       dataInMem_hi_1089 = {dataInMem_hi_hi_705, dataInMem_hi_lo_321};
  wire [47:0]       dataInMem_lo_898 = {dataInMem_lo_hi_514, dataRegroupBySew_0_1_52};
  wire [31:0]       dataInMem_hi_hi_706 = {dataRegroupBySew_6_1_52, dataRegroupBySew_5_1_52};
  wire [63:0]       dataInMem_hi_1090 = {dataInMem_hi_hi_706, dataInMem_hi_lo_322};
  wire [47:0]       dataInMem_lo_899 = {dataInMem_lo_hi_515, dataRegroupBySew_0_1_53};
  wire [31:0]       dataInMem_hi_hi_707 = {dataRegroupBySew_6_1_53, dataRegroupBySew_5_1_53};
  wire [63:0]       dataInMem_hi_1091 = {dataInMem_hi_hi_707, dataInMem_hi_lo_323};
  wire [47:0]       dataInMem_lo_900 = {dataInMem_lo_hi_516, dataRegroupBySew_0_1_54};
  wire [31:0]       dataInMem_hi_hi_708 = {dataRegroupBySew_6_1_54, dataRegroupBySew_5_1_54};
  wire [63:0]       dataInMem_hi_1092 = {dataInMem_hi_hi_708, dataInMem_hi_lo_324};
  wire [47:0]       dataInMem_lo_901 = {dataInMem_lo_hi_517, dataRegroupBySew_0_1_55};
  wire [31:0]       dataInMem_hi_hi_709 = {dataRegroupBySew_6_1_55, dataRegroupBySew_5_1_55};
  wire [63:0]       dataInMem_hi_1093 = {dataInMem_hi_hi_709, dataInMem_hi_lo_325};
  wire [47:0]       dataInMem_lo_902 = {dataInMem_lo_hi_518, dataRegroupBySew_0_1_56};
  wire [31:0]       dataInMem_hi_hi_710 = {dataRegroupBySew_6_1_56, dataRegroupBySew_5_1_56};
  wire [63:0]       dataInMem_hi_1094 = {dataInMem_hi_hi_710, dataInMem_hi_lo_326};
  wire [47:0]       dataInMem_lo_903 = {dataInMem_lo_hi_519, dataRegroupBySew_0_1_57};
  wire [31:0]       dataInMem_hi_hi_711 = {dataRegroupBySew_6_1_57, dataRegroupBySew_5_1_57};
  wire [63:0]       dataInMem_hi_1095 = {dataInMem_hi_hi_711, dataInMem_hi_lo_327};
  wire [47:0]       dataInMem_lo_904 = {dataInMem_lo_hi_520, dataRegroupBySew_0_1_58};
  wire [31:0]       dataInMem_hi_hi_712 = {dataRegroupBySew_6_1_58, dataRegroupBySew_5_1_58};
  wire [63:0]       dataInMem_hi_1096 = {dataInMem_hi_hi_712, dataInMem_hi_lo_328};
  wire [47:0]       dataInMem_lo_905 = {dataInMem_lo_hi_521, dataRegroupBySew_0_1_59};
  wire [31:0]       dataInMem_hi_hi_713 = {dataRegroupBySew_6_1_59, dataRegroupBySew_5_1_59};
  wire [63:0]       dataInMem_hi_1097 = {dataInMem_hi_hi_713, dataInMem_hi_lo_329};
  wire [47:0]       dataInMem_lo_906 = {dataInMem_lo_hi_522, dataRegroupBySew_0_1_60};
  wire [31:0]       dataInMem_hi_hi_714 = {dataRegroupBySew_6_1_60, dataRegroupBySew_5_1_60};
  wire [63:0]       dataInMem_hi_1098 = {dataInMem_hi_hi_714, dataInMem_hi_lo_330};
  wire [47:0]       dataInMem_lo_907 = {dataInMem_lo_hi_523, dataRegroupBySew_0_1_61};
  wire [31:0]       dataInMem_hi_hi_715 = {dataRegroupBySew_6_1_61, dataRegroupBySew_5_1_61};
  wire [63:0]       dataInMem_hi_1099 = {dataInMem_hi_hi_715, dataInMem_hi_lo_331};
  wire [47:0]       dataInMem_lo_908 = {dataInMem_lo_hi_524, dataRegroupBySew_0_1_62};
  wire [31:0]       dataInMem_hi_hi_716 = {dataRegroupBySew_6_1_62, dataRegroupBySew_5_1_62};
  wire [63:0]       dataInMem_hi_1100 = {dataInMem_hi_hi_716, dataInMem_hi_lo_332};
  wire [47:0]       dataInMem_lo_909 = {dataInMem_lo_hi_525, dataRegroupBySew_0_1_63};
  wire [31:0]       dataInMem_hi_hi_717 = {dataRegroupBySew_6_1_63, dataRegroupBySew_5_1_63};
  wire [63:0]       dataInMem_hi_1101 = {dataInMem_hi_hi_717, dataInMem_hi_lo_333};
  wire [223:0]      dataInMem_lo_lo_lo_lo_lo_14 = {dataInMem_hi_1039, dataInMem_lo_847, dataInMem_hi_1038, dataInMem_lo_846};
  wire [223:0]      dataInMem_lo_lo_lo_lo_hi_14 = {dataInMem_hi_1041, dataInMem_lo_849, dataInMem_hi_1040, dataInMem_lo_848};
  wire [447:0]      dataInMem_lo_lo_lo_lo_14 = {dataInMem_lo_lo_lo_lo_hi_14, dataInMem_lo_lo_lo_lo_lo_14};
  wire [223:0]      dataInMem_lo_lo_lo_hi_lo_14 = {dataInMem_hi_1043, dataInMem_lo_851, dataInMem_hi_1042, dataInMem_lo_850};
  wire [223:0]      dataInMem_lo_lo_lo_hi_hi_14 = {dataInMem_hi_1045, dataInMem_lo_853, dataInMem_hi_1044, dataInMem_lo_852};
  wire [447:0]      dataInMem_lo_lo_lo_hi_14 = {dataInMem_lo_lo_lo_hi_hi_14, dataInMem_lo_lo_lo_hi_lo_14};
  wire [895:0]      dataInMem_lo_lo_lo_14 = {dataInMem_lo_lo_lo_hi_14, dataInMem_lo_lo_lo_lo_14};
  wire [223:0]      dataInMem_lo_lo_hi_lo_lo_14 = {dataInMem_hi_1047, dataInMem_lo_855, dataInMem_hi_1046, dataInMem_lo_854};
  wire [223:0]      dataInMem_lo_lo_hi_lo_hi_14 = {dataInMem_hi_1049, dataInMem_lo_857, dataInMem_hi_1048, dataInMem_lo_856};
  wire [447:0]      dataInMem_lo_lo_hi_lo_14 = {dataInMem_lo_lo_hi_lo_hi_14, dataInMem_lo_lo_hi_lo_lo_14};
  wire [223:0]      dataInMem_lo_lo_hi_hi_lo_14 = {dataInMem_hi_1051, dataInMem_lo_859, dataInMem_hi_1050, dataInMem_lo_858};
  wire [223:0]      dataInMem_lo_lo_hi_hi_hi_14 = {dataInMem_hi_1053, dataInMem_lo_861, dataInMem_hi_1052, dataInMem_lo_860};
  wire [447:0]      dataInMem_lo_lo_hi_hi_14 = {dataInMem_lo_lo_hi_hi_hi_14, dataInMem_lo_lo_hi_hi_lo_14};
  wire [895:0]      dataInMem_lo_lo_hi_14 = {dataInMem_lo_lo_hi_hi_14, dataInMem_lo_lo_hi_lo_14};
  wire [1791:0]     dataInMem_lo_lo_142 = {dataInMem_lo_lo_hi_14, dataInMem_lo_lo_lo_14};
  wire [223:0]      dataInMem_lo_hi_lo_lo_lo_14 = {dataInMem_hi_1055, dataInMem_lo_863, dataInMem_hi_1054, dataInMem_lo_862};
  wire [223:0]      dataInMem_lo_hi_lo_lo_hi_14 = {dataInMem_hi_1057, dataInMem_lo_865, dataInMem_hi_1056, dataInMem_lo_864};
  wire [447:0]      dataInMem_lo_hi_lo_lo_14 = {dataInMem_lo_hi_lo_lo_hi_14, dataInMem_lo_hi_lo_lo_lo_14};
  wire [223:0]      dataInMem_lo_hi_lo_hi_lo_14 = {dataInMem_hi_1059, dataInMem_lo_867, dataInMem_hi_1058, dataInMem_lo_866};
  wire [223:0]      dataInMem_lo_hi_lo_hi_hi_14 = {dataInMem_hi_1061, dataInMem_lo_869, dataInMem_hi_1060, dataInMem_lo_868};
  wire [447:0]      dataInMem_lo_hi_lo_hi_14 = {dataInMem_lo_hi_lo_hi_hi_14, dataInMem_lo_hi_lo_hi_lo_14};
  wire [895:0]      dataInMem_lo_hi_lo_14 = {dataInMem_lo_hi_lo_hi_14, dataInMem_lo_hi_lo_lo_14};
  wire [223:0]      dataInMem_lo_hi_hi_lo_lo_14 = {dataInMem_hi_1063, dataInMem_lo_871, dataInMem_hi_1062, dataInMem_lo_870};
  wire [223:0]      dataInMem_lo_hi_hi_lo_hi_14 = {dataInMem_hi_1065, dataInMem_lo_873, dataInMem_hi_1064, dataInMem_lo_872};
  wire [447:0]      dataInMem_lo_hi_hi_lo_14 = {dataInMem_lo_hi_hi_lo_hi_14, dataInMem_lo_hi_hi_lo_lo_14};
  wire [223:0]      dataInMem_lo_hi_hi_hi_lo_14 = {dataInMem_hi_1067, dataInMem_lo_875, dataInMem_hi_1066, dataInMem_lo_874};
  wire [223:0]      dataInMem_lo_hi_hi_hi_hi_14 = {dataInMem_hi_1069, dataInMem_lo_877, dataInMem_hi_1068, dataInMem_lo_876};
  wire [447:0]      dataInMem_lo_hi_hi_hi_14 = {dataInMem_lo_hi_hi_hi_hi_14, dataInMem_lo_hi_hi_hi_lo_14};
  wire [895:0]      dataInMem_lo_hi_hi_14 = {dataInMem_lo_hi_hi_hi_14, dataInMem_lo_hi_hi_lo_14};
  wire [1791:0]     dataInMem_lo_hi_526 = {dataInMem_lo_hi_hi_14, dataInMem_lo_hi_lo_14};
  wire [3583:0]     dataInMem_lo_910 = {dataInMem_lo_hi_526, dataInMem_lo_lo_142};
  wire [223:0]      dataInMem_hi_lo_lo_lo_lo_14 = {dataInMem_hi_1071, dataInMem_lo_879, dataInMem_hi_1070, dataInMem_lo_878};
  wire [223:0]      dataInMem_hi_lo_lo_lo_hi_14 = {dataInMem_hi_1073, dataInMem_lo_881, dataInMem_hi_1072, dataInMem_lo_880};
  wire [447:0]      dataInMem_hi_lo_lo_lo_14 = {dataInMem_hi_lo_lo_lo_hi_14, dataInMem_hi_lo_lo_lo_lo_14};
  wire [223:0]      dataInMem_hi_lo_lo_hi_lo_14 = {dataInMem_hi_1075, dataInMem_lo_883, dataInMem_hi_1074, dataInMem_lo_882};
  wire [223:0]      dataInMem_hi_lo_lo_hi_hi_14 = {dataInMem_hi_1077, dataInMem_lo_885, dataInMem_hi_1076, dataInMem_lo_884};
  wire [447:0]      dataInMem_hi_lo_lo_hi_14 = {dataInMem_hi_lo_lo_hi_hi_14, dataInMem_hi_lo_lo_hi_lo_14};
  wire [895:0]      dataInMem_hi_lo_lo_14 = {dataInMem_hi_lo_lo_hi_14, dataInMem_hi_lo_lo_lo_14};
  wire [223:0]      dataInMem_hi_lo_hi_lo_lo_14 = {dataInMem_hi_1079, dataInMem_lo_887, dataInMem_hi_1078, dataInMem_lo_886};
  wire [223:0]      dataInMem_hi_lo_hi_lo_hi_14 = {dataInMem_hi_1081, dataInMem_lo_889, dataInMem_hi_1080, dataInMem_lo_888};
  wire [447:0]      dataInMem_hi_lo_hi_lo_14 = {dataInMem_hi_lo_hi_lo_hi_14, dataInMem_hi_lo_hi_lo_lo_14};
  wire [223:0]      dataInMem_hi_lo_hi_hi_lo_14 = {dataInMem_hi_1083, dataInMem_lo_891, dataInMem_hi_1082, dataInMem_lo_890};
  wire [223:0]      dataInMem_hi_lo_hi_hi_hi_14 = {dataInMem_hi_1085, dataInMem_lo_893, dataInMem_hi_1084, dataInMem_lo_892};
  wire [447:0]      dataInMem_hi_lo_hi_hi_14 = {dataInMem_hi_lo_hi_hi_hi_14, dataInMem_hi_lo_hi_hi_lo_14};
  wire [895:0]      dataInMem_hi_lo_hi_14 = {dataInMem_hi_lo_hi_hi_14, dataInMem_hi_lo_hi_lo_14};
  wire [1791:0]     dataInMem_hi_lo_334 = {dataInMem_hi_lo_hi_14, dataInMem_hi_lo_lo_14};
  wire [223:0]      dataInMem_hi_hi_lo_lo_lo_14 = {dataInMem_hi_1087, dataInMem_lo_895, dataInMem_hi_1086, dataInMem_lo_894};
  wire [223:0]      dataInMem_hi_hi_lo_lo_hi_14 = {dataInMem_hi_1089, dataInMem_lo_897, dataInMem_hi_1088, dataInMem_lo_896};
  wire [447:0]      dataInMem_hi_hi_lo_lo_14 = {dataInMem_hi_hi_lo_lo_hi_14, dataInMem_hi_hi_lo_lo_lo_14};
  wire [223:0]      dataInMem_hi_hi_lo_hi_lo_14 = {dataInMem_hi_1091, dataInMem_lo_899, dataInMem_hi_1090, dataInMem_lo_898};
  wire [223:0]      dataInMem_hi_hi_lo_hi_hi_14 = {dataInMem_hi_1093, dataInMem_lo_901, dataInMem_hi_1092, dataInMem_lo_900};
  wire [447:0]      dataInMem_hi_hi_lo_hi_14 = {dataInMem_hi_hi_lo_hi_hi_14, dataInMem_hi_hi_lo_hi_lo_14};
  wire [895:0]      dataInMem_hi_hi_lo_14 = {dataInMem_hi_hi_lo_hi_14, dataInMem_hi_hi_lo_lo_14};
  wire [223:0]      dataInMem_hi_hi_hi_lo_lo_14 = {dataInMem_hi_1095, dataInMem_lo_903, dataInMem_hi_1094, dataInMem_lo_902};
  wire [223:0]      dataInMem_hi_hi_hi_lo_hi_14 = {dataInMem_hi_1097, dataInMem_lo_905, dataInMem_hi_1096, dataInMem_lo_904};
  wire [447:0]      dataInMem_hi_hi_hi_lo_14 = {dataInMem_hi_hi_hi_lo_hi_14, dataInMem_hi_hi_hi_lo_lo_14};
  wire [223:0]      dataInMem_hi_hi_hi_hi_lo_14 = {dataInMem_hi_1099, dataInMem_lo_907, dataInMem_hi_1098, dataInMem_lo_906};
  wire [223:0]      dataInMem_hi_hi_hi_hi_hi_14 = {dataInMem_hi_1101, dataInMem_lo_909, dataInMem_hi_1100, dataInMem_lo_908};
  wire [447:0]      dataInMem_hi_hi_hi_hi_14 = {dataInMem_hi_hi_hi_hi_hi_14, dataInMem_hi_hi_hi_hi_lo_14};
  wire [895:0]      dataInMem_hi_hi_hi_14 = {dataInMem_hi_hi_hi_hi_14, dataInMem_hi_hi_hi_lo_14};
  wire [1791:0]     dataInMem_hi_hi_718 = {dataInMem_hi_hi_hi_14, dataInMem_hi_hi_lo_14};
  wire [3583:0]     dataInMem_hi_1102 = {dataInMem_hi_hi_718, dataInMem_hi_lo_334};
  wire [7167:0]     dataInMem_14 = {dataInMem_hi_1102, dataInMem_lo_910};
  wire [1023:0]     regroupCacheLine_14_0 = dataInMem_14[1023:0];
  wire [1023:0]     regroupCacheLine_14_1 = dataInMem_14[2047:1024];
  wire [1023:0]     regroupCacheLine_14_2 = dataInMem_14[3071:2048];
  wire [1023:0]     regroupCacheLine_14_3 = dataInMem_14[4095:3072];
  wire [1023:0]     regroupCacheLine_14_4 = dataInMem_14[5119:4096];
  wire [1023:0]     regroupCacheLine_14_5 = dataInMem_14[6143:5120];
  wire [1023:0]     regroupCacheLine_14_6 = dataInMem_14[7167:6144];
  wire [1023:0]     res_112 = regroupCacheLine_14_0;
  wire [1023:0]     res_113 = regroupCacheLine_14_1;
  wire [1023:0]     res_114 = regroupCacheLine_14_2;
  wire [1023:0]     res_115 = regroupCacheLine_14_3;
  wire [1023:0]     res_116 = regroupCacheLine_14_4;
  wire [1023:0]     res_117 = regroupCacheLine_14_5;
  wire [1023:0]     res_118 = regroupCacheLine_14_6;
  wire [2047:0]     lo_lo_14 = {res_113, res_112};
  wire [2047:0]     lo_hi_14 = {res_115, res_114};
  wire [4095:0]     lo_14 = {lo_hi_14, lo_lo_14};
  wire [2047:0]     hi_lo_14 = {res_117, res_116};
  wire [2047:0]     hi_hi_14 = {1024'h0, res_118};
  wire [4095:0]     hi_14 = {hi_hi_14, hi_lo_14};
  wire [8191:0]     regroupLoadData_1_6 = {hi_14, lo_14};
  wire [63:0]       dataInMem_lo_911 = {dataInMem_lo_hi_527, dataInMem_lo_lo_143};
  wire [31:0]       dataInMem_hi_hi_719 = {dataRegroupBySew_7_1_0, dataRegroupBySew_6_1_0};
  wire [63:0]       dataInMem_hi_1103 = {dataInMem_hi_hi_719, dataInMem_hi_lo_335};
  wire [63:0]       dataInMem_lo_912 = {dataInMem_lo_hi_528, dataInMem_lo_lo_144};
  wire [31:0]       dataInMem_hi_hi_720 = {dataRegroupBySew_7_1_1, dataRegroupBySew_6_1_1};
  wire [63:0]       dataInMem_hi_1104 = {dataInMem_hi_hi_720, dataInMem_hi_lo_336};
  wire [63:0]       dataInMem_lo_913 = {dataInMem_lo_hi_529, dataInMem_lo_lo_145};
  wire [31:0]       dataInMem_hi_hi_721 = {dataRegroupBySew_7_1_2, dataRegroupBySew_6_1_2};
  wire [63:0]       dataInMem_hi_1105 = {dataInMem_hi_hi_721, dataInMem_hi_lo_337};
  wire [63:0]       dataInMem_lo_914 = {dataInMem_lo_hi_530, dataInMem_lo_lo_146};
  wire [31:0]       dataInMem_hi_hi_722 = {dataRegroupBySew_7_1_3, dataRegroupBySew_6_1_3};
  wire [63:0]       dataInMem_hi_1106 = {dataInMem_hi_hi_722, dataInMem_hi_lo_338};
  wire [63:0]       dataInMem_lo_915 = {dataInMem_lo_hi_531, dataInMem_lo_lo_147};
  wire [31:0]       dataInMem_hi_hi_723 = {dataRegroupBySew_7_1_4, dataRegroupBySew_6_1_4};
  wire [63:0]       dataInMem_hi_1107 = {dataInMem_hi_hi_723, dataInMem_hi_lo_339};
  wire [63:0]       dataInMem_lo_916 = {dataInMem_lo_hi_532, dataInMem_lo_lo_148};
  wire [31:0]       dataInMem_hi_hi_724 = {dataRegroupBySew_7_1_5, dataRegroupBySew_6_1_5};
  wire [63:0]       dataInMem_hi_1108 = {dataInMem_hi_hi_724, dataInMem_hi_lo_340};
  wire [63:0]       dataInMem_lo_917 = {dataInMem_lo_hi_533, dataInMem_lo_lo_149};
  wire [31:0]       dataInMem_hi_hi_725 = {dataRegroupBySew_7_1_6, dataRegroupBySew_6_1_6};
  wire [63:0]       dataInMem_hi_1109 = {dataInMem_hi_hi_725, dataInMem_hi_lo_341};
  wire [63:0]       dataInMem_lo_918 = {dataInMem_lo_hi_534, dataInMem_lo_lo_150};
  wire [31:0]       dataInMem_hi_hi_726 = {dataRegroupBySew_7_1_7, dataRegroupBySew_6_1_7};
  wire [63:0]       dataInMem_hi_1110 = {dataInMem_hi_hi_726, dataInMem_hi_lo_342};
  wire [63:0]       dataInMem_lo_919 = {dataInMem_lo_hi_535, dataInMem_lo_lo_151};
  wire [31:0]       dataInMem_hi_hi_727 = {dataRegroupBySew_7_1_8, dataRegroupBySew_6_1_8};
  wire [63:0]       dataInMem_hi_1111 = {dataInMem_hi_hi_727, dataInMem_hi_lo_343};
  wire [63:0]       dataInMem_lo_920 = {dataInMem_lo_hi_536, dataInMem_lo_lo_152};
  wire [31:0]       dataInMem_hi_hi_728 = {dataRegroupBySew_7_1_9, dataRegroupBySew_6_1_9};
  wire [63:0]       dataInMem_hi_1112 = {dataInMem_hi_hi_728, dataInMem_hi_lo_344};
  wire [63:0]       dataInMem_lo_921 = {dataInMem_lo_hi_537, dataInMem_lo_lo_153};
  wire [31:0]       dataInMem_hi_hi_729 = {dataRegroupBySew_7_1_10, dataRegroupBySew_6_1_10};
  wire [63:0]       dataInMem_hi_1113 = {dataInMem_hi_hi_729, dataInMem_hi_lo_345};
  wire [63:0]       dataInMem_lo_922 = {dataInMem_lo_hi_538, dataInMem_lo_lo_154};
  wire [31:0]       dataInMem_hi_hi_730 = {dataRegroupBySew_7_1_11, dataRegroupBySew_6_1_11};
  wire [63:0]       dataInMem_hi_1114 = {dataInMem_hi_hi_730, dataInMem_hi_lo_346};
  wire [63:0]       dataInMem_lo_923 = {dataInMem_lo_hi_539, dataInMem_lo_lo_155};
  wire [31:0]       dataInMem_hi_hi_731 = {dataRegroupBySew_7_1_12, dataRegroupBySew_6_1_12};
  wire [63:0]       dataInMem_hi_1115 = {dataInMem_hi_hi_731, dataInMem_hi_lo_347};
  wire [63:0]       dataInMem_lo_924 = {dataInMem_lo_hi_540, dataInMem_lo_lo_156};
  wire [31:0]       dataInMem_hi_hi_732 = {dataRegroupBySew_7_1_13, dataRegroupBySew_6_1_13};
  wire [63:0]       dataInMem_hi_1116 = {dataInMem_hi_hi_732, dataInMem_hi_lo_348};
  wire [63:0]       dataInMem_lo_925 = {dataInMem_lo_hi_541, dataInMem_lo_lo_157};
  wire [31:0]       dataInMem_hi_hi_733 = {dataRegroupBySew_7_1_14, dataRegroupBySew_6_1_14};
  wire [63:0]       dataInMem_hi_1117 = {dataInMem_hi_hi_733, dataInMem_hi_lo_349};
  wire [63:0]       dataInMem_lo_926 = {dataInMem_lo_hi_542, dataInMem_lo_lo_158};
  wire [31:0]       dataInMem_hi_hi_734 = {dataRegroupBySew_7_1_15, dataRegroupBySew_6_1_15};
  wire [63:0]       dataInMem_hi_1118 = {dataInMem_hi_hi_734, dataInMem_hi_lo_350};
  wire [63:0]       dataInMem_lo_927 = {dataInMem_lo_hi_543, dataInMem_lo_lo_159};
  wire [31:0]       dataInMem_hi_hi_735 = {dataRegroupBySew_7_1_16, dataRegroupBySew_6_1_16};
  wire [63:0]       dataInMem_hi_1119 = {dataInMem_hi_hi_735, dataInMem_hi_lo_351};
  wire [63:0]       dataInMem_lo_928 = {dataInMem_lo_hi_544, dataInMem_lo_lo_160};
  wire [31:0]       dataInMem_hi_hi_736 = {dataRegroupBySew_7_1_17, dataRegroupBySew_6_1_17};
  wire [63:0]       dataInMem_hi_1120 = {dataInMem_hi_hi_736, dataInMem_hi_lo_352};
  wire [63:0]       dataInMem_lo_929 = {dataInMem_lo_hi_545, dataInMem_lo_lo_161};
  wire [31:0]       dataInMem_hi_hi_737 = {dataRegroupBySew_7_1_18, dataRegroupBySew_6_1_18};
  wire [63:0]       dataInMem_hi_1121 = {dataInMem_hi_hi_737, dataInMem_hi_lo_353};
  wire [63:0]       dataInMem_lo_930 = {dataInMem_lo_hi_546, dataInMem_lo_lo_162};
  wire [31:0]       dataInMem_hi_hi_738 = {dataRegroupBySew_7_1_19, dataRegroupBySew_6_1_19};
  wire [63:0]       dataInMem_hi_1122 = {dataInMem_hi_hi_738, dataInMem_hi_lo_354};
  wire [63:0]       dataInMem_lo_931 = {dataInMem_lo_hi_547, dataInMem_lo_lo_163};
  wire [31:0]       dataInMem_hi_hi_739 = {dataRegroupBySew_7_1_20, dataRegroupBySew_6_1_20};
  wire [63:0]       dataInMem_hi_1123 = {dataInMem_hi_hi_739, dataInMem_hi_lo_355};
  wire [63:0]       dataInMem_lo_932 = {dataInMem_lo_hi_548, dataInMem_lo_lo_164};
  wire [31:0]       dataInMem_hi_hi_740 = {dataRegroupBySew_7_1_21, dataRegroupBySew_6_1_21};
  wire [63:0]       dataInMem_hi_1124 = {dataInMem_hi_hi_740, dataInMem_hi_lo_356};
  wire [63:0]       dataInMem_lo_933 = {dataInMem_lo_hi_549, dataInMem_lo_lo_165};
  wire [31:0]       dataInMem_hi_hi_741 = {dataRegroupBySew_7_1_22, dataRegroupBySew_6_1_22};
  wire [63:0]       dataInMem_hi_1125 = {dataInMem_hi_hi_741, dataInMem_hi_lo_357};
  wire [63:0]       dataInMem_lo_934 = {dataInMem_lo_hi_550, dataInMem_lo_lo_166};
  wire [31:0]       dataInMem_hi_hi_742 = {dataRegroupBySew_7_1_23, dataRegroupBySew_6_1_23};
  wire [63:0]       dataInMem_hi_1126 = {dataInMem_hi_hi_742, dataInMem_hi_lo_358};
  wire [63:0]       dataInMem_lo_935 = {dataInMem_lo_hi_551, dataInMem_lo_lo_167};
  wire [31:0]       dataInMem_hi_hi_743 = {dataRegroupBySew_7_1_24, dataRegroupBySew_6_1_24};
  wire [63:0]       dataInMem_hi_1127 = {dataInMem_hi_hi_743, dataInMem_hi_lo_359};
  wire [63:0]       dataInMem_lo_936 = {dataInMem_lo_hi_552, dataInMem_lo_lo_168};
  wire [31:0]       dataInMem_hi_hi_744 = {dataRegroupBySew_7_1_25, dataRegroupBySew_6_1_25};
  wire [63:0]       dataInMem_hi_1128 = {dataInMem_hi_hi_744, dataInMem_hi_lo_360};
  wire [63:0]       dataInMem_lo_937 = {dataInMem_lo_hi_553, dataInMem_lo_lo_169};
  wire [31:0]       dataInMem_hi_hi_745 = {dataRegroupBySew_7_1_26, dataRegroupBySew_6_1_26};
  wire [63:0]       dataInMem_hi_1129 = {dataInMem_hi_hi_745, dataInMem_hi_lo_361};
  wire [63:0]       dataInMem_lo_938 = {dataInMem_lo_hi_554, dataInMem_lo_lo_170};
  wire [31:0]       dataInMem_hi_hi_746 = {dataRegroupBySew_7_1_27, dataRegroupBySew_6_1_27};
  wire [63:0]       dataInMem_hi_1130 = {dataInMem_hi_hi_746, dataInMem_hi_lo_362};
  wire [63:0]       dataInMem_lo_939 = {dataInMem_lo_hi_555, dataInMem_lo_lo_171};
  wire [31:0]       dataInMem_hi_hi_747 = {dataRegroupBySew_7_1_28, dataRegroupBySew_6_1_28};
  wire [63:0]       dataInMem_hi_1131 = {dataInMem_hi_hi_747, dataInMem_hi_lo_363};
  wire [63:0]       dataInMem_lo_940 = {dataInMem_lo_hi_556, dataInMem_lo_lo_172};
  wire [31:0]       dataInMem_hi_hi_748 = {dataRegroupBySew_7_1_29, dataRegroupBySew_6_1_29};
  wire [63:0]       dataInMem_hi_1132 = {dataInMem_hi_hi_748, dataInMem_hi_lo_364};
  wire [63:0]       dataInMem_lo_941 = {dataInMem_lo_hi_557, dataInMem_lo_lo_173};
  wire [31:0]       dataInMem_hi_hi_749 = {dataRegroupBySew_7_1_30, dataRegroupBySew_6_1_30};
  wire [63:0]       dataInMem_hi_1133 = {dataInMem_hi_hi_749, dataInMem_hi_lo_365};
  wire [63:0]       dataInMem_lo_942 = {dataInMem_lo_hi_558, dataInMem_lo_lo_174};
  wire [31:0]       dataInMem_hi_hi_750 = {dataRegroupBySew_7_1_31, dataRegroupBySew_6_1_31};
  wire [63:0]       dataInMem_hi_1134 = {dataInMem_hi_hi_750, dataInMem_hi_lo_366};
  wire [63:0]       dataInMem_lo_943 = {dataInMem_lo_hi_559, dataInMem_lo_lo_175};
  wire [31:0]       dataInMem_hi_hi_751 = {dataRegroupBySew_7_1_32, dataRegroupBySew_6_1_32};
  wire [63:0]       dataInMem_hi_1135 = {dataInMem_hi_hi_751, dataInMem_hi_lo_367};
  wire [63:0]       dataInMem_lo_944 = {dataInMem_lo_hi_560, dataInMem_lo_lo_176};
  wire [31:0]       dataInMem_hi_hi_752 = {dataRegroupBySew_7_1_33, dataRegroupBySew_6_1_33};
  wire [63:0]       dataInMem_hi_1136 = {dataInMem_hi_hi_752, dataInMem_hi_lo_368};
  wire [63:0]       dataInMem_lo_945 = {dataInMem_lo_hi_561, dataInMem_lo_lo_177};
  wire [31:0]       dataInMem_hi_hi_753 = {dataRegroupBySew_7_1_34, dataRegroupBySew_6_1_34};
  wire [63:0]       dataInMem_hi_1137 = {dataInMem_hi_hi_753, dataInMem_hi_lo_369};
  wire [63:0]       dataInMem_lo_946 = {dataInMem_lo_hi_562, dataInMem_lo_lo_178};
  wire [31:0]       dataInMem_hi_hi_754 = {dataRegroupBySew_7_1_35, dataRegroupBySew_6_1_35};
  wire [63:0]       dataInMem_hi_1138 = {dataInMem_hi_hi_754, dataInMem_hi_lo_370};
  wire [63:0]       dataInMem_lo_947 = {dataInMem_lo_hi_563, dataInMem_lo_lo_179};
  wire [31:0]       dataInMem_hi_hi_755 = {dataRegroupBySew_7_1_36, dataRegroupBySew_6_1_36};
  wire [63:0]       dataInMem_hi_1139 = {dataInMem_hi_hi_755, dataInMem_hi_lo_371};
  wire [63:0]       dataInMem_lo_948 = {dataInMem_lo_hi_564, dataInMem_lo_lo_180};
  wire [31:0]       dataInMem_hi_hi_756 = {dataRegroupBySew_7_1_37, dataRegroupBySew_6_1_37};
  wire [63:0]       dataInMem_hi_1140 = {dataInMem_hi_hi_756, dataInMem_hi_lo_372};
  wire [63:0]       dataInMem_lo_949 = {dataInMem_lo_hi_565, dataInMem_lo_lo_181};
  wire [31:0]       dataInMem_hi_hi_757 = {dataRegroupBySew_7_1_38, dataRegroupBySew_6_1_38};
  wire [63:0]       dataInMem_hi_1141 = {dataInMem_hi_hi_757, dataInMem_hi_lo_373};
  wire [63:0]       dataInMem_lo_950 = {dataInMem_lo_hi_566, dataInMem_lo_lo_182};
  wire [31:0]       dataInMem_hi_hi_758 = {dataRegroupBySew_7_1_39, dataRegroupBySew_6_1_39};
  wire [63:0]       dataInMem_hi_1142 = {dataInMem_hi_hi_758, dataInMem_hi_lo_374};
  wire [63:0]       dataInMem_lo_951 = {dataInMem_lo_hi_567, dataInMem_lo_lo_183};
  wire [31:0]       dataInMem_hi_hi_759 = {dataRegroupBySew_7_1_40, dataRegroupBySew_6_1_40};
  wire [63:0]       dataInMem_hi_1143 = {dataInMem_hi_hi_759, dataInMem_hi_lo_375};
  wire [63:0]       dataInMem_lo_952 = {dataInMem_lo_hi_568, dataInMem_lo_lo_184};
  wire [31:0]       dataInMem_hi_hi_760 = {dataRegroupBySew_7_1_41, dataRegroupBySew_6_1_41};
  wire [63:0]       dataInMem_hi_1144 = {dataInMem_hi_hi_760, dataInMem_hi_lo_376};
  wire [63:0]       dataInMem_lo_953 = {dataInMem_lo_hi_569, dataInMem_lo_lo_185};
  wire [31:0]       dataInMem_hi_hi_761 = {dataRegroupBySew_7_1_42, dataRegroupBySew_6_1_42};
  wire [63:0]       dataInMem_hi_1145 = {dataInMem_hi_hi_761, dataInMem_hi_lo_377};
  wire [63:0]       dataInMem_lo_954 = {dataInMem_lo_hi_570, dataInMem_lo_lo_186};
  wire [31:0]       dataInMem_hi_hi_762 = {dataRegroupBySew_7_1_43, dataRegroupBySew_6_1_43};
  wire [63:0]       dataInMem_hi_1146 = {dataInMem_hi_hi_762, dataInMem_hi_lo_378};
  wire [63:0]       dataInMem_lo_955 = {dataInMem_lo_hi_571, dataInMem_lo_lo_187};
  wire [31:0]       dataInMem_hi_hi_763 = {dataRegroupBySew_7_1_44, dataRegroupBySew_6_1_44};
  wire [63:0]       dataInMem_hi_1147 = {dataInMem_hi_hi_763, dataInMem_hi_lo_379};
  wire [63:0]       dataInMem_lo_956 = {dataInMem_lo_hi_572, dataInMem_lo_lo_188};
  wire [31:0]       dataInMem_hi_hi_764 = {dataRegroupBySew_7_1_45, dataRegroupBySew_6_1_45};
  wire [63:0]       dataInMem_hi_1148 = {dataInMem_hi_hi_764, dataInMem_hi_lo_380};
  wire [63:0]       dataInMem_lo_957 = {dataInMem_lo_hi_573, dataInMem_lo_lo_189};
  wire [31:0]       dataInMem_hi_hi_765 = {dataRegroupBySew_7_1_46, dataRegroupBySew_6_1_46};
  wire [63:0]       dataInMem_hi_1149 = {dataInMem_hi_hi_765, dataInMem_hi_lo_381};
  wire [63:0]       dataInMem_lo_958 = {dataInMem_lo_hi_574, dataInMem_lo_lo_190};
  wire [31:0]       dataInMem_hi_hi_766 = {dataRegroupBySew_7_1_47, dataRegroupBySew_6_1_47};
  wire [63:0]       dataInMem_hi_1150 = {dataInMem_hi_hi_766, dataInMem_hi_lo_382};
  wire [63:0]       dataInMem_lo_959 = {dataInMem_lo_hi_575, dataInMem_lo_lo_191};
  wire [31:0]       dataInMem_hi_hi_767 = {dataRegroupBySew_7_1_48, dataRegroupBySew_6_1_48};
  wire [63:0]       dataInMem_hi_1151 = {dataInMem_hi_hi_767, dataInMem_hi_lo_383};
  wire [63:0]       dataInMem_lo_960 = {dataInMem_lo_hi_576, dataInMem_lo_lo_192};
  wire [31:0]       dataInMem_hi_hi_768 = {dataRegroupBySew_7_1_49, dataRegroupBySew_6_1_49};
  wire [63:0]       dataInMem_hi_1152 = {dataInMem_hi_hi_768, dataInMem_hi_lo_384};
  wire [63:0]       dataInMem_lo_961 = {dataInMem_lo_hi_577, dataInMem_lo_lo_193};
  wire [31:0]       dataInMem_hi_hi_769 = {dataRegroupBySew_7_1_50, dataRegroupBySew_6_1_50};
  wire [63:0]       dataInMem_hi_1153 = {dataInMem_hi_hi_769, dataInMem_hi_lo_385};
  wire [63:0]       dataInMem_lo_962 = {dataInMem_lo_hi_578, dataInMem_lo_lo_194};
  wire [31:0]       dataInMem_hi_hi_770 = {dataRegroupBySew_7_1_51, dataRegroupBySew_6_1_51};
  wire [63:0]       dataInMem_hi_1154 = {dataInMem_hi_hi_770, dataInMem_hi_lo_386};
  wire [63:0]       dataInMem_lo_963 = {dataInMem_lo_hi_579, dataInMem_lo_lo_195};
  wire [31:0]       dataInMem_hi_hi_771 = {dataRegroupBySew_7_1_52, dataRegroupBySew_6_1_52};
  wire [63:0]       dataInMem_hi_1155 = {dataInMem_hi_hi_771, dataInMem_hi_lo_387};
  wire [63:0]       dataInMem_lo_964 = {dataInMem_lo_hi_580, dataInMem_lo_lo_196};
  wire [31:0]       dataInMem_hi_hi_772 = {dataRegroupBySew_7_1_53, dataRegroupBySew_6_1_53};
  wire [63:0]       dataInMem_hi_1156 = {dataInMem_hi_hi_772, dataInMem_hi_lo_388};
  wire [63:0]       dataInMem_lo_965 = {dataInMem_lo_hi_581, dataInMem_lo_lo_197};
  wire [31:0]       dataInMem_hi_hi_773 = {dataRegroupBySew_7_1_54, dataRegroupBySew_6_1_54};
  wire [63:0]       dataInMem_hi_1157 = {dataInMem_hi_hi_773, dataInMem_hi_lo_389};
  wire [63:0]       dataInMem_lo_966 = {dataInMem_lo_hi_582, dataInMem_lo_lo_198};
  wire [31:0]       dataInMem_hi_hi_774 = {dataRegroupBySew_7_1_55, dataRegroupBySew_6_1_55};
  wire [63:0]       dataInMem_hi_1158 = {dataInMem_hi_hi_774, dataInMem_hi_lo_390};
  wire [63:0]       dataInMem_lo_967 = {dataInMem_lo_hi_583, dataInMem_lo_lo_199};
  wire [31:0]       dataInMem_hi_hi_775 = {dataRegroupBySew_7_1_56, dataRegroupBySew_6_1_56};
  wire [63:0]       dataInMem_hi_1159 = {dataInMem_hi_hi_775, dataInMem_hi_lo_391};
  wire [63:0]       dataInMem_lo_968 = {dataInMem_lo_hi_584, dataInMem_lo_lo_200};
  wire [31:0]       dataInMem_hi_hi_776 = {dataRegroupBySew_7_1_57, dataRegroupBySew_6_1_57};
  wire [63:0]       dataInMem_hi_1160 = {dataInMem_hi_hi_776, dataInMem_hi_lo_392};
  wire [63:0]       dataInMem_lo_969 = {dataInMem_lo_hi_585, dataInMem_lo_lo_201};
  wire [31:0]       dataInMem_hi_hi_777 = {dataRegroupBySew_7_1_58, dataRegroupBySew_6_1_58};
  wire [63:0]       dataInMem_hi_1161 = {dataInMem_hi_hi_777, dataInMem_hi_lo_393};
  wire [63:0]       dataInMem_lo_970 = {dataInMem_lo_hi_586, dataInMem_lo_lo_202};
  wire [31:0]       dataInMem_hi_hi_778 = {dataRegroupBySew_7_1_59, dataRegroupBySew_6_1_59};
  wire [63:0]       dataInMem_hi_1162 = {dataInMem_hi_hi_778, dataInMem_hi_lo_394};
  wire [63:0]       dataInMem_lo_971 = {dataInMem_lo_hi_587, dataInMem_lo_lo_203};
  wire [31:0]       dataInMem_hi_hi_779 = {dataRegroupBySew_7_1_60, dataRegroupBySew_6_1_60};
  wire [63:0]       dataInMem_hi_1163 = {dataInMem_hi_hi_779, dataInMem_hi_lo_395};
  wire [63:0]       dataInMem_lo_972 = {dataInMem_lo_hi_588, dataInMem_lo_lo_204};
  wire [31:0]       dataInMem_hi_hi_780 = {dataRegroupBySew_7_1_61, dataRegroupBySew_6_1_61};
  wire [63:0]       dataInMem_hi_1164 = {dataInMem_hi_hi_780, dataInMem_hi_lo_396};
  wire [63:0]       dataInMem_lo_973 = {dataInMem_lo_hi_589, dataInMem_lo_lo_205};
  wire [31:0]       dataInMem_hi_hi_781 = {dataRegroupBySew_7_1_62, dataRegroupBySew_6_1_62};
  wire [63:0]       dataInMem_hi_1165 = {dataInMem_hi_hi_781, dataInMem_hi_lo_397};
  wire [63:0]       dataInMem_lo_974 = {dataInMem_lo_hi_590, dataInMem_lo_lo_206};
  wire [31:0]       dataInMem_hi_hi_782 = {dataRegroupBySew_7_1_63, dataRegroupBySew_6_1_63};
  wire [63:0]       dataInMem_hi_1166 = {dataInMem_hi_hi_782, dataInMem_hi_lo_398};
  wire [255:0]      dataInMem_lo_lo_lo_lo_lo_15 = {dataInMem_hi_1104, dataInMem_lo_912, dataInMem_hi_1103, dataInMem_lo_911};
  wire [255:0]      dataInMem_lo_lo_lo_lo_hi_15 = {dataInMem_hi_1106, dataInMem_lo_914, dataInMem_hi_1105, dataInMem_lo_913};
  wire [511:0]      dataInMem_lo_lo_lo_lo_15 = {dataInMem_lo_lo_lo_lo_hi_15, dataInMem_lo_lo_lo_lo_lo_15};
  wire [255:0]      dataInMem_lo_lo_lo_hi_lo_15 = {dataInMem_hi_1108, dataInMem_lo_916, dataInMem_hi_1107, dataInMem_lo_915};
  wire [255:0]      dataInMem_lo_lo_lo_hi_hi_15 = {dataInMem_hi_1110, dataInMem_lo_918, dataInMem_hi_1109, dataInMem_lo_917};
  wire [511:0]      dataInMem_lo_lo_lo_hi_15 = {dataInMem_lo_lo_lo_hi_hi_15, dataInMem_lo_lo_lo_hi_lo_15};
  wire [1023:0]     dataInMem_lo_lo_lo_15 = {dataInMem_lo_lo_lo_hi_15, dataInMem_lo_lo_lo_lo_15};
  wire [255:0]      dataInMem_lo_lo_hi_lo_lo_15 = {dataInMem_hi_1112, dataInMem_lo_920, dataInMem_hi_1111, dataInMem_lo_919};
  wire [255:0]      dataInMem_lo_lo_hi_lo_hi_15 = {dataInMem_hi_1114, dataInMem_lo_922, dataInMem_hi_1113, dataInMem_lo_921};
  wire [511:0]      dataInMem_lo_lo_hi_lo_15 = {dataInMem_lo_lo_hi_lo_hi_15, dataInMem_lo_lo_hi_lo_lo_15};
  wire [255:0]      dataInMem_lo_lo_hi_hi_lo_15 = {dataInMem_hi_1116, dataInMem_lo_924, dataInMem_hi_1115, dataInMem_lo_923};
  wire [255:0]      dataInMem_lo_lo_hi_hi_hi_15 = {dataInMem_hi_1118, dataInMem_lo_926, dataInMem_hi_1117, dataInMem_lo_925};
  wire [511:0]      dataInMem_lo_lo_hi_hi_15 = {dataInMem_lo_lo_hi_hi_hi_15, dataInMem_lo_lo_hi_hi_lo_15};
  wire [1023:0]     dataInMem_lo_lo_hi_15 = {dataInMem_lo_lo_hi_hi_15, dataInMem_lo_lo_hi_lo_15};
  wire [2047:0]     dataInMem_lo_lo_207 = {dataInMem_lo_lo_hi_15, dataInMem_lo_lo_lo_15};
  wire [255:0]      dataInMem_lo_hi_lo_lo_lo_15 = {dataInMem_hi_1120, dataInMem_lo_928, dataInMem_hi_1119, dataInMem_lo_927};
  wire [255:0]      dataInMem_lo_hi_lo_lo_hi_15 = {dataInMem_hi_1122, dataInMem_lo_930, dataInMem_hi_1121, dataInMem_lo_929};
  wire [511:0]      dataInMem_lo_hi_lo_lo_15 = {dataInMem_lo_hi_lo_lo_hi_15, dataInMem_lo_hi_lo_lo_lo_15};
  wire [255:0]      dataInMem_lo_hi_lo_hi_lo_15 = {dataInMem_hi_1124, dataInMem_lo_932, dataInMem_hi_1123, dataInMem_lo_931};
  wire [255:0]      dataInMem_lo_hi_lo_hi_hi_15 = {dataInMem_hi_1126, dataInMem_lo_934, dataInMem_hi_1125, dataInMem_lo_933};
  wire [511:0]      dataInMem_lo_hi_lo_hi_15 = {dataInMem_lo_hi_lo_hi_hi_15, dataInMem_lo_hi_lo_hi_lo_15};
  wire [1023:0]     dataInMem_lo_hi_lo_15 = {dataInMem_lo_hi_lo_hi_15, dataInMem_lo_hi_lo_lo_15};
  wire [255:0]      dataInMem_lo_hi_hi_lo_lo_15 = {dataInMem_hi_1128, dataInMem_lo_936, dataInMem_hi_1127, dataInMem_lo_935};
  wire [255:0]      dataInMem_lo_hi_hi_lo_hi_15 = {dataInMem_hi_1130, dataInMem_lo_938, dataInMem_hi_1129, dataInMem_lo_937};
  wire [511:0]      dataInMem_lo_hi_hi_lo_15 = {dataInMem_lo_hi_hi_lo_hi_15, dataInMem_lo_hi_hi_lo_lo_15};
  wire [255:0]      dataInMem_lo_hi_hi_hi_lo_15 = {dataInMem_hi_1132, dataInMem_lo_940, dataInMem_hi_1131, dataInMem_lo_939};
  wire [255:0]      dataInMem_lo_hi_hi_hi_hi_15 = {dataInMem_hi_1134, dataInMem_lo_942, dataInMem_hi_1133, dataInMem_lo_941};
  wire [511:0]      dataInMem_lo_hi_hi_hi_15 = {dataInMem_lo_hi_hi_hi_hi_15, dataInMem_lo_hi_hi_hi_lo_15};
  wire [1023:0]     dataInMem_lo_hi_hi_15 = {dataInMem_lo_hi_hi_hi_15, dataInMem_lo_hi_hi_lo_15};
  wire [2047:0]     dataInMem_lo_hi_591 = {dataInMem_lo_hi_hi_15, dataInMem_lo_hi_lo_15};
  wire [4095:0]     dataInMem_lo_975 = {dataInMem_lo_hi_591, dataInMem_lo_lo_207};
  wire [255:0]      dataInMem_hi_lo_lo_lo_lo_15 = {dataInMem_hi_1136, dataInMem_lo_944, dataInMem_hi_1135, dataInMem_lo_943};
  wire [255:0]      dataInMem_hi_lo_lo_lo_hi_15 = {dataInMem_hi_1138, dataInMem_lo_946, dataInMem_hi_1137, dataInMem_lo_945};
  wire [511:0]      dataInMem_hi_lo_lo_lo_15 = {dataInMem_hi_lo_lo_lo_hi_15, dataInMem_hi_lo_lo_lo_lo_15};
  wire [255:0]      dataInMem_hi_lo_lo_hi_lo_15 = {dataInMem_hi_1140, dataInMem_lo_948, dataInMem_hi_1139, dataInMem_lo_947};
  wire [255:0]      dataInMem_hi_lo_lo_hi_hi_15 = {dataInMem_hi_1142, dataInMem_lo_950, dataInMem_hi_1141, dataInMem_lo_949};
  wire [511:0]      dataInMem_hi_lo_lo_hi_15 = {dataInMem_hi_lo_lo_hi_hi_15, dataInMem_hi_lo_lo_hi_lo_15};
  wire [1023:0]     dataInMem_hi_lo_lo_15 = {dataInMem_hi_lo_lo_hi_15, dataInMem_hi_lo_lo_lo_15};
  wire [255:0]      dataInMem_hi_lo_hi_lo_lo_15 = {dataInMem_hi_1144, dataInMem_lo_952, dataInMem_hi_1143, dataInMem_lo_951};
  wire [255:0]      dataInMem_hi_lo_hi_lo_hi_15 = {dataInMem_hi_1146, dataInMem_lo_954, dataInMem_hi_1145, dataInMem_lo_953};
  wire [511:0]      dataInMem_hi_lo_hi_lo_15 = {dataInMem_hi_lo_hi_lo_hi_15, dataInMem_hi_lo_hi_lo_lo_15};
  wire [255:0]      dataInMem_hi_lo_hi_hi_lo_15 = {dataInMem_hi_1148, dataInMem_lo_956, dataInMem_hi_1147, dataInMem_lo_955};
  wire [255:0]      dataInMem_hi_lo_hi_hi_hi_15 = {dataInMem_hi_1150, dataInMem_lo_958, dataInMem_hi_1149, dataInMem_lo_957};
  wire [511:0]      dataInMem_hi_lo_hi_hi_15 = {dataInMem_hi_lo_hi_hi_hi_15, dataInMem_hi_lo_hi_hi_lo_15};
  wire [1023:0]     dataInMem_hi_lo_hi_15 = {dataInMem_hi_lo_hi_hi_15, dataInMem_hi_lo_hi_lo_15};
  wire [2047:0]     dataInMem_hi_lo_399 = {dataInMem_hi_lo_hi_15, dataInMem_hi_lo_lo_15};
  wire [255:0]      dataInMem_hi_hi_lo_lo_lo_15 = {dataInMem_hi_1152, dataInMem_lo_960, dataInMem_hi_1151, dataInMem_lo_959};
  wire [255:0]      dataInMem_hi_hi_lo_lo_hi_15 = {dataInMem_hi_1154, dataInMem_lo_962, dataInMem_hi_1153, dataInMem_lo_961};
  wire [511:0]      dataInMem_hi_hi_lo_lo_15 = {dataInMem_hi_hi_lo_lo_hi_15, dataInMem_hi_hi_lo_lo_lo_15};
  wire [255:0]      dataInMem_hi_hi_lo_hi_lo_15 = {dataInMem_hi_1156, dataInMem_lo_964, dataInMem_hi_1155, dataInMem_lo_963};
  wire [255:0]      dataInMem_hi_hi_lo_hi_hi_15 = {dataInMem_hi_1158, dataInMem_lo_966, dataInMem_hi_1157, dataInMem_lo_965};
  wire [511:0]      dataInMem_hi_hi_lo_hi_15 = {dataInMem_hi_hi_lo_hi_hi_15, dataInMem_hi_hi_lo_hi_lo_15};
  wire [1023:0]     dataInMem_hi_hi_lo_15 = {dataInMem_hi_hi_lo_hi_15, dataInMem_hi_hi_lo_lo_15};
  wire [255:0]      dataInMem_hi_hi_hi_lo_lo_15 = {dataInMem_hi_1160, dataInMem_lo_968, dataInMem_hi_1159, dataInMem_lo_967};
  wire [255:0]      dataInMem_hi_hi_hi_lo_hi_15 = {dataInMem_hi_1162, dataInMem_lo_970, dataInMem_hi_1161, dataInMem_lo_969};
  wire [511:0]      dataInMem_hi_hi_hi_lo_15 = {dataInMem_hi_hi_hi_lo_hi_15, dataInMem_hi_hi_hi_lo_lo_15};
  wire [255:0]      dataInMem_hi_hi_hi_hi_lo_15 = {dataInMem_hi_1164, dataInMem_lo_972, dataInMem_hi_1163, dataInMem_lo_971};
  wire [255:0]      dataInMem_hi_hi_hi_hi_hi_15 = {dataInMem_hi_1166, dataInMem_lo_974, dataInMem_hi_1165, dataInMem_lo_973};
  wire [511:0]      dataInMem_hi_hi_hi_hi_15 = {dataInMem_hi_hi_hi_hi_hi_15, dataInMem_hi_hi_hi_hi_lo_15};
  wire [1023:0]     dataInMem_hi_hi_hi_15 = {dataInMem_hi_hi_hi_hi_15, dataInMem_hi_hi_hi_lo_15};
  wire [2047:0]     dataInMem_hi_hi_783 = {dataInMem_hi_hi_hi_15, dataInMem_hi_hi_lo_15};
  wire [4095:0]     dataInMem_hi_1167 = {dataInMem_hi_hi_783, dataInMem_hi_lo_399};
  wire [8191:0]     dataInMem_15 = {dataInMem_hi_1167, dataInMem_lo_975};
  wire [1023:0]     regroupCacheLine_15_0 = dataInMem_15[1023:0];
  wire [1023:0]     regroupCacheLine_15_1 = dataInMem_15[2047:1024];
  wire [1023:0]     regroupCacheLine_15_2 = dataInMem_15[3071:2048];
  wire [1023:0]     regroupCacheLine_15_3 = dataInMem_15[4095:3072];
  wire [1023:0]     regroupCacheLine_15_4 = dataInMem_15[5119:4096];
  wire [1023:0]     regroupCacheLine_15_5 = dataInMem_15[6143:5120];
  wire [1023:0]     regroupCacheLine_15_6 = dataInMem_15[7167:6144];
  wire [1023:0]     regroupCacheLine_15_7 = dataInMem_15[8191:7168];
  wire [1023:0]     res_120 = regroupCacheLine_15_0;
  wire [1023:0]     res_121 = regroupCacheLine_15_1;
  wire [1023:0]     res_122 = regroupCacheLine_15_2;
  wire [1023:0]     res_123 = regroupCacheLine_15_3;
  wire [1023:0]     res_124 = regroupCacheLine_15_4;
  wire [1023:0]     res_125 = regroupCacheLine_15_5;
  wire [1023:0]     res_126 = regroupCacheLine_15_6;
  wire [1023:0]     res_127 = regroupCacheLine_15_7;
  wire [2047:0]     lo_lo_15 = {res_121, res_120};
  wire [2047:0]     lo_hi_15 = {res_123, res_122};
  wire [4095:0]     lo_15 = {lo_hi_15, lo_lo_15};
  wire [2047:0]     hi_lo_15 = {res_125, res_124};
  wire [2047:0]     hi_hi_15 = {res_127, res_126};
  wire [4095:0]     hi_15 = {hi_hi_15, hi_lo_15};
  wire [8191:0]     regroupLoadData_1_7 = {hi_15, lo_15};
  wire [31:0]       dataRegroupBySew_0_2_0 = bufferStageEnqueueData_0[31:0];
  wire [31:0]       dataRegroupBySew_0_2_1 = bufferStageEnqueueData_0[63:32];
  wire [31:0]       dataRegroupBySew_0_2_2 = bufferStageEnqueueData_0[95:64];
  wire [31:0]       dataRegroupBySew_0_2_3 = bufferStageEnqueueData_0[127:96];
  wire [31:0]       dataRegroupBySew_0_2_4 = bufferStageEnqueueData_0[159:128];
  wire [31:0]       dataRegroupBySew_0_2_5 = bufferStageEnqueueData_0[191:160];
  wire [31:0]       dataRegroupBySew_0_2_6 = bufferStageEnqueueData_0[223:192];
  wire [31:0]       dataRegroupBySew_0_2_7 = bufferStageEnqueueData_0[255:224];
  wire [31:0]       dataRegroupBySew_0_2_8 = bufferStageEnqueueData_0[287:256];
  wire [31:0]       dataRegroupBySew_0_2_9 = bufferStageEnqueueData_0[319:288];
  wire [31:0]       dataRegroupBySew_0_2_10 = bufferStageEnqueueData_0[351:320];
  wire [31:0]       dataRegroupBySew_0_2_11 = bufferStageEnqueueData_0[383:352];
  wire [31:0]       dataRegroupBySew_0_2_12 = bufferStageEnqueueData_0[415:384];
  wire [31:0]       dataRegroupBySew_0_2_13 = bufferStageEnqueueData_0[447:416];
  wire [31:0]       dataRegroupBySew_0_2_14 = bufferStageEnqueueData_0[479:448];
  wire [31:0]       dataRegroupBySew_0_2_15 = bufferStageEnqueueData_0[511:480];
  wire [31:0]       dataRegroupBySew_0_2_16 = bufferStageEnqueueData_0[543:512];
  wire [31:0]       dataRegroupBySew_0_2_17 = bufferStageEnqueueData_0[575:544];
  wire [31:0]       dataRegroupBySew_0_2_18 = bufferStageEnqueueData_0[607:576];
  wire [31:0]       dataRegroupBySew_0_2_19 = bufferStageEnqueueData_0[639:608];
  wire [31:0]       dataRegroupBySew_0_2_20 = bufferStageEnqueueData_0[671:640];
  wire [31:0]       dataRegroupBySew_0_2_21 = bufferStageEnqueueData_0[703:672];
  wire [31:0]       dataRegroupBySew_0_2_22 = bufferStageEnqueueData_0[735:704];
  wire [31:0]       dataRegroupBySew_0_2_23 = bufferStageEnqueueData_0[767:736];
  wire [31:0]       dataRegroupBySew_0_2_24 = bufferStageEnqueueData_0[799:768];
  wire [31:0]       dataRegroupBySew_0_2_25 = bufferStageEnqueueData_0[831:800];
  wire [31:0]       dataRegroupBySew_0_2_26 = bufferStageEnqueueData_0[863:832];
  wire [31:0]       dataRegroupBySew_0_2_27 = bufferStageEnqueueData_0[895:864];
  wire [31:0]       dataRegroupBySew_0_2_28 = bufferStageEnqueueData_0[927:896];
  wire [31:0]       dataRegroupBySew_0_2_29 = bufferStageEnqueueData_0[959:928];
  wire [31:0]       dataRegroupBySew_0_2_30 = bufferStageEnqueueData_0[991:960];
  wire [31:0]       dataRegroupBySew_0_2_31 = bufferStageEnqueueData_0[1023:992];
  wire [31:0]       dataRegroupBySew_1_2_0 = bufferStageEnqueueData_1[31:0];
  wire [31:0]       dataRegroupBySew_1_2_1 = bufferStageEnqueueData_1[63:32];
  wire [31:0]       dataRegroupBySew_1_2_2 = bufferStageEnqueueData_1[95:64];
  wire [31:0]       dataRegroupBySew_1_2_3 = bufferStageEnqueueData_1[127:96];
  wire [31:0]       dataRegroupBySew_1_2_4 = bufferStageEnqueueData_1[159:128];
  wire [31:0]       dataRegroupBySew_1_2_5 = bufferStageEnqueueData_1[191:160];
  wire [31:0]       dataRegroupBySew_1_2_6 = bufferStageEnqueueData_1[223:192];
  wire [31:0]       dataRegroupBySew_1_2_7 = bufferStageEnqueueData_1[255:224];
  wire [31:0]       dataRegroupBySew_1_2_8 = bufferStageEnqueueData_1[287:256];
  wire [31:0]       dataRegroupBySew_1_2_9 = bufferStageEnqueueData_1[319:288];
  wire [31:0]       dataRegroupBySew_1_2_10 = bufferStageEnqueueData_1[351:320];
  wire [31:0]       dataRegroupBySew_1_2_11 = bufferStageEnqueueData_1[383:352];
  wire [31:0]       dataRegroupBySew_1_2_12 = bufferStageEnqueueData_1[415:384];
  wire [31:0]       dataRegroupBySew_1_2_13 = bufferStageEnqueueData_1[447:416];
  wire [31:0]       dataRegroupBySew_1_2_14 = bufferStageEnqueueData_1[479:448];
  wire [31:0]       dataRegroupBySew_1_2_15 = bufferStageEnqueueData_1[511:480];
  wire [31:0]       dataRegroupBySew_1_2_16 = bufferStageEnqueueData_1[543:512];
  wire [31:0]       dataRegroupBySew_1_2_17 = bufferStageEnqueueData_1[575:544];
  wire [31:0]       dataRegroupBySew_1_2_18 = bufferStageEnqueueData_1[607:576];
  wire [31:0]       dataRegroupBySew_1_2_19 = bufferStageEnqueueData_1[639:608];
  wire [31:0]       dataRegroupBySew_1_2_20 = bufferStageEnqueueData_1[671:640];
  wire [31:0]       dataRegroupBySew_1_2_21 = bufferStageEnqueueData_1[703:672];
  wire [31:0]       dataRegroupBySew_1_2_22 = bufferStageEnqueueData_1[735:704];
  wire [31:0]       dataRegroupBySew_1_2_23 = bufferStageEnqueueData_1[767:736];
  wire [31:0]       dataRegroupBySew_1_2_24 = bufferStageEnqueueData_1[799:768];
  wire [31:0]       dataRegroupBySew_1_2_25 = bufferStageEnqueueData_1[831:800];
  wire [31:0]       dataRegroupBySew_1_2_26 = bufferStageEnqueueData_1[863:832];
  wire [31:0]       dataRegroupBySew_1_2_27 = bufferStageEnqueueData_1[895:864];
  wire [31:0]       dataRegroupBySew_1_2_28 = bufferStageEnqueueData_1[927:896];
  wire [31:0]       dataRegroupBySew_1_2_29 = bufferStageEnqueueData_1[959:928];
  wire [31:0]       dataRegroupBySew_1_2_30 = bufferStageEnqueueData_1[991:960];
  wire [31:0]       dataRegroupBySew_1_2_31 = bufferStageEnqueueData_1[1023:992];
  wire [31:0]       dataRegroupBySew_2_2_0 = bufferStageEnqueueData_2[31:0];
  wire [31:0]       dataRegroupBySew_2_2_1 = bufferStageEnqueueData_2[63:32];
  wire [31:0]       dataRegroupBySew_2_2_2 = bufferStageEnqueueData_2[95:64];
  wire [31:0]       dataRegroupBySew_2_2_3 = bufferStageEnqueueData_2[127:96];
  wire [31:0]       dataRegroupBySew_2_2_4 = bufferStageEnqueueData_2[159:128];
  wire [31:0]       dataRegroupBySew_2_2_5 = bufferStageEnqueueData_2[191:160];
  wire [31:0]       dataRegroupBySew_2_2_6 = bufferStageEnqueueData_2[223:192];
  wire [31:0]       dataRegroupBySew_2_2_7 = bufferStageEnqueueData_2[255:224];
  wire [31:0]       dataRegroupBySew_2_2_8 = bufferStageEnqueueData_2[287:256];
  wire [31:0]       dataRegroupBySew_2_2_9 = bufferStageEnqueueData_2[319:288];
  wire [31:0]       dataRegroupBySew_2_2_10 = bufferStageEnqueueData_2[351:320];
  wire [31:0]       dataRegroupBySew_2_2_11 = bufferStageEnqueueData_2[383:352];
  wire [31:0]       dataRegroupBySew_2_2_12 = bufferStageEnqueueData_2[415:384];
  wire [31:0]       dataRegroupBySew_2_2_13 = bufferStageEnqueueData_2[447:416];
  wire [31:0]       dataRegroupBySew_2_2_14 = bufferStageEnqueueData_2[479:448];
  wire [31:0]       dataRegroupBySew_2_2_15 = bufferStageEnqueueData_2[511:480];
  wire [31:0]       dataRegroupBySew_2_2_16 = bufferStageEnqueueData_2[543:512];
  wire [31:0]       dataRegroupBySew_2_2_17 = bufferStageEnqueueData_2[575:544];
  wire [31:0]       dataRegroupBySew_2_2_18 = bufferStageEnqueueData_2[607:576];
  wire [31:0]       dataRegroupBySew_2_2_19 = bufferStageEnqueueData_2[639:608];
  wire [31:0]       dataRegroupBySew_2_2_20 = bufferStageEnqueueData_2[671:640];
  wire [31:0]       dataRegroupBySew_2_2_21 = bufferStageEnqueueData_2[703:672];
  wire [31:0]       dataRegroupBySew_2_2_22 = bufferStageEnqueueData_2[735:704];
  wire [31:0]       dataRegroupBySew_2_2_23 = bufferStageEnqueueData_2[767:736];
  wire [31:0]       dataRegroupBySew_2_2_24 = bufferStageEnqueueData_2[799:768];
  wire [31:0]       dataRegroupBySew_2_2_25 = bufferStageEnqueueData_2[831:800];
  wire [31:0]       dataRegroupBySew_2_2_26 = bufferStageEnqueueData_2[863:832];
  wire [31:0]       dataRegroupBySew_2_2_27 = bufferStageEnqueueData_2[895:864];
  wire [31:0]       dataRegroupBySew_2_2_28 = bufferStageEnqueueData_2[927:896];
  wire [31:0]       dataRegroupBySew_2_2_29 = bufferStageEnqueueData_2[959:928];
  wire [31:0]       dataRegroupBySew_2_2_30 = bufferStageEnqueueData_2[991:960];
  wire [31:0]       dataRegroupBySew_2_2_31 = bufferStageEnqueueData_2[1023:992];
  wire [31:0]       dataRegroupBySew_3_2_0 = bufferStageEnqueueData_3[31:0];
  wire [31:0]       dataRegroupBySew_3_2_1 = bufferStageEnqueueData_3[63:32];
  wire [31:0]       dataRegroupBySew_3_2_2 = bufferStageEnqueueData_3[95:64];
  wire [31:0]       dataRegroupBySew_3_2_3 = bufferStageEnqueueData_3[127:96];
  wire [31:0]       dataRegroupBySew_3_2_4 = bufferStageEnqueueData_3[159:128];
  wire [31:0]       dataRegroupBySew_3_2_5 = bufferStageEnqueueData_3[191:160];
  wire [31:0]       dataRegroupBySew_3_2_6 = bufferStageEnqueueData_3[223:192];
  wire [31:0]       dataRegroupBySew_3_2_7 = bufferStageEnqueueData_3[255:224];
  wire [31:0]       dataRegroupBySew_3_2_8 = bufferStageEnqueueData_3[287:256];
  wire [31:0]       dataRegroupBySew_3_2_9 = bufferStageEnqueueData_3[319:288];
  wire [31:0]       dataRegroupBySew_3_2_10 = bufferStageEnqueueData_3[351:320];
  wire [31:0]       dataRegroupBySew_3_2_11 = bufferStageEnqueueData_3[383:352];
  wire [31:0]       dataRegroupBySew_3_2_12 = bufferStageEnqueueData_3[415:384];
  wire [31:0]       dataRegroupBySew_3_2_13 = bufferStageEnqueueData_3[447:416];
  wire [31:0]       dataRegroupBySew_3_2_14 = bufferStageEnqueueData_3[479:448];
  wire [31:0]       dataRegroupBySew_3_2_15 = bufferStageEnqueueData_3[511:480];
  wire [31:0]       dataRegroupBySew_3_2_16 = bufferStageEnqueueData_3[543:512];
  wire [31:0]       dataRegroupBySew_3_2_17 = bufferStageEnqueueData_3[575:544];
  wire [31:0]       dataRegroupBySew_3_2_18 = bufferStageEnqueueData_3[607:576];
  wire [31:0]       dataRegroupBySew_3_2_19 = bufferStageEnqueueData_3[639:608];
  wire [31:0]       dataRegroupBySew_3_2_20 = bufferStageEnqueueData_3[671:640];
  wire [31:0]       dataRegroupBySew_3_2_21 = bufferStageEnqueueData_3[703:672];
  wire [31:0]       dataRegroupBySew_3_2_22 = bufferStageEnqueueData_3[735:704];
  wire [31:0]       dataRegroupBySew_3_2_23 = bufferStageEnqueueData_3[767:736];
  wire [31:0]       dataRegroupBySew_3_2_24 = bufferStageEnqueueData_3[799:768];
  wire [31:0]       dataRegroupBySew_3_2_25 = bufferStageEnqueueData_3[831:800];
  wire [31:0]       dataRegroupBySew_3_2_26 = bufferStageEnqueueData_3[863:832];
  wire [31:0]       dataRegroupBySew_3_2_27 = bufferStageEnqueueData_3[895:864];
  wire [31:0]       dataRegroupBySew_3_2_28 = bufferStageEnqueueData_3[927:896];
  wire [31:0]       dataRegroupBySew_3_2_29 = bufferStageEnqueueData_3[959:928];
  wire [31:0]       dataRegroupBySew_3_2_30 = bufferStageEnqueueData_3[991:960];
  wire [31:0]       dataRegroupBySew_3_2_31 = bufferStageEnqueueData_3[1023:992];
  wire [31:0]       dataRegroupBySew_4_2_0 = bufferStageEnqueueData_4[31:0];
  wire [31:0]       dataRegroupBySew_4_2_1 = bufferStageEnqueueData_4[63:32];
  wire [31:0]       dataRegroupBySew_4_2_2 = bufferStageEnqueueData_4[95:64];
  wire [31:0]       dataRegroupBySew_4_2_3 = bufferStageEnqueueData_4[127:96];
  wire [31:0]       dataRegroupBySew_4_2_4 = bufferStageEnqueueData_4[159:128];
  wire [31:0]       dataRegroupBySew_4_2_5 = bufferStageEnqueueData_4[191:160];
  wire [31:0]       dataRegroupBySew_4_2_6 = bufferStageEnqueueData_4[223:192];
  wire [31:0]       dataRegroupBySew_4_2_7 = bufferStageEnqueueData_4[255:224];
  wire [31:0]       dataRegroupBySew_4_2_8 = bufferStageEnqueueData_4[287:256];
  wire [31:0]       dataRegroupBySew_4_2_9 = bufferStageEnqueueData_4[319:288];
  wire [31:0]       dataRegroupBySew_4_2_10 = bufferStageEnqueueData_4[351:320];
  wire [31:0]       dataRegroupBySew_4_2_11 = bufferStageEnqueueData_4[383:352];
  wire [31:0]       dataRegroupBySew_4_2_12 = bufferStageEnqueueData_4[415:384];
  wire [31:0]       dataRegroupBySew_4_2_13 = bufferStageEnqueueData_4[447:416];
  wire [31:0]       dataRegroupBySew_4_2_14 = bufferStageEnqueueData_4[479:448];
  wire [31:0]       dataRegroupBySew_4_2_15 = bufferStageEnqueueData_4[511:480];
  wire [31:0]       dataRegroupBySew_4_2_16 = bufferStageEnqueueData_4[543:512];
  wire [31:0]       dataRegroupBySew_4_2_17 = bufferStageEnqueueData_4[575:544];
  wire [31:0]       dataRegroupBySew_4_2_18 = bufferStageEnqueueData_4[607:576];
  wire [31:0]       dataRegroupBySew_4_2_19 = bufferStageEnqueueData_4[639:608];
  wire [31:0]       dataRegroupBySew_4_2_20 = bufferStageEnqueueData_4[671:640];
  wire [31:0]       dataRegroupBySew_4_2_21 = bufferStageEnqueueData_4[703:672];
  wire [31:0]       dataRegroupBySew_4_2_22 = bufferStageEnqueueData_4[735:704];
  wire [31:0]       dataRegroupBySew_4_2_23 = bufferStageEnqueueData_4[767:736];
  wire [31:0]       dataRegroupBySew_4_2_24 = bufferStageEnqueueData_4[799:768];
  wire [31:0]       dataRegroupBySew_4_2_25 = bufferStageEnqueueData_4[831:800];
  wire [31:0]       dataRegroupBySew_4_2_26 = bufferStageEnqueueData_4[863:832];
  wire [31:0]       dataRegroupBySew_4_2_27 = bufferStageEnqueueData_4[895:864];
  wire [31:0]       dataRegroupBySew_4_2_28 = bufferStageEnqueueData_4[927:896];
  wire [31:0]       dataRegroupBySew_4_2_29 = bufferStageEnqueueData_4[959:928];
  wire [31:0]       dataRegroupBySew_4_2_30 = bufferStageEnqueueData_4[991:960];
  wire [31:0]       dataRegroupBySew_4_2_31 = bufferStageEnqueueData_4[1023:992];
  wire [31:0]       dataRegroupBySew_5_2_0 = bufferStageEnqueueData_5[31:0];
  wire [31:0]       dataRegroupBySew_5_2_1 = bufferStageEnqueueData_5[63:32];
  wire [31:0]       dataRegroupBySew_5_2_2 = bufferStageEnqueueData_5[95:64];
  wire [31:0]       dataRegroupBySew_5_2_3 = bufferStageEnqueueData_5[127:96];
  wire [31:0]       dataRegroupBySew_5_2_4 = bufferStageEnqueueData_5[159:128];
  wire [31:0]       dataRegroupBySew_5_2_5 = bufferStageEnqueueData_5[191:160];
  wire [31:0]       dataRegroupBySew_5_2_6 = bufferStageEnqueueData_5[223:192];
  wire [31:0]       dataRegroupBySew_5_2_7 = bufferStageEnqueueData_5[255:224];
  wire [31:0]       dataRegroupBySew_5_2_8 = bufferStageEnqueueData_5[287:256];
  wire [31:0]       dataRegroupBySew_5_2_9 = bufferStageEnqueueData_5[319:288];
  wire [31:0]       dataRegroupBySew_5_2_10 = bufferStageEnqueueData_5[351:320];
  wire [31:0]       dataRegroupBySew_5_2_11 = bufferStageEnqueueData_5[383:352];
  wire [31:0]       dataRegroupBySew_5_2_12 = bufferStageEnqueueData_5[415:384];
  wire [31:0]       dataRegroupBySew_5_2_13 = bufferStageEnqueueData_5[447:416];
  wire [31:0]       dataRegroupBySew_5_2_14 = bufferStageEnqueueData_5[479:448];
  wire [31:0]       dataRegroupBySew_5_2_15 = bufferStageEnqueueData_5[511:480];
  wire [31:0]       dataRegroupBySew_5_2_16 = bufferStageEnqueueData_5[543:512];
  wire [31:0]       dataRegroupBySew_5_2_17 = bufferStageEnqueueData_5[575:544];
  wire [31:0]       dataRegroupBySew_5_2_18 = bufferStageEnqueueData_5[607:576];
  wire [31:0]       dataRegroupBySew_5_2_19 = bufferStageEnqueueData_5[639:608];
  wire [31:0]       dataRegroupBySew_5_2_20 = bufferStageEnqueueData_5[671:640];
  wire [31:0]       dataRegroupBySew_5_2_21 = bufferStageEnqueueData_5[703:672];
  wire [31:0]       dataRegroupBySew_5_2_22 = bufferStageEnqueueData_5[735:704];
  wire [31:0]       dataRegroupBySew_5_2_23 = bufferStageEnqueueData_5[767:736];
  wire [31:0]       dataRegroupBySew_5_2_24 = bufferStageEnqueueData_5[799:768];
  wire [31:0]       dataRegroupBySew_5_2_25 = bufferStageEnqueueData_5[831:800];
  wire [31:0]       dataRegroupBySew_5_2_26 = bufferStageEnqueueData_5[863:832];
  wire [31:0]       dataRegroupBySew_5_2_27 = bufferStageEnqueueData_5[895:864];
  wire [31:0]       dataRegroupBySew_5_2_28 = bufferStageEnqueueData_5[927:896];
  wire [31:0]       dataRegroupBySew_5_2_29 = bufferStageEnqueueData_5[959:928];
  wire [31:0]       dataRegroupBySew_5_2_30 = bufferStageEnqueueData_5[991:960];
  wire [31:0]       dataRegroupBySew_5_2_31 = bufferStageEnqueueData_5[1023:992];
  wire [31:0]       dataRegroupBySew_6_2_0 = bufferStageEnqueueData_6[31:0];
  wire [31:0]       dataRegroupBySew_6_2_1 = bufferStageEnqueueData_6[63:32];
  wire [31:0]       dataRegroupBySew_6_2_2 = bufferStageEnqueueData_6[95:64];
  wire [31:0]       dataRegroupBySew_6_2_3 = bufferStageEnqueueData_6[127:96];
  wire [31:0]       dataRegroupBySew_6_2_4 = bufferStageEnqueueData_6[159:128];
  wire [31:0]       dataRegroupBySew_6_2_5 = bufferStageEnqueueData_6[191:160];
  wire [31:0]       dataRegroupBySew_6_2_6 = bufferStageEnqueueData_6[223:192];
  wire [31:0]       dataRegroupBySew_6_2_7 = bufferStageEnqueueData_6[255:224];
  wire [31:0]       dataRegroupBySew_6_2_8 = bufferStageEnqueueData_6[287:256];
  wire [31:0]       dataRegroupBySew_6_2_9 = bufferStageEnqueueData_6[319:288];
  wire [31:0]       dataRegroupBySew_6_2_10 = bufferStageEnqueueData_6[351:320];
  wire [31:0]       dataRegroupBySew_6_2_11 = bufferStageEnqueueData_6[383:352];
  wire [31:0]       dataRegroupBySew_6_2_12 = bufferStageEnqueueData_6[415:384];
  wire [31:0]       dataRegroupBySew_6_2_13 = bufferStageEnqueueData_6[447:416];
  wire [31:0]       dataRegroupBySew_6_2_14 = bufferStageEnqueueData_6[479:448];
  wire [31:0]       dataRegroupBySew_6_2_15 = bufferStageEnqueueData_6[511:480];
  wire [31:0]       dataRegroupBySew_6_2_16 = bufferStageEnqueueData_6[543:512];
  wire [31:0]       dataRegroupBySew_6_2_17 = bufferStageEnqueueData_6[575:544];
  wire [31:0]       dataRegroupBySew_6_2_18 = bufferStageEnqueueData_6[607:576];
  wire [31:0]       dataRegroupBySew_6_2_19 = bufferStageEnqueueData_6[639:608];
  wire [31:0]       dataRegroupBySew_6_2_20 = bufferStageEnqueueData_6[671:640];
  wire [31:0]       dataRegroupBySew_6_2_21 = bufferStageEnqueueData_6[703:672];
  wire [31:0]       dataRegroupBySew_6_2_22 = bufferStageEnqueueData_6[735:704];
  wire [31:0]       dataRegroupBySew_6_2_23 = bufferStageEnqueueData_6[767:736];
  wire [31:0]       dataRegroupBySew_6_2_24 = bufferStageEnqueueData_6[799:768];
  wire [31:0]       dataRegroupBySew_6_2_25 = bufferStageEnqueueData_6[831:800];
  wire [31:0]       dataRegroupBySew_6_2_26 = bufferStageEnqueueData_6[863:832];
  wire [31:0]       dataRegroupBySew_6_2_27 = bufferStageEnqueueData_6[895:864];
  wire [31:0]       dataRegroupBySew_6_2_28 = bufferStageEnqueueData_6[927:896];
  wire [31:0]       dataRegroupBySew_6_2_29 = bufferStageEnqueueData_6[959:928];
  wire [31:0]       dataRegroupBySew_6_2_30 = bufferStageEnqueueData_6[991:960];
  wire [31:0]       dataRegroupBySew_6_2_31 = bufferStageEnqueueData_6[1023:992];
  wire [31:0]       dataRegroupBySew_7_2_0 = bufferStageEnqueueData_7[31:0];
  wire [31:0]       dataRegroupBySew_7_2_1 = bufferStageEnqueueData_7[63:32];
  wire [31:0]       dataRegroupBySew_7_2_2 = bufferStageEnqueueData_7[95:64];
  wire [31:0]       dataRegroupBySew_7_2_3 = bufferStageEnqueueData_7[127:96];
  wire [31:0]       dataRegroupBySew_7_2_4 = bufferStageEnqueueData_7[159:128];
  wire [31:0]       dataRegroupBySew_7_2_5 = bufferStageEnqueueData_7[191:160];
  wire [31:0]       dataRegroupBySew_7_2_6 = bufferStageEnqueueData_7[223:192];
  wire [31:0]       dataRegroupBySew_7_2_7 = bufferStageEnqueueData_7[255:224];
  wire [31:0]       dataRegroupBySew_7_2_8 = bufferStageEnqueueData_7[287:256];
  wire [31:0]       dataRegroupBySew_7_2_9 = bufferStageEnqueueData_7[319:288];
  wire [31:0]       dataRegroupBySew_7_2_10 = bufferStageEnqueueData_7[351:320];
  wire [31:0]       dataRegroupBySew_7_2_11 = bufferStageEnqueueData_7[383:352];
  wire [31:0]       dataRegroupBySew_7_2_12 = bufferStageEnqueueData_7[415:384];
  wire [31:0]       dataRegroupBySew_7_2_13 = bufferStageEnqueueData_7[447:416];
  wire [31:0]       dataRegroupBySew_7_2_14 = bufferStageEnqueueData_7[479:448];
  wire [31:0]       dataRegroupBySew_7_2_15 = bufferStageEnqueueData_7[511:480];
  wire [31:0]       dataRegroupBySew_7_2_16 = bufferStageEnqueueData_7[543:512];
  wire [31:0]       dataRegroupBySew_7_2_17 = bufferStageEnqueueData_7[575:544];
  wire [31:0]       dataRegroupBySew_7_2_18 = bufferStageEnqueueData_7[607:576];
  wire [31:0]       dataRegroupBySew_7_2_19 = bufferStageEnqueueData_7[639:608];
  wire [31:0]       dataRegroupBySew_7_2_20 = bufferStageEnqueueData_7[671:640];
  wire [31:0]       dataRegroupBySew_7_2_21 = bufferStageEnqueueData_7[703:672];
  wire [31:0]       dataRegroupBySew_7_2_22 = bufferStageEnqueueData_7[735:704];
  wire [31:0]       dataRegroupBySew_7_2_23 = bufferStageEnqueueData_7[767:736];
  wire [31:0]       dataRegroupBySew_7_2_24 = bufferStageEnqueueData_7[799:768];
  wire [31:0]       dataRegroupBySew_7_2_25 = bufferStageEnqueueData_7[831:800];
  wire [31:0]       dataRegroupBySew_7_2_26 = bufferStageEnqueueData_7[863:832];
  wire [31:0]       dataRegroupBySew_7_2_27 = bufferStageEnqueueData_7[895:864];
  wire [31:0]       dataRegroupBySew_7_2_28 = bufferStageEnqueueData_7[927:896];
  wire [31:0]       dataRegroupBySew_7_2_29 = bufferStageEnqueueData_7[959:928];
  wire [31:0]       dataRegroupBySew_7_2_30 = bufferStageEnqueueData_7[991:960];
  wire [31:0]       dataRegroupBySew_7_2_31 = bufferStageEnqueueData_7[1023:992];
  wire [63:0]       dataInMem_lo_lo_lo_lo_16 = {dataRegroupBySew_0_2_1, dataRegroupBySew_0_2_0};
  wire [63:0]       dataInMem_lo_lo_lo_hi_16 = {dataRegroupBySew_0_2_3, dataRegroupBySew_0_2_2};
  wire [127:0]      dataInMem_lo_lo_lo_16 = {dataInMem_lo_lo_lo_hi_16, dataInMem_lo_lo_lo_lo_16};
  wire [63:0]       dataInMem_lo_lo_hi_lo_16 = {dataRegroupBySew_0_2_5, dataRegroupBySew_0_2_4};
  wire [63:0]       dataInMem_lo_lo_hi_hi_16 = {dataRegroupBySew_0_2_7, dataRegroupBySew_0_2_6};
  wire [127:0]      dataInMem_lo_lo_hi_16 = {dataInMem_lo_lo_hi_hi_16, dataInMem_lo_lo_hi_lo_16};
  wire [255:0]      dataInMem_lo_lo_208 = {dataInMem_lo_lo_hi_16, dataInMem_lo_lo_lo_16};
  wire [63:0]       dataInMem_lo_hi_lo_lo_16 = {dataRegroupBySew_0_2_9, dataRegroupBySew_0_2_8};
  wire [63:0]       dataInMem_lo_hi_lo_hi_16 = {dataRegroupBySew_0_2_11, dataRegroupBySew_0_2_10};
  wire [127:0]      dataInMem_lo_hi_lo_16 = {dataInMem_lo_hi_lo_hi_16, dataInMem_lo_hi_lo_lo_16};
  wire [63:0]       dataInMem_lo_hi_hi_lo_16 = {dataRegroupBySew_0_2_13, dataRegroupBySew_0_2_12};
  wire [63:0]       dataInMem_lo_hi_hi_hi_16 = {dataRegroupBySew_0_2_15, dataRegroupBySew_0_2_14};
  wire [127:0]      dataInMem_lo_hi_hi_16 = {dataInMem_lo_hi_hi_hi_16, dataInMem_lo_hi_hi_lo_16};
  wire [255:0]      dataInMem_lo_hi_592 = {dataInMem_lo_hi_hi_16, dataInMem_lo_hi_lo_16};
  wire [511:0]      dataInMem_lo_976 = {dataInMem_lo_hi_592, dataInMem_lo_lo_208};
  wire [63:0]       dataInMem_hi_lo_lo_lo_16 = {dataRegroupBySew_0_2_17, dataRegroupBySew_0_2_16};
  wire [63:0]       dataInMem_hi_lo_lo_hi_16 = {dataRegroupBySew_0_2_19, dataRegroupBySew_0_2_18};
  wire [127:0]      dataInMem_hi_lo_lo_16 = {dataInMem_hi_lo_lo_hi_16, dataInMem_hi_lo_lo_lo_16};
  wire [63:0]       dataInMem_hi_lo_hi_lo_16 = {dataRegroupBySew_0_2_21, dataRegroupBySew_0_2_20};
  wire [63:0]       dataInMem_hi_lo_hi_hi_16 = {dataRegroupBySew_0_2_23, dataRegroupBySew_0_2_22};
  wire [127:0]      dataInMem_hi_lo_hi_16 = {dataInMem_hi_lo_hi_hi_16, dataInMem_hi_lo_hi_lo_16};
  wire [255:0]      dataInMem_hi_lo_400 = {dataInMem_hi_lo_hi_16, dataInMem_hi_lo_lo_16};
  wire [63:0]       dataInMem_hi_hi_lo_lo_16 = {dataRegroupBySew_0_2_25, dataRegroupBySew_0_2_24};
  wire [63:0]       dataInMem_hi_hi_lo_hi_16 = {dataRegroupBySew_0_2_27, dataRegroupBySew_0_2_26};
  wire [127:0]      dataInMem_hi_hi_lo_16 = {dataInMem_hi_hi_lo_hi_16, dataInMem_hi_hi_lo_lo_16};
  wire [63:0]       dataInMem_hi_hi_hi_lo_16 = {dataRegroupBySew_0_2_29, dataRegroupBySew_0_2_28};
  wire [63:0]       dataInMem_hi_hi_hi_hi_16 = {dataRegroupBySew_0_2_31, dataRegroupBySew_0_2_30};
  wire [127:0]      dataInMem_hi_hi_hi_16 = {dataInMem_hi_hi_hi_hi_16, dataInMem_hi_hi_hi_lo_16};
  wire [255:0]      dataInMem_hi_hi_784 = {dataInMem_hi_hi_hi_16, dataInMem_hi_hi_lo_16};
  wire [511:0]      dataInMem_hi_1168 = {dataInMem_hi_hi_784, dataInMem_hi_lo_400};
  wire [1023:0]     dataInMem_16 = {dataInMem_hi_1168, dataInMem_lo_976};
  wire [1023:0]     regroupCacheLine_16_0 = dataInMem_16;
  wire [1023:0]     res_128 = regroupCacheLine_16_0;
  wire [2047:0]     lo_lo_16 = {1024'h0, res_128};
  wire [4095:0]     lo_16 = {2048'h0, lo_lo_16};
  wire [8191:0]     regroupLoadData_2_0 = {4096'h0, lo_16};
  wire [127:0]      dataInMem_lo_lo_lo_lo_17 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1, dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [127:0]      dataInMem_lo_lo_lo_hi_17 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3, dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [255:0]      dataInMem_lo_lo_lo_17 = {dataInMem_lo_lo_lo_hi_17, dataInMem_lo_lo_lo_lo_17};
  wire [127:0]      dataInMem_lo_lo_hi_lo_17 = {dataRegroupBySew_1_2_5, dataRegroupBySew_0_2_5, dataRegroupBySew_1_2_4, dataRegroupBySew_0_2_4};
  wire [127:0]      dataInMem_lo_lo_hi_hi_17 = {dataRegroupBySew_1_2_7, dataRegroupBySew_0_2_7, dataRegroupBySew_1_2_6, dataRegroupBySew_0_2_6};
  wire [255:0]      dataInMem_lo_lo_hi_17 = {dataInMem_lo_lo_hi_hi_17, dataInMem_lo_lo_hi_lo_17};
  wire [511:0]      dataInMem_lo_lo_209 = {dataInMem_lo_lo_hi_17, dataInMem_lo_lo_lo_17};
  wire [127:0]      dataInMem_lo_hi_lo_lo_17 = {dataRegroupBySew_1_2_9, dataRegroupBySew_0_2_9, dataRegroupBySew_1_2_8, dataRegroupBySew_0_2_8};
  wire [127:0]      dataInMem_lo_hi_lo_hi_17 = {dataRegroupBySew_1_2_11, dataRegroupBySew_0_2_11, dataRegroupBySew_1_2_10, dataRegroupBySew_0_2_10};
  wire [255:0]      dataInMem_lo_hi_lo_17 = {dataInMem_lo_hi_lo_hi_17, dataInMem_lo_hi_lo_lo_17};
  wire [127:0]      dataInMem_lo_hi_hi_lo_17 = {dataRegroupBySew_1_2_13, dataRegroupBySew_0_2_13, dataRegroupBySew_1_2_12, dataRegroupBySew_0_2_12};
  wire [127:0]      dataInMem_lo_hi_hi_hi_17 = {dataRegroupBySew_1_2_15, dataRegroupBySew_0_2_15, dataRegroupBySew_1_2_14, dataRegroupBySew_0_2_14};
  wire [255:0]      dataInMem_lo_hi_hi_17 = {dataInMem_lo_hi_hi_hi_17, dataInMem_lo_hi_hi_lo_17};
  wire [511:0]      dataInMem_lo_hi_593 = {dataInMem_lo_hi_hi_17, dataInMem_lo_hi_lo_17};
  wire [1023:0]     dataInMem_lo_977 = {dataInMem_lo_hi_593, dataInMem_lo_lo_209};
  wire [127:0]      dataInMem_hi_lo_lo_lo_17 = {dataRegroupBySew_1_2_17, dataRegroupBySew_0_2_17, dataRegroupBySew_1_2_16, dataRegroupBySew_0_2_16};
  wire [127:0]      dataInMem_hi_lo_lo_hi_17 = {dataRegroupBySew_1_2_19, dataRegroupBySew_0_2_19, dataRegroupBySew_1_2_18, dataRegroupBySew_0_2_18};
  wire [255:0]      dataInMem_hi_lo_lo_17 = {dataInMem_hi_lo_lo_hi_17, dataInMem_hi_lo_lo_lo_17};
  wire [127:0]      dataInMem_hi_lo_hi_lo_17 = {dataRegroupBySew_1_2_21, dataRegroupBySew_0_2_21, dataRegroupBySew_1_2_20, dataRegroupBySew_0_2_20};
  wire [127:0]      dataInMem_hi_lo_hi_hi_17 = {dataRegroupBySew_1_2_23, dataRegroupBySew_0_2_23, dataRegroupBySew_1_2_22, dataRegroupBySew_0_2_22};
  wire [255:0]      dataInMem_hi_lo_hi_17 = {dataInMem_hi_lo_hi_hi_17, dataInMem_hi_lo_hi_lo_17};
  wire [511:0]      dataInMem_hi_lo_401 = {dataInMem_hi_lo_hi_17, dataInMem_hi_lo_lo_17};
  wire [127:0]      dataInMem_hi_hi_lo_lo_17 = {dataRegroupBySew_1_2_25, dataRegroupBySew_0_2_25, dataRegroupBySew_1_2_24, dataRegroupBySew_0_2_24};
  wire [127:0]      dataInMem_hi_hi_lo_hi_17 = {dataRegroupBySew_1_2_27, dataRegroupBySew_0_2_27, dataRegroupBySew_1_2_26, dataRegroupBySew_0_2_26};
  wire [255:0]      dataInMem_hi_hi_lo_17 = {dataInMem_hi_hi_lo_hi_17, dataInMem_hi_hi_lo_lo_17};
  wire [127:0]      dataInMem_hi_hi_hi_lo_17 = {dataRegroupBySew_1_2_29, dataRegroupBySew_0_2_29, dataRegroupBySew_1_2_28, dataRegroupBySew_0_2_28};
  wire [127:0]      dataInMem_hi_hi_hi_hi_17 = {dataRegroupBySew_1_2_31, dataRegroupBySew_0_2_31, dataRegroupBySew_1_2_30, dataRegroupBySew_0_2_30};
  wire [255:0]      dataInMem_hi_hi_hi_17 = {dataInMem_hi_hi_hi_hi_17, dataInMem_hi_hi_hi_lo_17};
  wire [511:0]      dataInMem_hi_hi_785 = {dataInMem_hi_hi_hi_17, dataInMem_hi_hi_lo_17};
  wire [1023:0]     dataInMem_hi_1169 = {dataInMem_hi_hi_785, dataInMem_hi_lo_401};
  wire [2047:0]     dataInMem_17 = {dataInMem_hi_1169, dataInMem_lo_977};
  wire [1023:0]     regroupCacheLine_17_0 = dataInMem_17[1023:0];
  wire [1023:0]     regroupCacheLine_17_1 = dataInMem_17[2047:1024];
  wire [1023:0]     res_136 = regroupCacheLine_17_0;
  wire [1023:0]     res_137 = regroupCacheLine_17_1;
  wire [2047:0]     lo_lo_17 = {res_137, res_136};
  wire [4095:0]     lo_17 = {2048'h0, lo_lo_17};
  wire [8191:0]     regroupLoadData_2_1 = {4096'h0, lo_17};
  wire [63:0]       _GEN_966 = {dataRegroupBySew_2_2_0, dataRegroupBySew_1_2_0};
  wire [63:0]       dataInMem_hi_1170;
  assign dataInMem_hi_1170 = _GEN_966;
  wire [63:0]       dataInMem_lo_hi_597;
  assign dataInMem_lo_hi_597 = _GEN_966;
  wire [63:0]       dataInMem_lo_hi_630;
  assign dataInMem_lo_hi_630 = _GEN_966;
  wire [63:0]       _GEN_967 = {dataRegroupBySew_2_2_1, dataRegroupBySew_1_2_1};
  wire [63:0]       dataInMem_hi_1171;
  assign dataInMem_hi_1171 = _GEN_967;
  wire [63:0]       dataInMem_lo_hi_598;
  assign dataInMem_lo_hi_598 = _GEN_967;
  wire [63:0]       dataInMem_lo_hi_631;
  assign dataInMem_lo_hi_631 = _GEN_967;
  wire [63:0]       _GEN_968 = {dataRegroupBySew_2_2_2, dataRegroupBySew_1_2_2};
  wire [63:0]       dataInMem_hi_1172;
  assign dataInMem_hi_1172 = _GEN_968;
  wire [63:0]       dataInMem_lo_hi_599;
  assign dataInMem_lo_hi_599 = _GEN_968;
  wire [63:0]       dataInMem_lo_hi_632;
  assign dataInMem_lo_hi_632 = _GEN_968;
  wire [63:0]       _GEN_969 = {dataRegroupBySew_2_2_3, dataRegroupBySew_1_2_3};
  wire [63:0]       dataInMem_hi_1173;
  assign dataInMem_hi_1173 = _GEN_969;
  wire [63:0]       dataInMem_lo_hi_600;
  assign dataInMem_lo_hi_600 = _GEN_969;
  wire [63:0]       dataInMem_lo_hi_633;
  assign dataInMem_lo_hi_633 = _GEN_969;
  wire [63:0]       _GEN_970 = {dataRegroupBySew_2_2_4, dataRegroupBySew_1_2_4};
  wire [63:0]       dataInMem_hi_1174;
  assign dataInMem_hi_1174 = _GEN_970;
  wire [63:0]       dataInMem_lo_hi_601;
  assign dataInMem_lo_hi_601 = _GEN_970;
  wire [63:0]       dataInMem_lo_hi_634;
  assign dataInMem_lo_hi_634 = _GEN_970;
  wire [63:0]       _GEN_971 = {dataRegroupBySew_2_2_5, dataRegroupBySew_1_2_5};
  wire [63:0]       dataInMem_hi_1175;
  assign dataInMem_hi_1175 = _GEN_971;
  wire [63:0]       dataInMem_lo_hi_602;
  assign dataInMem_lo_hi_602 = _GEN_971;
  wire [63:0]       dataInMem_lo_hi_635;
  assign dataInMem_lo_hi_635 = _GEN_971;
  wire [63:0]       _GEN_972 = {dataRegroupBySew_2_2_6, dataRegroupBySew_1_2_6};
  wire [63:0]       dataInMem_hi_1176;
  assign dataInMem_hi_1176 = _GEN_972;
  wire [63:0]       dataInMem_lo_hi_603;
  assign dataInMem_lo_hi_603 = _GEN_972;
  wire [63:0]       dataInMem_lo_hi_636;
  assign dataInMem_lo_hi_636 = _GEN_972;
  wire [63:0]       _GEN_973 = {dataRegroupBySew_2_2_7, dataRegroupBySew_1_2_7};
  wire [63:0]       dataInMem_hi_1177;
  assign dataInMem_hi_1177 = _GEN_973;
  wire [63:0]       dataInMem_lo_hi_604;
  assign dataInMem_lo_hi_604 = _GEN_973;
  wire [63:0]       dataInMem_lo_hi_637;
  assign dataInMem_lo_hi_637 = _GEN_973;
  wire [63:0]       _GEN_974 = {dataRegroupBySew_2_2_8, dataRegroupBySew_1_2_8};
  wire [63:0]       dataInMem_hi_1178;
  assign dataInMem_hi_1178 = _GEN_974;
  wire [63:0]       dataInMem_lo_hi_605;
  assign dataInMem_lo_hi_605 = _GEN_974;
  wire [63:0]       dataInMem_lo_hi_638;
  assign dataInMem_lo_hi_638 = _GEN_974;
  wire [63:0]       _GEN_975 = {dataRegroupBySew_2_2_9, dataRegroupBySew_1_2_9};
  wire [63:0]       dataInMem_hi_1179;
  assign dataInMem_hi_1179 = _GEN_975;
  wire [63:0]       dataInMem_lo_hi_606;
  assign dataInMem_lo_hi_606 = _GEN_975;
  wire [63:0]       dataInMem_lo_hi_639;
  assign dataInMem_lo_hi_639 = _GEN_975;
  wire [63:0]       _GEN_976 = {dataRegroupBySew_2_2_10, dataRegroupBySew_1_2_10};
  wire [63:0]       dataInMem_hi_1180;
  assign dataInMem_hi_1180 = _GEN_976;
  wire [63:0]       dataInMem_lo_hi_607;
  assign dataInMem_lo_hi_607 = _GEN_976;
  wire [63:0]       dataInMem_lo_hi_640;
  assign dataInMem_lo_hi_640 = _GEN_976;
  wire [63:0]       _GEN_977 = {dataRegroupBySew_2_2_11, dataRegroupBySew_1_2_11};
  wire [63:0]       dataInMem_hi_1181;
  assign dataInMem_hi_1181 = _GEN_977;
  wire [63:0]       dataInMem_lo_hi_608;
  assign dataInMem_lo_hi_608 = _GEN_977;
  wire [63:0]       dataInMem_lo_hi_641;
  assign dataInMem_lo_hi_641 = _GEN_977;
  wire [63:0]       _GEN_978 = {dataRegroupBySew_2_2_12, dataRegroupBySew_1_2_12};
  wire [63:0]       dataInMem_hi_1182;
  assign dataInMem_hi_1182 = _GEN_978;
  wire [63:0]       dataInMem_lo_hi_609;
  assign dataInMem_lo_hi_609 = _GEN_978;
  wire [63:0]       dataInMem_lo_hi_642;
  assign dataInMem_lo_hi_642 = _GEN_978;
  wire [63:0]       _GEN_979 = {dataRegroupBySew_2_2_13, dataRegroupBySew_1_2_13};
  wire [63:0]       dataInMem_hi_1183;
  assign dataInMem_hi_1183 = _GEN_979;
  wire [63:0]       dataInMem_lo_hi_610;
  assign dataInMem_lo_hi_610 = _GEN_979;
  wire [63:0]       dataInMem_lo_hi_643;
  assign dataInMem_lo_hi_643 = _GEN_979;
  wire [63:0]       _GEN_980 = {dataRegroupBySew_2_2_14, dataRegroupBySew_1_2_14};
  wire [63:0]       dataInMem_hi_1184;
  assign dataInMem_hi_1184 = _GEN_980;
  wire [63:0]       dataInMem_lo_hi_611;
  assign dataInMem_lo_hi_611 = _GEN_980;
  wire [63:0]       dataInMem_lo_hi_644;
  assign dataInMem_lo_hi_644 = _GEN_980;
  wire [63:0]       _GEN_981 = {dataRegroupBySew_2_2_15, dataRegroupBySew_1_2_15};
  wire [63:0]       dataInMem_hi_1185;
  assign dataInMem_hi_1185 = _GEN_981;
  wire [63:0]       dataInMem_lo_hi_612;
  assign dataInMem_lo_hi_612 = _GEN_981;
  wire [63:0]       dataInMem_lo_hi_645;
  assign dataInMem_lo_hi_645 = _GEN_981;
  wire [63:0]       _GEN_982 = {dataRegroupBySew_2_2_16, dataRegroupBySew_1_2_16};
  wire [63:0]       dataInMem_hi_1186;
  assign dataInMem_hi_1186 = _GEN_982;
  wire [63:0]       dataInMem_lo_hi_613;
  assign dataInMem_lo_hi_613 = _GEN_982;
  wire [63:0]       dataInMem_lo_hi_646;
  assign dataInMem_lo_hi_646 = _GEN_982;
  wire [63:0]       _GEN_983 = {dataRegroupBySew_2_2_17, dataRegroupBySew_1_2_17};
  wire [63:0]       dataInMem_hi_1187;
  assign dataInMem_hi_1187 = _GEN_983;
  wire [63:0]       dataInMem_lo_hi_614;
  assign dataInMem_lo_hi_614 = _GEN_983;
  wire [63:0]       dataInMem_lo_hi_647;
  assign dataInMem_lo_hi_647 = _GEN_983;
  wire [63:0]       _GEN_984 = {dataRegroupBySew_2_2_18, dataRegroupBySew_1_2_18};
  wire [63:0]       dataInMem_hi_1188;
  assign dataInMem_hi_1188 = _GEN_984;
  wire [63:0]       dataInMem_lo_hi_615;
  assign dataInMem_lo_hi_615 = _GEN_984;
  wire [63:0]       dataInMem_lo_hi_648;
  assign dataInMem_lo_hi_648 = _GEN_984;
  wire [63:0]       _GEN_985 = {dataRegroupBySew_2_2_19, dataRegroupBySew_1_2_19};
  wire [63:0]       dataInMem_hi_1189;
  assign dataInMem_hi_1189 = _GEN_985;
  wire [63:0]       dataInMem_lo_hi_616;
  assign dataInMem_lo_hi_616 = _GEN_985;
  wire [63:0]       dataInMem_lo_hi_649;
  assign dataInMem_lo_hi_649 = _GEN_985;
  wire [63:0]       _GEN_986 = {dataRegroupBySew_2_2_20, dataRegroupBySew_1_2_20};
  wire [63:0]       dataInMem_hi_1190;
  assign dataInMem_hi_1190 = _GEN_986;
  wire [63:0]       dataInMem_lo_hi_617;
  assign dataInMem_lo_hi_617 = _GEN_986;
  wire [63:0]       dataInMem_lo_hi_650;
  assign dataInMem_lo_hi_650 = _GEN_986;
  wire [63:0]       _GEN_987 = {dataRegroupBySew_2_2_21, dataRegroupBySew_1_2_21};
  wire [63:0]       dataInMem_hi_1191;
  assign dataInMem_hi_1191 = _GEN_987;
  wire [63:0]       dataInMem_lo_hi_618;
  assign dataInMem_lo_hi_618 = _GEN_987;
  wire [63:0]       dataInMem_lo_hi_651;
  assign dataInMem_lo_hi_651 = _GEN_987;
  wire [63:0]       _GEN_988 = {dataRegroupBySew_2_2_22, dataRegroupBySew_1_2_22};
  wire [63:0]       dataInMem_hi_1192;
  assign dataInMem_hi_1192 = _GEN_988;
  wire [63:0]       dataInMem_lo_hi_619;
  assign dataInMem_lo_hi_619 = _GEN_988;
  wire [63:0]       dataInMem_lo_hi_652;
  assign dataInMem_lo_hi_652 = _GEN_988;
  wire [63:0]       _GEN_989 = {dataRegroupBySew_2_2_23, dataRegroupBySew_1_2_23};
  wire [63:0]       dataInMem_hi_1193;
  assign dataInMem_hi_1193 = _GEN_989;
  wire [63:0]       dataInMem_lo_hi_620;
  assign dataInMem_lo_hi_620 = _GEN_989;
  wire [63:0]       dataInMem_lo_hi_653;
  assign dataInMem_lo_hi_653 = _GEN_989;
  wire [63:0]       _GEN_990 = {dataRegroupBySew_2_2_24, dataRegroupBySew_1_2_24};
  wire [63:0]       dataInMem_hi_1194;
  assign dataInMem_hi_1194 = _GEN_990;
  wire [63:0]       dataInMem_lo_hi_621;
  assign dataInMem_lo_hi_621 = _GEN_990;
  wire [63:0]       dataInMem_lo_hi_654;
  assign dataInMem_lo_hi_654 = _GEN_990;
  wire [63:0]       _GEN_991 = {dataRegroupBySew_2_2_25, dataRegroupBySew_1_2_25};
  wire [63:0]       dataInMem_hi_1195;
  assign dataInMem_hi_1195 = _GEN_991;
  wire [63:0]       dataInMem_lo_hi_622;
  assign dataInMem_lo_hi_622 = _GEN_991;
  wire [63:0]       dataInMem_lo_hi_655;
  assign dataInMem_lo_hi_655 = _GEN_991;
  wire [63:0]       _GEN_992 = {dataRegroupBySew_2_2_26, dataRegroupBySew_1_2_26};
  wire [63:0]       dataInMem_hi_1196;
  assign dataInMem_hi_1196 = _GEN_992;
  wire [63:0]       dataInMem_lo_hi_623;
  assign dataInMem_lo_hi_623 = _GEN_992;
  wire [63:0]       dataInMem_lo_hi_656;
  assign dataInMem_lo_hi_656 = _GEN_992;
  wire [63:0]       _GEN_993 = {dataRegroupBySew_2_2_27, dataRegroupBySew_1_2_27};
  wire [63:0]       dataInMem_hi_1197;
  assign dataInMem_hi_1197 = _GEN_993;
  wire [63:0]       dataInMem_lo_hi_624;
  assign dataInMem_lo_hi_624 = _GEN_993;
  wire [63:0]       dataInMem_lo_hi_657;
  assign dataInMem_lo_hi_657 = _GEN_993;
  wire [63:0]       _GEN_994 = {dataRegroupBySew_2_2_28, dataRegroupBySew_1_2_28};
  wire [63:0]       dataInMem_hi_1198;
  assign dataInMem_hi_1198 = _GEN_994;
  wire [63:0]       dataInMem_lo_hi_625;
  assign dataInMem_lo_hi_625 = _GEN_994;
  wire [63:0]       dataInMem_lo_hi_658;
  assign dataInMem_lo_hi_658 = _GEN_994;
  wire [63:0]       _GEN_995 = {dataRegroupBySew_2_2_29, dataRegroupBySew_1_2_29};
  wire [63:0]       dataInMem_hi_1199;
  assign dataInMem_hi_1199 = _GEN_995;
  wire [63:0]       dataInMem_lo_hi_626;
  assign dataInMem_lo_hi_626 = _GEN_995;
  wire [63:0]       dataInMem_lo_hi_659;
  assign dataInMem_lo_hi_659 = _GEN_995;
  wire [63:0]       _GEN_996 = {dataRegroupBySew_2_2_30, dataRegroupBySew_1_2_30};
  wire [63:0]       dataInMem_hi_1200;
  assign dataInMem_hi_1200 = _GEN_996;
  wire [63:0]       dataInMem_lo_hi_627;
  assign dataInMem_lo_hi_627 = _GEN_996;
  wire [63:0]       dataInMem_lo_hi_660;
  assign dataInMem_lo_hi_660 = _GEN_996;
  wire [63:0]       _GEN_997 = {dataRegroupBySew_2_2_31, dataRegroupBySew_1_2_31};
  wire [63:0]       dataInMem_hi_1201;
  assign dataInMem_hi_1201 = _GEN_997;
  wire [63:0]       dataInMem_lo_hi_628;
  assign dataInMem_lo_hi_628 = _GEN_997;
  wire [63:0]       dataInMem_lo_hi_661;
  assign dataInMem_lo_hi_661 = _GEN_997;
  wire [191:0]      dataInMem_lo_lo_lo_lo_18 = {dataInMem_hi_1171, dataRegroupBySew_0_2_1, dataInMem_hi_1170, dataRegroupBySew_0_2_0};
  wire [191:0]      dataInMem_lo_lo_lo_hi_18 = {dataInMem_hi_1173, dataRegroupBySew_0_2_3, dataInMem_hi_1172, dataRegroupBySew_0_2_2};
  wire [383:0]      dataInMem_lo_lo_lo_18 = {dataInMem_lo_lo_lo_hi_18, dataInMem_lo_lo_lo_lo_18};
  wire [191:0]      dataInMem_lo_lo_hi_lo_18 = {dataInMem_hi_1175, dataRegroupBySew_0_2_5, dataInMem_hi_1174, dataRegroupBySew_0_2_4};
  wire [191:0]      dataInMem_lo_lo_hi_hi_18 = {dataInMem_hi_1177, dataRegroupBySew_0_2_7, dataInMem_hi_1176, dataRegroupBySew_0_2_6};
  wire [383:0]      dataInMem_lo_lo_hi_18 = {dataInMem_lo_lo_hi_hi_18, dataInMem_lo_lo_hi_lo_18};
  wire [767:0]      dataInMem_lo_lo_210 = {dataInMem_lo_lo_hi_18, dataInMem_lo_lo_lo_18};
  wire [191:0]      dataInMem_lo_hi_lo_lo_18 = {dataInMem_hi_1179, dataRegroupBySew_0_2_9, dataInMem_hi_1178, dataRegroupBySew_0_2_8};
  wire [191:0]      dataInMem_lo_hi_lo_hi_18 = {dataInMem_hi_1181, dataRegroupBySew_0_2_11, dataInMem_hi_1180, dataRegroupBySew_0_2_10};
  wire [383:0]      dataInMem_lo_hi_lo_18 = {dataInMem_lo_hi_lo_hi_18, dataInMem_lo_hi_lo_lo_18};
  wire [191:0]      dataInMem_lo_hi_hi_lo_18 = {dataInMem_hi_1183, dataRegroupBySew_0_2_13, dataInMem_hi_1182, dataRegroupBySew_0_2_12};
  wire [191:0]      dataInMem_lo_hi_hi_hi_18 = {dataInMem_hi_1185, dataRegroupBySew_0_2_15, dataInMem_hi_1184, dataRegroupBySew_0_2_14};
  wire [383:0]      dataInMem_lo_hi_hi_18 = {dataInMem_lo_hi_hi_hi_18, dataInMem_lo_hi_hi_lo_18};
  wire [767:0]      dataInMem_lo_hi_594 = {dataInMem_lo_hi_hi_18, dataInMem_lo_hi_lo_18};
  wire [1535:0]     dataInMem_lo_978 = {dataInMem_lo_hi_594, dataInMem_lo_lo_210};
  wire [191:0]      dataInMem_hi_lo_lo_lo_18 = {dataInMem_hi_1187, dataRegroupBySew_0_2_17, dataInMem_hi_1186, dataRegroupBySew_0_2_16};
  wire [191:0]      dataInMem_hi_lo_lo_hi_18 = {dataInMem_hi_1189, dataRegroupBySew_0_2_19, dataInMem_hi_1188, dataRegroupBySew_0_2_18};
  wire [383:0]      dataInMem_hi_lo_lo_18 = {dataInMem_hi_lo_lo_hi_18, dataInMem_hi_lo_lo_lo_18};
  wire [191:0]      dataInMem_hi_lo_hi_lo_18 = {dataInMem_hi_1191, dataRegroupBySew_0_2_21, dataInMem_hi_1190, dataRegroupBySew_0_2_20};
  wire [191:0]      dataInMem_hi_lo_hi_hi_18 = {dataInMem_hi_1193, dataRegroupBySew_0_2_23, dataInMem_hi_1192, dataRegroupBySew_0_2_22};
  wire [383:0]      dataInMem_hi_lo_hi_18 = {dataInMem_hi_lo_hi_hi_18, dataInMem_hi_lo_hi_lo_18};
  wire [767:0]      dataInMem_hi_lo_402 = {dataInMem_hi_lo_hi_18, dataInMem_hi_lo_lo_18};
  wire [191:0]      dataInMem_hi_hi_lo_lo_18 = {dataInMem_hi_1195, dataRegroupBySew_0_2_25, dataInMem_hi_1194, dataRegroupBySew_0_2_24};
  wire [191:0]      dataInMem_hi_hi_lo_hi_18 = {dataInMem_hi_1197, dataRegroupBySew_0_2_27, dataInMem_hi_1196, dataRegroupBySew_0_2_26};
  wire [383:0]      dataInMem_hi_hi_lo_18 = {dataInMem_hi_hi_lo_hi_18, dataInMem_hi_hi_lo_lo_18};
  wire [191:0]      dataInMem_hi_hi_hi_lo_18 = {dataInMem_hi_1199, dataRegroupBySew_0_2_29, dataInMem_hi_1198, dataRegroupBySew_0_2_28};
  wire [191:0]      dataInMem_hi_hi_hi_hi_18 = {dataInMem_hi_1201, dataRegroupBySew_0_2_31, dataInMem_hi_1200, dataRegroupBySew_0_2_30};
  wire [383:0]      dataInMem_hi_hi_hi_18 = {dataInMem_hi_hi_hi_hi_18, dataInMem_hi_hi_hi_lo_18};
  wire [767:0]      dataInMem_hi_hi_786 = {dataInMem_hi_hi_hi_18, dataInMem_hi_hi_lo_18};
  wire [1535:0]     dataInMem_hi_1202 = {dataInMem_hi_hi_786, dataInMem_hi_lo_402};
  wire [3071:0]     dataInMem_18 = {dataInMem_hi_1202, dataInMem_lo_978};
  wire [1023:0]     regroupCacheLine_18_0 = dataInMem_18[1023:0];
  wire [1023:0]     regroupCacheLine_18_1 = dataInMem_18[2047:1024];
  wire [1023:0]     regroupCacheLine_18_2 = dataInMem_18[3071:2048];
  wire [1023:0]     res_144 = regroupCacheLine_18_0;
  wire [1023:0]     res_145 = regroupCacheLine_18_1;
  wire [1023:0]     res_146 = regroupCacheLine_18_2;
  wire [2047:0]     lo_lo_18 = {res_145, res_144};
  wire [2047:0]     lo_hi_18 = {1024'h0, res_146};
  wire [4095:0]     lo_18 = {lo_hi_18, lo_lo_18};
  wire [8191:0]     regroupLoadData_2_2 = {4096'h0, lo_18};
  wire [63:0]       _GEN_998 = {dataRegroupBySew_1_2_0, dataRegroupBySew_0_2_0};
  wire [63:0]       dataInMem_lo_979;
  assign dataInMem_lo_979 = _GEN_998;
  wire [63:0]       dataInMem_lo_1012;
  assign dataInMem_lo_1012 = _GEN_998;
  wire [63:0]       dataInMem_lo_lo_215;
  assign dataInMem_lo_lo_215 = _GEN_998;
  wire [63:0]       _GEN_999 = {dataRegroupBySew_3_2_0, dataRegroupBySew_2_2_0};
  wire [63:0]       dataInMem_hi_1203;
  assign dataInMem_hi_1203 = _GEN_999;
  wire [63:0]       dataInMem_lo_hi_663;
  assign dataInMem_lo_hi_663 = _GEN_999;
  wire [63:0]       _GEN_1000 = {dataRegroupBySew_1_2_1, dataRegroupBySew_0_2_1};
  wire [63:0]       dataInMem_lo_980;
  assign dataInMem_lo_980 = _GEN_1000;
  wire [63:0]       dataInMem_lo_1013;
  assign dataInMem_lo_1013 = _GEN_1000;
  wire [63:0]       dataInMem_lo_lo_216;
  assign dataInMem_lo_lo_216 = _GEN_1000;
  wire [63:0]       _GEN_1001 = {dataRegroupBySew_3_2_1, dataRegroupBySew_2_2_1};
  wire [63:0]       dataInMem_hi_1204;
  assign dataInMem_hi_1204 = _GEN_1001;
  wire [63:0]       dataInMem_lo_hi_664;
  assign dataInMem_lo_hi_664 = _GEN_1001;
  wire [63:0]       _GEN_1002 = {dataRegroupBySew_1_2_2, dataRegroupBySew_0_2_2};
  wire [63:0]       dataInMem_lo_981;
  assign dataInMem_lo_981 = _GEN_1002;
  wire [63:0]       dataInMem_lo_1014;
  assign dataInMem_lo_1014 = _GEN_1002;
  wire [63:0]       dataInMem_lo_lo_217;
  assign dataInMem_lo_lo_217 = _GEN_1002;
  wire [63:0]       _GEN_1003 = {dataRegroupBySew_3_2_2, dataRegroupBySew_2_2_2};
  wire [63:0]       dataInMem_hi_1205;
  assign dataInMem_hi_1205 = _GEN_1003;
  wire [63:0]       dataInMem_lo_hi_665;
  assign dataInMem_lo_hi_665 = _GEN_1003;
  wire [63:0]       _GEN_1004 = {dataRegroupBySew_1_2_3, dataRegroupBySew_0_2_3};
  wire [63:0]       dataInMem_lo_982;
  assign dataInMem_lo_982 = _GEN_1004;
  wire [63:0]       dataInMem_lo_1015;
  assign dataInMem_lo_1015 = _GEN_1004;
  wire [63:0]       dataInMem_lo_lo_218;
  assign dataInMem_lo_lo_218 = _GEN_1004;
  wire [63:0]       _GEN_1005 = {dataRegroupBySew_3_2_3, dataRegroupBySew_2_2_3};
  wire [63:0]       dataInMem_hi_1206;
  assign dataInMem_hi_1206 = _GEN_1005;
  wire [63:0]       dataInMem_lo_hi_666;
  assign dataInMem_lo_hi_666 = _GEN_1005;
  wire [63:0]       _GEN_1006 = {dataRegroupBySew_1_2_4, dataRegroupBySew_0_2_4};
  wire [63:0]       dataInMem_lo_983;
  assign dataInMem_lo_983 = _GEN_1006;
  wire [63:0]       dataInMem_lo_1016;
  assign dataInMem_lo_1016 = _GEN_1006;
  wire [63:0]       dataInMem_lo_lo_219;
  assign dataInMem_lo_lo_219 = _GEN_1006;
  wire [63:0]       _GEN_1007 = {dataRegroupBySew_3_2_4, dataRegroupBySew_2_2_4};
  wire [63:0]       dataInMem_hi_1207;
  assign dataInMem_hi_1207 = _GEN_1007;
  wire [63:0]       dataInMem_lo_hi_667;
  assign dataInMem_lo_hi_667 = _GEN_1007;
  wire [63:0]       _GEN_1008 = {dataRegroupBySew_1_2_5, dataRegroupBySew_0_2_5};
  wire [63:0]       dataInMem_lo_984;
  assign dataInMem_lo_984 = _GEN_1008;
  wire [63:0]       dataInMem_lo_1017;
  assign dataInMem_lo_1017 = _GEN_1008;
  wire [63:0]       dataInMem_lo_lo_220;
  assign dataInMem_lo_lo_220 = _GEN_1008;
  wire [63:0]       _GEN_1009 = {dataRegroupBySew_3_2_5, dataRegroupBySew_2_2_5};
  wire [63:0]       dataInMem_hi_1208;
  assign dataInMem_hi_1208 = _GEN_1009;
  wire [63:0]       dataInMem_lo_hi_668;
  assign dataInMem_lo_hi_668 = _GEN_1009;
  wire [63:0]       _GEN_1010 = {dataRegroupBySew_1_2_6, dataRegroupBySew_0_2_6};
  wire [63:0]       dataInMem_lo_985;
  assign dataInMem_lo_985 = _GEN_1010;
  wire [63:0]       dataInMem_lo_1018;
  assign dataInMem_lo_1018 = _GEN_1010;
  wire [63:0]       dataInMem_lo_lo_221;
  assign dataInMem_lo_lo_221 = _GEN_1010;
  wire [63:0]       _GEN_1011 = {dataRegroupBySew_3_2_6, dataRegroupBySew_2_2_6};
  wire [63:0]       dataInMem_hi_1209;
  assign dataInMem_hi_1209 = _GEN_1011;
  wire [63:0]       dataInMem_lo_hi_669;
  assign dataInMem_lo_hi_669 = _GEN_1011;
  wire [63:0]       _GEN_1012 = {dataRegroupBySew_1_2_7, dataRegroupBySew_0_2_7};
  wire [63:0]       dataInMem_lo_986;
  assign dataInMem_lo_986 = _GEN_1012;
  wire [63:0]       dataInMem_lo_1019;
  assign dataInMem_lo_1019 = _GEN_1012;
  wire [63:0]       dataInMem_lo_lo_222;
  assign dataInMem_lo_lo_222 = _GEN_1012;
  wire [63:0]       _GEN_1013 = {dataRegroupBySew_3_2_7, dataRegroupBySew_2_2_7};
  wire [63:0]       dataInMem_hi_1210;
  assign dataInMem_hi_1210 = _GEN_1013;
  wire [63:0]       dataInMem_lo_hi_670;
  assign dataInMem_lo_hi_670 = _GEN_1013;
  wire [63:0]       _GEN_1014 = {dataRegroupBySew_1_2_8, dataRegroupBySew_0_2_8};
  wire [63:0]       dataInMem_lo_987;
  assign dataInMem_lo_987 = _GEN_1014;
  wire [63:0]       dataInMem_lo_1020;
  assign dataInMem_lo_1020 = _GEN_1014;
  wire [63:0]       dataInMem_lo_lo_223;
  assign dataInMem_lo_lo_223 = _GEN_1014;
  wire [63:0]       _GEN_1015 = {dataRegroupBySew_3_2_8, dataRegroupBySew_2_2_8};
  wire [63:0]       dataInMem_hi_1211;
  assign dataInMem_hi_1211 = _GEN_1015;
  wire [63:0]       dataInMem_lo_hi_671;
  assign dataInMem_lo_hi_671 = _GEN_1015;
  wire [63:0]       _GEN_1016 = {dataRegroupBySew_1_2_9, dataRegroupBySew_0_2_9};
  wire [63:0]       dataInMem_lo_988;
  assign dataInMem_lo_988 = _GEN_1016;
  wire [63:0]       dataInMem_lo_1021;
  assign dataInMem_lo_1021 = _GEN_1016;
  wire [63:0]       dataInMem_lo_lo_224;
  assign dataInMem_lo_lo_224 = _GEN_1016;
  wire [63:0]       _GEN_1017 = {dataRegroupBySew_3_2_9, dataRegroupBySew_2_2_9};
  wire [63:0]       dataInMem_hi_1212;
  assign dataInMem_hi_1212 = _GEN_1017;
  wire [63:0]       dataInMem_lo_hi_672;
  assign dataInMem_lo_hi_672 = _GEN_1017;
  wire [63:0]       _GEN_1018 = {dataRegroupBySew_1_2_10, dataRegroupBySew_0_2_10};
  wire [63:0]       dataInMem_lo_989;
  assign dataInMem_lo_989 = _GEN_1018;
  wire [63:0]       dataInMem_lo_1022;
  assign dataInMem_lo_1022 = _GEN_1018;
  wire [63:0]       dataInMem_lo_lo_225;
  assign dataInMem_lo_lo_225 = _GEN_1018;
  wire [63:0]       _GEN_1019 = {dataRegroupBySew_3_2_10, dataRegroupBySew_2_2_10};
  wire [63:0]       dataInMem_hi_1213;
  assign dataInMem_hi_1213 = _GEN_1019;
  wire [63:0]       dataInMem_lo_hi_673;
  assign dataInMem_lo_hi_673 = _GEN_1019;
  wire [63:0]       _GEN_1020 = {dataRegroupBySew_1_2_11, dataRegroupBySew_0_2_11};
  wire [63:0]       dataInMem_lo_990;
  assign dataInMem_lo_990 = _GEN_1020;
  wire [63:0]       dataInMem_lo_1023;
  assign dataInMem_lo_1023 = _GEN_1020;
  wire [63:0]       dataInMem_lo_lo_226;
  assign dataInMem_lo_lo_226 = _GEN_1020;
  wire [63:0]       _GEN_1021 = {dataRegroupBySew_3_2_11, dataRegroupBySew_2_2_11};
  wire [63:0]       dataInMem_hi_1214;
  assign dataInMem_hi_1214 = _GEN_1021;
  wire [63:0]       dataInMem_lo_hi_674;
  assign dataInMem_lo_hi_674 = _GEN_1021;
  wire [63:0]       _GEN_1022 = {dataRegroupBySew_1_2_12, dataRegroupBySew_0_2_12};
  wire [63:0]       dataInMem_lo_991;
  assign dataInMem_lo_991 = _GEN_1022;
  wire [63:0]       dataInMem_lo_1024;
  assign dataInMem_lo_1024 = _GEN_1022;
  wire [63:0]       dataInMem_lo_lo_227;
  assign dataInMem_lo_lo_227 = _GEN_1022;
  wire [63:0]       _GEN_1023 = {dataRegroupBySew_3_2_12, dataRegroupBySew_2_2_12};
  wire [63:0]       dataInMem_hi_1215;
  assign dataInMem_hi_1215 = _GEN_1023;
  wire [63:0]       dataInMem_lo_hi_675;
  assign dataInMem_lo_hi_675 = _GEN_1023;
  wire [63:0]       _GEN_1024 = {dataRegroupBySew_1_2_13, dataRegroupBySew_0_2_13};
  wire [63:0]       dataInMem_lo_992;
  assign dataInMem_lo_992 = _GEN_1024;
  wire [63:0]       dataInMem_lo_1025;
  assign dataInMem_lo_1025 = _GEN_1024;
  wire [63:0]       dataInMem_lo_lo_228;
  assign dataInMem_lo_lo_228 = _GEN_1024;
  wire [63:0]       _GEN_1025 = {dataRegroupBySew_3_2_13, dataRegroupBySew_2_2_13};
  wire [63:0]       dataInMem_hi_1216;
  assign dataInMem_hi_1216 = _GEN_1025;
  wire [63:0]       dataInMem_lo_hi_676;
  assign dataInMem_lo_hi_676 = _GEN_1025;
  wire [63:0]       _GEN_1026 = {dataRegroupBySew_1_2_14, dataRegroupBySew_0_2_14};
  wire [63:0]       dataInMem_lo_993;
  assign dataInMem_lo_993 = _GEN_1026;
  wire [63:0]       dataInMem_lo_1026;
  assign dataInMem_lo_1026 = _GEN_1026;
  wire [63:0]       dataInMem_lo_lo_229;
  assign dataInMem_lo_lo_229 = _GEN_1026;
  wire [63:0]       _GEN_1027 = {dataRegroupBySew_3_2_14, dataRegroupBySew_2_2_14};
  wire [63:0]       dataInMem_hi_1217;
  assign dataInMem_hi_1217 = _GEN_1027;
  wire [63:0]       dataInMem_lo_hi_677;
  assign dataInMem_lo_hi_677 = _GEN_1027;
  wire [63:0]       _GEN_1028 = {dataRegroupBySew_1_2_15, dataRegroupBySew_0_2_15};
  wire [63:0]       dataInMem_lo_994;
  assign dataInMem_lo_994 = _GEN_1028;
  wire [63:0]       dataInMem_lo_1027;
  assign dataInMem_lo_1027 = _GEN_1028;
  wire [63:0]       dataInMem_lo_lo_230;
  assign dataInMem_lo_lo_230 = _GEN_1028;
  wire [63:0]       _GEN_1029 = {dataRegroupBySew_3_2_15, dataRegroupBySew_2_2_15};
  wire [63:0]       dataInMem_hi_1218;
  assign dataInMem_hi_1218 = _GEN_1029;
  wire [63:0]       dataInMem_lo_hi_678;
  assign dataInMem_lo_hi_678 = _GEN_1029;
  wire [63:0]       _GEN_1030 = {dataRegroupBySew_1_2_16, dataRegroupBySew_0_2_16};
  wire [63:0]       dataInMem_lo_995;
  assign dataInMem_lo_995 = _GEN_1030;
  wire [63:0]       dataInMem_lo_1028;
  assign dataInMem_lo_1028 = _GEN_1030;
  wire [63:0]       dataInMem_lo_lo_231;
  assign dataInMem_lo_lo_231 = _GEN_1030;
  wire [63:0]       _GEN_1031 = {dataRegroupBySew_3_2_16, dataRegroupBySew_2_2_16};
  wire [63:0]       dataInMem_hi_1219;
  assign dataInMem_hi_1219 = _GEN_1031;
  wire [63:0]       dataInMem_lo_hi_679;
  assign dataInMem_lo_hi_679 = _GEN_1031;
  wire [63:0]       _GEN_1032 = {dataRegroupBySew_1_2_17, dataRegroupBySew_0_2_17};
  wire [63:0]       dataInMem_lo_996;
  assign dataInMem_lo_996 = _GEN_1032;
  wire [63:0]       dataInMem_lo_1029;
  assign dataInMem_lo_1029 = _GEN_1032;
  wire [63:0]       dataInMem_lo_lo_232;
  assign dataInMem_lo_lo_232 = _GEN_1032;
  wire [63:0]       _GEN_1033 = {dataRegroupBySew_3_2_17, dataRegroupBySew_2_2_17};
  wire [63:0]       dataInMem_hi_1220;
  assign dataInMem_hi_1220 = _GEN_1033;
  wire [63:0]       dataInMem_lo_hi_680;
  assign dataInMem_lo_hi_680 = _GEN_1033;
  wire [63:0]       _GEN_1034 = {dataRegroupBySew_1_2_18, dataRegroupBySew_0_2_18};
  wire [63:0]       dataInMem_lo_997;
  assign dataInMem_lo_997 = _GEN_1034;
  wire [63:0]       dataInMem_lo_1030;
  assign dataInMem_lo_1030 = _GEN_1034;
  wire [63:0]       dataInMem_lo_lo_233;
  assign dataInMem_lo_lo_233 = _GEN_1034;
  wire [63:0]       _GEN_1035 = {dataRegroupBySew_3_2_18, dataRegroupBySew_2_2_18};
  wire [63:0]       dataInMem_hi_1221;
  assign dataInMem_hi_1221 = _GEN_1035;
  wire [63:0]       dataInMem_lo_hi_681;
  assign dataInMem_lo_hi_681 = _GEN_1035;
  wire [63:0]       _GEN_1036 = {dataRegroupBySew_1_2_19, dataRegroupBySew_0_2_19};
  wire [63:0]       dataInMem_lo_998;
  assign dataInMem_lo_998 = _GEN_1036;
  wire [63:0]       dataInMem_lo_1031;
  assign dataInMem_lo_1031 = _GEN_1036;
  wire [63:0]       dataInMem_lo_lo_234;
  assign dataInMem_lo_lo_234 = _GEN_1036;
  wire [63:0]       _GEN_1037 = {dataRegroupBySew_3_2_19, dataRegroupBySew_2_2_19};
  wire [63:0]       dataInMem_hi_1222;
  assign dataInMem_hi_1222 = _GEN_1037;
  wire [63:0]       dataInMem_lo_hi_682;
  assign dataInMem_lo_hi_682 = _GEN_1037;
  wire [63:0]       _GEN_1038 = {dataRegroupBySew_1_2_20, dataRegroupBySew_0_2_20};
  wire [63:0]       dataInMem_lo_999;
  assign dataInMem_lo_999 = _GEN_1038;
  wire [63:0]       dataInMem_lo_1032;
  assign dataInMem_lo_1032 = _GEN_1038;
  wire [63:0]       dataInMem_lo_lo_235;
  assign dataInMem_lo_lo_235 = _GEN_1038;
  wire [63:0]       _GEN_1039 = {dataRegroupBySew_3_2_20, dataRegroupBySew_2_2_20};
  wire [63:0]       dataInMem_hi_1223;
  assign dataInMem_hi_1223 = _GEN_1039;
  wire [63:0]       dataInMem_lo_hi_683;
  assign dataInMem_lo_hi_683 = _GEN_1039;
  wire [63:0]       _GEN_1040 = {dataRegroupBySew_1_2_21, dataRegroupBySew_0_2_21};
  wire [63:0]       dataInMem_lo_1000;
  assign dataInMem_lo_1000 = _GEN_1040;
  wire [63:0]       dataInMem_lo_1033;
  assign dataInMem_lo_1033 = _GEN_1040;
  wire [63:0]       dataInMem_lo_lo_236;
  assign dataInMem_lo_lo_236 = _GEN_1040;
  wire [63:0]       _GEN_1041 = {dataRegroupBySew_3_2_21, dataRegroupBySew_2_2_21};
  wire [63:0]       dataInMem_hi_1224;
  assign dataInMem_hi_1224 = _GEN_1041;
  wire [63:0]       dataInMem_lo_hi_684;
  assign dataInMem_lo_hi_684 = _GEN_1041;
  wire [63:0]       _GEN_1042 = {dataRegroupBySew_1_2_22, dataRegroupBySew_0_2_22};
  wire [63:0]       dataInMem_lo_1001;
  assign dataInMem_lo_1001 = _GEN_1042;
  wire [63:0]       dataInMem_lo_1034;
  assign dataInMem_lo_1034 = _GEN_1042;
  wire [63:0]       dataInMem_lo_lo_237;
  assign dataInMem_lo_lo_237 = _GEN_1042;
  wire [63:0]       _GEN_1043 = {dataRegroupBySew_3_2_22, dataRegroupBySew_2_2_22};
  wire [63:0]       dataInMem_hi_1225;
  assign dataInMem_hi_1225 = _GEN_1043;
  wire [63:0]       dataInMem_lo_hi_685;
  assign dataInMem_lo_hi_685 = _GEN_1043;
  wire [63:0]       _GEN_1044 = {dataRegroupBySew_1_2_23, dataRegroupBySew_0_2_23};
  wire [63:0]       dataInMem_lo_1002;
  assign dataInMem_lo_1002 = _GEN_1044;
  wire [63:0]       dataInMem_lo_1035;
  assign dataInMem_lo_1035 = _GEN_1044;
  wire [63:0]       dataInMem_lo_lo_238;
  assign dataInMem_lo_lo_238 = _GEN_1044;
  wire [63:0]       _GEN_1045 = {dataRegroupBySew_3_2_23, dataRegroupBySew_2_2_23};
  wire [63:0]       dataInMem_hi_1226;
  assign dataInMem_hi_1226 = _GEN_1045;
  wire [63:0]       dataInMem_lo_hi_686;
  assign dataInMem_lo_hi_686 = _GEN_1045;
  wire [63:0]       _GEN_1046 = {dataRegroupBySew_1_2_24, dataRegroupBySew_0_2_24};
  wire [63:0]       dataInMem_lo_1003;
  assign dataInMem_lo_1003 = _GEN_1046;
  wire [63:0]       dataInMem_lo_1036;
  assign dataInMem_lo_1036 = _GEN_1046;
  wire [63:0]       dataInMem_lo_lo_239;
  assign dataInMem_lo_lo_239 = _GEN_1046;
  wire [63:0]       _GEN_1047 = {dataRegroupBySew_3_2_24, dataRegroupBySew_2_2_24};
  wire [63:0]       dataInMem_hi_1227;
  assign dataInMem_hi_1227 = _GEN_1047;
  wire [63:0]       dataInMem_lo_hi_687;
  assign dataInMem_lo_hi_687 = _GEN_1047;
  wire [63:0]       _GEN_1048 = {dataRegroupBySew_1_2_25, dataRegroupBySew_0_2_25};
  wire [63:0]       dataInMem_lo_1004;
  assign dataInMem_lo_1004 = _GEN_1048;
  wire [63:0]       dataInMem_lo_1037;
  assign dataInMem_lo_1037 = _GEN_1048;
  wire [63:0]       dataInMem_lo_lo_240;
  assign dataInMem_lo_lo_240 = _GEN_1048;
  wire [63:0]       _GEN_1049 = {dataRegroupBySew_3_2_25, dataRegroupBySew_2_2_25};
  wire [63:0]       dataInMem_hi_1228;
  assign dataInMem_hi_1228 = _GEN_1049;
  wire [63:0]       dataInMem_lo_hi_688;
  assign dataInMem_lo_hi_688 = _GEN_1049;
  wire [63:0]       _GEN_1050 = {dataRegroupBySew_1_2_26, dataRegroupBySew_0_2_26};
  wire [63:0]       dataInMem_lo_1005;
  assign dataInMem_lo_1005 = _GEN_1050;
  wire [63:0]       dataInMem_lo_1038;
  assign dataInMem_lo_1038 = _GEN_1050;
  wire [63:0]       dataInMem_lo_lo_241;
  assign dataInMem_lo_lo_241 = _GEN_1050;
  wire [63:0]       _GEN_1051 = {dataRegroupBySew_3_2_26, dataRegroupBySew_2_2_26};
  wire [63:0]       dataInMem_hi_1229;
  assign dataInMem_hi_1229 = _GEN_1051;
  wire [63:0]       dataInMem_lo_hi_689;
  assign dataInMem_lo_hi_689 = _GEN_1051;
  wire [63:0]       _GEN_1052 = {dataRegroupBySew_1_2_27, dataRegroupBySew_0_2_27};
  wire [63:0]       dataInMem_lo_1006;
  assign dataInMem_lo_1006 = _GEN_1052;
  wire [63:0]       dataInMem_lo_1039;
  assign dataInMem_lo_1039 = _GEN_1052;
  wire [63:0]       dataInMem_lo_lo_242;
  assign dataInMem_lo_lo_242 = _GEN_1052;
  wire [63:0]       _GEN_1053 = {dataRegroupBySew_3_2_27, dataRegroupBySew_2_2_27};
  wire [63:0]       dataInMem_hi_1230;
  assign dataInMem_hi_1230 = _GEN_1053;
  wire [63:0]       dataInMem_lo_hi_690;
  assign dataInMem_lo_hi_690 = _GEN_1053;
  wire [63:0]       _GEN_1054 = {dataRegroupBySew_1_2_28, dataRegroupBySew_0_2_28};
  wire [63:0]       dataInMem_lo_1007;
  assign dataInMem_lo_1007 = _GEN_1054;
  wire [63:0]       dataInMem_lo_1040;
  assign dataInMem_lo_1040 = _GEN_1054;
  wire [63:0]       dataInMem_lo_lo_243;
  assign dataInMem_lo_lo_243 = _GEN_1054;
  wire [63:0]       _GEN_1055 = {dataRegroupBySew_3_2_28, dataRegroupBySew_2_2_28};
  wire [63:0]       dataInMem_hi_1231;
  assign dataInMem_hi_1231 = _GEN_1055;
  wire [63:0]       dataInMem_lo_hi_691;
  assign dataInMem_lo_hi_691 = _GEN_1055;
  wire [63:0]       _GEN_1056 = {dataRegroupBySew_1_2_29, dataRegroupBySew_0_2_29};
  wire [63:0]       dataInMem_lo_1008;
  assign dataInMem_lo_1008 = _GEN_1056;
  wire [63:0]       dataInMem_lo_1041;
  assign dataInMem_lo_1041 = _GEN_1056;
  wire [63:0]       dataInMem_lo_lo_244;
  assign dataInMem_lo_lo_244 = _GEN_1056;
  wire [63:0]       _GEN_1057 = {dataRegroupBySew_3_2_29, dataRegroupBySew_2_2_29};
  wire [63:0]       dataInMem_hi_1232;
  assign dataInMem_hi_1232 = _GEN_1057;
  wire [63:0]       dataInMem_lo_hi_692;
  assign dataInMem_lo_hi_692 = _GEN_1057;
  wire [63:0]       _GEN_1058 = {dataRegroupBySew_1_2_30, dataRegroupBySew_0_2_30};
  wire [63:0]       dataInMem_lo_1009;
  assign dataInMem_lo_1009 = _GEN_1058;
  wire [63:0]       dataInMem_lo_1042;
  assign dataInMem_lo_1042 = _GEN_1058;
  wire [63:0]       dataInMem_lo_lo_245;
  assign dataInMem_lo_lo_245 = _GEN_1058;
  wire [63:0]       _GEN_1059 = {dataRegroupBySew_3_2_30, dataRegroupBySew_2_2_30};
  wire [63:0]       dataInMem_hi_1233;
  assign dataInMem_hi_1233 = _GEN_1059;
  wire [63:0]       dataInMem_lo_hi_693;
  assign dataInMem_lo_hi_693 = _GEN_1059;
  wire [63:0]       _GEN_1060 = {dataRegroupBySew_1_2_31, dataRegroupBySew_0_2_31};
  wire [63:0]       dataInMem_lo_1010;
  assign dataInMem_lo_1010 = _GEN_1060;
  wire [63:0]       dataInMem_lo_1043;
  assign dataInMem_lo_1043 = _GEN_1060;
  wire [63:0]       dataInMem_lo_lo_246;
  assign dataInMem_lo_lo_246 = _GEN_1060;
  wire [63:0]       _GEN_1061 = {dataRegroupBySew_3_2_31, dataRegroupBySew_2_2_31};
  wire [63:0]       dataInMem_hi_1234;
  assign dataInMem_hi_1234 = _GEN_1061;
  wire [63:0]       dataInMem_lo_hi_694;
  assign dataInMem_lo_hi_694 = _GEN_1061;
  wire [255:0]      dataInMem_lo_lo_lo_lo_19 = {dataInMem_hi_1204, dataInMem_lo_980, dataInMem_hi_1203, dataInMem_lo_979};
  wire [255:0]      dataInMem_lo_lo_lo_hi_19 = {dataInMem_hi_1206, dataInMem_lo_982, dataInMem_hi_1205, dataInMem_lo_981};
  wire [511:0]      dataInMem_lo_lo_lo_19 = {dataInMem_lo_lo_lo_hi_19, dataInMem_lo_lo_lo_lo_19};
  wire [255:0]      dataInMem_lo_lo_hi_lo_19 = {dataInMem_hi_1208, dataInMem_lo_984, dataInMem_hi_1207, dataInMem_lo_983};
  wire [255:0]      dataInMem_lo_lo_hi_hi_19 = {dataInMem_hi_1210, dataInMem_lo_986, dataInMem_hi_1209, dataInMem_lo_985};
  wire [511:0]      dataInMem_lo_lo_hi_19 = {dataInMem_lo_lo_hi_hi_19, dataInMem_lo_lo_hi_lo_19};
  wire [1023:0]     dataInMem_lo_lo_211 = {dataInMem_lo_lo_hi_19, dataInMem_lo_lo_lo_19};
  wire [255:0]      dataInMem_lo_hi_lo_lo_19 = {dataInMem_hi_1212, dataInMem_lo_988, dataInMem_hi_1211, dataInMem_lo_987};
  wire [255:0]      dataInMem_lo_hi_lo_hi_19 = {dataInMem_hi_1214, dataInMem_lo_990, dataInMem_hi_1213, dataInMem_lo_989};
  wire [511:0]      dataInMem_lo_hi_lo_19 = {dataInMem_lo_hi_lo_hi_19, dataInMem_lo_hi_lo_lo_19};
  wire [255:0]      dataInMem_lo_hi_hi_lo_19 = {dataInMem_hi_1216, dataInMem_lo_992, dataInMem_hi_1215, dataInMem_lo_991};
  wire [255:0]      dataInMem_lo_hi_hi_hi_19 = {dataInMem_hi_1218, dataInMem_lo_994, dataInMem_hi_1217, dataInMem_lo_993};
  wire [511:0]      dataInMem_lo_hi_hi_19 = {dataInMem_lo_hi_hi_hi_19, dataInMem_lo_hi_hi_lo_19};
  wire [1023:0]     dataInMem_lo_hi_595 = {dataInMem_lo_hi_hi_19, dataInMem_lo_hi_lo_19};
  wire [2047:0]     dataInMem_lo_1011 = {dataInMem_lo_hi_595, dataInMem_lo_lo_211};
  wire [255:0]      dataInMem_hi_lo_lo_lo_19 = {dataInMem_hi_1220, dataInMem_lo_996, dataInMem_hi_1219, dataInMem_lo_995};
  wire [255:0]      dataInMem_hi_lo_lo_hi_19 = {dataInMem_hi_1222, dataInMem_lo_998, dataInMem_hi_1221, dataInMem_lo_997};
  wire [511:0]      dataInMem_hi_lo_lo_19 = {dataInMem_hi_lo_lo_hi_19, dataInMem_hi_lo_lo_lo_19};
  wire [255:0]      dataInMem_hi_lo_hi_lo_19 = {dataInMem_hi_1224, dataInMem_lo_1000, dataInMem_hi_1223, dataInMem_lo_999};
  wire [255:0]      dataInMem_hi_lo_hi_hi_19 = {dataInMem_hi_1226, dataInMem_lo_1002, dataInMem_hi_1225, dataInMem_lo_1001};
  wire [511:0]      dataInMem_hi_lo_hi_19 = {dataInMem_hi_lo_hi_hi_19, dataInMem_hi_lo_hi_lo_19};
  wire [1023:0]     dataInMem_hi_lo_403 = {dataInMem_hi_lo_hi_19, dataInMem_hi_lo_lo_19};
  wire [255:0]      dataInMem_hi_hi_lo_lo_19 = {dataInMem_hi_1228, dataInMem_lo_1004, dataInMem_hi_1227, dataInMem_lo_1003};
  wire [255:0]      dataInMem_hi_hi_lo_hi_19 = {dataInMem_hi_1230, dataInMem_lo_1006, dataInMem_hi_1229, dataInMem_lo_1005};
  wire [511:0]      dataInMem_hi_hi_lo_19 = {dataInMem_hi_hi_lo_hi_19, dataInMem_hi_hi_lo_lo_19};
  wire [255:0]      dataInMem_hi_hi_hi_lo_19 = {dataInMem_hi_1232, dataInMem_lo_1008, dataInMem_hi_1231, dataInMem_lo_1007};
  wire [255:0]      dataInMem_hi_hi_hi_hi_19 = {dataInMem_hi_1234, dataInMem_lo_1010, dataInMem_hi_1233, dataInMem_lo_1009};
  wire [511:0]      dataInMem_hi_hi_hi_19 = {dataInMem_hi_hi_hi_hi_19, dataInMem_hi_hi_hi_lo_19};
  wire [1023:0]     dataInMem_hi_hi_787 = {dataInMem_hi_hi_hi_19, dataInMem_hi_hi_lo_19};
  wire [2047:0]     dataInMem_hi_1235 = {dataInMem_hi_hi_787, dataInMem_hi_lo_403};
  wire [4095:0]     dataInMem_19 = {dataInMem_hi_1235, dataInMem_lo_1011};
  wire [1023:0]     regroupCacheLine_19_0 = dataInMem_19[1023:0];
  wire [1023:0]     regroupCacheLine_19_1 = dataInMem_19[2047:1024];
  wire [1023:0]     regroupCacheLine_19_2 = dataInMem_19[3071:2048];
  wire [1023:0]     regroupCacheLine_19_3 = dataInMem_19[4095:3072];
  wire [1023:0]     res_152 = regroupCacheLine_19_0;
  wire [1023:0]     res_153 = regroupCacheLine_19_1;
  wire [1023:0]     res_154 = regroupCacheLine_19_2;
  wire [1023:0]     res_155 = regroupCacheLine_19_3;
  wire [2047:0]     lo_lo_19 = {res_153, res_152};
  wire [2047:0]     lo_hi_19 = {res_155, res_154};
  wire [4095:0]     lo_19 = {lo_hi_19, lo_lo_19};
  wire [8191:0]     regroupLoadData_2_3 = {4096'h0, lo_19};
  wire [63:0]       _GEN_1062 = {dataRegroupBySew_4_2_0, dataRegroupBySew_3_2_0};
  wire [63:0]       dataInMem_hi_hi_788;
  assign dataInMem_hi_hi_788 = _GEN_1062;
  wire [63:0]       dataInMem_hi_lo_406;
  assign dataInMem_hi_lo_406 = _GEN_1062;
  wire [95:0]       dataInMem_hi_1236 = {dataInMem_hi_hi_788, dataRegroupBySew_2_2_0};
  wire [63:0]       _GEN_1063 = {dataRegroupBySew_4_2_1, dataRegroupBySew_3_2_1};
  wire [63:0]       dataInMem_hi_hi_789;
  assign dataInMem_hi_hi_789 = _GEN_1063;
  wire [63:0]       dataInMem_hi_lo_407;
  assign dataInMem_hi_lo_407 = _GEN_1063;
  wire [95:0]       dataInMem_hi_1237 = {dataInMem_hi_hi_789, dataRegroupBySew_2_2_1};
  wire [63:0]       _GEN_1064 = {dataRegroupBySew_4_2_2, dataRegroupBySew_3_2_2};
  wire [63:0]       dataInMem_hi_hi_790;
  assign dataInMem_hi_hi_790 = _GEN_1064;
  wire [63:0]       dataInMem_hi_lo_408;
  assign dataInMem_hi_lo_408 = _GEN_1064;
  wire [95:0]       dataInMem_hi_1238 = {dataInMem_hi_hi_790, dataRegroupBySew_2_2_2};
  wire [63:0]       _GEN_1065 = {dataRegroupBySew_4_2_3, dataRegroupBySew_3_2_3};
  wire [63:0]       dataInMem_hi_hi_791;
  assign dataInMem_hi_hi_791 = _GEN_1065;
  wire [63:0]       dataInMem_hi_lo_409;
  assign dataInMem_hi_lo_409 = _GEN_1065;
  wire [95:0]       dataInMem_hi_1239 = {dataInMem_hi_hi_791, dataRegroupBySew_2_2_3};
  wire [63:0]       _GEN_1066 = {dataRegroupBySew_4_2_4, dataRegroupBySew_3_2_4};
  wire [63:0]       dataInMem_hi_hi_792;
  assign dataInMem_hi_hi_792 = _GEN_1066;
  wire [63:0]       dataInMem_hi_lo_410;
  assign dataInMem_hi_lo_410 = _GEN_1066;
  wire [95:0]       dataInMem_hi_1240 = {dataInMem_hi_hi_792, dataRegroupBySew_2_2_4};
  wire [63:0]       _GEN_1067 = {dataRegroupBySew_4_2_5, dataRegroupBySew_3_2_5};
  wire [63:0]       dataInMem_hi_hi_793;
  assign dataInMem_hi_hi_793 = _GEN_1067;
  wire [63:0]       dataInMem_hi_lo_411;
  assign dataInMem_hi_lo_411 = _GEN_1067;
  wire [95:0]       dataInMem_hi_1241 = {dataInMem_hi_hi_793, dataRegroupBySew_2_2_5};
  wire [63:0]       _GEN_1068 = {dataRegroupBySew_4_2_6, dataRegroupBySew_3_2_6};
  wire [63:0]       dataInMem_hi_hi_794;
  assign dataInMem_hi_hi_794 = _GEN_1068;
  wire [63:0]       dataInMem_hi_lo_412;
  assign dataInMem_hi_lo_412 = _GEN_1068;
  wire [95:0]       dataInMem_hi_1242 = {dataInMem_hi_hi_794, dataRegroupBySew_2_2_6};
  wire [63:0]       _GEN_1069 = {dataRegroupBySew_4_2_7, dataRegroupBySew_3_2_7};
  wire [63:0]       dataInMem_hi_hi_795;
  assign dataInMem_hi_hi_795 = _GEN_1069;
  wire [63:0]       dataInMem_hi_lo_413;
  assign dataInMem_hi_lo_413 = _GEN_1069;
  wire [95:0]       dataInMem_hi_1243 = {dataInMem_hi_hi_795, dataRegroupBySew_2_2_7};
  wire [63:0]       _GEN_1070 = {dataRegroupBySew_4_2_8, dataRegroupBySew_3_2_8};
  wire [63:0]       dataInMem_hi_hi_796;
  assign dataInMem_hi_hi_796 = _GEN_1070;
  wire [63:0]       dataInMem_hi_lo_414;
  assign dataInMem_hi_lo_414 = _GEN_1070;
  wire [95:0]       dataInMem_hi_1244 = {dataInMem_hi_hi_796, dataRegroupBySew_2_2_8};
  wire [63:0]       _GEN_1071 = {dataRegroupBySew_4_2_9, dataRegroupBySew_3_2_9};
  wire [63:0]       dataInMem_hi_hi_797;
  assign dataInMem_hi_hi_797 = _GEN_1071;
  wire [63:0]       dataInMem_hi_lo_415;
  assign dataInMem_hi_lo_415 = _GEN_1071;
  wire [95:0]       dataInMem_hi_1245 = {dataInMem_hi_hi_797, dataRegroupBySew_2_2_9};
  wire [63:0]       _GEN_1072 = {dataRegroupBySew_4_2_10, dataRegroupBySew_3_2_10};
  wire [63:0]       dataInMem_hi_hi_798;
  assign dataInMem_hi_hi_798 = _GEN_1072;
  wire [63:0]       dataInMem_hi_lo_416;
  assign dataInMem_hi_lo_416 = _GEN_1072;
  wire [95:0]       dataInMem_hi_1246 = {dataInMem_hi_hi_798, dataRegroupBySew_2_2_10};
  wire [63:0]       _GEN_1073 = {dataRegroupBySew_4_2_11, dataRegroupBySew_3_2_11};
  wire [63:0]       dataInMem_hi_hi_799;
  assign dataInMem_hi_hi_799 = _GEN_1073;
  wire [63:0]       dataInMem_hi_lo_417;
  assign dataInMem_hi_lo_417 = _GEN_1073;
  wire [95:0]       dataInMem_hi_1247 = {dataInMem_hi_hi_799, dataRegroupBySew_2_2_11};
  wire [63:0]       _GEN_1074 = {dataRegroupBySew_4_2_12, dataRegroupBySew_3_2_12};
  wire [63:0]       dataInMem_hi_hi_800;
  assign dataInMem_hi_hi_800 = _GEN_1074;
  wire [63:0]       dataInMem_hi_lo_418;
  assign dataInMem_hi_lo_418 = _GEN_1074;
  wire [95:0]       dataInMem_hi_1248 = {dataInMem_hi_hi_800, dataRegroupBySew_2_2_12};
  wire [63:0]       _GEN_1075 = {dataRegroupBySew_4_2_13, dataRegroupBySew_3_2_13};
  wire [63:0]       dataInMem_hi_hi_801;
  assign dataInMem_hi_hi_801 = _GEN_1075;
  wire [63:0]       dataInMem_hi_lo_419;
  assign dataInMem_hi_lo_419 = _GEN_1075;
  wire [95:0]       dataInMem_hi_1249 = {dataInMem_hi_hi_801, dataRegroupBySew_2_2_13};
  wire [63:0]       _GEN_1076 = {dataRegroupBySew_4_2_14, dataRegroupBySew_3_2_14};
  wire [63:0]       dataInMem_hi_hi_802;
  assign dataInMem_hi_hi_802 = _GEN_1076;
  wire [63:0]       dataInMem_hi_lo_420;
  assign dataInMem_hi_lo_420 = _GEN_1076;
  wire [95:0]       dataInMem_hi_1250 = {dataInMem_hi_hi_802, dataRegroupBySew_2_2_14};
  wire [63:0]       _GEN_1077 = {dataRegroupBySew_4_2_15, dataRegroupBySew_3_2_15};
  wire [63:0]       dataInMem_hi_hi_803;
  assign dataInMem_hi_hi_803 = _GEN_1077;
  wire [63:0]       dataInMem_hi_lo_421;
  assign dataInMem_hi_lo_421 = _GEN_1077;
  wire [95:0]       dataInMem_hi_1251 = {dataInMem_hi_hi_803, dataRegroupBySew_2_2_15};
  wire [63:0]       _GEN_1078 = {dataRegroupBySew_4_2_16, dataRegroupBySew_3_2_16};
  wire [63:0]       dataInMem_hi_hi_804;
  assign dataInMem_hi_hi_804 = _GEN_1078;
  wire [63:0]       dataInMem_hi_lo_422;
  assign dataInMem_hi_lo_422 = _GEN_1078;
  wire [95:0]       dataInMem_hi_1252 = {dataInMem_hi_hi_804, dataRegroupBySew_2_2_16};
  wire [63:0]       _GEN_1079 = {dataRegroupBySew_4_2_17, dataRegroupBySew_3_2_17};
  wire [63:0]       dataInMem_hi_hi_805;
  assign dataInMem_hi_hi_805 = _GEN_1079;
  wire [63:0]       dataInMem_hi_lo_423;
  assign dataInMem_hi_lo_423 = _GEN_1079;
  wire [95:0]       dataInMem_hi_1253 = {dataInMem_hi_hi_805, dataRegroupBySew_2_2_17};
  wire [63:0]       _GEN_1080 = {dataRegroupBySew_4_2_18, dataRegroupBySew_3_2_18};
  wire [63:0]       dataInMem_hi_hi_806;
  assign dataInMem_hi_hi_806 = _GEN_1080;
  wire [63:0]       dataInMem_hi_lo_424;
  assign dataInMem_hi_lo_424 = _GEN_1080;
  wire [95:0]       dataInMem_hi_1254 = {dataInMem_hi_hi_806, dataRegroupBySew_2_2_18};
  wire [63:0]       _GEN_1081 = {dataRegroupBySew_4_2_19, dataRegroupBySew_3_2_19};
  wire [63:0]       dataInMem_hi_hi_807;
  assign dataInMem_hi_hi_807 = _GEN_1081;
  wire [63:0]       dataInMem_hi_lo_425;
  assign dataInMem_hi_lo_425 = _GEN_1081;
  wire [95:0]       dataInMem_hi_1255 = {dataInMem_hi_hi_807, dataRegroupBySew_2_2_19};
  wire [63:0]       _GEN_1082 = {dataRegroupBySew_4_2_20, dataRegroupBySew_3_2_20};
  wire [63:0]       dataInMem_hi_hi_808;
  assign dataInMem_hi_hi_808 = _GEN_1082;
  wire [63:0]       dataInMem_hi_lo_426;
  assign dataInMem_hi_lo_426 = _GEN_1082;
  wire [95:0]       dataInMem_hi_1256 = {dataInMem_hi_hi_808, dataRegroupBySew_2_2_20};
  wire [63:0]       _GEN_1083 = {dataRegroupBySew_4_2_21, dataRegroupBySew_3_2_21};
  wire [63:0]       dataInMem_hi_hi_809;
  assign dataInMem_hi_hi_809 = _GEN_1083;
  wire [63:0]       dataInMem_hi_lo_427;
  assign dataInMem_hi_lo_427 = _GEN_1083;
  wire [95:0]       dataInMem_hi_1257 = {dataInMem_hi_hi_809, dataRegroupBySew_2_2_21};
  wire [63:0]       _GEN_1084 = {dataRegroupBySew_4_2_22, dataRegroupBySew_3_2_22};
  wire [63:0]       dataInMem_hi_hi_810;
  assign dataInMem_hi_hi_810 = _GEN_1084;
  wire [63:0]       dataInMem_hi_lo_428;
  assign dataInMem_hi_lo_428 = _GEN_1084;
  wire [95:0]       dataInMem_hi_1258 = {dataInMem_hi_hi_810, dataRegroupBySew_2_2_22};
  wire [63:0]       _GEN_1085 = {dataRegroupBySew_4_2_23, dataRegroupBySew_3_2_23};
  wire [63:0]       dataInMem_hi_hi_811;
  assign dataInMem_hi_hi_811 = _GEN_1085;
  wire [63:0]       dataInMem_hi_lo_429;
  assign dataInMem_hi_lo_429 = _GEN_1085;
  wire [95:0]       dataInMem_hi_1259 = {dataInMem_hi_hi_811, dataRegroupBySew_2_2_23};
  wire [63:0]       _GEN_1086 = {dataRegroupBySew_4_2_24, dataRegroupBySew_3_2_24};
  wire [63:0]       dataInMem_hi_hi_812;
  assign dataInMem_hi_hi_812 = _GEN_1086;
  wire [63:0]       dataInMem_hi_lo_430;
  assign dataInMem_hi_lo_430 = _GEN_1086;
  wire [95:0]       dataInMem_hi_1260 = {dataInMem_hi_hi_812, dataRegroupBySew_2_2_24};
  wire [63:0]       _GEN_1087 = {dataRegroupBySew_4_2_25, dataRegroupBySew_3_2_25};
  wire [63:0]       dataInMem_hi_hi_813;
  assign dataInMem_hi_hi_813 = _GEN_1087;
  wire [63:0]       dataInMem_hi_lo_431;
  assign dataInMem_hi_lo_431 = _GEN_1087;
  wire [95:0]       dataInMem_hi_1261 = {dataInMem_hi_hi_813, dataRegroupBySew_2_2_25};
  wire [63:0]       _GEN_1088 = {dataRegroupBySew_4_2_26, dataRegroupBySew_3_2_26};
  wire [63:0]       dataInMem_hi_hi_814;
  assign dataInMem_hi_hi_814 = _GEN_1088;
  wire [63:0]       dataInMem_hi_lo_432;
  assign dataInMem_hi_lo_432 = _GEN_1088;
  wire [95:0]       dataInMem_hi_1262 = {dataInMem_hi_hi_814, dataRegroupBySew_2_2_26};
  wire [63:0]       _GEN_1089 = {dataRegroupBySew_4_2_27, dataRegroupBySew_3_2_27};
  wire [63:0]       dataInMem_hi_hi_815;
  assign dataInMem_hi_hi_815 = _GEN_1089;
  wire [63:0]       dataInMem_hi_lo_433;
  assign dataInMem_hi_lo_433 = _GEN_1089;
  wire [95:0]       dataInMem_hi_1263 = {dataInMem_hi_hi_815, dataRegroupBySew_2_2_27};
  wire [63:0]       _GEN_1090 = {dataRegroupBySew_4_2_28, dataRegroupBySew_3_2_28};
  wire [63:0]       dataInMem_hi_hi_816;
  assign dataInMem_hi_hi_816 = _GEN_1090;
  wire [63:0]       dataInMem_hi_lo_434;
  assign dataInMem_hi_lo_434 = _GEN_1090;
  wire [95:0]       dataInMem_hi_1264 = {dataInMem_hi_hi_816, dataRegroupBySew_2_2_28};
  wire [63:0]       _GEN_1091 = {dataRegroupBySew_4_2_29, dataRegroupBySew_3_2_29};
  wire [63:0]       dataInMem_hi_hi_817;
  assign dataInMem_hi_hi_817 = _GEN_1091;
  wire [63:0]       dataInMem_hi_lo_435;
  assign dataInMem_hi_lo_435 = _GEN_1091;
  wire [95:0]       dataInMem_hi_1265 = {dataInMem_hi_hi_817, dataRegroupBySew_2_2_29};
  wire [63:0]       _GEN_1092 = {dataRegroupBySew_4_2_30, dataRegroupBySew_3_2_30};
  wire [63:0]       dataInMem_hi_hi_818;
  assign dataInMem_hi_hi_818 = _GEN_1092;
  wire [63:0]       dataInMem_hi_lo_436;
  assign dataInMem_hi_lo_436 = _GEN_1092;
  wire [95:0]       dataInMem_hi_1266 = {dataInMem_hi_hi_818, dataRegroupBySew_2_2_30};
  wire [63:0]       _GEN_1093 = {dataRegroupBySew_4_2_31, dataRegroupBySew_3_2_31};
  wire [63:0]       dataInMem_hi_hi_819;
  assign dataInMem_hi_hi_819 = _GEN_1093;
  wire [63:0]       dataInMem_hi_lo_437;
  assign dataInMem_hi_lo_437 = _GEN_1093;
  wire [95:0]       dataInMem_hi_1267 = {dataInMem_hi_hi_819, dataRegroupBySew_2_2_31};
  wire [319:0]      dataInMem_lo_lo_lo_lo_20 = {dataInMem_hi_1237, dataInMem_lo_1013, dataInMem_hi_1236, dataInMem_lo_1012};
  wire [319:0]      dataInMem_lo_lo_lo_hi_20 = {dataInMem_hi_1239, dataInMem_lo_1015, dataInMem_hi_1238, dataInMem_lo_1014};
  wire [639:0]      dataInMem_lo_lo_lo_20 = {dataInMem_lo_lo_lo_hi_20, dataInMem_lo_lo_lo_lo_20};
  wire [319:0]      dataInMem_lo_lo_hi_lo_20 = {dataInMem_hi_1241, dataInMem_lo_1017, dataInMem_hi_1240, dataInMem_lo_1016};
  wire [319:0]      dataInMem_lo_lo_hi_hi_20 = {dataInMem_hi_1243, dataInMem_lo_1019, dataInMem_hi_1242, dataInMem_lo_1018};
  wire [639:0]      dataInMem_lo_lo_hi_20 = {dataInMem_lo_lo_hi_hi_20, dataInMem_lo_lo_hi_lo_20};
  wire [1279:0]     dataInMem_lo_lo_212 = {dataInMem_lo_lo_hi_20, dataInMem_lo_lo_lo_20};
  wire [319:0]      dataInMem_lo_hi_lo_lo_20 = {dataInMem_hi_1245, dataInMem_lo_1021, dataInMem_hi_1244, dataInMem_lo_1020};
  wire [319:0]      dataInMem_lo_hi_lo_hi_20 = {dataInMem_hi_1247, dataInMem_lo_1023, dataInMem_hi_1246, dataInMem_lo_1022};
  wire [639:0]      dataInMem_lo_hi_lo_20 = {dataInMem_lo_hi_lo_hi_20, dataInMem_lo_hi_lo_lo_20};
  wire [319:0]      dataInMem_lo_hi_hi_lo_20 = {dataInMem_hi_1249, dataInMem_lo_1025, dataInMem_hi_1248, dataInMem_lo_1024};
  wire [319:0]      dataInMem_lo_hi_hi_hi_20 = {dataInMem_hi_1251, dataInMem_lo_1027, dataInMem_hi_1250, dataInMem_lo_1026};
  wire [639:0]      dataInMem_lo_hi_hi_20 = {dataInMem_lo_hi_hi_hi_20, dataInMem_lo_hi_hi_lo_20};
  wire [1279:0]     dataInMem_lo_hi_596 = {dataInMem_lo_hi_hi_20, dataInMem_lo_hi_lo_20};
  wire [2559:0]     dataInMem_lo_1044 = {dataInMem_lo_hi_596, dataInMem_lo_lo_212};
  wire [319:0]      dataInMem_hi_lo_lo_lo_20 = {dataInMem_hi_1253, dataInMem_lo_1029, dataInMem_hi_1252, dataInMem_lo_1028};
  wire [319:0]      dataInMem_hi_lo_lo_hi_20 = {dataInMem_hi_1255, dataInMem_lo_1031, dataInMem_hi_1254, dataInMem_lo_1030};
  wire [639:0]      dataInMem_hi_lo_lo_20 = {dataInMem_hi_lo_lo_hi_20, dataInMem_hi_lo_lo_lo_20};
  wire [319:0]      dataInMem_hi_lo_hi_lo_20 = {dataInMem_hi_1257, dataInMem_lo_1033, dataInMem_hi_1256, dataInMem_lo_1032};
  wire [319:0]      dataInMem_hi_lo_hi_hi_20 = {dataInMem_hi_1259, dataInMem_lo_1035, dataInMem_hi_1258, dataInMem_lo_1034};
  wire [639:0]      dataInMem_hi_lo_hi_20 = {dataInMem_hi_lo_hi_hi_20, dataInMem_hi_lo_hi_lo_20};
  wire [1279:0]     dataInMem_hi_lo_404 = {dataInMem_hi_lo_hi_20, dataInMem_hi_lo_lo_20};
  wire [319:0]      dataInMem_hi_hi_lo_lo_20 = {dataInMem_hi_1261, dataInMem_lo_1037, dataInMem_hi_1260, dataInMem_lo_1036};
  wire [319:0]      dataInMem_hi_hi_lo_hi_20 = {dataInMem_hi_1263, dataInMem_lo_1039, dataInMem_hi_1262, dataInMem_lo_1038};
  wire [639:0]      dataInMem_hi_hi_lo_20 = {dataInMem_hi_hi_lo_hi_20, dataInMem_hi_hi_lo_lo_20};
  wire [319:0]      dataInMem_hi_hi_hi_lo_20 = {dataInMem_hi_1265, dataInMem_lo_1041, dataInMem_hi_1264, dataInMem_lo_1040};
  wire [319:0]      dataInMem_hi_hi_hi_hi_20 = {dataInMem_hi_1267, dataInMem_lo_1043, dataInMem_hi_1266, dataInMem_lo_1042};
  wire [639:0]      dataInMem_hi_hi_hi_20 = {dataInMem_hi_hi_hi_hi_20, dataInMem_hi_hi_hi_lo_20};
  wire [1279:0]     dataInMem_hi_hi_820 = {dataInMem_hi_hi_hi_20, dataInMem_hi_hi_lo_20};
  wire [2559:0]     dataInMem_hi_1268 = {dataInMem_hi_hi_820, dataInMem_hi_lo_404};
  wire [5119:0]     dataInMem_20 = {dataInMem_hi_1268, dataInMem_lo_1044};
  wire [1023:0]     regroupCacheLine_20_0 = dataInMem_20[1023:0];
  wire [1023:0]     regroupCacheLine_20_1 = dataInMem_20[2047:1024];
  wire [1023:0]     regroupCacheLine_20_2 = dataInMem_20[3071:2048];
  wire [1023:0]     regroupCacheLine_20_3 = dataInMem_20[4095:3072];
  wire [1023:0]     regroupCacheLine_20_4 = dataInMem_20[5119:4096];
  wire [1023:0]     res_160 = regroupCacheLine_20_0;
  wire [1023:0]     res_161 = regroupCacheLine_20_1;
  wire [1023:0]     res_162 = regroupCacheLine_20_2;
  wire [1023:0]     res_163 = regroupCacheLine_20_3;
  wire [1023:0]     res_164 = regroupCacheLine_20_4;
  wire [2047:0]     lo_lo_20 = {res_161, res_160};
  wire [2047:0]     lo_hi_20 = {res_163, res_162};
  wire [4095:0]     lo_20 = {lo_hi_20, lo_lo_20};
  wire [2047:0]     hi_lo_20 = {1024'h0, res_164};
  wire [4095:0]     hi_20 = {2048'h0, hi_lo_20};
  wire [8191:0]     regroupLoadData_2_4 = {hi_20, lo_20};
  wire [95:0]       dataInMem_lo_1045 = {dataInMem_lo_hi_597, dataRegroupBySew_0_2_0};
  wire [63:0]       _GEN_1094 = {dataRegroupBySew_5_2_0, dataRegroupBySew_4_2_0};
  wire [63:0]       dataInMem_hi_hi_821;
  assign dataInMem_hi_hi_821 = _GEN_1094;
  wire [63:0]       dataInMem_hi_lo_439;
  assign dataInMem_hi_lo_439 = _GEN_1094;
  wire [95:0]       dataInMem_hi_1269 = {dataInMem_hi_hi_821, dataRegroupBySew_3_2_0};
  wire [95:0]       dataInMem_lo_1046 = {dataInMem_lo_hi_598, dataRegroupBySew_0_2_1};
  wire [63:0]       _GEN_1095 = {dataRegroupBySew_5_2_1, dataRegroupBySew_4_2_1};
  wire [63:0]       dataInMem_hi_hi_822;
  assign dataInMem_hi_hi_822 = _GEN_1095;
  wire [63:0]       dataInMem_hi_lo_440;
  assign dataInMem_hi_lo_440 = _GEN_1095;
  wire [95:0]       dataInMem_hi_1270 = {dataInMem_hi_hi_822, dataRegroupBySew_3_2_1};
  wire [95:0]       dataInMem_lo_1047 = {dataInMem_lo_hi_599, dataRegroupBySew_0_2_2};
  wire [63:0]       _GEN_1096 = {dataRegroupBySew_5_2_2, dataRegroupBySew_4_2_2};
  wire [63:0]       dataInMem_hi_hi_823;
  assign dataInMem_hi_hi_823 = _GEN_1096;
  wire [63:0]       dataInMem_hi_lo_441;
  assign dataInMem_hi_lo_441 = _GEN_1096;
  wire [95:0]       dataInMem_hi_1271 = {dataInMem_hi_hi_823, dataRegroupBySew_3_2_2};
  wire [95:0]       dataInMem_lo_1048 = {dataInMem_lo_hi_600, dataRegroupBySew_0_2_3};
  wire [63:0]       _GEN_1097 = {dataRegroupBySew_5_2_3, dataRegroupBySew_4_2_3};
  wire [63:0]       dataInMem_hi_hi_824;
  assign dataInMem_hi_hi_824 = _GEN_1097;
  wire [63:0]       dataInMem_hi_lo_442;
  assign dataInMem_hi_lo_442 = _GEN_1097;
  wire [95:0]       dataInMem_hi_1272 = {dataInMem_hi_hi_824, dataRegroupBySew_3_2_3};
  wire [95:0]       dataInMem_lo_1049 = {dataInMem_lo_hi_601, dataRegroupBySew_0_2_4};
  wire [63:0]       _GEN_1098 = {dataRegroupBySew_5_2_4, dataRegroupBySew_4_2_4};
  wire [63:0]       dataInMem_hi_hi_825;
  assign dataInMem_hi_hi_825 = _GEN_1098;
  wire [63:0]       dataInMem_hi_lo_443;
  assign dataInMem_hi_lo_443 = _GEN_1098;
  wire [95:0]       dataInMem_hi_1273 = {dataInMem_hi_hi_825, dataRegroupBySew_3_2_4};
  wire [95:0]       dataInMem_lo_1050 = {dataInMem_lo_hi_602, dataRegroupBySew_0_2_5};
  wire [63:0]       _GEN_1099 = {dataRegroupBySew_5_2_5, dataRegroupBySew_4_2_5};
  wire [63:0]       dataInMem_hi_hi_826;
  assign dataInMem_hi_hi_826 = _GEN_1099;
  wire [63:0]       dataInMem_hi_lo_444;
  assign dataInMem_hi_lo_444 = _GEN_1099;
  wire [95:0]       dataInMem_hi_1274 = {dataInMem_hi_hi_826, dataRegroupBySew_3_2_5};
  wire [95:0]       dataInMem_lo_1051 = {dataInMem_lo_hi_603, dataRegroupBySew_0_2_6};
  wire [63:0]       _GEN_1100 = {dataRegroupBySew_5_2_6, dataRegroupBySew_4_2_6};
  wire [63:0]       dataInMem_hi_hi_827;
  assign dataInMem_hi_hi_827 = _GEN_1100;
  wire [63:0]       dataInMem_hi_lo_445;
  assign dataInMem_hi_lo_445 = _GEN_1100;
  wire [95:0]       dataInMem_hi_1275 = {dataInMem_hi_hi_827, dataRegroupBySew_3_2_6};
  wire [95:0]       dataInMem_lo_1052 = {dataInMem_lo_hi_604, dataRegroupBySew_0_2_7};
  wire [63:0]       _GEN_1101 = {dataRegroupBySew_5_2_7, dataRegroupBySew_4_2_7};
  wire [63:0]       dataInMem_hi_hi_828;
  assign dataInMem_hi_hi_828 = _GEN_1101;
  wire [63:0]       dataInMem_hi_lo_446;
  assign dataInMem_hi_lo_446 = _GEN_1101;
  wire [95:0]       dataInMem_hi_1276 = {dataInMem_hi_hi_828, dataRegroupBySew_3_2_7};
  wire [95:0]       dataInMem_lo_1053 = {dataInMem_lo_hi_605, dataRegroupBySew_0_2_8};
  wire [63:0]       _GEN_1102 = {dataRegroupBySew_5_2_8, dataRegroupBySew_4_2_8};
  wire [63:0]       dataInMem_hi_hi_829;
  assign dataInMem_hi_hi_829 = _GEN_1102;
  wire [63:0]       dataInMem_hi_lo_447;
  assign dataInMem_hi_lo_447 = _GEN_1102;
  wire [95:0]       dataInMem_hi_1277 = {dataInMem_hi_hi_829, dataRegroupBySew_3_2_8};
  wire [95:0]       dataInMem_lo_1054 = {dataInMem_lo_hi_606, dataRegroupBySew_0_2_9};
  wire [63:0]       _GEN_1103 = {dataRegroupBySew_5_2_9, dataRegroupBySew_4_2_9};
  wire [63:0]       dataInMem_hi_hi_830;
  assign dataInMem_hi_hi_830 = _GEN_1103;
  wire [63:0]       dataInMem_hi_lo_448;
  assign dataInMem_hi_lo_448 = _GEN_1103;
  wire [95:0]       dataInMem_hi_1278 = {dataInMem_hi_hi_830, dataRegroupBySew_3_2_9};
  wire [95:0]       dataInMem_lo_1055 = {dataInMem_lo_hi_607, dataRegroupBySew_0_2_10};
  wire [63:0]       _GEN_1104 = {dataRegroupBySew_5_2_10, dataRegroupBySew_4_2_10};
  wire [63:0]       dataInMem_hi_hi_831;
  assign dataInMem_hi_hi_831 = _GEN_1104;
  wire [63:0]       dataInMem_hi_lo_449;
  assign dataInMem_hi_lo_449 = _GEN_1104;
  wire [95:0]       dataInMem_hi_1279 = {dataInMem_hi_hi_831, dataRegroupBySew_3_2_10};
  wire [95:0]       dataInMem_lo_1056 = {dataInMem_lo_hi_608, dataRegroupBySew_0_2_11};
  wire [63:0]       _GEN_1105 = {dataRegroupBySew_5_2_11, dataRegroupBySew_4_2_11};
  wire [63:0]       dataInMem_hi_hi_832;
  assign dataInMem_hi_hi_832 = _GEN_1105;
  wire [63:0]       dataInMem_hi_lo_450;
  assign dataInMem_hi_lo_450 = _GEN_1105;
  wire [95:0]       dataInMem_hi_1280 = {dataInMem_hi_hi_832, dataRegroupBySew_3_2_11};
  wire [95:0]       dataInMem_lo_1057 = {dataInMem_lo_hi_609, dataRegroupBySew_0_2_12};
  wire [63:0]       _GEN_1106 = {dataRegroupBySew_5_2_12, dataRegroupBySew_4_2_12};
  wire [63:0]       dataInMem_hi_hi_833;
  assign dataInMem_hi_hi_833 = _GEN_1106;
  wire [63:0]       dataInMem_hi_lo_451;
  assign dataInMem_hi_lo_451 = _GEN_1106;
  wire [95:0]       dataInMem_hi_1281 = {dataInMem_hi_hi_833, dataRegroupBySew_3_2_12};
  wire [95:0]       dataInMem_lo_1058 = {dataInMem_lo_hi_610, dataRegroupBySew_0_2_13};
  wire [63:0]       _GEN_1107 = {dataRegroupBySew_5_2_13, dataRegroupBySew_4_2_13};
  wire [63:0]       dataInMem_hi_hi_834;
  assign dataInMem_hi_hi_834 = _GEN_1107;
  wire [63:0]       dataInMem_hi_lo_452;
  assign dataInMem_hi_lo_452 = _GEN_1107;
  wire [95:0]       dataInMem_hi_1282 = {dataInMem_hi_hi_834, dataRegroupBySew_3_2_13};
  wire [95:0]       dataInMem_lo_1059 = {dataInMem_lo_hi_611, dataRegroupBySew_0_2_14};
  wire [63:0]       _GEN_1108 = {dataRegroupBySew_5_2_14, dataRegroupBySew_4_2_14};
  wire [63:0]       dataInMem_hi_hi_835;
  assign dataInMem_hi_hi_835 = _GEN_1108;
  wire [63:0]       dataInMem_hi_lo_453;
  assign dataInMem_hi_lo_453 = _GEN_1108;
  wire [95:0]       dataInMem_hi_1283 = {dataInMem_hi_hi_835, dataRegroupBySew_3_2_14};
  wire [95:0]       dataInMem_lo_1060 = {dataInMem_lo_hi_612, dataRegroupBySew_0_2_15};
  wire [63:0]       _GEN_1109 = {dataRegroupBySew_5_2_15, dataRegroupBySew_4_2_15};
  wire [63:0]       dataInMem_hi_hi_836;
  assign dataInMem_hi_hi_836 = _GEN_1109;
  wire [63:0]       dataInMem_hi_lo_454;
  assign dataInMem_hi_lo_454 = _GEN_1109;
  wire [95:0]       dataInMem_hi_1284 = {dataInMem_hi_hi_836, dataRegroupBySew_3_2_15};
  wire [95:0]       dataInMem_lo_1061 = {dataInMem_lo_hi_613, dataRegroupBySew_0_2_16};
  wire [63:0]       _GEN_1110 = {dataRegroupBySew_5_2_16, dataRegroupBySew_4_2_16};
  wire [63:0]       dataInMem_hi_hi_837;
  assign dataInMem_hi_hi_837 = _GEN_1110;
  wire [63:0]       dataInMem_hi_lo_455;
  assign dataInMem_hi_lo_455 = _GEN_1110;
  wire [95:0]       dataInMem_hi_1285 = {dataInMem_hi_hi_837, dataRegroupBySew_3_2_16};
  wire [95:0]       dataInMem_lo_1062 = {dataInMem_lo_hi_614, dataRegroupBySew_0_2_17};
  wire [63:0]       _GEN_1111 = {dataRegroupBySew_5_2_17, dataRegroupBySew_4_2_17};
  wire [63:0]       dataInMem_hi_hi_838;
  assign dataInMem_hi_hi_838 = _GEN_1111;
  wire [63:0]       dataInMem_hi_lo_456;
  assign dataInMem_hi_lo_456 = _GEN_1111;
  wire [95:0]       dataInMem_hi_1286 = {dataInMem_hi_hi_838, dataRegroupBySew_3_2_17};
  wire [95:0]       dataInMem_lo_1063 = {dataInMem_lo_hi_615, dataRegroupBySew_0_2_18};
  wire [63:0]       _GEN_1112 = {dataRegroupBySew_5_2_18, dataRegroupBySew_4_2_18};
  wire [63:0]       dataInMem_hi_hi_839;
  assign dataInMem_hi_hi_839 = _GEN_1112;
  wire [63:0]       dataInMem_hi_lo_457;
  assign dataInMem_hi_lo_457 = _GEN_1112;
  wire [95:0]       dataInMem_hi_1287 = {dataInMem_hi_hi_839, dataRegroupBySew_3_2_18};
  wire [95:0]       dataInMem_lo_1064 = {dataInMem_lo_hi_616, dataRegroupBySew_0_2_19};
  wire [63:0]       _GEN_1113 = {dataRegroupBySew_5_2_19, dataRegroupBySew_4_2_19};
  wire [63:0]       dataInMem_hi_hi_840;
  assign dataInMem_hi_hi_840 = _GEN_1113;
  wire [63:0]       dataInMem_hi_lo_458;
  assign dataInMem_hi_lo_458 = _GEN_1113;
  wire [95:0]       dataInMem_hi_1288 = {dataInMem_hi_hi_840, dataRegroupBySew_3_2_19};
  wire [95:0]       dataInMem_lo_1065 = {dataInMem_lo_hi_617, dataRegroupBySew_0_2_20};
  wire [63:0]       _GEN_1114 = {dataRegroupBySew_5_2_20, dataRegroupBySew_4_2_20};
  wire [63:0]       dataInMem_hi_hi_841;
  assign dataInMem_hi_hi_841 = _GEN_1114;
  wire [63:0]       dataInMem_hi_lo_459;
  assign dataInMem_hi_lo_459 = _GEN_1114;
  wire [95:0]       dataInMem_hi_1289 = {dataInMem_hi_hi_841, dataRegroupBySew_3_2_20};
  wire [95:0]       dataInMem_lo_1066 = {dataInMem_lo_hi_618, dataRegroupBySew_0_2_21};
  wire [63:0]       _GEN_1115 = {dataRegroupBySew_5_2_21, dataRegroupBySew_4_2_21};
  wire [63:0]       dataInMem_hi_hi_842;
  assign dataInMem_hi_hi_842 = _GEN_1115;
  wire [63:0]       dataInMem_hi_lo_460;
  assign dataInMem_hi_lo_460 = _GEN_1115;
  wire [95:0]       dataInMem_hi_1290 = {dataInMem_hi_hi_842, dataRegroupBySew_3_2_21};
  wire [95:0]       dataInMem_lo_1067 = {dataInMem_lo_hi_619, dataRegroupBySew_0_2_22};
  wire [63:0]       _GEN_1116 = {dataRegroupBySew_5_2_22, dataRegroupBySew_4_2_22};
  wire [63:0]       dataInMem_hi_hi_843;
  assign dataInMem_hi_hi_843 = _GEN_1116;
  wire [63:0]       dataInMem_hi_lo_461;
  assign dataInMem_hi_lo_461 = _GEN_1116;
  wire [95:0]       dataInMem_hi_1291 = {dataInMem_hi_hi_843, dataRegroupBySew_3_2_22};
  wire [95:0]       dataInMem_lo_1068 = {dataInMem_lo_hi_620, dataRegroupBySew_0_2_23};
  wire [63:0]       _GEN_1117 = {dataRegroupBySew_5_2_23, dataRegroupBySew_4_2_23};
  wire [63:0]       dataInMem_hi_hi_844;
  assign dataInMem_hi_hi_844 = _GEN_1117;
  wire [63:0]       dataInMem_hi_lo_462;
  assign dataInMem_hi_lo_462 = _GEN_1117;
  wire [95:0]       dataInMem_hi_1292 = {dataInMem_hi_hi_844, dataRegroupBySew_3_2_23};
  wire [95:0]       dataInMem_lo_1069 = {dataInMem_lo_hi_621, dataRegroupBySew_0_2_24};
  wire [63:0]       _GEN_1118 = {dataRegroupBySew_5_2_24, dataRegroupBySew_4_2_24};
  wire [63:0]       dataInMem_hi_hi_845;
  assign dataInMem_hi_hi_845 = _GEN_1118;
  wire [63:0]       dataInMem_hi_lo_463;
  assign dataInMem_hi_lo_463 = _GEN_1118;
  wire [95:0]       dataInMem_hi_1293 = {dataInMem_hi_hi_845, dataRegroupBySew_3_2_24};
  wire [95:0]       dataInMem_lo_1070 = {dataInMem_lo_hi_622, dataRegroupBySew_0_2_25};
  wire [63:0]       _GEN_1119 = {dataRegroupBySew_5_2_25, dataRegroupBySew_4_2_25};
  wire [63:0]       dataInMem_hi_hi_846;
  assign dataInMem_hi_hi_846 = _GEN_1119;
  wire [63:0]       dataInMem_hi_lo_464;
  assign dataInMem_hi_lo_464 = _GEN_1119;
  wire [95:0]       dataInMem_hi_1294 = {dataInMem_hi_hi_846, dataRegroupBySew_3_2_25};
  wire [95:0]       dataInMem_lo_1071 = {dataInMem_lo_hi_623, dataRegroupBySew_0_2_26};
  wire [63:0]       _GEN_1120 = {dataRegroupBySew_5_2_26, dataRegroupBySew_4_2_26};
  wire [63:0]       dataInMem_hi_hi_847;
  assign dataInMem_hi_hi_847 = _GEN_1120;
  wire [63:0]       dataInMem_hi_lo_465;
  assign dataInMem_hi_lo_465 = _GEN_1120;
  wire [95:0]       dataInMem_hi_1295 = {dataInMem_hi_hi_847, dataRegroupBySew_3_2_26};
  wire [95:0]       dataInMem_lo_1072 = {dataInMem_lo_hi_624, dataRegroupBySew_0_2_27};
  wire [63:0]       _GEN_1121 = {dataRegroupBySew_5_2_27, dataRegroupBySew_4_2_27};
  wire [63:0]       dataInMem_hi_hi_848;
  assign dataInMem_hi_hi_848 = _GEN_1121;
  wire [63:0]       dataInMem_hi_lo_466;
  assign dataInMem_hi_lo_466 = _GEN_1121;
  wire [95:0]       dataInMem_hi_1296 = {dataInMem_hi_hi_848, dataRegroupBySew_3_2_27};
  wire [95:0]       dataInMem_lo_1073 = {dataInMem_lo_hi_625, dataRegroupBySew_0_2_28};
  wire [63:0]       _GEN_1122 = {dataRegroupBySew_5_2_28, dataRegroupBySew_4_2_28};
  wire [63:0]       dataInMem_hi_hi_849;
  assign dataInMem_hi_hi_849 = _GEN_1122;
  wire [63:0]       dataInMem_hi_lo_467;
  assign dataInMem_hi_lo_467 = _GEN_1122;
  wire [95:0]       dataInMem_hi_1297 = {dataInMem_hi_hi_849, dataRegroupBySew_3_2_28};
  wire [95:0]       dataInMem_lo_1074 = {dataInMem_lo_hi_626, dataRegroupBySew_0_2_29};
  wire [63:0]       _GEN_1123 = {dataRegroupBySew_5_2_29, dataRegroupBySew_4_2_29};
  wire [63:0]       dataInMem_hi_hi_850;
  assign dataInMem_hi_hi_850 = _GEN_1123;
  wire [63:0]       dataInMem_hi_lo_468;
  assign dataInMem_hi_lo_468 = _GEN_1123;
  wire [95:0]       dataInMem_hi_1298 = {dataInMem_hi_hi_850, dataRegroupBySew_3_2_29};
  wire [95:0]       dataInMem_lo_1075 = {dataInMem_lo_hi_627, dataRegroupBySew_0_2_30};
  wire [63:0]       _GEN_1124 = {dataRegroupBySew_5_2_30, dataRegroupBySew_4_2_30};
  wire [63:0]       dataInMem_hi_hi_851;
  assign dataInMem_hi_hi_851 = _GEN_1124;
  wire [63:0]       dataInMem_hi_lo_469;
  assign dataInMem_hi_lo_469 = _GEN_1124;
  wire [95:0]       dataInMem_hi_1299 = {dataInMem_hi_hi_851, dataRegroupBySew_3_2_30};
  wire [95:0]       dataInMem_lo_1076 = {dataInMem_lo_hi_628, dataRegroupBySew_0_2_31};
  wire [63:0]       _GEN_1125 = {dataRegroupBySew_5_2_31, dataRegroupBySew_4_2_31};
  wire [63:0]       dataInMem_hi_hi_852;
  assign dataInMem_hi_hi_852 = _GEN_1125;
  wire [63:0]       dataInMem_hi_lo_470;
  assign dataInMem_hi_lo_470 = _GEN_1125;
  wire [95:0]       dataInMem_hi_1300 = {dataInMem_hi_hi_852, dataRegroupBySew_3_2_31};
  wire [383:0]      dataInMem_lo_lo_lo_lo_21 = {dataInMem_hi_1270, dataInMem_lo_1046, dataInMem_hi_1269, dataInMem_lo_1045};
  wire [383:0]      dataInMem_lo_lo_lo_hi_21 = {dataInMem_hi_1272, dataInMem_lo_1048, dataInMem_hi_1271, dataInMem_lo_1047};
  wire [767:0]      dataInMem_lo_lo_lo_21 = {dataInMem_lo_lo_lo_hi_21, dataInMem_lo_lo_lo_lo_21};
  wire [383:0]      dataInMem_lo_lo_hi_lo_21 = {dataInMem_hi_1274, dataInMem_lo_1050, dataInMem_hi_1273, dataInMem_lo_1049};
  wire [383:0]      dataInMem_lo_lo_hi_hi_21 = {dataInMem_hi_1276, dataInMem_lo_1052, dataInMem_hi_1275, dataInMem_lo_1051};
  wire [767:0]      dataInMem_lo_lo_hi_21 = {dataInMem_lo_lo_hi_hi_21, dataInMem_lo_lo_hi_lo_21};
  wire [1535:0]     dataInMem_lo_lo_213 = {dataInMem_lo_lo_hi_21, dataInMem_lo_lo_lo_21};
  wire [383:0]      dataInMem_lo_hi_lo_lo_21 = {dataInMem_hi_1278, dataInMem_lo_1054, dataInMem_hi_1277, dataInMem_lo_1053};
  wire [383:0]      dataInMem_lo_hi_lo_hi_21 = {dataInMem_hi_1280, dataInMem_lo_1056, dataInMem_hi_1279, dataInMem_lo_1055};
  wire [767:0]      dataInMem_lo_hi_lo_21 = {dataInMem_lo_hi_lo_hi_21, dataInMem_lo_hi_lo_lo_21};
  wire [383:0]      dataInMem_lo_hi_hi_lo_21 = {dataInMem_hi_1282, dataInMem_lo_1058, dataInMem_hi_1281, dataInMem_lo_1057};
  wire [383:0]      dataInMem_lo_hi_hi_hi_21 = {dataInMem_hi_1284, dataInMem_lo_1060, dataInMem_hi_1283, dataInMem_lo_1059};
  wire [767:0]      dataInMem_lo_hi_hi_21 = {dataInMem_lo_hi_hi_hi_21, dataInMem_lo_hi_hi_lo_21};
  wire [1535:0]     dataInMem_lo_hi_629 = {dataInMem_lo_hi_hi_21, dataInMem_lo_hi_lo_21};
  wire [3071:0]     dataInMem_lo_1077 = {dataInMem_lo_hi_629, dataInMem_lo_lo_213};
  wire [383:0]      dataInMem_hi_lo_lo_lo_21 = {dataInMem_hi_1286, dataInMem_lo_1062, dataInMem_hi_1285, dataInMem_lo_1061};
  wire [383:0]      dataInMem_hi_lo_lo_hi_21 = {dataInMem_hi_1288, dataInMem_lo_1064, dataInMem_hi_1287, dataInMem_lo_1063};
  wire [767:0]      dataInMem_hi_lo_lo_21 = {dataInMem_hi_lo_lo_hi_21, dataInMem_hi_lo_lo_lo_21};
  wire [383:0]      dataInMem_hi_lo_hi_lo_21 = {dataInMem_hi_1290, dataInMem_lo_1066, dataInMem_hi_1289, dataInMem_lo_1065};
  wire [383:0]      dataInMem_hi_lo_hi_hi_21 = {dataInMem_hi_1292, dataInMem_lo_1068, dataInMem_hi_1291, dataInMem_lo_1067};
  wire [767:0]      dataInMem_hi_lo_hi_21 = {dataInMem_hi_lo_hi_hi_21, dataInMem_hi_lo_hi_lo_21};
  wire [1535:0]     dataInMem_hi_lo_405 = {dataInMem_hi_lo_hi_21, dataInMem_hi_lo_lo_21};
  wire [383:0]      dataInMem_hi_hi_lo_lo_21 = {dataInMem_hi_1294, dataInMem_lo_1070, dataInMem_hi_1293, dataInMem_lo_1069};
  wire [383:0]      dataInMem_hi_hi_lo_hi_21 = {dataInMem_hi_1296, dataInMem_lo_1072, dataInMem_hi_1295, dataInMem_lo_1071};
  wire [767:0]      dataInMem_hi_hi_lo_21 = {dataInMem_hi_hi_lo_hi_21, dataInMem_hi_hi_lo_lo_21};
  wire [383:0]      dataInMem_hi_hi_hi_lo_21 = {dataInMem_hi_1298, dataInMem_lo_1074, dataInMem_hi_1297, dataInMem_lo_1073};
  wire [383:0]      dataInMem_hi_hi_hi_hi_21 = {dataInMem_hi_1300, dataInMem_lo_1076, dataInMem_hi_1299, dataInMem_lo_1075};
  wire [767:0]      dataInMem_hi_hi_hi_21 = {dataInMem_hi_hi_hi_hi_21, dataInMem_hi_hi_hi_lo_21};
  wire [1535:0]     dataInMem_hi_hi_853 = {dataInMem_hi_hi_hi_21, dataInMem_hi_hi_lo_21};
  wire [3071:0]     dataInMem_hi_1301 = {dataInMem_hi_hi_853, dataInMem_hi_lo_405};
  wire [6143:0]     dataInMem_21 = {dataInMem_hi_1301, dataInMem_lo_1077};
  wire [1023:0]     regroupCacheLine_21_0 = dataInMem_21[1023:0];
  wire [1023:0]     regroupCacheLine_21_1 = dataInMem_21[2047:1024];
  wire [1023:0]     regroupCacheLine_21_2 = dataInMem_21[3071:2048];
  wire [1023:0]     regroupCacheLine_21_3 = dataInMem_21[4095:3072];
  wire [1023:0]     regroupCacheLine_21_4 = dataInMem_21[5119:4096];
  wire [1023:0]     regroupCacheLine_21_5 = dataInMem_21[6143:5120];
  wire [1023:0]     res_168 = regroupCacheLine_21_0;
  wire [1023:0]     res_169 = regroupCacheLine_21_1;
  wire [1023:0]     res_170 = regroupCacheLine_21_2;
  wire [1023:0]     res_171 = regroupCacheLine_21_3;
  wire [1023:0]     res_172 = regroupCacheLine_21_4;
  wire [1023:0]     res_173 = regroupCacheLine_21_5;
  wire [2047:0]     lo_lo_21 = {res_169, res_168};
  wire [2047:0]     lo_hi_21 = {res_171, res_170};
  wire [4095:0]     lo_21 = {lo_hi_21, lo_lo_21};
  wire [2047:0]     hi_lo_21 = {res_173, res_172};
  wire [4095:0]     hi_21 = {2048'h0, hi_lo_21};
  wire [8191:0]     regroupLoadData_2_5 = {hi_21, lo_21};
  wire [95:0]       dataInMem_lo_1078 = {dataInMem_lo_hi_630, dataRegroupBySew_0_2_0};
  wire [63:0]       dataInMem_hi_hi_854 = {dataRegroupBySew_6_2_0, dataRegroupBySew_5_2_0};
  wire [127:0]      dataInMem_hi_1302 = {dataInMem_hi_hi_854, dataInMem_hi_lo_406};
  wire [95:0]       dataInMem_lo_1079 = {dataInMem_lo_hi_631, dataRegroupBySew_0_2_1};
  wire [63:0]       dataInMem_hi_hi_855 = {dataRegroupBySew_6_2_1, dataRegroupBySew_5_2_1};
  wire [127:0]      dataInMem_hi_1303 = {dataInMem_hi_hi_855, dataInMem_hi_lo_407};
  wire [95:0]       dataInMem_lo_1080 = {dataInMem_lo_hi_632, dataRegroupBySew_0_2_2};
  wire [63:0]       dataInMem_hi_hi_856 = {dataRegroupBySew_6_2_2, dataRegroupBySew_5_2_2};
  wire [127:0]      dataInMem_hi_1304 = {dataInMem_hi_hi_856, dataInMem_hi_lo_408};
  wire [95:0]       dataInMem_lo_1081 = {dataInMem_lo_hi_633, dataRegroupBySew_0_2_3};
  wire [63:0]       dataInMem_hi_hi_857 = {dataRegroupBySew_6_2_3, dataRegroupBySew_5_2_3};
  wire [127:0]      dataInMem_hi_1305 = {dataInMem_hi_hi_857, dataInMem_hi_lo_409};
  wire [95:0]       dataInMem_lo_1082 = {dataInMem_lo_hi_634, dataRegroupBySew_0_2_4};
  wire [63:0]       dataInMem_hi_hi_858 = {dataRegroupBySew_6_2_4, dataRegroupBySew_5_2_4};
  wire [127:0]      dataInMem_hi_1306 = {dataInMem_hi_hi_858, dataInMem_hi_lo_410};
  wire [95:0]       dataInMem_lo_1083 = {dataInMem_lo_hi_635, dataRegroupBySew_0_2_5};
  wire [63:0]       dataInMem_hi_hi_859 = {dataRegroupBySew_6_2_5, dataRegroupBySew_5_2_5};
  wire [127:0]      dataInMem_hi_1307 = {dataInMem_hi_hi_859, dataInMem_hi_lo_411};
  wire [95:0]       dataInMem_lo_1084 = {dataInMem_lo_hi_636, dataRegroupBySew_0_2_6};
  wire [63:0]       dataInMem_hi_hi_860 = {dataRegroupBySew_6_2_6, dataRegroupBySew_5_2_6};
  wire [127:0]      dataInMem_hi_1308 = {dataInMem_hi_hi_860, dataInMem_hi_lo_412};
  wire [95:0]       dataInMem_lo_1085 = {dataInMem_lo_hi_637, dataRegroupBySew_0_2_7};
  wire [63:0]       dataInMem_hi_hi_861 = {dataRegroupBySew_6_2_7, dataRegroupBySew_5_2_7};
  wire [127:0]      dataInMem_hi_1309 = {dataInMem_hi_hi_861, dataInMem_hi_lo_413};
  wire [95:0]       dataInMem_lo_1086 = {dataInMem_lo_hi_638, dataRegroupBySew_0_2_8};
  wire [63:0]       dataInMem_hi_hi_862 = {dataRegroupBySew_6_2_8, dataRegroupBySew_5_2_8};
  wire [127:0]      dataInMem_hi_1310 = {dataInMem_hi_hi_862, dataInMem_hi_lo_414};
  wire [95:0]       dataInMem_lo_1087 = {dataInMem_lo_hi_639, dataRegroupBySew_0_2_9};
  wire [63:0]       dataInMem_hi_hi_863 = {dataRegroupBySew_6_2_9, dataRegroupBySew_5_2_9};
  wire [127:0]      dataInMem_hi_1311 = {dataInMem_hi_hi_863, dataInMem_hi_lo_415};
  wire [95:0]       dataInMem_lo_1088 = {dataInMem_lo_hi_640, dataRegroupBySew_0_2_10};
  wire [63:0]       dataInMem_hi_hi_864 = {dataRegroupBySew_6_2_10, dataRegroupBySew_5_2_10};
  wire [127:0]      dataInMem_hi_1312 = {dataInMem_hi_hi_864, dataInMem_hi_lo_416};
  wire [95:0]       dataInMem_lo_1089 = {dataInMem_lo_hi_641, dataRegroupBySew_0_2_11};
  wire [63:0]       dataInMem_hi_hi_865 = {dataRegroupBySew_6_2_11, dataRegroupBySew_5_2_11};
  wire [127:0]      dataInMem_hi_1313 = {dataInMem_hi_hi_865, dataInMem_hi_lo_417};
  wire [95:0]       dataInMem_lo_1090 = {dataInMem_lo_hi_642, dataRegroupBySew_0_2_12};
  wire [63:0]       dataInMem_hi_hi_866 = {dataRegroupBySew_6_2_12, dataRegroupBySew_5_2_12};
  wire [127:0]      dataInMem_hi_1314 = {dataInMem_hi_hi_866, dataInMem_hi_lo_418};
  wire [95:0]       dataInMem_lo_1091 = {dataInMem_lo_hi_643, dataRegroupBySew_0_2_13};
  wire [63:0]       dataInMem_hi_hi_867 = {dataRegroupBySew_6_2_13, dataRegroupBySew_5_2_13};
  wire [127:0]      dataInMem_hi_1315 = {dataInMem_hi_hi_867, dataInMem_hi_lo_419};
  wire [95:0]       dataInMem_lo_1092 = {dataInMem_lo_hi_644, dataRegroupBySew_0_2_14};
  wire [63:0]       dataInMem_hi_hi_868 = {dataRegroupBySew_6_2_14, dataRegroupBySew_5_2_14};
  wire [127:0]      dataInMem_hi_1316 = {dataInMem_hi_hi_868, dataInMem_hi_lo_420};
  wire [95:0]       dataInMem_lo_1093 = {dataInMem_lo_hi_645, dataRegroupBySew_0_2_15};
  wire [63:0]       dataInMem_hi_hi_869 = {dataRegroupBySew_6_2_15, dataRegroupBySew_5_2_15};
  wire [127:0]      dataInMem_hi_1317 = {dataInMem_hi_hi_869, dataInMem_hi_lo_421};
  wire [95:0]       dataInMem_lo_1094 = {dataInMem_lo_hi_646, dataRegroupBySew_0_2_16};
  wire [63:0]       dataInMem_hi_hi_870 = {dataRegroupBySew_6_2_16, dataRegroupBySew_5_2_16};
  wire [127:0]      dataInMem_hi_1318 = {dataInMem_hi_hi_870, dataInMem_hi_lo_422};
  wire [95:0]       dataInMem_lo_1095 = {dataInMem_lo_hi_647, dataRegroupBySew_0_2_17};
  wire [63:0]       dataInMem_hi_hi_871 = {dataRegroupBySew_6_2_17, dataRegroupBySew_5_2_17};
  wire [127:0]      dataInMem_hi_1319 = {dataInMem_hi_hi_871, dataInMem_hi_lo_423};
  wire [95:0]       dataInMem_lo_1096 = {dataInMem_lo_hi_648, dataRegroupBySew_0_2_18};
  wire [63:0]       dataInMem_hi_hi_872 = {dataRegroupBySew_6_2_18, dataRegroupBySew_5_2_18};
  wire [127:0]      dataInMem_hi_1320 = {dataInMem_hi_hi_872, dataInMem_hi_lo_424};
  wire [95:0]       dataInMem_lo_1097 = {dataInMem_lo_hi_649, dataRegroupBySew_0_2_19};
  wire [63:0]       dataInMem_hi_hi_873 = {dataRegroupBySew_6_2_19, dataRegroupBySew_5_2_19};
  wire [127:0]      dataInMem_hi_1321 = {dataInMem_hi_hi_873, dataInMem_hi_lo_425};
  wire [95:0]       dataInMem_lo_1098 = {dataInMem_lo_hi_650, dataRegroupBySew_0_2_20};
  wire [63:0]       dataInMem_hi_hi_874 = {dataRegroupBySew_6_2_20, dataRegroupBySew_5_2_20};
  wire [127:0]      dataInMem_hi_1322 = {dataInMem_hi_hi_874, dataInMem_hi_lo_426};
  wire [95:0]       dataInMem_lo_1099 = {dataInMem_lo_hi_651, dataRegroupBySew_0_2_21};
  wire [63:0]       dataInMem_hi_hi_875 = {dataRegroupBySew_6_2_21, dataRegroupBySew_5_2_21};
  wire [127:0]      dataInMem_hi_1323 = {dataInMem_hi_hi_875, dataInMem_hi_lo_427};
  wire [95:0]       dataInMem_lo_1100 = {dataInMem_lo_hi_652, dataRegroupBySew_0_2_22};
  wire [63:0]       dataInMem_hi_hi_876 = {dataRegroupBySew_6_2_22, dataRegroupBySew_5_2_22};
  wire [127:0]      dataInMem_hi_1324 = {dataInMem_hi_hi_876, dataInMem_hi_lo_428};
  wire [95:0]       dataInMem_lo_1101 = {dataInMem_lo_hi_653, dataRegroupBySew_0_2_23};
  wire [63:0]       dataInMem_hi_hi_877 = {dataRegroupBySew_6_2_23, dataRegroupBySew_5_2_23};
  wire [127:0]      dataInMem_hi_1325 = {dataInMem_hi_hi_877, dataInMem_hi_lo_429};
  wire [95:0]       dataInMem_lo_1102 = {dataInMem_lo_hi_654, dataRegroupBySew_0_2_24};
  wire [63:0]       dataInMem_hi_hi_878 = {dataRegroupBySew_6_2_24, dataRegroupBySew_5_2_24};
  wire [127:0]      dataInMem_hi_1326 = {dataInMem_hi_hi_878, dataInMem_hi_lo_430};
  wire [95:0]       dataInMem_lo_1103 = {dataInMem_lo_hi_655, dataRegroupBySew_0_2_25};
  wire [63:0]       dataInMem_hi_hi_879 = {dataRegroupBySew_6_2_25, dataRegroupBySew_5_2_25};
  wire [127:0]      dataInMem_hi_1327 = {dataInMem_hi_hi_879, dataInMem_hi_lo_431};
  wire [95:0]       dataInMem_lo_1104 = {dataInMem_lo_hi_656, dataRegroupBySew_0_2_26};
  wire [63:0]       dataInMem_hi_hi_880 = {dataRegroupBySew_6_2_26, dataRegroupBySew_5_2_26};
  wire [127:0]      dataInMem_hi_1328 = {dataInMem_hi_hi_880, dataInMem_hi_lo_432};
  wire [95:0]       dataInMem_lo_1105 = {dataInMem_lo_hi_657, dataRegroupBySew_0_2_27};
  wire [63:0]       dataInMem_hi_hi_881 = {dataRegroupBySew_6_2_27, dataRegroupBySew_5_2_27};
  wire [127:0]      dataInMem_hi_1329 = {dataInMem_hi_hi_881, dataInMem_hi_lo_433};
  wire [95:0]       dataInMem_lo_1106 = {dataInMem_lo_hi_658, dataRegroupBySew_0_2_28};
  wire [63:0]       dataInMem_hi_hi_882 = {dataRegroupBySew_6_2_28, dataRegroupBySew_5_2_28};
  wire [127:0]      dataInMem_hi_1330 = {dataInMem_hi_hi_882, dataInMem_hi_lo_434};
  wire [95:0]       dataInMem_lo_1107 = {dataInMem_lo_hi_659, dataRegroupBySew_0_2_29};
  wire [63:0]       dataInMem_hi_hi_883 = {dataRegroupBySew_6_2_29, dataRegroupBySew_5_2_29};
  wire [127:0]      dataInMem_hi_1331 = {dataInMem_hi_hi_883, dataInMem_hi_lo_435};
  wire [95:0]       dataInMem_lo_1108 = {dataInMem_lo_hi_660, dataRegroupBySew_0_2_30};
  wire [63:0]       dataInMem_hi_hi_884 = {dataRegroupBySew_6_2_30, dataRegroupBySew_5_2_30};
  wire [127:0]      dataInMem_hi_1332 = {dataInMem_hi_hi_884, dataInMem_hi_lo_436};
  wire [95:0]       dataInMem_lo_1109 = {dataInMem_lo_hi_661, dataRegroupBySew_0_2_31};
  wire [63:0]       dataInMem_hi_hi_885 = {dataRegroupBySew_6_2_31, dataRegroupBySew_5_2_31};
  wire [127:0]      dataInMem_hi_1333 = {dataInMem_hi_hi_885, dataInMem_hi_lo_437};
  wire [447:0]      dataInMem_lo_lo_lo_lo_22 = {dataInMem_hi_1303, dataInMem_lo_1079, dataInMem_hi_1302, dataInMem_lo_1078};
  wire [447:0]      dataInMem_lo_lo_lo_hi_22 = {dataInMem_hi_1305, dataInMem_lo_1081, dataInMem_hi_1304, dataInMem_lo_1080};
  wire [895:0]      dataInMem_lo_lo_lo_22 = {dataInMem_lo_lo_lo_hi_22, dataInMem_lo_lo_lo_lo_22};
  wire [447:0]      dataInMem_lo_lo_hi_lo_22 = {dataInMem_hi_1307, dataInMem_lo_1083, dataInMem_hi_1306, dataInMem_lo_1082};
  wire [447:0]      dataInMem_lo_lo_hi_hi_22 = {dataInMem_hi_1309, dataInMem_lo_1085, dataInMem_hi_1308, dataInMem_lo_1084};
  wire [895:0]      dataInMem_lo_lo_hi_22 = {dataInMem_lo_lo_hi_hi_22, dataInMem_lo_lo_hi_lo_22};
  wire [1791:0]     dataInMem_lo_lo_214 = {dataInMem_lo_lo_hi_22, dataInMem_lo_lo_lo_22};
  wire [447:0]      dataInMem_lo_hi_lo_lo_22 = {dataInMem_hi_1311, dataInMem_lo_1087, dataInMem_hi_1310, dataInMem_lo_1086};
  wire [447:0]      dataInMem_lo_hi_lo_hi_22 = {dataInMem_hi_1313, dataInMem_lo_1089, dataInMem_hi_1312, dataInMem_lo_1088};
  wire [895:0]      dataInMem_lo_hi_lo_22 = {dataInMem_lo_hi_lo_hi_22, dataInMem_lo_hi_lo_lo_22};
  wire [447:0]      dataInMem_lo_hi_hi_lo_22 = {dataInMem_hi_1315, dataInMem_lo_1091, dataInMem_hi_1314, dataInMem_lo_1090};
  wire [447:0]      dataInMem_lo_hi_hi_hi_22 = {dataInMem_hi_1317, dataInMem_lo_1093, dataInMem_hi_1316, dataInMem_lo_1092};
  wire [895:0]      dataInMem_lo_hi_hi_22 = {dataInMem_lo_hi_hi_hi_22, dataInMem_lo_hi_hi_lo_22};
  wire [1791:0]     dataInMem_lo_hi_662 = {dataInMem_lo_hi_hi_22, dataInMem_lo_hi_lo_22};
  wire [3583:0]     dataInMem_lo_1110 = {dataInMem_lo_hi_662, dataInMem_lo_lo_214};
  wire [447:0]      dataInMem_hi_lo_lo_lo_22 = {dataInMem_hi_1319, dataInMem_lo_1095, dataInMem_hi_1318, dataInMem_lo_1094};
  wire [447:0]      dataInMem_hi_lo_lo_hi_22 = {dataInMem_hi_1321, dataInMem_lo_1097, dataInMem_hi_1320, dataInMem_lo_1096};
  wire [895:0]      dataInMem_hi_lo_lo_22 = {dataInMem_hi_lo_lo_hi_22, dataInMem_hi_lo_lo_lo_22};
  wire [447:0]      dataInMem_hi_lo_hi_lo_22 = {dataInMem_hi_1323, dataInMem_lo_1099, dataInMem_hi_1322, dataInMem_lo_1098};
  wire [447:0]      dataInMem_hi_lo_hi_hi_22 = {dataInMem_hi_1325, dataInMem_lo_1101, dataInMem_hi_1324, dataInMem_lo_1100};
  wire [895:0]      dataInMem_hi_lo_hi_22 = {dataInMem_hi_lo_hi_hi_22, dataInMem_hi_lo_hi_lo_22};
  wire [1791:0]     dataInMem_hi_lo_438 = {dataInMem_hi_lo_hi_22, dataInMem_hi_lo_lo_22};
  wire [447:0]      dataInMem_hi_hi_lo_lo_22 = {dataInMem_hi_1327, dataInMem_lo_1103, dataInMem_hi_1326, dataInMem_lo_1102};
  wire [447:0]      dataInMem_hi_hi_lo_hi_22 = {dataInMem_hi_1329, dataInMem_lo_1105, dataInMem_hi_1328, dataInMem_lo_1104};
  wire [895:0]      dataInMem_hi_hi_lo_22 = {dataInMem_hi_hi_lo_hi_22, dataInMem_hi_hi_lo_lo_22};
  wire [447:0]      dataInMem_hi_hi_hi_lo_22 = {dataInMem_hi_1331, dataInMem_lo_1107, dataInMem_hi_1330, dataInMem_lo_1106};
  wire [447:0]      dataInMem_hi_hi_hi_hi_22 = {dataInMem_hi_1333, dataInMem_lo_1109, dataInMem_hi_1332, dataInMem_lo_1108};
  wire [895:0]      dataInMem_hi_hi_hi_22 = {dataInMem_hi_hi_hi_hi_22, dataInMem_hi_hi_hi_lo_22};
  wire [1791:0]     dataInMem_hi_hi_886 = {dataInMem_hi_hi_hi_22, dataInMem_hi_hi_lo_22};
  wire [3583:0]     dataInMem_hi_1334 = {dataInMem_hi_hi_886, dataInMem_hi_lo_438};
  wire [7167:0]     dataInMem_22 = {dataInMem_hi_1334, dataInMem_lo_1110};
  wire [1023:0]     regroupCacheLine_22_0 = dataInMem_22[1023:0];
  wire [1023:0]     regroupCacheLine_22_1 = dataInMem_22[2047:1024];
  wire [1023:0]     regroupCacheLine_22_2 = dataInMem_22[3071:2048];
  wire [1023:0]     regroupCacheLine_22_3 = dataInMem_22[4095:3072];
  wire [1023:0]     regroupCacheLine_22_4 = dataInMem_22[5119:4096];
  wire [1023:0]     regroupCacheLine_22_5 = dataInMem_22[6143:5120];
  wire [1023:0]     regroupCacheLine_22_6 = dataInMem_22[7167:6144];
  wire [1023:0]     res_176 = regroupCacheLine_22_0;
  wire [1023:0]     res_177 = regroupCacheLine_22_1;
  wire [1023:0]     res_178 = regroupCacheLine_22_2;
  wire [1023:0]     res_179 = regroupCacheLine_22_3;
  wire [1023:0]     res_180 = regroupCacheLine_22_4;
  wire [1023:0]     res_181 = regroupCacheLine_22_5;
  wire [1023:0]     res_182 = regroupCacheLine_22_6;
  wire [2047:0]     lo_lo_22 = {res_177, res_176};
  wire [2047:0]     lo_hi_22 = {res_179, res_178};
  wire [4095:0]     lo_22 = {lo_hi_22, lo_lo_22};
  wire [2047:0]     hi_lo_22 = {res_181, res_180};
  wire [2047:0]     hi_hi_22 = {1024'h0, res_182};
  wire [4095:0]     hi_22 = {hi_hi_22, hi_lo_22};
  wire [8191:0]     regroupLoadData_2_6 = {hi_22, lo_22};
  wire [127:0]      dataInMem_lo_1111 = {dataInMem_lo_hi_663, dataInMem_lo_lo_215};
  wire [63:0]       dataInMem_hi_hi_887 = {dataRegroupBySew_7_2_0, dataRegroupBySew_6_2_0};
  wire [127:0]      dataInMem_hi_1335 = {dataInMem_hi_hi_887, dataInMem_hi_lo_439};
  wire [127:0]      dataInMem_lo_1112 = {dataInMem_lo_hi_664, dataInMem_lo_lo_216};
  wire [63:0]       dataInMem_hi_hi_888 = {dataRegroupBySew_7_2_1, dataRegroupBySew_6_2_1};
  wire [127:0]      dataInMem_hi_1336 = {dataInMem_hi_hi_888, dataInMem_hi_lo_440};
  wire [127:0]      dataInMem_lo_1113 = {dataInMem_lo_hi_665, dataInMem_lo_lo_217};
  wire [63:0]       dataInMem_hi_hi_889 = {dataRegroupBySew_7_2_2, dataRegroupBySew_6_2_2};
  wire [127:0]      dataInMem_hi_1337 = {dataInMem_hi_hi_889, dataInMem_hi_lo_441};
  wire [127:0]      dataInMem_lo_1114 = {dataInMem_lo_hi_666, dataInMem_lo_lo_218};
  wire [63:0]       dataInMem_hi_hi_890 = {dataRegroupBySew_7_2_3, dataRegroupBySew_6_2_3};
  wire [127:0]      dataInMem_hi_1338 = {dataInMem_hi_hi_890, dataInMem_hi_lo_442};
  wire [127:0]      dataInMem_lo_1115 = {dataInMem_lo_hi_667, dataInMem_lo_lo_219};
  wire [63:0]       dataInMem_hi_hi_891 = {dataRegroupBySew_7_2_4, dataRegroupBySew_6_2_4};
  wire [127:0]      dataInMem_hi_1339 = {dataInMem_hi_hi_891, dataInMem_hi_lo_443};
  wire [127:0]      dataInMem_lo_1116 = {dataInMem_lo_hi_668, dataInMem_lo_lo_220};
  wire [63:0]       dataInMem_hi_hi_892 = {dataRegroupBySew_7_2_5, dataRegroupBySew_6_2_5};
  wire [127:0]      dataInMem_hi_1340 = {dataInMem_hi_hi_892, dataInMem_hi_lo_444};
  wire [127:0]      dataInMem_lo_1117 = {dataInMem_lo_hi_669, dataInMem_lo_lo_221};
  wire [63:0]       dataInMem_hi_hi_893 = {dataRegroupBySew_7_2_6, dataRegroupBySew_6_2_6};
  wire [127:0]      dataInMem_hi_1341 = {dataInMem_hi_hi_893, dataInMem_hi_lo_445};
  wire [127:0]      dataInMem_lo_1118 = {dataInMem_lo_hi_670, dataInMem_lo_lo_222};
  wire [63:0]       dataInMem_hi_hi_894 = {dataRegroupBySew_7_2_7, dataRegroupBySew_6_2_7};
  wire [127:0]      dataInMem_hi_1342 = {dataInMem_hi_hi_894, dataInMem_hi_lo_446};
  wire [127:0]      dataInMem_lo_1119 = {dataInMem_lo_hi_671, dataInMem_lo_lo_223};
  wire [63:0]       dataInMem_hi_hi_895 = {dataRegroupBySew_7_2_8, dataRegroupBySew_6_2_8};
  wire [127:0]      dataInMem_hi_1343 = {dataInMem_hi_hi_895, dataInMem_hi_lo_447};
  wire [127:0]      dataInMem_lo_1120 = {dataInMem_lo_hi_672, dataInMem_lo_lo_224};
  wire [63:0]       dataInMem_hi_hi_896 = {dataRegroupBySew_7_2_9, dataRegroupBySew_6_2_9};
  wire [127:0]      dataInMem_hi_1344 = {dataInMem_hi_hi_896, dataInMem_hi_lo_448};
  wire [127:0]      dataInMem_lo_1121 = {dataInMem_lo_hi_673, dataInMem_lo_lo_225};
  wire [63:0]       dataInMem_hi_hi_897 = {dataRegroupBySew_7_2_10, dataRegroupBySew_6_2_10};
  wire [127:0]      dataInMem_hi_1345 = {dataInMem_hi_hi_897, dataInMem_hi_lo_449};
  wire [127:0]      dataInMem_lo_1122 = {dataInMem_lo_hi_674, dataInMem_lo_lo_226};
  wire [63:0]       dataInMem_hi_hi_898 = {dataRegroupBySew_7_2_11, dataRegroupBySew_6_2_11};
  wire [127:0]      dataInMem_hi_1346 = {dataInMem_hi_hi_898, dataInMem_hi_lo_450};
  wire [127:0]      dataInMem_lo_1123 = {dataInMem_lo_hi_675, dataInMem_lo_lo_227};
  wire [63:0]       dataInMem_hi_hi_899 = {dataRegroupBySew_7_2_12, dataRegroupBySew_6_2_12};
  wire [127:0]      dataInMem_hi_1347 = {dataInMem_hi_hi_899, dataInMem_hi_lo_451};
  wire [127:0]      dataInMem_lo_1124 = {dataInMem_lo_hi_676, dataInMem_lo_lo_228};
  wire [63:0]       dataInMem_hi_hi_900 = {dataRegroupBySew_7_2_13, dataRegroupBySew_6_2_13};
  wire [127:0]      dataInMem_hi_1348 = {dataInMem_hi_hi_900, dataInMem_hi_lo_452};
  wire [127:0]      dataInMem_lo_1125 = {dataInMem_lo_hi_677, dataInMem_lo_lo_229};
  wire [63:0]       dataInMem_hi_hi_901 = {dataRegroupBySew_7_2_14, dataRegroupBySew_6_2_14};
  wire [127:0]      dataInMem_hi_1349 = {dataInMem_hi_hi_901, dataInMem_hi_lo_453};
  wire [127:0]      dataInMem_lo_1126 = {dataInMem_lo_hi_678, dataInMem_lo_lo_230};
  wire [63:0]       dataInMem_hi_hi_902 = {dataRegroupBySew_7_2_15, dataRegroupBySew_6_2_15};
  wire [127:0]      dataInMem_hi_1350 = {dataInMem_hi_hi_902, dataInMem_hi_lo_454};
  wire [127:0]      dataInMem_lo_1127 = {dataInMem_lo_hi_679, dataInMem_lo_lo_231};
  wire [63:0]       dataInMem_hi_hi_903 = {dataRegroupBySew_7_2_16, dataRegroupBySew_6_2_16};
  wire [127:0]      dataInMem_hi_1351 = {dataInMem_hi_hi_903, dataInMem_hi_lo_455};
  wire [127:0]      dataInMem_lo_1128 = {dataInMem_lo_hi_680, dataInMem_lo_lo_232};
  wire [63:0]       dataInMem_hi_hi_904 = {dataRegroupBySew_7_2_17, dataRegroupBySew_6_2_17};
  wire [127:0]      dataInMem_hi_1352 = {dataInMem_hi_hi_904, dataInMem_hi_lo_456};
  wire [127:0]      dataInMem_lo_1129 = {dataInMem_lo_hi_681, dataInMem_lo_lo_233};
  wire [63:0]       dataInMem_hi_hi_905 = {dataRegroupBySew_7_2_18, dataRegroupBySew_6_2_18};
  wire [127:0]      dataInMem_hi_1353 = {dataInMem_hi_hi_905, dataInMem_hi_lo_457};
  wire [127:0]      dataInMem_lo_1130 = {dataInMem_lo_hi_682, dataInMem_lo_lo_234};
  wire [63:0]       dataInMem_hi_hi_906 = {dataRegroupBySew_7_2_19, dataRegroupBySew_6_2_19};
  wire [127:0]      dataInMem_hi_1354 = {dataInMem_hi_hi_906, dataInMem_hi_lo_458};
  wire [127:0]      dataInMem_lo_1131 = {dataInMem_lo_hi_683, dataInMem_lo_lo_235};
  wire [63:0]       dataInMem_hi_hi_907 = {dataRegroupBySew_7_2_20, dataRegroupBySew_6_2_20};
  wire [127:0]      dataInMem_hi_1355 = {dataInMem_hi_hi_907, dataInMem_hi_lo_459};
  wire [127:0]      dataInMem_lo_1132 = {dataInMem_lo_hi_684, dataInMem_lo_lo_236};
  wire [63:0]       dataInMem_hi_hi_908 = {dataRegroupBySew_7_2_21, dataRegroupBySew_6_2_21};
  wire [127:0]      dataInMem_hi_1356 = {dataInMem_hi_hi_908, dataInMem_hi_lo_460};
  wire [127:0]      dataInMem_lo_1133 = {dataInMem_lo_hi_685, dataInMem_lo_lo_237};
  wire [63:0]       dataInMem_hi_hi_909 = {dataRegroupBySew_7_2_22, dataRegroupBySew_6_2_22};
  wire [127:0]      dataInMem_hi_1357 = {dataInMem_hi_hi_909, dataInMem_hi_lo_461};
  wire [127:0]      dataInMem_lo_1134 = {dataInMem_lo_hi_686, dataInMem_lo_lo_238};
  wire [63:0]       dataInMem_hi_hi_910 = {dataRegroupBySew_7_2_23, dataRegroupBySew_6_2_23};
  wire [127:0]      dataInMem_hi_1358 = {dataInMem_hi_hi_910, dataInMem_hi_lo_462};
  wire [127:0]      dataInMem_lo_1135 = {dataInMem_lo_hi_687, dataInMem_lo_lo_239};
  wire [63:0]       dataInMem_hi_hi_911 = {dataRegroupBySew_7_2_24, dataRegroupBySew_6_2_24};
  wire [127:0]      dataInMem_hi_1359 = {dataInMem_hi_hi_911, dataInMem_hi_lo_463};
  wire [127:0]      dataInMem_lo_1136 = {dataInMem_lo_hi_688, dataInMem_lo_lo_240};
  wire [63:0]       dataInMem_hi_hi_912 = {dataRegroupBySew_7_2_25, dataRegroupBySew_6_2_25};
  wire [127:0]      dataInMem_hi_1360 = {dataInMem_hi_hi_912, dataInMem_hi_lo_464};
  wire [127:0]      dataInMem_lo_1137 = {dataInMem_lo_hi_689, dataInMem_lo_lo_241};
  wire [63:0]       dataInMem_hi_hi_913 = {dataRegroupBySew_7_2_26, dataRegroupBySew_6_2_26};
  wire [127:0]      dataInMem_hi_1361 = {dataInMem_hi_hi_913, dataInMem_hi_lo_465};
  wire [127:0]      dataInMem_lo_1138 = {dataInMem_lo_hi_690, dataInMem_lo_lo_242};
  wire [63:0]       dataInMem_hi_hi_914 = {dataRegroupBySew_7_2_27, dataRegroupBySew_6_2_27};
  wire [127:0]      dataInMem_hi_1362 = {dataInMem_hi_hi_914, dataInMem_hi_lo_466};
  wire [127:0]      dataInMem_lo_1139 = {dataInMem_lo_hi_691, dataInMem_lo_lo_243};
  wire [63:0]       dataInMem_hi_hi_915 = {dataRegroupBySew_7_2_28, dataRegroupBySew_6_2_28};
  wire [127:0]      dataInMem_hi_1363 = {dataInMem_hi_hi_915, dataInMem_hi_lo_467};
  wire [127:0]      dataInMem_lo_1140 = {dataInMem_lo_hi_692, dataInMem_lo_lo_244};
  wire [63:0]       dataInMem_hi_hi_916 = {dataRegroupBySew_7_2_29, dataRegroupBySew_6_2_29};
  wire [127:0]      dataInMem_hi_1364 = {dataInMem_hi_hi_916, dataInMem_hi_lo_468};
  wire [127:0]      dataInMem_lo_1141 = {dataInMem_lo_hi_693, dataInMem_lo_lo_245};
  wire [63:0]       dataInMem_hi_hi_917 = {dataRegroupBySew_7_2_30, dataRegroupBySew_6_2_30};
  wire [127:0]      dataInMem_hi_1365 = {dataInMem_hi_hi_917, dataInMem_hi_lo_469};
  wire [127:0]      dataInMem_lo_1142 = {dataInMem_lo_hi_694, dataInMem_lo_lo_246};
  wire [63:0]       dataInMem_hi_hi_918 = {dataRegroupBySew_7_2_31, dataRegroupBySew_6_2_31};
  wire [127:0]      dataInMem_hi_1366 = {dataInMem_hi_hi_918, dataInMem_hi_lo_470};
  wire [511:0]      dataInMem_lo_lo_lo_lo_23 = {dataInMem_hi_1336, dataInMem_lo_1112, dataInMem_hi_1335, dataInMem_lo_1111};
  wire [511:0]      dataInMem_lo_lo_lo_hi_23 = {dataInMem_hi_1338, dataInMem_lo_1114, dataInMem_hi_1337, dataInMem_lo_1113};
  wire [1023:0]     dataInMem_lo_lo_lo_23 = {dataInMem_lo_lo_lo_hi_23, dataInMem_lo_lo_lo_lo_23};
  wire [511:0]      dataInMem_lo_lo_hi_lo_23 = {dataInMem_hi_1340, dataInMem_lo_1116, dataInMem_hi_1339, dataInMem_lo_1115};
  wire [511:0]      dataInMem_lo_lo_hi_hi_23 = {dataInMem_hi_1342, dataInMem_lo_1118, dataInMem_hi_1341, dataInMem_lo_1117};
  wire [1023:0]     dataInMem_lo_lo_hi_23 = {dataInMem_lo_lo_hi_hi_23, dataInMem_lo_lo_hi_lo_23};
  wire [2047:0]     dataInMem_lo_lo_247 = {dataInMem_lo_lo_hi_23, dataInMem_lo_lo_lo_23};
  wire [511:0]      dataInMem_lo_hi_lo_lo_23 = {dataInMem_hi_1344, dataInMem_lo_1120, dataInMem_hi_1343, dataInMem_lo_1119};
  wire [511:0]      dataInMem_lo_hi_lo_hi_23 = {dataInMem_hi_1346, dataInMem_lo_1122, dataInMem_hi_1345, dataInMem_lo_1121};
  wire [1023:0]     dataInMem_lo_hi_lo_23 = {dataInMem_lo_hi_lo_hi_23, dataInMem_lo_hi_lo_lo_23};
  wire [511:0]      dataInMem_lo_hi_hi_lo_23 = {dataInMem_hi_1348, dataInMem_lo_1124, dataInMem_hi_1347, dataInMem_lo_1123};
  wire [511:0]      dataInMem_lo_hi_hi_hi_23 = {dataInMem_hi_1350, dataInMem_lo_1126, dataInMem_hi_1349, dataInMem_lo_1125};
  wire [1023:0]     dataInMem_lo_hi_hi_23 = {dataInMem_lo_hi_hi_hi_23, dataInMem_lo_hi_hi_lo_23};
  wire [2047:0]     dataInMem_lo_hi_695 = {dataInMem_lo_hi_hi_23, dataInMem_lo_hi_lo_23};
  wire [4095:0]     dataInMem_lo_1143 = {dataInMem_lo_hi_695, dataInMem_lo_lo_247};
  wire [511:0]      dataInMem_hi_lo_lo_lo_23 = {dataInMem_hi_1352, dataInMem_lo_1128, dataInMem_hi_1351, dataInMem_lo_1127};
  wire [511:0]      dataInMem_hi_lo_lo_hi_23 = {dataInMem_hi_1354, dataInMem_lo_1130, dataInMem_hi_1353, dataInMem_lo_1129};
  wire [1023:0]     dataInMem_hi_lo_lo_23 = {dataInMem_hi_lo_lo_hi_23, dataInMem_hi_lo_lo_lo_23};
  wire [511:0]      dataInMem_hi_lo_hi_lo_23 = {dataInMem_hi_1356, dataInMem_lo_1132, dataInMem_hi_1355, dataInMem_lo_1131};
  wire [511:0]      dataInMem_hi_lo_hi_hi_23 = {dataInMem_hi_1358, dataInMem_lo_1134, dataInMem_hi_1357, dataInMem_lo_1133};
  wire [1023:0]     dataInMem_hi_lo_hi_23 = {dataInMem_hi_lo_hi_hi_23, dataInMem_hi_lo_hi_lo_23};
  wire [2047:0]     dataInMem_hi_lo_471 = {dataInMem_hi_lo_hi_23, dataInMem_hi_lo_lo_23};
  wire [511:0]      dataInMem_hi_hi_lo_lo_23 = {dataInMem_hi_1360, dataInMem_lo_1136, dataInMem_hi_1359, dataInMem_lo_1135};
  wire [511:0]      dataInMem_hi_hi_lo_hi_23 = {dataInMem_hi_1362, dataInMem_lo_1138, dataInMem_hi_1361, dataInMem_lo_1137};
  wire [1023:0]     dataInMem_hi_hi_lo_23 = {dataInMem_hi_hi_lo_hi_23, dataInMem_hi_hi_lo_lo_23};
  wire [511:0]      dataInMem_hi_hi_hi_lo_23 = {dataInMem_hi_1364, dataInMem_lo_1140, dataInMem_hi_1363, dataInMem_lo_1139};
  wire [511:0]      dataInMem_hi_hi_hi_hi_23 = {dataInMem_hi_1366, dataInMem_lo_1142, dataInMem_hi_1365, dataInMem_lo_1141};
  wire [1023:0]     dataInMem_hi_hi_hi_23 = {dataInMem_hi_hi_hi_hi_23, dataInMem_hi_hi_hi_lo_23};
  wire [2047:0]     dataInMem_hi_hi_919 = {dataInMem_hi_hi_hi_23, dataInMem_hi_hi_lo_23};
  wire [4095:0]     dataInMem_hi_1367 = {dataInMem_hi_hi_919, dataInMem_hi_lo_471};
  wire [8191:0]     dataInMem_23 = {dataInMem_hi_1367, dataInMem_lo_1143};
  wire [1023:0]     regroupCacheLine_23_0 = dataInMem_23[1023:0];
  wire [1023:0]     regroupCacheLine_23_1 = dataInMem_23[2047:1024];
  wire [1023:0]     regroupCacheLine_23_2 = dataInMem_23[3071:2048];
  wire [1023:0]     regroupCacheLine_23_3 = dataInMem_23[4095:3072];
  wire [1023:0]     regroupCacheLine_23_4 = dataInMem_23[5119:4096];
  wire [1023:0]     regroupCacheLine_23_5 = dataInMem_23[6143:5120];
  wire [1023:0]     regroupCacheLine_23_6 = dataInMem_23[7167:6144];
  wire [1023:0]     regroupCacheLine_23_7 = dataInMem_23[8191:7168];
  wire [1023:0]     res_184 = regroupCacheLine_23_0;
  wire [1023:0]     res_185 = regroupCacheLine_23_1;
  wire [1023:0]     res_186 = regroupCacheLine_23_2;
  wire [1023:0]     res_187 = regroupCacheLine_23_3;
  wire [1023:0]     res_188 = regroupCacheLine_23_4;
  wire [1023:0]     res_189 = regroupCacheLine_23_5;
  wire [1023:0]     res_190 = regroupCacheLine_23_6;
  wire [1023:0]     res_191 = regroupCacheLine_23_7;
  wire [2047:0]     lo_lo_23 = {res_185, res_184};
  wire [2047:0]     lo_hi_23 = {res_187, res_186};
  wire [4095:0]     lo_23 = {lo_hi_23, lo_lo_23};
  wire [2047:0]     hi_lo_23 = {res_189, res_188};
  wire [2047:0]     hi_hi_23 = {res_191, res_190};
  wire [4095:0]     hi_23 = {hi_hi_23, hi_lo_23};
  wire [8191:0]     regroupLoadData_2_7 = {hi_23, lo_23};
  wire              _GEN_1126 = lsuRequest_valid | accessBufferDequeueFire;
  wire              _GEN_1127 = isLastDataGroup & ~isLastMaskGroup;
  wire              _maskSelect_valid_output = _GEN_1126 & _GEN_1127;
  wire [7:0][127:0] _GEN_1128 = {{maskForBufferData_7}, {maskForBufferData_6}, {maskForBufferData_5}, {maskForBufferData_4}, {maskForBufferData_3}, {maskForBufferData_2}, {maskForBufferData_1}, {maskForBufferData_0}};
  wire [127:0]      _GEN_1129 = _GEN_1128[cacheLineIndexInBuffer];
  wire              needSendTail = {7'h0, bufferBaseCacheLineIndex} == cacheLineNumberReg;
  assign memRequest_valid_0 = (bufferValid | canSendTail & needSendTail) & addressQueueFree;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo = {cacheLineTemp[8], cacheLineTemp[0]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi = {cacheLineTemp[24], cacheLineTemp[16]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo = {cacheLineTemp[40], cacheLineTemp[32]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi = {cacheLineTemp[56], cacheLineTemp[48]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo = {cacheLineTemp[72], cacheLineTemp[64]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi = {cacheLineTemp[88], cacheLineTemp[80]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo = {cacheLineTemp[104], cacheLineTemp[96]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi = {cacheLineTemp[120], cacheLineTemp[112]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi = {memRequest_bits_data_lo_lo_lo_lo_hi_hi, memRequest_bits_data_lo_lo_lo_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo = {cacheLineTemp[136], cacheLineTemp[128]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi = {cacheLineTemp[152], cacheLineTemp[144]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo = {cacheLineTemp[168], cacheLineTemp[160]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi = {cacheLineTemp[184], cacheLineTemp[176]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo = {memRequest_bits_data_lo_lo_lo_hi_lo_hi, memRequest_bits_data_lo_lo_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo = {cacheLineTemp[200], cacheLineTemp[192]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi = {cacheLineTemp[216], cacheLineTemp[208]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo = {cacheLineTemp[232], cacheLineTemp[224]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi = {cacheLineTemp[248], cacheLineTemp[240]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi = {memRequest_bits_data_lo_lo_lo_hi_hi_hi, memRequest_bits_data_lo_lo_lo_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi = {memRequest_bits_data_lo_lo_lo_hi_hi, memRequest_bits_data_lo_lo_lo_hi_lo};
  wire [31:0]       memRequest_bits_data_lo_lo_lo = {memRequest_bits_data_lo_lo_lo_hi, memRequest_bits_data_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo = {cacheLineTemp[264], cacheLineTemp[256]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi = {cacheLineTemp[280], cacheLineTemp[272]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo = {cacheLineTemp[296], cacheLineTemp[288]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi = {cacheLineTemp[312], cacheLineTemp[304]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo = {memRequest_bits_data_lo_lo_hi_lo_lo_hi, memRequest_bits_data_lo_lo_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo = {cacheLineTemp[328], cacheLineTemp[320]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi = {cacheLineTemp[344], cacheLineTemp[336]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo = {cacheLineTemp[360], cacheLineTemp[352]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi = {cacheLineTemp[376], cacheLineTemp[368]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi = {memRequest_bits_data_lo_lo_hi_lo_hi_hi, memRequest_bits_data_lo_lo_hi_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo = {memRequest_bits_data_lo_lo_hi_lo_hi, memRequest_bits_data_lo_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo = {cacheLineTemp[392], cacheLineTemp[384]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi = {cacheLineTemp[408], cacheLineTemp[400]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo = {cacheLineTemp[424], cacheLineTemp[416]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi = {cacheLineTemp[440], cacheLineTemp[432]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo = {memRequest_bits_data_lo_lo_hi_hi_lo_hi, memRequest_bits_data_lo_lo_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo = {cacheLineTemp[456], cacheLineTemp[448]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi = {cacheLineTemp[472], cacheLineTemp[464]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo = {cacheLineTemp[488], cacheLineTemp[480]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi = {cacheLineTemp[504], cacheLineTemp[496]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi = {memRequest_bits_data_lo_lo_hi_hi_hi_hi, memRequest_bits_data_lo_lo_hi_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi = {memRequest_bits_data_lo_lo_hi_hi_hi, memRequest_bits_data_lo_lo_hi_hi_lo};
  wire [31:0]       memRequest_bits_data_lo_lo_hi = {memRequest_bits_data_lo_lo_hi_hi, memRequest_bits_data_lo_lo_hi_lo};
  wire [63:0]       memRequest_bits_data_lo_lo = {memRequest_bits_data_lo_lo_hi, memRequest_bits_data_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo = {cacheLineTemp[520], cacheLineTemp[512]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi = {cacheLineTemp[536], cacheLineTemp[528]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo = {cacheLineTemp[552], cacheLineTemp[544]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi = {cacheLineTemp[568], cacheLineTemp[560]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo = {memRequest_bits_data_lo_hi_lo_lo_lo_hi, memRequest_bits_data_lo_hi_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo = {cacheLineTemp[584], cacheLineTemp[576]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi = {cacheLineTemp[600], cacheLineTemp[592]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo = {cacheLineTemp[616], cacheLineTemp[608]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi = {cacheLineTemp[632], cacheLineTemp[624]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi = {memRequest_bits_data_lo_hi_lo_lo_hi_hi, memRequest_bits_data_lo_hi_lo_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo = {memRequest_bits_data_lo_hi_lo_lo_hi, memRequest_bits_data_lo_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo = {cacheLineTemp[648], cacheLineTemp[640]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi = {cacheLineTemp[664], cacheLineTemp[656]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo = {cacheLineTemp[680], cacheLineTemp[672]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi = {cacheLineTemp[696], cacheLineTemp[688]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo = {memRequest_bits_data_lo_hi_lo_hi_lo_hi, memRequest_bits_data_lo_hi_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo = {cacheLineTemp[712], cacheLineTemp[704]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi = {cacheLineTemp[728], cacheLineTemp[720]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo = {cacheLineTemp[744], cacheLineTemp[736]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi = {cacheLineTemp[760], cacheLineTemp[752]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi = {memRequest_bits_data_lo_hi_lo_hi_hi_hi, memRequest_bits_data_lo_hi_lo_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi = {memRequest_bits_data_lo_hi_lo_hi_hi, memRequest_bits_data_lo_hi_lo_hi_lo};
  wire [31:0]       memRequest_bits_data_lo_hi_lo = {memRequest_bits_data_lo_hi_lo_hi, memRequest_bits_data_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo = {cacheLineTemp[776], cacheLineTemp[768]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi = {cacheLineTemp[792], cacheLineTemp[784]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo = {cacheLineTemp[808], cacheLineTemp[800]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi = {cacheLineTemp[824], cacheLineTemp[816]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo = {memRequest_bits_data_lo_hi_hi_lo_lo_hi, memRequest_bits_data_lo_hi_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo = {cacheLineTemp[840], cacheLineTemp[832]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi = {cacheLineTemp[856], cacheLineTemp[848]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo = {cacheLineTemp[872], cacheLineTemp[864]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi = {cacheLineTemp[888], cacheLineTemp[880]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi = {memRequest_bits_data_lo_hi_hi_lo_hi_hi, memRequest_bits_data_lo_hi_hi_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo = {memRequest_bits_data_lo_hi_hi_lo_hi, memRequest_bits_data_lo_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo = {cacheLineTemp[904], cacheLineTemp[896]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi = {cacheLineTemp[920], cacheLineTemp[912]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo = {cacheLineTemp[936], cacheLineTemp[928]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi = {cacheLineTemp[952], cacheLineTemp[944]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo = {memRequest_bits_data_lo_hi_hi_hi_lo_hi, memRequest_bits_data_lo_hi_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo = {cacheLineTemp[968], cacheLineTemp[960]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi = {cacheLineTemp[984], cacheLineTemp[976]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo = {cacheLineTemp[1000], cacheLineTemp[992]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi = {cacheLineTemp[1016], cacheLineTemp[1008]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi = {memRequest_bits_data_lo_hi_hi_hi_hi_hi, memRequest_bits_data_lo_hi_hi_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi = {memRequest_bits_data_lo_hi_hi_hi_hi, memRequest_bits_data_lo_hi_hi_hi_lo};
  wire [31:0]       memRequest_bits_data_lo_hi_hi = {memRequest_bits_data_lo_hi_hi_hi, memRequest_bits_data_lo_hi_hi_lo};
  wire [63:0]       memRequest_bits_data_lo_hi = {memRequest_bits_data_lo_hi_hi, memRequest_bits_data_lo_hi_lo};
  wire [127:0]      memRequest_bits_data_lo = {memRequest_bits_data_lo_hi, memRequest_bits_data_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo = {dataBuffer_0[8], dataBuffer_0[0]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi = {dataBuffer_0[24], dataBuffer_0[16]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo = {dataBuffer_0[40], dataBuffer_0[32]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi = {dataBuffer_0[56], dataBuffer_0[48]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo = {memRequest_bits_data_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo = {dataBuffer_0[72], dataBuffer_0[64]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi = {dataBuffer_0[88], dataBuffer_0[80]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo = {dataBuffer_0[104], dataBuffer_0[96]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi = {dataBuffer_0[120], dataBuffer_0[112]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_lo_lo_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo = {memRequest_bits_data_hi_lo_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo = {dataBuffer_0[136], dataBuffer_0[128]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi = {dataBuffer_0[152], dataBuffer_0[144]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo = {dataBuffer_0[168], dataBuffer_0[160]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi = {dataBuffer_0[184], dataBuffer_0[176]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo = {memRequest_bits_data_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_lo_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo = {dataBuffer_0[200], dataBuffer_0[192]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi = {dataBuffer_0[216], dataBuffer_0[208]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo = {dataBuffer_0[232], dataBuffer_0[224]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi = {dataBuffer_0[248], dataBuffer_0[240]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_lo_lo_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi = {memRequest_bits_data_hi_lo_lo_hi_hi, memRequest_bits_data_hi_lo_lo_hi_lo};
  wire [31:0]       memRequest_bits_data_hi_lo_lo = {memRequest_bits_data_hi_lo_lo_hi, memRequest_bits_data_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo = {dataBuffer_0[264], dataBuffer_0[256]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi = {dataBuffer_0[280], dataBuffer_0[272]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo = {dataBuffer_0[296], dataBuffer_0[288]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi = {dataBuffer_0[312], dataBuffer_0[304]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo = {memRequest_bits_data_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_lo_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo = {dataBuffer_0[328], dataBuffer_0[320]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi = {dataBuffer_0[344], dataBuffer_0[336]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo = {dataBuffer_0[360], dataBuffer_0[352]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi = {dataBuffer_0[376], dataBuffer_0[368]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_lo_hi_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo = {memRequest_bits_data_hi_lo_hi_lo_hi, memRequest_bits_data_hi_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo = {dataBuffer_0[392], dataBuffer_0[384]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi = {dataBuffer_0[408], dataBuffer_0[400]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo = {dataBuffer_0[424], dataBuffer_0[416]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi = {dataBuffer_0[440], dataBuffer_0[432]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo = {memRequest_bits_data_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_lo_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo = {dataBuffer_0[456], dataBuffer_0[448]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi = {dataBuffer_0[472], dataBuffer_0[464]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo = {dataBuffer_0[488], dataBuffer_0[480]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi = {dataBuffer_0[504], dataBuffer_0[496]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_lo_hi_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi = {memRequest_bits_data_hi_lo_hi_hi_hi, memRequest_bits_data_hi_lo_hi_hi_lo};
  wire [31:0]       memRequest_bits_data_hi_lo_hi = {memRequest_bits_data_hi_lo_hi_hi, memRequest_bits_data_hi_lo_hi_lo};
  wire [63:0]       memRequest_bits_data_hi_lo = {memRequest_bits_data_hi_lo_hi, memRequest_bits_data_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo = {dataBuffer_0[520], dataBuffer_0[512]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi = {dataBuffer_0[536], dataBuffer_0[528]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo = {dataBuffer_0[552], dataBuffer_0[544]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi = {dataBuffer_0[568], dataBuffer_0[560]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo = {memRequest_bits_data_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_hi_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo = {dataBuffer_0[584], dataBuffer_0[576]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi = {dataBuffer_0[600], dataBuffer_0[592]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo = {dataBuffer_0[616], dataBuffer_0[608]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi = {dataBuffer_0[632], dataBuffer_0[624]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_hi_lo_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo = {memRequest_bits_data_hi_hi_lo_lo_hi, memRequest_bits_data_hi_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo = {dataBuffer_0[648], dataBuffer_0[640]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi = {dataBuffer_0[664], dataBuffer_0[656]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo = {dataBuffer_0[680], dataBuffer_0[672]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi = {dataBuffer_0[696], dataBuffer_0[688]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo = {memRequest_bits_data_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_hi_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo = {dataBuffer_0[712], dataBuffer_0[704]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi = {dataBuffer_0[728], dataBuffer_0[720]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo = {dataBuffer_0[744], dataBuffer_0[736]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi = {dataBuffer_0[760], dataBuffer_0[752]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_hi_lo_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi = {memRequest_bits_data_hi_hi_lo_hi_hi, memRequest_bits_data_hi_hi_lo_hi_lo};
  wire [31:0]       memRequest_bits_data_hi_hi_lo = {memRequest_bits_data_hi_hi_lo_hi, memRequest_bits_data_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo = {dataBuffer_0[776], dataBuffer_0[768]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi = {dataBuffer_0[792], dataBuffer_0[784]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo = {dataBuffer_0[808], dataBuffer_0[800]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi = {dataBuffer_0[824], dataBuffer_0[816]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo = {memRequest_bits_data_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_hi_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo = {dataBuffer_0[840], dataBuffer_0[832]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi = {dataBuffer_0[856], dataBuffer_0[848]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo = {dataBuffer_0[872], dataBuffer_0[864]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi = {dataBuffer_0[888], dataBuffer_0[880]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_hi_hi_lo_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo = {memRequest_bits_data_hi_hi_hi_lo_hi, memRequest_bits_data_hi_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo = {dataBuffer_0[904], dataBuffer_0[896]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi = {dataBuffer_0[920], dataBuffer_0[912]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo = {dataBuffer_0[936], dataBuffer_0[928]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi = {dataBuffer_0[952], dataBuffer_0[944]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo = {memRequest_bits_data_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_hi_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo = {dataBuffer_0[968], dataBuffer_0[960]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi = {dataBuffer_0[984], dataBuffer_0[976]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo = {dataBuffer_0[1000], dataBuffer_0[992]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi = {dataBuffer_0[1016], dataBuffer_0[1008]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_hi_hi_lo};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_hi_lo};
  wire [31:0]       memRequest_bits_data_hi_hi_hi = {memRequest_bits_data_hi_hi_hi_hi, memRequest_bits_data_hi_hi_hi_lo};
  wire [63:0]       memRequest_bits_data_hi_hi = {memRequest_bits_data_hi_hi_hi, memRequest_bits_data_hi_hi_lo};
  wire [127:0]      memRequest_bits_data_hi = {memRequest_bits_data_hi_hi, memRequest_bits_data_hi_lo};
  wire [382:0]      _GEN_1130 = {376'h0, initOffset};
  wire [382:0]      _memRequest_bits_data_T_2050 = {127'h0, memRequest_bits_data_hi, memRequest_bits_data_lo} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_1 = {cacheLineTemp[9], cacheLineTemp[1]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_1 = {cacheLineTemp[25], cacheLineTemp[17]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_1 = {cacheLineTemp[41], cacheLineTemp[33]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_1 = {cacheLineTemp[57], cacheLineTemp[49]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_1 = {cacheLineTemp[73], cacheLineTemp[65]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_1 = {cacheLineTemp[89], cacheLineTemp[81]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_1 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_1 = {cacheLineTemp[105], cacheLineTemp[97]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_1 = {cacheLineTemp[121], cacheLineTemp[113]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_1 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_1, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_lo_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_1 = {cacheLineTemp[137], cacheLineTemp[129]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_1 = {cacheLineTemp[153], cacheLineTemp[145]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_1 = {cacheLineTemp[169], cacheLineTemp[161]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_1 = {cacheLineTemp[185], cacheLineTemp[177]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_1 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_1, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_1, memRequest_bits_data_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_1 = {cacheLineTemp[201], cacheLineTemp[193]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_1 = {cacheLineTemp[217], cacheLineTemp[209]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_1, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_1 = {cacheLineTemp[233], cacheLineTemp[225]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_1 = {cacheLineTemp[249], cacheLineTemp[241]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_1 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_1, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi_1 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_1, memRequest_bits_data_lo_lo_lo_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_lo_hi_lo_1};
  wire [31:0]       memRequest_bits_data_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_1 = {cacheLineTemp[265], cacheLineTemp[257]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_1 = {cacheLineTemp[281], cacheLineTemp[273]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_1, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_1 = {cacheLineTemp[297], cacheLineTemp[289]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_1 = {cacheLineTemp[313], cacheLineTemp[305]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_1, memRequest_bits_data_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_1 = {cacheLineTemp[329], cacheLineTemp[321]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_1 = {cacheLineTemp[345], cacheLineTemp[337]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_1 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_1, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_1 = {cacheLineTemp[361], cacheLineTemp[353]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_1 = {cacheLineTemp[377], cacheLineTemp[369]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_1 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_1 = {memRequest_bits_data_lo_lo_hi_lo_hi_1, memRequest_bits_data_lo_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_1 = {cacheLineTemp[393], cacheLineTemp[385]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_1 = {cacheLineTemp[409], cacheLineTemp[401]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_1, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_1 = {cacheLineTemp[425], cacheLineTemp[417]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_1 = {cacheLineTemp[441], cacheLineTemp[433]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo_1 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_1, memRequest_bits_data_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_1 = {cacheLineTemp[457], cacheLineTemp[449]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_1 = {cacheLineTemp[473], cacheLineTemp[465]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_1 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_1, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_1 = {cacheLineTemp[489], cacheLineTemp[481]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_1 = {cacheLineTemp[505], cacheLineTemp[497]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_1, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_1, memRequest_bits_data_lo_lo_hi_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_hi_1, memRequest_bits_data_lo_lo_hi_hi_lo_1};
  wire [31:0]       memRequest_bits_data_lo_lo_hi_1 = {memRequest_bits_data_lo_lo_hi_hi_1, memRequest_bits_data_lo_lo_hi_lo_1};
  wire [63:0]       memRequest_bits_data_lo_lo_1 = {memRequest_bits_data_lo_lo_hi_1, memRequest_bits_data_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_1 = {cacheLineTemp[521], cacheLineTemp[513]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_1 = {cacheLineTemp[537], cacheLineTemp[529]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_1 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_1 = {cacheLineTemp[553], cacheLineTemp[545]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_1 = {cacheLineTemp[569], cacheLineTemp[561]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_1 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo_1 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_1 = {cacheLineTemp[585], cacheLineTemp[577]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_1 = {cacheLineTemp[601], cacheLineTemp[593]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_1 = {cacheLineTemp[617], cacheLineTemp[609]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_1 = {cacheLineTemp[633], cacheLineTemp[625]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi_1 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_1 = {memRequest_bits_data_lo_hi_lo_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_1 = {cacheLineTemp[649], cacheLineTemp[641]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_1 = {cacheLineTemp[665], cacheLineTemp[657]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_1, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_1 = {cacheLineTemp[681], cacheLineTemp[673]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_1 = {cacheLineTemp[697], cacheLineTemp[689]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_1 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_1 = {cacheLineTemp[713], cacheLineTemp[705]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_1 = {cacheLineTemp[729], cacheLineTemp[721]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_1 = {cacheLineTemp[745], cacheLineTemp[737]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_1 = {cacheLineTemp[761], cacheLineTemp[753]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_1 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_1, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_lo_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_1 = {memRequest_bits_data_lo_hi_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_hi_lo_1};
  wire [31:0]       memRequest_bits_data_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_1 = {cacheLineTemp[777], cacheLineTemp[769]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_1 = {cacheLineTemp[793], cacheLineTemp[785]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_1 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_1, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_1 = {cacheLineTemp[809], cacheLineTemp[801]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_1 = {cacheLineTemp[825], cacheLineTemp[817]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo_1 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_1, memRequest_bits_data_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_1 = {cacheLineTemp[841], cacheLineTemp[833]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_1 = {cacheLineTemp[857], cacheLineTemp[849]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_1 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_1, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_1 = {cacheLineTemp[873], cacheLineTemp[865]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_1 = {cacheLineTemp[889], cacheLineTemp[881]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_1 = {memRequest_bits_data_lo_hi_hi_lo_hi_1, memRequest_bits_data_lo_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_1 = {cacheLineTemp[905], cacheLineTemp[897]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_1 = {cacheLineTemp[921], cacheLineTemp[913]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_1 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_1, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_1 = {cacheLineTemp[937], cacheLineTemp[929]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_1 = {cacheLineTemp[953], cacheLineTemp[945]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_1, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo_1 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_1, memRequest_bits_data_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_1 = {cacheLineTemp[969], cacheLineTemp[961]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_1 = {cacheLineTemp[985], cacheLineTemp[977]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_1 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_1, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_1 = {cacheLineTemp[1001], cacheLineTemp[993]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_1 = {cacheLineTemp[1017], cacheLineTemp[1009]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_hi_lo_1};
  wire [31:0]       memRequest_bits_data_lo_hi_hi_1 = {memRequest_bits_data_lo_hi_hi_hi_1, memRequest_bits_data_lo_hi_hi_lo_1};
  wire [63:0]       memRequest_bits_data_lo_hi_1 = {memRequest_bits_data_lo_hi_hi_1, memRequest_bits_data_lo_hi_lo_1};
  wire [127:0]      memRequest_bits_data_lo_1 = {memRequest_bits_data_lo_hi_1, memRequest_bits_data_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_1 = {dataBuffer_0[9], dataBuffer_0[1]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_1 = {dataBuffer_0[25], dataBuffer_0[17]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_1 = {dataBuffer_0[41], dataBuffer_0[33]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_1 = {dataBuffer_0[57], dataBuffer_0[49]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_1 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_1, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_1 = {dataBuffer_0[73], dataBuffer_0[65]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_1 = {dataBuffer_0[89], dataBuffer_0[81]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_1 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_1 = {dataBuffer_0[105], dataBuffer_0[97]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_1 = {dataBuffer_0[121], dataBuffer_0[113]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_1 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_1, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi_1 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_1, memRequest_bits_data_hi_lo_lo_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_1 = {dataBuffer_0[137], dataBuffer_0[129]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_1 = {dataBuffer_0[153], dataBuffer_0[145]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_1 = {dataBuffer_0[169], dataBuffer_0[161]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_1 = {dataBuffer_0[185], dataBuffer_0[177]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_1 = {dataBuffer_0[201], dataBuffer_0[193]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_1 = {dataBuffer_0[217], dataBuffer_0[209]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_1 = {dataBuffer_0[233], dataBuffer_0[225]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_1 = {dataBuffer_0[249], dataBuffer_0[241]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_1 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_1, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi_1 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_1, memRequest_bits_data_hi_lo_lo_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_1 = {memRequest_bits_data_hi_lo_lo_hi_hi_1, memRequest_bits_data_hi_lo_lo_hi_lo_1};
  wire [31:0]       memRequest_bits_data_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_1 = {dataBuffer_0[265], dataBuffer_0[257]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_1 = {dataBuffer_0[281], dataBuffer_0[273]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_1 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_1, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_1 = {dataBuffer_0[297], dataBuffer_0[289]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_1 = {dataBuffer_0[313], dataBuffer_0[305]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_1 = {dataBuffer_0[329], dataBuffer_0[321]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_1 = {dataBuffer_0[345], dataBuffer_0[337]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_1, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_1 = {dataBuffer_0[361], dataBuffer_0[353]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_1 = {dataBuffer_0[377], dataBuffer_0[369]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_1 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_lo_hi_1, memRequest_bits_data_hi_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_1 = {dataBuffer_0[393], dataBuffer_0[385]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_1 = {dataBuffer_0[409], dataBuffer_0[401]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_1 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_1, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_1 = {dataBuffer_0[425], dataBuffer_0[417]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_1 = {dataBuffer_0[441], dataBuffer_0[433]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_1, memRequest_bits_data_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_1 = {dataBuffer_0[457], dataBuffer_0[449]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_1 = {dataBuffer_0[473], dataBuffer_0[465]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_1, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_1 = {dataBuffer_0[489], dataBuffer_0[481]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_1 = {dataBuffer_0[505], dataBuffer_0[497]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_1, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_1, memRequest_bits_data_hi_lo_hi_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_hi_1, memRequest_bits_data_hi_lo_hi_hi_lo_1};
  wire [31:0]       memRequest_bits_data_hi_lo_hi_1 = {memRequest_bits_data_hi_lo_hi_hi_1, memRequest_bits_data_hi_lo_hi_lo_1};
  wire [63:0]       memRequest_bits_data_hi_lo_1 = {memRequest_bits_data_hi_lo_hi_1, memRequest_bits_data_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_1 = {dataBuffer_0[521], dataBuffer_0[513]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_1 = {dataBuffer_0[537], dataBuffer_0[529]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_1 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_1 = {dataBuffer_0[553], dataBuffer_0[545]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_1 = {dataBuffer_0[569], dataBuffer_0[561]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_1 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_1, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo_1 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_1 = {dataBuffer_0[585], dataBuffer_0[577]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_1 = {dataBuffer_0[601], dataBuffer_0[593]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_1 = {dataBuffer_0[617], dataBuffer_0[609]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_1 = {dataBuffer_0[633], dataBuffer_0[625]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_1 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi_1 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_1, memRequest_bits_data_hi_hi_lo_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_1 = {memRequest_bits_data_hi_hi_lo_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_1 = {dataBuffer_0[649], dataBuffer_0[641]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_1 = {dataBuffer_0[665], dataBuffer_0[657]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_1, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_1 = {dataBuffer_0[681], dataBuffer_0[673]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_1 = {dataBuffer_0[697], dataBuffer_0[689]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_1 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_1, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_1 = {dataBuffer_0[713], dataBuffer_0[705]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_1 = {dataBuffer_0[729], dataBuffer_0[721]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_1 = {dataBuffer_0[745], dataBuffer_0[737]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_1 = {dataBuffer_0[761], dataBuffer_0[753]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi_1 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_1 = {memRequest_bits_data_hi_hi_lo_hi_hi_1, memRequest_bits_data_hi_hi_lo_hi_lo_1};
  wire [31:0]       memRequest_bits_data_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_1 = {dataBuffer_0[777], dataBuffer_0[769]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_1 = {dataBuffer_0[793], dataBuffer_0[785]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_1 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_1, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_1 = {dataBuffer_0[809], dataBuffer_0[801]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_1 = {dataBuffer_0[825], dataBuffer_0[817]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_1 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo_1 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_1, memRequest_bits_data_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_1 = {dataBuffer_0[841], dataBuffer_0[833]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_1 = {dataBuffer_0[857], dataBuffer_0[849]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_1 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_1, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_1 = {dataBuffer_0[873], dataBuffer_0[865]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_1 = {dataBuffer_0[889], dataBuffer_0[881]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi_1 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_1 = {dataBuffer_0[905], dataBuffer_0[897]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_1 = {dataBuffer_0[921], dataBuffer_0[913]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_1 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_1, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_1 = {dataBuffer_0[937], dataBuffer_0[929]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_1 = {dataBuffer_0[953], dataBuffer_0[945]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_1, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_1 = {dataBuffer_0[969], dataBuffer_0[961]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_1 = {dataBuffer_0[985], dataBuffer_0[977]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_1 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_1, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_1};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_1 = {dataBuffer_0[1001], dataBuffer_0[993]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_1 = {dataBuffer_0[1017], dataBuffer_0[1009]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_1};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_hi_hi_lo_1};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_hi_lo_1};
  wire [31:0]       memRequest_bits_data_hi_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_hi_1, memRequest_bits_data_hi_hi_hi_lo_1};
  wire [63:0]       memRequest_bits_data_hi_hi_1 = {memRequest_bits_data_hi_hi_hi_1, memRequest_bits_data_hi_hi_lo_1};
  wire [127:0]      memRequest_bits_data_hi_1 = {memRequest_bits_data_hi_hi_1, memRequest_bits_data_hi_lo_1};
  wire [382:0]      _memRequest_bits_data_T_2435 = {127'h0, memRequest_bits_data_hi_1, memRequest_bits_data_lo_1} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_2 = {cacheLineTemp[10], cacheLineTemp[2]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_2 = {cacheLineTemp[26], cacheLineTemp[18]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_2 = {cacheLineTemp[42], cacheLineTemp[34]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_2 = {cacheLineTemp[58], cacheLineTemp[50]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_2 = {cacheLineTemp[74], cacheLineTemp[66]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_2 = {cacheLineTemp[90], cacheLineTemp[82]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_2 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_2 = {cacheLineTemp[106], cacheLineTemp[98]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_2 = {cacheLineTemp[122], cacheLineTemp[114]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_2 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_2, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_lo_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_2 = {cacheLineTemp[138], cacheLineTemp[130]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_2 = {cacheLineTemp[154], cacheLineTemp[146]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_2 = {cacheLineTemp[170], cacheLineTemp[162]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_2 = {cacheLineTemp[186], cacheLineTemp[178]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_2 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_2, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_2, memRequest_bits_data_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_2 = {cacheLineTemp[202], cacheLineTemp[194]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_2 = {cacheLineTemp[218], cacheLineTemp[210]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_2, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_2 = {cacheLineTemp[234], cacheLineTemp[226]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_2 = {cacheLineTemp[250], cacheLineTemp[242]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_2 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_2, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi_2 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_2, memRequest_bits_data_lo_lo_lo_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_lo_hi_lo_2};
  wire [31:0]       memRequest_bits_data_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_2 = {cacheLineTemp[266], cacheLineTemp[258]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_2 = {cacheLineTemp[282], cacheLineTemp[274]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_2, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_2 = {cacheLineTemp[298], cacheLineTemp[290]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_2 = {cacheLineTemp[314], cacheLineTemp[306]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_2, memRequest_bits_data_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_2 = {cacheLineTemp[330], cacheLineTemp[322]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_2 = {cacheLineTemp[346], cacheLineTemp[338]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_2 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_2, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_2 = {cacheLineTemp[362], cacheLineTemp[354]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_2 = {cacheLineTemp[378], cacheLineTemp[370]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_2 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_2 = {memRequest_bits_data_lo_lo_hi_lo_hi_2, memRequest_bits_data_lo_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_2 = {cacheLineTemp[394], cacheLineTemp[386]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_2 = {cacheLineTemp[410], cacheLineTemp[402]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_2, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_2 = {cacheLineTemp[426], cacheLineTemp[418]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_2 = {cacheLineTemp[442], cacheLineTemp[434]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo_2 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_2, memRequest_bits_data_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_2 = {cacheLineTemp[458], cacheLineTemp[450]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_2 = {cacheLineTemp[474], cacheLineTemp[466]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_2 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_2, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_2 = {cacheLineTemp[490], cacheLineTemp[482]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_2 = {cacheLineTemp[506], cacheLineTemp[498]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_2, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_2, memRequest_bits_data_lo_lo_hi_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_hi_2, memRequest_bits_data_lo_lo_hi_hi_lo_2};
  wire [31:0]       memRequest_bits_data_lo_lo_hi_2 = {memRequest_bits_data_lo_lo_hi_hi_2, memRequest_bits_data_lo_lo_hi_lo_2};
  wire [63:0]       memRequest_bits_data_lo_lo_2 = {memRequest_bits_data_lo_lo_hi_2, memRequest_bits_data_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_2 = {cacheLineTemp[522], cacheLineTemp[514]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_2 = {cacheLineTemp[538], cacheLineTemp[530]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_2 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_2 = {cacheLineTemp[554], cacheLineTemp[546]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_2 = {cacheLineTemp[570], cacheLineTemp[562]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_2 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo_2 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_2 = {cacheLineTemp[586], cacheLineTemp[578]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_2 = {cacheLineTemp[602], cacheLineTemp[594]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_2 = {cacheLineTemp[618], cacheLineTemp[610]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_2 = {cacheLineTemp[634], cacheLineTemp[626]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi_2 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_2 = {memRequest_bits_data_lo_hi_lo_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_2 = {cacheLineTemp[650], cacheLineTemp[642]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_2 = {cacheLineTemp[666], cacheLineTemp[658]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_2, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_2 = {cacheLineTemp[682], cacheLineTemp[674]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_2 = {cacheLineTemp[698], cacheLineTemp[690]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_2 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_2 = {cacheLineTemp[714], cacheLineTemp[706]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_2 = {cacheLineTemp[730], cacheLineTemp[722]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_2 = {cacheLineTemp[746], cacheLineTemp[738]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_2 = {cacheLineTemp[762], cacheLineTemp[754]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_2 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_2, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_lo_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_2 = {memRequest_bits_data_lo_hi_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_hi_lo_2};
  wire [31:0]       memRequest_bits_data_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_2 = {cacheLineTemp[778], cacheLineTemp[770]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_2 = {cacheLineTemp[794], cacheLineTemp[786]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_2 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_2, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_2 = {cacheLineTemp[810], cacheLineTemp[802]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_2 = {cacheLineTemp[826], cacheLineTemp[818]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo_2 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_2, memRequest_bits_data_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_2 = {cacheLineTemp[842], cacheLineTemp[834]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_2 = {cacheLineTemp[858], cacheLineTemp[850]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_2 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_2, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_2 = {cacheLineTemp[874], cacheLineTemp[866]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_2 = {cacheLineTemp[890], cacheLineTemp[882]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_2 = {memRequest_bits_data_lo_hi_hi_lo_hi_2, memRequest_bits_data_lo_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_2 = {cacheLineTemp[906], cacheLineTemp[898]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_2 = {cacheLineTemp[922], cacheLineTemp[914]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_2 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_2, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_2 = {cacheLineTemp[938], cacheLineTemp[930]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_2 = {cacheLineTemp[954], cacheLineTemp[946]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_2, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo_2 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_2, memRequest_bits_data_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_2 = {cacheLineTemp[970], cacheLineTemp[962]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_2 = {cacheLineTemp[986], cacheLineTemp[978]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_2 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_2, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_2 = {cacheLineTemp[1002], cacheLineTemp[994]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_2 = {cacheLineTemp[1018], cacheLineTemp[1010]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_hi_lo_2};
  wire [31:0]       memRequest_bits_data_lo_hi_hi_2 = {memRequest_bits_data_lo_hi_hi_hi_2, memRequest_bits_data_lo_hi_hi_lo_2};
  wire [63:0]       memRequest_bits_data_lo_hi_2 = {memRequest_bits_data_lo_hi_hi_2, memRequest_bits_data_lo_hi_lo_2};
  wire [127:0]      memRequest_bits_data_lo_2 = {memRequest_bits_data_lo_hi_2, memRequest_bits_data_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_2 = {dataBuffer_0[10], dataBuffer_0[2]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_2 = {dataBuffer_0[26], dataBuffer_0[18]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_2 = {dataBuffer_0[42], dataBuffer_0[34]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_2 = {dataBuffer_0[58], dataBuffer_0[50]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_2 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_2, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_2 = {dataBuffer_0[74], dataBuffer_0[66]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_2 = {dataBuffer_0[90], dataBuffer_0[82]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_2 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_2 = {dataBuffer_0[106], dataBuffer_0[98]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_2 = {dataBuffer_0[122], dataBuffer_0[114]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_2 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_2, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi_2 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_2, memRequest_bits_data_hi_lo_lo_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_2 = {dataBuffer_0[138], dataBuffer_0[130]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_2 = {dataBuffer_0[154], dataBuffer_0[146]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_2 = {dataBuffer_0[170], dataBuffer_0[162]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_2 = {dataBuffer_0[186], dataBuffer_0[178]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_2 = {dataBuffer_0[202], dataBuffer_0[194]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_2 = {dataBuffer_0[218], dataBuffer_0[210]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_2 = {dataBuffer_0[234], dataBuffer_0[226]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_2 = {dataBuffer_0[250], dataBuffer_0[242]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_2 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_2, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi_2 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_2, memRequest_bits_data_hi_lo_lo_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_2 = {memRequest_bits_data_hi_lo_lo_hi_hi_2, memRequest_bits_data_hi_lo_lo_hi_lo_2};
  wire [31:0]       memRequest_bits_data_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_2 = {dataBuffer_0[266], dataBuffer_0[258]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_2 = {dataBuffer_0[282], dataBuffer_0[274]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_2 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_2, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_2 = {dataBuffer_0[298], dataBuffer_0[290]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_2 = {dataBuffer_0[314], dataBuffer_0[306]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_2 = {dataBuffer_0[330], dataBuffer_0[322]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_2 = {dataBuffer_0[346], dataBuffer_0[338]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_2, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_2 = {dataBuffer_0[362], dataBuffer_0[354]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_2 = {dataBuffer_0[378], dataBuffer_0[370]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_2 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_lo_hi_2, memRequest_bits_data_hi_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_2 = {dataBuffer_0[394], dataBuffer_0[386]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_2 = {dataBuffer_0[410], dataBuffer_0[402]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_2 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_2, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_2 = {dataBuffer_0[426], dataBuffer_0[418]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_2 = {dataBuffer_0[442], dataBuffer_0[434]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_2, memRequest_bits_data_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_2 = {dataBuffer_0[458], dataBuffer_0[450]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_2 = {dataBuffer_0[474], dataBuffer_0[466]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_2, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_2 = {dataBuffer_0[490], dataBuffer_0[482]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_2 = {dataBuffer_0[506], dataBuffer_0[498]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_2, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_2, memRequest_bits_data_hi_lo_hi_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_hi_2, memRequest_bits_data_hi_lo_hi_hi_lo_2};
  wire [31:0]       memRequest_bits_data_hi_lo_hi_2 = {memRequest_bits_data_hi_lo_hi_hi_2, memRequest_bits_data_hi_lo_hi_lo_2};
  wire [63:0]       memRequest_bits_data_hi_lo_2 = {memRequest_bits_data_hi_lo_hi_2, memRequest_bits_data_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_2 = {dataBuffer_0[522], dataBuffer_0[514]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_2 = {dataBuffer_0[538], dataBuffer_0[530]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_2 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_2 = {dataBuffer_0[554], dataBuffer_0[546]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_2 = {dataBuffer_0[570], dataBuffer_0[562]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_2 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_2, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo_2 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_2 = {dataBuffer_0[586], dataBuffer_0[578]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_2 = {dataBuffer_0[602], dataBuffer_0[594]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_2 = {dataBuffer_0[618], dataBuffer_0[610]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_2 = {dataBuffer_0[634], dataBuffer_0[626]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_2 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi_2 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_2, memRequest_bits_data_hi_hi_lo_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_2 = {memRequest_bits_data_hi_hi_lo_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_2 = {dataBuffer_0[650], dataBuffer_0[642]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_2 = {dataBuffer_0[666], dataBuffer_0[658]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_2, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_2 = {dataBuffer_0[682], dataBuffer_0[674]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_2 = {dataBuffer_0[698], dataBuffer_0[690]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_2 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_2, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_2 = {dataBuffer_0[714], dataBuffer_0[706]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_2 = {dataBuffer_0[730], dataBuffer_0[722]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_2 = {dataBuffer_0[746], dataBuffer_0[738]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_2 = {dataBuffer_0[762], dataBuffer_0[754]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi_2 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_2 = {memRequest_bits_data_hi_hi_lo_hi_hi_2, memRequest_bits_data_hi_hi_lo_hi_lo_2};
  wire [31:0]       memRequest_bits_data_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_2 = {dataBuffer_0[778], dataBuffer_0[770]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_2 = {dataBuffer_0[794], dataBuffer_0[786]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_2 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_2, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_2 = {dataBuffer_0[810], dataBuffer_0[802]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_2 = {dataBuffer_0[826], dataBuffer_0[818]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_2 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo_2 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_2, memRequest_bits_data_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_2 = {dataBuffer_0[842], dataBuffer_0[834]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_2 = {dataBuffer_0[858], dataBuffer_0[850]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_2 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_2, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_2 = {dataBuffer_0[874], dataBuffer_0[866]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_2 = {dataBuffer_0[890], dataBuffer_0[882]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi_2 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_2 = {dataBuffer_0[906], dataBuffer_0[898]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_2 = {dataBuffer_0[922], dataBuffer_0[914]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_2 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_2, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_2 = {dataBuffer_0[938], dataBuffer_0[930]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_2 = {dataBuffer_0[954], dataBuffer_0[946]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_2, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_2 = {dataBuffer_0[970], dataBuffer_0[962]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_2 = {dataBuffer_0[986], dataBuffer_0[978]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_2 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_2, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_2};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_2 = {dataBuffer_0[1002], dataBuffer_0[994]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_2 = {dataBuffer_0[1018], dataBuffer_0[1010]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_2};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_hi_hi_lo_2};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_hi_lo_2};
  wire [31:0]       memRequest_bits_data_hi_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_hi_2, memRequest_bits_data_hi_hi_hi_lo_2};
  wire [63:0]       memRequest_bits_data_hi_hi_2 = {memRequest_bits_data_hi_hi_hi_2, memRequest_bits_data_hi_hi_lo_2};
  wire [127:0]      memRequest_bits_data_hi_2 = {memRequest_bits_data_hi_hi_2, memRequest_bits_data_hi_lo_2};
  wire [382:0]      _memRequest_bits_data_T_2820 = {127'h0, memRequest_bits_data_hi_2, memRequest_bits_data_lo_2} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_3 = {cacheLineTemp[11], cacheLineTemp[3]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_3 = {cacheLineTemp[27], cacheLineTemp[19]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_3 = {cacheLineTemp[43], cacheLineTemp[35]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_3 = {cacheLineTemp[59], cacheLineTemp[51]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_3 = {cacheLineTemp[75], cacheLineTemp[67]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_3 = {cacheLineTemp[91], cacheLineTemp[83]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_3 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_3 = {cacheLineTemp[107], cacheLineTemp[99]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_3 = {cacheLineTemp[123], cacheLineTemp[115]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_3 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_3, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_lo_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_3 = {cacheLineTemp[139], cacheLineTemp[131]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_3 = {cacheLineTemp[155], cacheLineTemp[147]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_3 = {cacheLineTemp[171], cacheLineTemp[163]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_3 = {cacheLineTemp[187], cacheLineTemp[179]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_3 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_3, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_3, memRequest_bits_data_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_3 = {cacheLineTemp[203], cacheLineTemp[195]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_3 = {cacheLineTemp[219], cacheLineTemp[211]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_3, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_3 = {cacheLineTemp[235], cacheLineTemp[227]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_3 = {cacheLineTemp[251], cacheLineTemp[243]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_3 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_3, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi_3 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_3, memRequest_bits_data_lo_lo_lo_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_lo_hi_lo_3};
  wire [31:0]       memRequest_bits_data_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_3 = {cacheLineTemp[267], cacheLineTemp[259]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_3 = {cacheLineTemp[283], cacheLineTemp[275]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_3, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_3 = {cacheLineTemp[299], cacheLineTemp[291]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_3 = {cacheLineTemp[315], cacheLineTemp[307]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_3, memRequest_bits_data_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_3 = {cacheLineTemp[331], cacheLineTemp[323]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_3 = {cacheLineTemp[347], cacheLineTemp[339]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_3 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_3, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_3 = {cacheLineTemp[363], cacheLineTemp[355]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_3 = {cacheLineTemp[379], cacheLineTemp[371]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_3 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_3 = {memRequest_bits_data_lo_lo_hi_lo_hi_3, memRequest_bits_data_lo_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_3 = {cacheLineTemp[395], cacheLineTemp[387]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_3 = {cacheLineTemp[411], cacheLineTemp[403]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_3, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_3 = {cacheLineTemp[427], cacheLineTemp[419]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_3 = {cacheLineTemp[443], cacheLineTemp[435]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo_3 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_3, memRequest_bits_data_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_3 = {cacheLineTemp[459], cacheLineTemp[451]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_3 = {cacheLineTemp[475], cacheLineTemp[467]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_3 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_3, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_3 = {cacheLineTemp[491], cacheLineTemp[483]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_3 = {cacheLineTemp[507], cacheLineTemp[499]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_3, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_3, memRequest_bits_data_lo_lo_hi_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_hi_3, memRequest_bits_data_lo_lo_hi_hi_lo_3};
  wire [31:0]       memRequest_bits_data_lo_lo_hi_3 = {memRequest_bits_data_lo_lo_hi_hi_3, memRequest_bits_data_lo_lo_hi_lo_3};
  wire [63:0]       memRequest_bits_data_lo_lo_3 = {memRequest_bits_data_lo_lo_hi_3, memRequest_bits_data_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_3 = {cacheLineTemp[523], cacheLineTemp[515]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_3 = {cacheLineTemp[539], cacheLineTemp[531]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_3 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_3 = {cacheLineTemp[555], cacheLineTemp[547]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_3 = {cacheLineTemp[571], cacheLineTemp[563]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_3 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo_3 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_3 = {cacheLineTemp[587], cacheLineTemp[579]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_3 = {cacheLineTemp[603], cacheLineTemp[595]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_3 = {cacheLineTemp[619], cacheLineTemp[611]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_3 = {cacheLineTemp[635], cacheLineTemp[627]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi_3 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_3 = {memRequest_bits_data_lo_hi_lo_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_3 = {cacheLineTemp[651], cacheLineTemp[643]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_3 = {cacheLineTemp[667], cacheLineTemp[659]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_3, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_3 = {cacheLineTemp[683], cacheLineTemp[675]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_3 = {cacheLineTemp[699], cacheLineTemp[691]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_3 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_3 = {cacheLineTemp[715], cacheLineTemp[707]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_3 = {cacheLineTemp[731], cacheLineTemp[723]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_3 = {cacheLineTemp[747], cacheLineTemp[739]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_3 = {cacheLineTemp[763], cacheLineTemp[755]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_3 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_3, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_lo_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_3 = {memRequest_bits_data_lo_hi_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_hi_lo_3};
  wire [31:0]       memRequest_bits_data_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_3 = {cacheLineTemp[779], cacheLineTemp[771]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_3 = {cacheLineTemp[795], cacheLineTemp[787]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_3 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_3, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_3 = {cacheLineTemp[811], cacheLineTemp[803]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_3 = {cacheLineTemp[827], cacheLineTemp[819]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo_3 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_3, memRequest_bits_data_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_3 = {cacheLineTemp[843], cacheLineTemp[835]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_3 = {cacheLineTemp[859], cacheLineTemp[851]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_3 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_3, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_3 = {cacheLineTemp[875], cacheLineTemp[867]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_3 = {cacheLineTemp[891], cacheLineTemp[883]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_3 = {memRequest_bits_data_lo_hi_hi_lo_hi_3, memRequest_bits_data_lo_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_3 = {cacheLineTemp[907], cacheLineTemp[899]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_3 = {cacheLineTemp[923], cacheLineTemp[915]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_3 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_3, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_3 = {cacheLineTemp[939], cacheLineTemp[931]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_3 = {cacheLineTemp[955], cacheLineTemp[947]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_3, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo_3 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_3, memRequest_bits_data_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_3 = {cacheLineTemp[971], cacheLineTemp[963]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_3 = {cacheLineTemp[987], cacheLineTemp[979]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_3 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_3, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_3 = {cacheLineTemp[1003], cacheLineTemp[995]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_3 = {cacheLineTemp[1019], cacheLineTemp[1011]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_hi_lo_3};
  wire [31:0]       memRequest_bits_data_lo_hi_hi_3 = {memRequest_bits_data_lo_hi_hi_hi_3, memRequest_bits_data_lo_hi_hi_lo_3};
  wire [63:0]       memRequest_bits_data_lo_hi_3 = {memRequest_bits_data_lo_hi_hi_3, memRequest_bits_data_lo_hi_lo_3};
  wire [127:0]      memRequest_bits_data_lo_3 = {memRequest_bits_data_lo_hi_3, memRequest_bits_data_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_3 = {dataBuffer_0[11], dataBuffer_0[3]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_3 = {dataBuffer_0[27], dataBuffer_0[19]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_3 = {dataBuffer_0[43], dataBuffer_0[35]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_3 = {dataBuffer_0[59], dataBuffer_0[51]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_3 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_3, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_3 = {dataBuffer_0[75], dataBuffer_0[67]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_3 = {dataBuffer_0[91], dataBuffer_0[83]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_3 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_3 = {dataBuffer_0[107], dataBuffer_0[99]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_3 = {dataBuffer_0[123], dataBuffer_0[115]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_3 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_3, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi_3 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_3, memRequest_bits_data_hi_lo_lo_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_3 = {dataBuffer_0[139], dataBuffer_0[131]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_3 = {dataBuffer_0[155], dataBuffer_0[147]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_3 = {dataBuffer_0[171], dataBuffer_0[163]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_3 = {dataBuffer_0[187], dataBuffer_0[179]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_3 = {dataBuffer_0[203], dataBuffer_0[195]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_3 = {dataBuffer_0[219], dataBuffer_0[211]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_3 = {dataBuffer_0[235], dataBuffer_0[227]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_3 = {dataBuffer_0[251], dataBuffer_0[243]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_3 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_3, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi_3 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_3, memRequest_bits_data_hi_lo_lo_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_3 = {memRequest_bits_data_hi_lo_lo_hi_hi_3, memRequest_bits_data_hi_lo_lo_hi_lo_3};
  wire [31:0]       memRequest_bits_data_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_3 = {dataBuffer_0[267], dataBuffer_0[259]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_3 = {dataBuffer_0[283], dataBuffer_0[275]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_3 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_3, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_3 = {dataBuffer_0[299], dataBuffer_0[291]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_3 = {dataBuffer_0[315], dataBuffer_0[307]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_3 = {dataBuffer_0[331], dataBuffer_0[323]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_3 = {dataBuffer_0[347], dataBuffer_0[339]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_3, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_3 = {dataBuffer_0[363], dataBuffer_0[355]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_3 = {dataBuffer_0[379], dataBuffer_0[371]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_3 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_lo_hi_3, memRequest_bits_data_hi_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_3 = {dataBuffer_0[395], dataBuffer_0[387]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_3 = {dataBuffer_0[411], dataBuffer_0[403]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_3 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_3, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_3 = {dataBuffer_0[427], dataBuffer_0[419]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_3 = {dataBuffer_0[443], dataBuffer_0[435]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_3, memRequest_bits_data_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_3 = {dataBuffer_0[459], dataBuffer_0[451]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_3 = {dataBuffer_0[475], dataBuffer_0[467]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_3, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_3 = {dataBuffer_0[491], dataBuffer_0[483]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_3 = {dataBuffer_0[507], dataBuffer_0[499]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_3, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_3, memRequest_bits_data_hi_lo_hi_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_hi_3, memRequest_bits_data_hi_lo_hi_hi_lo_3};
  wire [31:0]       memRequest_bits_data_hi_lo_hi_3 = {memRequest_bits_data_hi_lo_hi_hi_3, memRequest_bits_data_hi_lo_hi_lo_3};
  wire [63:0]       memRequest_bits_data_hi_lo_3 = {memRequest_bits_data_hi_lo_hi_3, memRequest_bits_data_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_3 = {dataBuffer_0[523], dataBuffer_0[515]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_3 = {dataBuffer_0[539], dataBuffer_0[531]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_3 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_3 = {dataBuffer_0[555], dataBuffer_0[547]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_3 = {dataBuffer_0[571], dataBuffer_0[563]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_3 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_3, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo_3 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_3 = {dataBuffer_0[587], dataBuffer_0[579]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_3 = {dataBuffer_0[603], dataBuffer_0[595]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_3 = {dataBuffer_0[619], dataBuffer_0[611]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_3 = {dataBuffer_0[635], dataBuffer_0[627]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_3 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi_3 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_3, memRequest_bits_data_hi_hi_lo_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_3 = {memRequest_bits_data_hi_hi_lo_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_3 = {dataBuffer_0[651], dataBuffer_0[643]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_3 = {dataBuffer_0[667], dataBuffer_0[659]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_3, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_3 = {dataBuffer_0[683], dataBuffer_0[675]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_3 = {dataBuffer_0[699], dataBuffer_0[691]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_3 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_3, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_3 = {dataBuffer_0[715], dataBuffer_0[707]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_3 = {dataBuffer_0[731], dataBuffer_0[723]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_3 = {dataBuffer_0[747], dataBuffer_0[739]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_3 = {dataBuffer_0[763], dataBuffer_0[755]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi_3 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_3 = {memRequest_bits_data_hi_hi_lo_hi_hi_3, memRequest_bits_data_hi_hi_lo_hi_lo_3};
  wire [31:0]       memRequest_bits_data_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_3 = {dataBuffer_0[779], dataBuffer_0[771]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_3 = {dataBuffer_0[795], dataBuffer_0[787]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_3 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_3, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_3 = {dataBuffer_0[811], dataBuffer_0[803]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_3 = {dataBuffer_0[827], dataBuffer_0[819]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_3 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo_3 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_3, memRequest_bits_data_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_3 = {dataBuffer_0[843], dataBuffer_0[835]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_3 = {dataBuffer_0[859], dataBuffer_0[851]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_3 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_3, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_3 = {dataBuffer_0[875], dataBuffer_0[867]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_3 = {dataBuffer_0[891], dataBuffer_0[883]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi_3 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_3 = {dataBuffer_0[907], dataBuffer_0[899]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_3 = {dataBuffer_0[923], dataBuffer_0[915]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_3 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_3, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_3 = {dataBuffer_0[939], dataBuffer_0[931]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_3 = {dataBuffer_0[955], dataBuffer_0[947]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_3, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_3 = {dataBuffer_0[971], dataBuffer_0[963]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_3 = {dataBuffer_0[987], dataBuffer_0[979]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_3 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_3, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_3};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_3 = {dataBuffer_0[1003], dataBuffer_0[995]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_3 = {dataBuffer_0[1019], dataBuffer_0[1011]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_3};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_hi_hi_lo_3};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_hi_lo_3};
  wire [31:0]       memRequest_bits_data_hi_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_hi_3, memRequest_bits_data_hi_hi_hi_lo_3};
  wire [63:0]       memRequest_bits_data_hi_hi_3 = {memRequest_bits_data_hi_hi_hi_3, memRequest_bits_data_hi_hi_lo_3};
  wire [127:0]      memRequest_bits_data_hi_3 = {memRequest_bits_data_hi_hi_3, memRequest_bits_data_hi_lo_3};
  wire [382:0]      _memRequest_bits_data_T_3205 = {127'h0, memRequest_bits_data_hi_3, memRequest_bits_data_lo_3} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_4 = {cacheLineTemp[12], cacheLineTemp[4]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_4 = {cacheLineTemp[28], cacheLineTemp[20]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_4 = {cacheLineTemp[44], cacheLineTemp[36]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_4 = {cacheLineTemp[60], cacheLineTemp[52]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_4 = {cacheLineTemp[76], cacheLineTemp[68]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_4 = {cacheLineTemp[92], cacheLineTemp[84]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_4 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_4 = {cacheLineTemp[108], cacheLineTemp[100]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_4 = {cacheLineTemp[124], cacheLineTemp[116]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_4 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_4, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_lo_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_4 = {cacheLineTemp[140], cacheLineTemp[132]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_4 = {cacheLineTemp[156], cacheLineTemp[148]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_4 = {cacheLineTemp[172], cacheLineTemp[164]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_4 = {cacheLineTemp[188], cacheLineTemp[180]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_4 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_4, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_4, memRequest_bits_data_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_4 = {cacheLineTemp[204], cacheLineTemp[196]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_4 = {cacheLineTemp[220], cacheLineTemp[212]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_4, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_4 = {cacheLineTemp[236], cacheLineTemp[228]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_4 = {cacheLineTemp[252], cacheLineTemp[244]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_4 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_4, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi_4 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_4, memRequest_bits_data_lo_lo_lo_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_lo_hi_lo_4};
  wire [31:0]       memRequest_bits_data_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_4 = {cacheLineTemp[268], cacheLineTemp[260]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_4 = {cacheLineTemp[284], cacheLineTemp[276]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_4, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_4 = {cacheLineTemp[300], cacheLineTemp[292]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_4 = {cacheLineTemp[316], cacheLineTemp[308]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_4, memRequest_bits_data_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_4 = {cacheLineTemp[332], cacheLineTemp[324]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_4 = {cacheLineTemp[348], cacheLineTemp[340]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_4 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_4, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_4 = {cacheLineTemp[364], cacheLineTemp[356]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_4 = {cacheLineTemp[380], cacheLineTemp[372]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_4 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_4 = {memRequest_bits_data_lo_lo_hi_lo_hi_4, memRequest_bits_data_lo_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_4 = {cacheLineTemp[396], cacheLineTemp[388]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_4 = {cacheLineTemp[412], cacheLineTemp[404]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_4, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_4 = {cacheLineTemp[428], cacheLineTemp[420]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_4 = {cacheLineTemp[444], cacheLineTemp[436]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo_4 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_4, memRequest_bits_data_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_4 = {cacheLineTemp[460], cacheLineTemp[452]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_4 = {cacheLineTemp[476], cacheLineTemp[468]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_4 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_4, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_4 = {cacheLineTemp[492], cacheLineTemp[484]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_4 = {cacheLineTemp[508], cacheLineTemp[500]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_4, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_4, memRequest_bits_data_lo_lo_hi_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_hi_4, memRequest_bits_data_lo_lo_hi_hi_lo_4};
  wire [31:0]       memRequest_bits_data_lo_lo_hi_4 = {memRequest_bits_data_lo_lo_hi_hi_4, memRequest_bits_data_lo_lo_hi_lo_4};
  wire [63:0]       memRequest_bits_data_lo_lo_4 = {memRequest_bits_data_lo_lo_hi_4, memRequest_bits_data_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_4 = {cacheLineTemp[524], cacheLineTemp[516]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_4 = {cacheLineTemp[540], cacheLineTemp[532]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_4 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_4 = {cacheLineTemp[556], cacheLineTemp[548]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_4 = {cacheLineTemp[572], cacheLineTemp[564]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_4 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo_4 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_4 = {cacheLineTemp[588], cacheLineTemp[580]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_4 = {cacheLineTemp[604], cacheLineTemp[596]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_4 = {cacheLineTemp[620], cacheLineTemp[612]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_4 = {cacheLineTemp[636], cacheLineTemp[628]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi_4 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_4 = {memRequest_bits_data_lo_hi_lo_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_4 = {cacheLineTemp[652], cacheLineTemp[644]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_4 = {cacheLineTemp[668], cacheLineTemp[660]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_4, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_4 = {cacheLineTemp[684], cacheLineTemp[676]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_4 = {cacheLineTemp[700], cacheLineTemp[692]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_4 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_4 = {cacheLineTemp[716], cacheLineTemp[708]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_4 = {cacheLineTemp[732], cacheLineTemp[724]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_4 = {cacheLineTemp[748], cacheLineTemp[740]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_4 = {cacheLineTemp[764], cacheLineTemp[756]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_4 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_4, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_lo_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_4 = {memRequest_bits_data_lo_hi_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_hi_lo_4};
  wire [31:0]       memRequest_bits_data_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_4 = {cacheLineTemp[780], cacheLineTemp[772]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_4 = {cacheLineTemp[796], cacheLineTemp[788]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_4 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_4, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_4 = {cacheLineTemp[812], cacheLineTemp[804]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_4 = {cacheLineTemp[828], cacheLineTemp[820]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo_4 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_4, memRequest_bits_data_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_4 = {cacheLineTemp[844], cacheLineTemp[836]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_4 = {cacheLineTemp[860], cacheLineTemp[852]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_4 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_4, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_4 = {cacheLineTemp[876], cacheLineTemp[868]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_4 = {cacheLineTemp[892], cacheLineTemp[884]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_4 = {memRequest_bits_data_lo_hi_hi_lo_hi_4, memRequest_bits_data_lo_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_4 = {cacheLineTemp[908], cacheLineTemp[900]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_4 = {cacheLineTemp[924], cacheLineTemp[916]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_4 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_4, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_4 = {cacheLineTemp[940], cacheLineTemp[932]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_4 = {cacheLineTemp[956], cacheLineTemp[948]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_4, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo_4 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_4, memRequest_bits_data_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_4 = {cacheLineTemp[972], cacheLineTemp[964]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_4 = {cacheLineTemp[988], cacheLineTemp[980]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_4 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_4, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_4 = {cacheLineTemp[1004], cacheLineTemp[996]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_4 = {cacheLineTemp[1020], cacheLineTemp[1012]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_hi_lo_4};
  wire [31:0]       memRequest_bits_data_lo_hi_hi_4 = {memRequest_bits_data_lo_hi_hi_hi_4, memRequest_bits_data_lo_hi_hi_lo_4};
  wire [63:0]       memRequest_bits_data_lo_hi_4 = {memRequest_bits_data_lo_hi_hi_4, memRequest_bits_data_lo_hi_lo_4};
  wire [127:0]      memRequest_bits_data_lo_4 = {memRequest_bits_data_lo_hi_4, memRequest_bits_data_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_4 = {dataBuffer_0[12], dataBuffer_0[4]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_4 = {dataBuffer_0[28], dataBuffer_0[20]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_4 = {dataBuffer_0[44], dataBuffer_0[36]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_4 = {dataBuffer_0[60], dataBuffer_0[52]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_4 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_4, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_4 = {dataBuffer_0[76], dataBuffer_0[68]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_4 = {dataBuffer_0[92], dataBuffer_0[84]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_4 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_4 = {dataBuffer_0[108], dataBuffer_0[100]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_4 = {dataBuffer_0[124], dataBuffer_0[116]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_4 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_4, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi_4 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_4, memRequest_bits_data_hi_lo_lo_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_4 = {dataBuffer_0[140], dataBuffer_0[132]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_4 = {dataBuffer_0[156], dataBuffer_0[148]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_4 = {dataBuffer_0[172], dataBuffer_0[164]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_4 = {dataBuffer_0[188], dataBuffer_0[180]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_4 = {dataBuffer_0[204], dataBuffer_0[196]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_4 = {dataBuffer_0[220], dataBuffer_0[212]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_4 = {dataBuffer_0[236], dataBuffer_0[228]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_4 = {dataBuffer_0[252], dataBuffer_0[244]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_4 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_4, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi_4 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_4, memRequest_bits_data_hi_lo_lo_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_4 = {memRequest_bits_data_hi_lo_lo_hi_hi_4, memRequest_bits_data_hi_lo_lo_hi_lo_4};
  wire [31:0]       memRequest_bits_data_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_4 = {dataBuffer_0[268], dataBuffer_0[260]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_4 = {dataBuffer_0[284], dataBuffer_0[276]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_4 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_4, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_4 = {dataBuffer_0[300], dataBuffer_0[292]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_4 = {dataBuffer_0[316], dataBuffer_0[308]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_4 = {dataBuffer_0[332], dataBuffer_0[324]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_4 = {dataBuffer_0[348], dataBuffer_0[340]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_4, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_4 = {dataBuffer_0[364], dataBuffer_0[356]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_4 = {dataBuffer_0[380], dataBuffer_0[372]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_4 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_lo_hi_4, memRequest_bits_data_hi_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_4 = {dataBuffer_0[396], dataBuffer_0[388]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_4 = {dataBuffer_0[412], dataBuffer_0[404]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_4 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_4, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_4 = {dataBuffer_0[428], dataBuffer_0[420]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_4 = {dataBuffer_0[444], dataBuffer_0[436]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_4, memRequest_bits_data_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_4 = {dataBuffer_0[460], dataBuffer_0[452]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_4 = {dataBuffer_0[476], dataBuffer_0[468]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_4, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_4 = {dataBuffer_0[492], dataBuffer_0[484]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_4 = {dataBuffer_0[508], dataBuffer_0[500]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_4, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_4, memRequest_bits_data_hi_lo_hi_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_hi_4, memRequest_bits_data_hi_lo_hi_hi_lo_4};
  wire [31:0]       memRequest_bits_data_hi_lo_hi_4 = {memRequest_bits_data_hi_lo_hi_hi_4, memRequest_bits_data_hi_lo_hi_lo_4};
  wire [63:0]       memRequest_bits_data_hi_lo_4 = {memRequest_bits_data_hi_lo_hi_4, memRequest_bits_data_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_4 = {dataBuffer_0[524], dataBuffer_0[516]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_4 = {dataBuffer_0[540], dataBuffer_0[532]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_4 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_4 = {dataBuffer_0[556], dataBuffer_0[548]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_4 = {dataBuffer_0[572], dataBuffer_0[564]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_4 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_4, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo_4 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_4 = {dataBuffer_0[588], dataBuffer_0[580]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_4 = {dataBuffer_0[604], dataBuffer_0[596]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_4 = {dataBuffer_0[620], dataBuffer_0[612]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_4 = {dataBuffer_0[636], dataBuffer_0[628]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_4 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi_4 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_4, memRequest_bits_data_hi_hi_lo_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_4 = {memRequest_bits_data_hi_hi_lo_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_4 = {dataBuffer_0[652], dataBuffer_0[644]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_4 = {dataBuffer_0[668], dataBuffer_0[660]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_4, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_4 = {dataBuffer_0[684], dataBuffer_0[676]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_4 = {dataBuffer_0[700], dataBuffer_0[692]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_4 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_4, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_4 = {dataBuffer_0[716], dataBuffer_0[708]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_4 = {dataBuffer_0[732], dataBuffer_0[724]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_4 = {dataBuffer_0[748], dataBuffer_0[740]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_4 = {dataBuffer_0[764], dataBuffer_0[756]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi_4 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_4 = {memRequest_bits_data_hi_hi_lo_hi_hi_4, memRequest_bits_data_hi_hi_lo_hi_lo_4};
  wire [31:0]       memRequest_bits_data_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_4 = {dataBuffer_0[780], dataBuffer_0[772]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_4 = {dataBuffer_0[796], dataBuffer_0[788]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_4 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_4, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_4 = {dataBuffer_0[812], dataBuffer_0[804]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_4 = {dataBuffer_0[828], dataBuffer_0[820]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_4 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo_4 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_4, memRequest_bits_data_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_4 = {dataBuffer_0[844], dataBuffer_0[836]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_4 = {dataBuffer_0[860], dataBuffer_0[852]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_4 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_4, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_4 = {dataBuffer_0[876], dataBuffer_0[868]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_4 = {dataBuffer_0[892], dataBuffer_0[884]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi_4 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_4 = {dataBuffer_0[908], dataBuffer_0[900]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_4 = {dataBuffer_0[924], dataBuffer_0[916]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_4 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_4, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_4 = {dataBuffer_0[940], dataBuffer_0[932]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_4 = {dataBuffer_0[956], dataBuffer_0[948]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_4, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_4 = {dataBuffer_0[972], dataBuffer_0[964]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_4 = {dataBuffer_0[988], dataBuffer_0[980]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_4 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_4, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_4};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_4 = {dataBuffer_0[1004], dataBuffer_0[996]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_4 = {dataBuffer_0[1020], dataBuffer_0[1012]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_4};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_hi_hi_lo_4};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_hi_lo_4};
  wire [31:0]       memRequest_bits_data_hi_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_hi_4, memRequest_bits_data_hi_hi_hi_lo_4};
  wire [63:0]       memRequest_bits_data_hi_hi_4 = {memRequest_bits_data_hi_hi_hi_4, memRequest_bits_data_hi_hi_lo_4};
  wire [127:0]      memRequest_bits_data_hi_4 = {memRequest_bits_data_hi_hi_4, memRequest_bits_data_hi_lo_4};
  wire [382:0]      _memRequest_bits_data_T_3590 = {127'h0, memRequest_bits_data_hi_4, memRequest_bits_data_lo_4} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_5 = {cacheLineTemp[13], cacheLineTemp[5]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_5 = {cacheLineTemp[29], cacheLineTemp[21]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_5 = {cacheLineTemp[45], cacheLineTemp[37]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_5 = {cacheLineTemp[61], cacheLineTemp[53]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_5 = {cacheLineTemp[77], cacheLineTemp[69]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_5 = {cacheLineTemp[93], cacheLineTemp[85]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_5 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_5 = {cacheLineTemp[109], cacheLineTemp[101]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_5 = {cacheLineTemp[125], cacheLineTemp[117]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_5 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_5, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_lo_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_5 = {cacheLineTemp[141], cacheLineTemp[133]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_5 = {cacheLineTemp[157], cacheLineTemp[149]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_5 = {cacheLineTemp[173], cacheLineTemp[165]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_5 = {cacheLineTemp[189], cacheLineTemp[181]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_5 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_5, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_5, memRequest_bits_data_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_5 = {cacheLineTemp[205], cacheLineTemp[197]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_5 = {cacheLineTemp[221], cacheLineTemp[213]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_5, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_5 = {cacheLineTemp[237], cacheLineTemp[229]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_5 = {cacheLineTemp[253], cacheLineTemp[245]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_5 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_5, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi_5 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_5, memRequest_bits_data_lo_lo_lo_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_lo_hi_lo_5};
  wire [31:0]       memRequest_bits_data_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_5 = {cacheLineTemp[269], cacheLineTemp[261]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_5 = {cacheLineTemp[285], cacheLineTemp[277]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_5, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_5 = {cacheLineTemp[301], cacheLineTemp[293]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_5 = {cacheLineTemp[317], cacheLineTemp[309]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_5, memRequest_bits_data_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_5 = {cacheLineTemp[333], cacheLineTemp[325]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_5 = {cacheLineTemp[349], cacheLineTemp[341]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_5 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_5, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_5 = {cacheLineTemp[365], cacheLineTemp[357]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_5 = {cacheLineTemp[381], cacheLineTemp[373]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_5 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_5 = {memRequest_bits_data_lo_lo_hi_lo_hi_5, memRequest_bits_data_lo_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_5 = {cacheLineTemp[397], cacheLineTemp[389]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_5 = {cacheLineTemp[413], cacheLineTemp[405]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_5, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_5 = {cacheLineTemp[429], cacheLineTemp[421]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_5 = {cacheLineTemp[445], cacheLineTemp[437]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo_5 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_5, memRequest_bits_data_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_5 = {cacheLineTemp[461], cacheLineTemp[453]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_5 = {cacheLineTemp[477], cacheLineTemp[469]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_5 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_5, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_5 = {cacheLineTemp[493], cacheLineTemp[485]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_5 = {cacheLineTemp[509], cacheLineTemp[501]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_5, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_5, memRequest_bits_data_lo_lo_hi_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_hi_5, memRequest_bits_data_lo_lo_hi_hi_lo_5};
  wire [31:0]       memRequest_bits_data_lo_lo_hi_5 = {memRequest_bits_data_lo_lo_hi_hi_5, memRequest_bits_data_lo_lo_hi_lo_5};
  wire [63:0]       memRequest_bits_data_lo_lo_5 = {memRequest_bits_data_lo_lo_hi_5, memRequest_bits_data_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_5 = {cacheLineTemp[525], cacheLineTemp[517]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_5 = {cacheLineTemp[541], cacheLineTemp[533]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_5 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_5 = {cacheLineTemp[557], cacheLineTemp[549]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_5 = {cacheLineTemp[573], cacheLineTemp[565]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_5 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo_5 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_5 = {cacheLineTemp[589], cacheLineTemp[581]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_5 = {cacheLineTemp[605], cacheLineTemp[597]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_5 = {cacheLineTemp[621], cacheLineTemp[613]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_5 = {cacheLineTemp[637], cacheLineTemp[629]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi_5 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_5 = {memRequest_bits_data_lo_hi_lo_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_5 = {cacheLineTemp[653], cacheLineTemp[645]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_5 = {cacheLineTemp[669], cacheLineTemp[661]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_5, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_5 = {cacheLineTemp[685], cacheLineTemp[677]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_5 = {cacheLineTemp[701], cacheLineTemp[693]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_5 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_5 = {cacheLineTemp[717], cacheLineTemp[709]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_5 = {cacheLineTemp[733], cacheLineTemp[725]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_5 = {cacheLineTemp[749], cacheLineTemp[741]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_5 = {cacheLineTemp[765], cacheLineTemp[757]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_5 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_5, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_lo_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_5 = {memRequest_bits_data_lo_hi_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_hi_lo_5};
  wire [31:0]       memRequest_bits_data_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_5 = {cacheLineTemp[781], cacheLineTemp[773]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_5 = {cacheLineTemp[797], cacheLineTemp[789]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_5 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_5, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_5 = {cacheLineTemp[813], cacheLineTemp[805]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_5 = {cacheLineTemp[829], cacheLineTemp[821]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo_5 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_5, memRequest_bits_data_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_5 = {cacheLineTemp[845], cacheLineTemp[837]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_5 = {cacheLineTemp[861], cacheLineTemp[853]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_5 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_5, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_5 = {cacheLineTemp[877], cacheLineTemp[869]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_5 = {cacheLineTemp[893], cacheLineTemp[885]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_5 = {memRequest_bits_data_lo_hi_hi_lo_hi_5, memRequest_bits_data_lo_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_5 = {cacheLineTemp[909], cacheLineTemp[901]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_5 = {cacheLineTemp[925], cacheLineTemp[917]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_5 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_5, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_5 = {cacheLineTemp[941], cacheLineTemp[933]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_5 = {cacheLineTemp[957], cacheLineTemp[949]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_5, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo_5 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_5, memRequest_bits_data_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_5 = {cacheLineTemp[973], cacheLineTemp[965]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_5 = {cacheLineTemp[989], cacheLineTemp[981]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_5 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_5, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_5 = {cacheLineTemp[1005], cacheLineTemp[997]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_5 = {cacheLineTemp[1021], cacheLineTemp[1013]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_hi_lo_5};
  wire [31:0]       memRequest_bits_data_lo_hi_hi_5 = {memRequest_bits_data_lo_hi_hi_hi_5, memRequest_bits_data_lo_hi_hi_lo_5};
  wire [63:0]       memRequest_bits_data_lo_hi_5 = {memRequest_bits_data_lo_hi_hi_5, memRequest_bits_data_lo_hi_lo_5};
  wire [127:0]      memRequest_bits_data_lo_5 = {memRequest_bits_data_lo_hi_5, memRequest_bits_data_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_5 = {dataBuffer_0[13], dataBuffer_0[5]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_5 = {dataBuffer_0[29], dataBuffer_0[21]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_5 = {dataBuffer_0[45], dataBuffer_0[37]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_5 = {dataBuffer_0[61], dataBuffer_0[53]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_5 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_5, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_5 = {dataBuffer_0[77], dataBuffer_0[69]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_5 = {dataBuffer_0[93], dataBuffer_0[85]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_5 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_5 = {dataBuffer_0[109], dataBuffer_0[101]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_5 = {dataBuffer_0[125], dataBuffer_0[117]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_5 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_5, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi_5 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_5, memRequest_bits_data_hi_lo_lo_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_5 = {dataBuffer_0[141], dataBuffer_0[133]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_5 = {dataBuffer_0[157], dataBuffer_0[149]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_5 = {dataBuffer_0[173], dataBuffer_0[165]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_5 = {dataBuffer_0[189], dataBuffer_0[181]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_5 = {dataBuffer_0[205], dataBuffer_0[197]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_5 = {dataBuffer_0[221], dataBuffer_0[213]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_5 = {dataBuffer_0[237], dataBuffer_0[229]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_5 = {dataBuffer_0[253], dataBuffer_0[245]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_5 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_5, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi_5 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_5, memRequest_bits_data_hi_lo_lo_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_5 = {memRequest_bits_data_hi_lo_lo_hi_hi_5, memRequest_bits_data_hi_lo_lo_hi_lo_5};
  wire [31:0]       memRequest_bits_data_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_5 = {dataBuffer_0[269], dataBuffer_0[261]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_5 = {dataBuffer_0[285], dataBuffer_0[277]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_5 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_5, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_5 = {dataBuffer_0[301], dataBuffer_0[293]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_5 = {dataBuffer_0[317], dataBuffer_0[309]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_5 = {dataBuffer_0[333], dataBuffer_0[325]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_5 = {dataBuffer_0[349], dataBuffer_0[341]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_5, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_5 = {dataBuffer_0[365], dataBuffer_0[357]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_5 = {dataBuffer_0[381], dataBuffer_0[373]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_5 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_lo_hi_5, memRequest_bits_data_hi_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_5 = {dataBuffer_0[397], dataBuffer_0[389]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_5 = {dataBuffer_0[413], dataBuffer_0[405]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_5 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_5, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_5 = {dataBuffer_0[429], dataBuffer_0[421]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_5 = {dataBuffer_0[445], dataBuffer_0[437]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_5, memRequest_bits_data_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_5 = {dataBuffer_0[461], dataBuffer_0[453]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_5 = {dataBuffer_0[477], dataBuffer_0[469]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_5, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_5 = {dataBuffer_0[493], dataBuffer_0[485]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_5 = {dataBuffer_0[509], dataBuffer_0[501]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_5, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_5, memRequest_bits_data_hi_lo_hi_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_hi_5, memRequest_bits_data_hi_lo_hi_hi_lo_5};
  wire [31:0]       memRequest_bits_data_hi_lo_hi_5 = {memRequest_bits_data_hi_lo_hi_hi_5, memRequest_bits_data_hi_lo_hi_lo_5};
  wire [63:0]       memRequest_bits_data_hi_lo_5 = {memRequest_bits_data_hi_lo_hi_5, memRequest_bits_data_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_5 = {dataBuffer_0[525], dataBuffer_0[517]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_5 = {dataBuffer_0[541], dataBuffer_0[533]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_5 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_5 = {dataBuffer_0[557], dataBuffer_0[549]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_5 = {dataBuffer_0[573], dataBuffer_0[565]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_5 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_5, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo_5 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_5 = {dataBuffer_0[589], dataBuffer_0[581]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_5 = {dataBuffer_0[605], dataBuffer_0[597]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_5 = {dataBuffer_0[621], dataBuffer_0[613]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_5 = {dataBuffer_0[637], dataBuffer_0[629]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_5 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi_5 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_5, memRequest_bits_data_hi_hi_lo_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_5 = {memRequest_bits_data_hi_hi_lo_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_5 = {dataBuffer_0[653], dataBuffer_0[645]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_5 = {dataBuffer_0[669], dataBuffer_0[661]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_5, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_5 = {dataBuffer_0[685], dataBuffer_0[677]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_5 = {dataBuffer_0[701], dataBuffer_0[693]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_5 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_5, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_5 = {dataBuffer_0[717], dataBuffer_0[709]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_5 = {dataBuffer_0[733], dataBuffer_0[725]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_5 = {dataBuffer_0[749], dataBuffer_0[741]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_5 = {dataBuffer_0[765], dataBuffer_0[757]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi_5 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_5 = {memRequest_bits_data_hi_hi_lo_hi_hi_5, memRequest_bits_data_hi_hi_lo_hi_lo_5};
  wire [31:0]       memRequest_bits_data_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_5 = {dataBuffer_0[781], dataBuffer_0[773]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_5 = {dataBuffer_0[797], dataBuffer_0[789]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_5 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_5, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_5 = {dataBuffer_0[813], dataBuffer_0[805]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_5 = {dataBuffer_0[829], dataBuffer_0[821]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_5 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo_5 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_5, memRequest_bits_data_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_5 = {dataBuffer_0[845], dataBuffer_0[837]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_5 = {dataBuffer_0[861], dataBuffer_0[853]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_5 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_5, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_5 = {dataBuffer_0[877], dataBuffer_0[869]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_5 = {dataBuffer_0[893], dataBuffer_0[885]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi_5 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_5 = {dataBuffer_0[909], dataBuffer_0[901]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_5 = {dataBuffer_0[925], dataBuffer_0[917]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_5 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_5, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_5 = {dataBuffer_0[941], dataBuffer_0[933]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_5 = {dataBuffer_0[957], dataBuffer_0[949]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_5, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_5 = {dataBuffer_0[973], dataBuffer_0[965]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_5 = {dataBuffer_0[989], dataBuffer_0[981]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_5 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_5, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_5};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_5 = {dataBuffer_0[1005], dataBuffer_0[997]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_5 = {dataBuffer_0[1021], dataBuffer_0[1013]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_5};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_hi_hi_lo_5};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_hi_lo_5};
  wire [31:0]       memRequest_bits_data_hi_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_hi_5, memRequest_bits_data_hi_hi_hi_lo_5};
  wire [63:0]       memRequest_bits_data_hi_hi_5 = {memRequest_bits_data_hi_hi_hi_5, memRequest_bits_data_hi_hi_lo_5};
  wire [127:0]      memRequest_bits_data_hi_5 = {memRequest_bits_data_hi_hi_5, memRequest_bits_data_hi_lo_5};
  wire [382:0]      _memRequest_bits_data_T_3975 = {127'h0, memRequest_bits_data_hi_5, memRequest_bits_data_lo_5} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_6 = {cacheLineTemp[14], cacheLineTemp[6]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_6 = {cacheLineTemp[30], cacheLineTemp[22]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_6 = {cacheLineTemp[46], cacheLineTemp[38]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_6 = {cacheLineTemp[62], cacheLineTemp[54]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_6 = {cacheLineTemp[78], cacheLineTemp[70]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_6 = {cacheLineTemp[94], cacheLineTemp[86]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_6 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_6 = {cacheLineTemp[110], cacheLineTemp[102]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_6 = {cacheLineTemp[126], cacheLineTemp[118]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_6 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_6, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_lo_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_6 = {cacheLineTemp[142], cacheLineTemp[134]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_6 = {cacheLineTemp[158], cacheLineTemp[150]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_6 = {cacheLineTemp[174], cacheLineTemp[166]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_6 = {cacheLineTemp[190], cacheLineTemp[182]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_6 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_6, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_6, memRequest_bits_data_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_6 = {cacheLineTemp[206], cacheLineTemp[198]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_6 = {cacheLineTemp[222], cacheLineTemp[214]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_6, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_6 = {cacheLineTemp[238], cacheLineTemp[230]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_6 = {cacheLineTemp[254], cacheLineTemp[246]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_6 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_6, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi_6 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_6, memRequest_bits_data_lo_lo_lo_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_lo_hi_lo_6};
  wire [31:0]       memRequest_bits_data_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_6 = {cacheLineTemp[270], cacheLineTemp[262]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_6 = {cacheLineTemp[286], cacheLineTemp[278]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_6, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_6 = {cacheLineTemp[302], cacheLineTemp[294]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_6 = {cacheLineTemp[318], cacheLineTemp[310]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_6, memRequest_bits_data_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_6 = {cacheLineTemp[334], cacheLineTemp[326]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_6 = {cacheLineTemp[350], cacheLineTemp[342]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_6 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_6, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_6 = {cacheLineTemp[366], cacheLineTemp[358]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_6 = {cacheLineTemp[382], cacheLineTemp[374]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_6 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_6 = {memRequest_bits_data_lo_lo_hi_lo_hi_6, memRequest_bits_data_lo_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_6 = {cacheLineTemp[398], cacheLineTemp[390]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_6 = {cacheLineTemp[414], cacheLineTemp[406]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_6, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_6 = {cacheLineTemp[430], cacheLineTemp[422]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_6 = {cacheLineTemp[446], cacheLineTemp[438]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo_6 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_6, memRequest_bits_data_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_6 = {cacheLineTemp[462], cacheLineTemp[454]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_6 = {cacheLineTemp[478], cacheLineTemp[470]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_6 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_6, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_6 = {cacheLineTemp[494], cacheLineTemp[486]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_6 = {cacheLineTemp[510], cacheLineTemp[502]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_6, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_6, memRequest_bits_data_lo_lo_hi_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_hi_6, memRequest_bits_data_lo_lo_hi_hi_lo_6};
  wire [31:0]       memRequest_bits_data_lo_lo_hi_6 = {memRequest_bits_data_lo_lo_hi_hi_6, memRequest_bits_data_lo_lo_hi_lo_6};
  wire [63:0]       memRequest_bits_data_lo_lo_6 = {memRequest_bits_data_lo_lo_hi_6, memRequest_bits_data_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_6 = {cacheLineTemp[526], cacheLineTemp[518]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_6 = {cacheLineTemp[542], cacheLineTemp[534]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_6 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_6 = {cacheLineTemp[558], cacheLineTemp[550]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_6 = {cacheLineTemp[574], cacheLineTemp[566]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_6 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo_6 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_6 = {cacheLineTemp[590], cacheLineTemp[582]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_6 = {cacheLineTemp[606], cacheLineTemp[598]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_6 = {cacheLineTemp[622], cacheLineTemp[614]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_6 = {cacheLineTemp[638], cacheLineTemp[630]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi_6 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_6 = {memRequest_bits_data_lo_hi_lo_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_6 = {cacheLineTemp[654], cacheLineTemp[646]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_6 = {cacheLineTemp[670], cacheLineTemp[662]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_6, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_6 = {cacheLineTemp[686], cacheLineTemp[678]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_6 = {cacheLineTemp[702], cacheLineTemp[694]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_6 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_6 = {cacheLineTemp[718], cacheLineTemp[710]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_6 = {cacheLineTemp[734], cacheLineTemp[726]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_6 = {cacheLineTemp[750], cacheLineTemp[742]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_6 = {cacheLineTemp[766], cacheLineTemp[758]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_6 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_6, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_lo_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_6 = {memRequest_bits_data_lo_hi_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_hi_lo_6};
  wire [31:0]       memRequest_bits_data_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_6 = {cacheLineTemp[782], cacheLineTemp[774]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_6 = {cacheLineTemp[798], cacheLineTemp[790]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_6 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_6, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_6 = {cacheLineTemp[814], cacheLineTemp[806]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_6 = {cacheLineTemp[830], cacheLineTemp[822]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo_6 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_6, memRequest_bits_data_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_6 = {cacheLineTemp[846], cacheLineTemp[838]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_6 = {cacheLineTemp[862], cacheLineTemp[854]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_6 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_6, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_6 = {cacheLineTemp[878], cacheLineTemp[870]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_6 = {cacheLineTemp[894], cacheLineTemp[886]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_6 = {memRequest_bits_data_lo_hi_hi_lo_hi_6, memRequest_bits_data_lo_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_6 = {cacheLineTemp[910], cacheLineTemp[902]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_6 = {cacheLineTemp[926], cacheLineTemp[918]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_6 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_6, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_6 = {cacheLineTemp[942], cacheLineTemp[934]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_6 = {cacheLineTemp[958], cacheLineTemp[950]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_6, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo_6 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_6, memRequest_bits_data_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_6 = {cacheLineTemp[974], cacheLineTemp[966]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_6 = {cacheLineTemp[990], cacheLineTemp[982]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_6 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_6, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_6 = {cacheLineTemp[1006], cacheLineTemp[998]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_6 = {cacheLineTemp[1022], cacheLineTemp[1014]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_hi_lo_6};
  wire [31:0]       memRequest_bits_data_lo_hi_hi_6 = {memRequest_bits_data_lo_hi_hi_hi_6, memRequest_bits_data_lo_hi_hi_lo_6};
  wire [63:0]       memRequest_bits_data_lo_hi_6 = {memRequest_bits_data_lo_hi_hi_6, memRequest_bits_data_lo_hi_lo_6};
  wire [127:0]      memRequest_bits_data_lo_6 = {memRequest_bits_data_lo_hi_6, memRequest_bits_data_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_6 = {dataBuffer_0[14], dataBuffer_0[6]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_6 = {dataBuffer_0[30], dataBuffer_0[22]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_6 = {dataBuffer_0[46], dataBuffer_0[38]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_6 = {dataBuffer_0[62], dataBuffer_0[54]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_6 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_6, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_6 = {dataBuffer_0[78], dataBuffer_0[70]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_6 = {dataBuffer_0[94], dataBuffer_0[86]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_6 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_6 = {dataBuffer_0[110], dataBuffer_0[102]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_6 = {dataBuffer_0[126], dataBuffer_0[118]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_6 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_6, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi_6 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_6, memRequest_bits_data_hi_lo_lo_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_6 = {dataBuffer_0[142], dataBuffer_0[134]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_6 = {dataBuffer_0[158], dataBuffer_0[150]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_6 = {dataBuffer_0[174], dataBuffer_0[166]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_6 = {dataBuffer_0[190], dataBuffer_0[182]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_6 = {dataBuffer_0[206], dataBuffer_0[198]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_6 = {dataBuffer_0[222], dataBuffer_0[214]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_6 = {dataBuffer_0[238], dataBuffer_0[230]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_6 = {dataBuffer_0[254], dataBuffer_0[246]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_6 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_6, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi_6 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_6, memRequest_bits_data_hi_lo_lo_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_6 = {memRequest_bits_data_hi_lo_lo_hi_hi_6, memRequest_bits_data_hi_lo_lo_hi_lo_6};
  wire [31:0]       memRequest_bits_data_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_6 = {dataBuffer_0[270], dataBuffer_0[262]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_6 = {dataBuffer_0[286], dataBuffer_0[278]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_6 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_6, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_6 = {dataBuffer_0[302], dataBuffer_0[294]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_6 = {dataBuffer_0[318], dataBuffer_0[310]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_6 = {dataBuffer_0[334], dataBuffer_0[326]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_6 = {dataBuffer_0[350], dataBuffer_0[342]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_6, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_6 = {dataBuffer_0[366], dataBuffer_0[358]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_6 = {dataBuffer_0[382], dataBuffer_0[374]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_6 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_lo_hi_6, memRequest_bits_data_hi_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_6 = {dataBuffer_0[398], dataBuffer_0[390]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_6 = {dataBuffer_0[414], dataBuffer_0[406]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_6 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_6, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_6 = {dataBuffer_0[430], dataBuffer_0[422]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_6 = {dataBuffer_0[446], dataBuffer_0[438]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_6, memRequest_bits_data_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_6 = {dataBuffer_0[462], dataBuffer_0[454]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_6 = {dataBuffer_0[478], dataBuffer_0[470]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_6, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_6 = {dataBuffer_0[494], dataBuffer_0[486]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_6 = {dataBuffer_0[510], dataBuffer_0[502]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_6, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_6, memRequest_bits_data_hi_lo_hi_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_hi_6, memRequest_bits_data_hi_lo_hi_hi_lo_6};
  wire [31:0]       memRequest_bits_data_hi_lo_hi_6 = {memRequest_bits_data_hi_lo_hi_hi_6, memRequest_bits_data_hi_lo_hi_lo_6};
  wire [63:0]       memRequest_bits_data_hi_lo_6 = {memRequest_bits_data_hi_lo_hi_6, memRequest_bits_data_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_6 = {dataBuffer_0[526], dataBuffer_0[518]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_6 = {dataBuffer_0[542], dataBuffer_0[534]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_6 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_6 = {dataBuffer_0[558], dataBuffer_0[550]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_6 = {dataBuffer_0[574], dataBuffer_0[566]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_6 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_6, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo_6 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_6 = {dataBuffer_0[590], dataBuffer_0[582]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_6 = {dataBuffer_0[606], dataBuffer_0[598]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_6 = {dataBuffer_0[622], dataBuffer_0[614]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_6 = {dataBuffer_0[638], dataBuffer_0[630]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_6 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi_6 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_6, memRequest_bits_data_hi_hi_lo_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_6 = {memRequest_bits_data_hi_hi_lo_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_6 = {dataBuffer_0[654], dataBuffer_0[646]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_6 = {dataBuffer_0[670], dataBuffer_0[662]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_6, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_6 = {dataBuffer_0[686], dataBuffer_0[678]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_6 = {dataBuffer_0[702], dataBuffer_0[694]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_6 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_6, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_6 = {dataBuffer_0[718], dataBuffer_0[710]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_6 = {dataBuffer_0[734], dataBuffer_0[726]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_6 = {dataBuffer_0[750], dataBuffer_0[742]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_6 = {dataBuffer_0[766], dataBuffer_0[758]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi_6 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_6 = {memRequest_bits_data_hi_hi_lo_hi_hi_6, memRequest_bits_data_hi_hi_lo_hi_lo_6};
  wire [31:0]       memRequest_bits_data_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_6 = {dataBuffer_0[782], dataBuffer_0[774]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_6 = {dataBuffer_0[798], dataBuffer_0[790]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_6 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_6, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_6 = {dataBuffer_0[814], dataBuffer_0[806]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_6 = {dataBuffer_0[830], dataBuffer_0[822]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_6 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo_6 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_6, memRequest_bits_data_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_6 = {dataBuffer_0[846], dataBuffer_0[838]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_6 = {dataBuffer_0[862], dataBuffer_0[854]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_6 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_6, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_6 = {dataBuffer_0[878], dataBuffer_0[870]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_6 = {dataBuffer_0[894], dataBuffer_0[886]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi_6 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_6 = {dataBuffer_0[910], dataBuffer_0[902]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_6 = {dataBuffer_0[926], dataBuffer_0[918]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_6 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_6, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_6 = {dataBuffer_0[942], dataBuffer_0[934]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_6 = {dataBuffer_0[958], dataBuffer_0[950]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_6, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_6 = {dataBuffer_0[974], dataBuffer_0[966]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_6 = {dataBuffer_0[990], dataBuffer_0[982]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_6 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_6, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_6};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_6 = {dataBuffer_0[1006], dataBuffer_0[998]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_6 = {dataBuffer_0[1022], dataBuffer_0[1014]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_6};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_hi_hi_lo_6};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_hi_lo_6};
  wire [31:0]       memRequest_bits_data_hi_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_hi_6, memRequest_bits_data_hi_hi_hi_lo_6};
  wire [63:0]       memRequest_bits_data_hi_hi_6 = {memRequest_bits_data_hi_hi_hi_6, memRequest_bits_data_hi_hi_lo_6};
  wire [127:0]      memRequest_bits_data_hi_6 = {memRequest_bits_data_hi_hi_6, memRequest_bits_data_hi_lo_6};
  wire [382:0]      _memRequest_bits_data_T_4360 = {127'h0, memRequest_bits_data_hi_6, memRequest_bits_data_lo_6} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_7 = {cacheLineTemp[15], cacheLineTemp[7]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_7 = {cacheLineTemp[31], cacheLineTemp[23]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_7 = {cacheLineTemp[47], cacheLineTemp[39]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_7 = {cacheLineTemp[63], cacheLineTemp[55]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_7 = {cacheLineTemp[79], cacheLineTemp[71]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_7 = {cacheLineTemp[95], cacheLineTemp[87]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_lo_7 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_7 = {cacheLineTemp[111], cacheLineTemp[103]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_7 = {cacheLineTemp[127], cacheLineTemp[119]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_lo_hi_hi_7 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_7, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_lo_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_7 = {cacheLineTemp[143], cacheLineTemp[135]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_7 = {cacheLineTemp[159], cacheLineTemp[151]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_7 = {cacheLineTemp[175], cacheLineTemp[167]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_7 = {cacheLineTemp[191], cacheLineTemp[183]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_lo_hi_7 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_7, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_7, memRequest_bits_data_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_7 = {cacheLineTemp[207], cacheLineTemp[199]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_7 = {cacheLineTemp[223], cacheLineTemp[215]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_7, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_7 = {cacheLineTemp[239], cacheLineTemp[231]};
  wire [1:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_7 = {cacheLineTemp[255], cacheLineTemp[247]};
  wire [3:0]        memRequest_bits_data_lo_lo_lo_hi_hi_hi_7 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_7, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_lo_hi_hi_7 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_7, memRequest_bits_data_lo_lo_lo_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_lo_hi_lo_7};
  wire [31:0]       memRequest_bits_data_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_7 = {cacheLineTemp[271], cacheLineTemp[263]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_7 = {cacheLineTemp[287], cacheLineTemp[279]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_7, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_7 = {cacheLineTemp[303], cacheLineTemp[295]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_7 = {cacheLineTemp[319], cacheLineTemp[311]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_7, memRequest_bits_data_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_7 = {cacheLineTemp[335], cacheLineTemp[327]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_7 = {cacheLineTemp[351], cacheLineTemp[343]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_lo_7 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_7, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_7 = {cacheLineTemp[367], cacheLineTemp[359]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_7 = {cacheLineTemp[383], cacheLineTemp[375]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_lo_hi_hi_7 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_7 = {memRequest_bits_data_lo_lo_hi_lo_hi_7, memRequest_bits_data_lo_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_7 = {cacheLineTemp[399], cacheLineTemp[391]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_7 = {cacheLineTemp[415], cacheLineTemp[407]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_7, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_7 = {cacheLineTemp[431], cacheLineTemp[423]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_7 = {cacheLineTemp[447], cacheLineTemp[439]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_lo_7 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_7, memRequest_bits_data_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_7 = {cacheLineTemp[463], cacheLineTemp[455]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_7 = {cacheLineTemp[479], cacheLineTemp[471]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_lo_7 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_7, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_7 = {cacheLineTemp[495], cacheLineTemp[487]};
  wire [1:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_7 = {cacheLineTemp[511], cacheLineTemp[503]};
  wire [3:0]        memRequest_bits_data_lo_lo_hi_hi_hi_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_7, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_lo_hi_hi_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_7, memRequest_bits_data_lo_lo_hi_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_hi_7, memRequest_bits_data_lo_lo_hi_hi_lo_7};
  wire [31:0]       memRequest_bits_data_lo_lo_hi_7 = {memRequest_bits_data_lo_lo_hi_hi_7, memRequest_bits_data_lo_lo_hi_lo_7};
  wire [63:0]       memRequest_bits_data_lo_lo_7 = {memRequest_bits_data_lo_lo_hi_7, memRequest_bits_data_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_7 = {cacheLineTemp[527], cacheLineTemp[519]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_7 = {cacheLineTemp[543], cacheLineTemp[535]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_lo_7 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_7 = {cacheLineTemp[559], cacheLineTemp[551]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_7 = {cacheLineTemp[575], cacheLineTemp[567]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_lo_hi_7 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_lo_7 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_7 = {cacheLineTemp[591], cacheLineTemp[583]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_7 = {cacheLineTemp[607], cacheLineTemp[599]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_7 = {cacheLineTemp[623], cacheLineTemp[615]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_7 = {cacheLineTemp[639], cacheLineTemp[631]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_lo_hi_7 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_7 = {memRequest_bits_data_lo_hi_lo_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_7 = {cacheLineTemp[655], cacheLineTemp[647]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_7 = {cacheLineTemp[671], cacheLineTemp[663]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_7, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_7 = {cacheLineTemp[687], cacheLineTemp[679]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_7 = {cacheLineTemp[703], cacheLineTemp[695]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_lo_hi_7 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_7 = {cacheLineTemp[719], cacheLineTemp[711]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_7 = {cacheLineTemp[735], cacheLineTemp[727]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_7 = {cacheLineTemp[751], cacheLineTemp[743]};
  wire [1:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_7 = {cacheLineTemp[767], cacheLineTemp[759]};
  wire [3:0]        memRequest_bits_data_lo_hi_lo_hi_hi_hi_7 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_7, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_lo_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_7 = {memRequest_bits_data_lo_hi_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_hi_lo_7};
  wire [31:0]       memRequest_bits_data_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_7 = {cacheLineTemp[783], cacheLineTemp[775]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_7 = {cacheLineTemp[799], cacheLineTemp[791]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_lo_7 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_7, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_7 = {cacheLineTemp[815], cacheLineTemp[807]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_7 = {cacheLineTemp[831], cacheLineTemp[823]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_lo_7 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_7, memRequest_bits_data_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_7 = {cacheLineTemp[847], cacheLineTemp[839]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_7 = {cacheLineTemp[863], cacheLineTemp[855]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_lo_7 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_7, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_7 = {cacheLineTemp[879], cacheLineTemp[871]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_7 = {cacheLineTemp[895], cacheLineTemp[887]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_7 = {memRequest_bits_data_lo_hi_hi_lo_hi_7, memRequest_bits_data_lo_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_7 = {cacheLineTemp[911], cacheLineTemp[903]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_7 = {cacheLineTemp[927], cacheLineTemp[919]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_lo_7 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_7, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_7 = {cacheLineTemp[943], cacheLineTemp[935]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_7 = {cacheLineTemp[959], cacheLineTemp[951]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_7, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_lo_7 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_7, memRequest_bits_data_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_7 = {cacheLineTemp[975], cacheLineTemp[967]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_7 = {cacheLineTemp[991], cacheLineTemp[983]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_lo_7 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_7, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_7 = {cacheLineTemp[1007], cacheLineTemp[999]};
  wire [1:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_7 = {cacheLineTemp[1023], cacheLineTemp[1015]};
  wire [3:0]        memRequest_bits_data_lo_hi_hi_hi_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_lo_hi_hi_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_hi_lo_7};
  wire [31:0]       memRequest_bits_data_lo_hi_hi_7 = {memRequest_bits_data_lo_hi_hi_hi_7, memRequest_bits_data_lo_hi_hi_lo_7};
  wire [63:0]       memRequest_bits_data_lo_hi_7 = {memRequest_bits_data_lo_hi_hi_7, memRequest_bits_data_lo_hi_lo_7};
  wire [127:0]      memRequest_bits_data_lo_7 = {memRequest_bits_data_lo_hi_7, memRequest_bits_data_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_7 = {dataBuffer_0[15], dataBuffer_0[7]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_7 = {dataBuffer_0[31], dataBuffer_0[23]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_7 = {dataBuffer_0[47], dataBuffer_0[39]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_7 = {dataBuffer_0[63], dataBuffer_0[55]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_lo_hi_7 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_7, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_7 = {dataBuffer_0[79], dataBuffer_0[71]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_7 = {dataBuffer_0[95], dataBuffer_0[87]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_lo_7 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_7 = {dataBuffer_0[111], dataBuffer_0[103]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_7 = {dataBuffer_0[127], dataBuffer_0[119]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_lo_hi_hi_7 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_7, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_lo_hi_7 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_7, memRequest_bits_data_hi_lo_lo_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_7 = {dataBuffer_0[143], dataBuffer_0[135]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_7 = {dataBuffer_0[159], dataBuffer_0[151]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_7 = {dataBuffer_0[175], dataBuffer_0[167]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_7 = {dataBuffer_0[191], dataBuffer_0[183]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_7 = {dataBuffer_0[207], dataBuffer_0[199]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_7 = {dataBuffer_0[223], dataBuffer_0[215]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_7 = {dataBuffer_0[239], dataBuffer_0[231]};
  wire [1:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_7 = {dataBuffer_0[255], dataBuffer_0[247]};
  wire [3:0]        memRequest_bits_data_hi_lo_lo_hi_hi_hi_7 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_7, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_lo_hi_hi_7 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_7, memRequest_bits_data_hi_lo_lo_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_7 = {memRequest_bits_data_hi_lo_lo_hi_hi_7, memRequest_bits_data_hi_lo_lo_hi_lo_7};
  wire [31:0]       memRequest_bits_data_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_7 = {dataBuffer_0[271], dataBuffer_0[263]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_7 = {dataBuffer_0[287], dataBuffer_0[279]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_lo_7 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_7, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_7 = {dataBuffer_0[303], dataBuffer_0[295]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_7 = {dataBuffer_0[319], dataBuffer_0[311]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_7 = {dataBuffer_0[335], dataBuffer_0[327]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_7 = {dataBuffer_0[351], dataBuffer_0[343]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_7, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_7 = {dataBuffer_0[367], dataBuffer_0[359]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_7 = {dataBuffer_0[383], dataBuffer_0[375]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_lo_hi_hi_7 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_lo_hi_7, memRequest_bits_data_hi_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_7 = {dataBuffer_0[399], dataBuffer_0[391]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_7 = {dataBuffer_0[415], dataBuffer_0[407]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_lo_7 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_7, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_7 = {dataBuffer_0[431], dataBuffer_0[423]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_7 = {dataBuffer_0[447], dataBuffer_0[439]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_7, memRequest_bits_data_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_7 = {dataBuffer_0[463], dataBuffer_0[455]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_7 = {dataBuffer_0[479], dataBuffer_0[471]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_7, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_7 = {dataBuffer_0[495], dataBuffer_0[487]};
  wire [1:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_7 = {dataBuffer_0[511], dataBuffer_0[503]};
  wire [3:0]        memRequest_bits_data_hi_lo_hi_hi_hi_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_7, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_lo_hi_hi_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_7, memRequest_bits_data_hi_lo_hi_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_hi_7, memRequest_bits_data_hi_lo_hi_hi_lo_7};
  wire [31:0]       memRequest_bits_data_hi_lo_hi_7 = {memRequest_bits_data_hi_lo_hi_hi_7, memRequest_bits_data_hi_lo_hi_lo_7};
  wire [63:0]       memRequest_bits_data_hi_lo_7 = {memRequest_bits_data_hi_lo_hi_7, memRequest_bits_data_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_7 = {dataBuffer_0[527], dataBuffer_0[519]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_7 = {dataBuffer_0[543], dataBuffer_0[535]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_lo_7 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_7 = {dataBuffer_0[559], dataBuffer_0[551]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_7 = {dataBuffer_0[575], dataBuffer_0[567]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_lo_hi_7 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_7, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_lo_7 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_7 = {dataBuffer_0[591], dataBuffer_0[583]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_7 = {dataBuffer_0[607], dataBuffer_0[599]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_7 = {dataBuffer_0[623], dataBuffer_0[615]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_7 = {dataBuffer_0[639], dataBuffer_0[631]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_lo_hi_hi_7 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_lo_hi_7 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_7, memRequest_bits_data_hi_hi_lo_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_7 = {memRequest_bits_data_hi_hi_lo_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_7 = {dataBuffer_0[655], dataBuffer_0[647]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_7 = {dataBuffer_0[671], dataBuffer_0[663]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_7, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_7 = {dataBuffer_0[687], dataBuffer_0[679]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_7 = {dataBuffer_0[703], dataBuffer_0[695]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_lo_hi_7 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_7, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_7 = {dataBuffer_0[719], dataBuffer_0[711]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_7 = {dataBuffer_0[735], dataBuffer_0[727]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_7 = {dataBuffer_0[751], dataBuffer_0[743]};
  wire [1:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_7 = {dataBuffer_0[767], dataBuffer_0[759]};
  wire [3:0]        memRequest_bits_data_hi_hi_lo_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_lo_hi_hi_7 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_7 = {memRequest_bits_data_hi_hi_lo_hi_hi_7, memRequest_bits_data_hi_hi_lo_hi_lo_7};
  wire [31:0]       memRequest_bits_data_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_7 = {dataBuffer_0[783], dataBuffer_0[775]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_7 = {dataBuffer_0[799], dataBuffer_0[791]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_lo_7 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_7, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_7 = {dataBuffer_0[815], dataBuffer_0[807]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_7 = {dataBuffer_0[831], dataBuffer_0[823]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_lo_hi_7 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_lo_7 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_7, memRequest_bits_data_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_7 = {dataBuffer_0[847], dataBuffer_0[839]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_7 = {dataBuffer_0[863], dataBuffer_0[855]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_lo_7 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_7, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_7 = {dataBuffer_0[879], dataBuffer_0[871]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_7 = {dataBuffer_0[895], dataBuffer_0[887]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_lo_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_lo_hi_7 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_7 = {dataBuffer_0[911], dataBuffer_0[903]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_7 = {dataBuffer_0[927], dataBuffer_0[919]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_lo_7 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_7, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_7 = {dataBuffer_0[943], dataBuffer_0[935]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_7 = {dataBuffer_0[959], dataBuffer_0[951]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_lo_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_7, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_7 = {dataBuffer_0[975], dataBuffer_0[967]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_7 = {dataBuffer_0[991], dataBuffer_0[983]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_lo_7 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_7, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_7};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_7 = {dataBuffer_0[1007], dataBuffer_0[999]};
  wire [1:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_7 = {dataBuffer_0[1023], dataBuffer_0[1015]};
  wire [3:0]        memRequest_bits_data_hi_hi_hi_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_7};
  wire [7:0]        memRequest_bits_data_hi_hi_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_hi_hi_lo_7};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_hi_lo_7};
  wire [31:0]       memRequest_bits_data_hi_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_hi_7, memRequest_bits_data_hi_hi_hi_lo_7};
  wire [63:0]       memRequest_bits_data_hi_hi_7 = {memRequest_bits_data_hi_hi_hi_7, memRequest_bits_data_hi_hi_lo_7};
  wire [127:0]      memRequest_bits_data_hi_7 = {memRequest_bits_data_hi_hi_7, memRequest_bits_data_hi_lo_7};
  wire [382:0]      _memRequest_bits_data_T_4745 = {127'h0, memRequest_bits_data_hi_7, memRequest_bits_data_lo_7} << _GEN_1130;
  wire [1:0]        memRequest_bits_data_lo_lo_8 = {_memRequest_bits_data_T_2435[0], _memRequest_bits_data_T_2050[0]};
  wire [1:0]        memRequest_bits_data_lo_hi_8 = {_memRequest_bits_data_T_3205[0], _memRequest_bits_data_T_2820[0]};
  wire [3:0]        memRequest_bits_data_lo_8 = {memRequest_bits_data_lo_hi_8, memRequest_bits_data_lo_lo_8};
  wire [1:0]        memRequest_bits_data_hi_lo_8 = {_memRequest_bits_data_T_3975[0], _memRequest_bits_data_T_3590[0]};
  wire [1:0]        memRequest_bits_data_hi_hi_8 = {_memRequest_bits_data_T_4745[0], _memRequest_bits_data_T_4360[0]};
  wire [3:0]        memRequest_bits_data_hi_8 = {memRequest_bits_data_hi_hi_8, memRequest_bits_data_hi_lo_8};
  wire [1:0]        memRequest_bits_data_lo_lo_9 = {_memRequest_bits_data_T_2435[1], _memRequest_bits_data_T_2050[1]};
  wire [1:0]        memRequest_bits_data_lo_hi_9 = {_memRequest_bits_data_T_3205[1], _memRequest_bits_data_T_2820[1]};
  wire [3:0]        memRequest_bits_data_lo_9 = {memRequest_bits_data_lo_hi_9, memRequest_bits_data_lo_lo_9};
  wire [1:0]        memRequest_bits_data_hi_lo_9 = {_memRequest_bits_data_T_3975[1], _memRequest_bits_data_T_3590[1]};
  wire [1:0]        memRequest_bits_data_hi_hi_9 = {_memRequest_bits_data_T_4745[1], _memRequest_bits_data_T_4360[1]};
  wire [3:0]        memRequest_bits_data_hi_9 = {memRequest_bits_data_hi_hi_9, memRequest_bits_data_hi_lo_9};
  wire [1:0]        memRequest_bits_data_lo_lo_10 = {_memRequest_bits_data_T_2435[2], _memRequest_bits_data_T_2050[2]};
  wire [1:0]        memRequest_bits_data_lo_hi_10 = {_memRequest_bits_data_T_3205[2], _memRequest_bits_data_T_2820[2]};
  wire [3:0]        memRequest_bits_data_lo_10 = {memRequest_bits_data_lo_hi_10, memRequest_bits_data_lo_lo_10};
  wire [1:0]        memRequest_bits_data_hi_lo_10 = {_memRequest_bits_data_T_3975[2], _memRequest_bits_data_T_3590[2]};
  wire [1:0]        memRequest_bits_data_hi_hi_10 = {_memRequest_bits_data_T_4745[2], _memRequest_bits_data_T_4360[2]};
  wire [3:0]        memRequest_bits_data_hi_10 = {memRequest_bits_data_hi_hi_10, memRequest_bits_data_hi_lo_10};
  wire [1:0]        memRequest_bits_data_lo_lo_11 = {_memRequest_bits_data_T_2435[3], _memRequest_bits_data_T_2050[3]};
  wire [1:0]        memRequest_bits_data_lo_hi_11 = {_memRequest_bits_data_T_3205[3], _memRequest_bits_data_T_2820[3]};
  wire [3:0]        memRequest_bits_data_lo_11 = {memRequest_bits_data_lo_hi_11, memRequest_bits_data_lo_lo_11};
  wire [1:0]        memRequest_bits_data_hi_lo_11 = {_memRequest_bits_data_T_3975[3], _memRequest_bits_data_T_3590[3]};
  wire [1:0]        memRequest_bits_data_hi_hi_11 = {_memRequest_bits_data_T_4745[3], _memRequest_bits_data_T_4360[3]};
  wire [3:0]        memRequest_bits_data_hi_11 = {memRequest_bits_data_hi_hi_11, memRequest_bits_data_hi_lo_11};
  wire [1:0]        memRequest_bits_data_lo_lo_12 = {_memRequest_bits_data_T_2435[4], _memRequest_bits_data_T_2050[4]};
  wire [1:0]        memRequest_bits_data_lo_hi_12 = {_memRequest_bits_data_T_3205[4], _memRequest_bits_data_T_2820[4]};
  wire [3:0]        memRequest_bits_data_lo_12 = {memRequest_bits_data_lo_hi_12, memRequest_bits_data_lo_lo_12};
  wire [1:0]        memRequest_bits_data_hi_lo_12 = {_memRequest_bits_data_T_3975[4], _memRequest_bits_data_T_3590[4]};
  wire [1:0]        memRequest_bits_data_hi_hi_12 = {_memRequest_bits_data_T_4745[4], _memRequest_bits_data_T_4360[4]};
  wire [3:0]        memRequest_bits_data_hi_12 = {memRequest_bits_data_hi_hi_12, memRequest_bits_data_hi_lo_12};
  wire [1:0]        memRequest_bits_data_lo_lo_13 = {_memRequest_bits_data_T_2435[5], _memRequest_bits_data_T_2050[5]};
  wire [1:0]        memRequest_bits_data_lo_hi_13 = {_memRequest_bits_data_T_3205[5], _memRequest_bits_data_T_2820[5]};
  wire [3:0]        memRequest_bits_data_lo_13 = {memRequest_bits_data_lo_hi_13, memRequest_bits_data_lo_lo_13};
  wire [1:0]        memRequest_bits_data_hi_lo_13 = {_memRequest_bits_data_T_3975[5], _memRequest_bits_data_T_3590[5]};
  wire [1:0]        memRequest_bits_data_hi_hi_13 = {_memRequest_bits_data_T_4745[5], _memRequest_bits_data_T_4360[5]};
  wire [3:0]        memRequest_bits_data_hi_13 = {memRequest_bits_data_hi_hi_13, memRequest_bits_data_hi_lo_13};
  wire [1:0]        memRequest_bits_data_lo_lo_14 = {_memRequest_bits_data_T_2435[6], _memRequest_bits_data_T_2050[6]};
  wire [1:0]        memRequest_bits_data_lo_hi_14 = {_memRequest_bits_data_T_3205[6], _memRequest_bits_data_T_2820[6]};
  wire [3:0]        memRequest_bits_data_lo_14 = {memRequest_bits_data_lo_hi_14, memRequest_bits_data_lo_lo_14};
  wire [1:0]        memRequest_bits_data_hi_lo_14 = {_memRequest_bits_data_T_3975[6], _memRequest_bits_data_T_3590[6]};
  wire [1:0]        memRequest_bits_data_hi_hi_14 = {_memRequest_bits_data_T_4745[6], _memRequest_bits_data_T_4360[6]};
  wire [3:0]        memRequest_bits_data_hi_14 = {memRequest_bits_data_hi_hi_14, memRequest_bits_data_hi_lo_14};
  wire [1:0]        memRequest_bits_data_lo_lo_15 = {_memRequest_bits_data_T_2435[7], _memRequest_bits_data_T_2050[7]};
  wire [1:0]        memRequest_bits_data_lo_hi_15 = {_memRequest_bits_data_T_3205[7], _memRequest_bits_data_T_2820[7]};
  wire [3:0]        memRequest_bits_data_lo_15 = {memRequest_bits_data_lo_hi_15, memRequest_bits_data_lo_lo_15};
  wire [1:0]        memRequest_bits_data_hi_lo_15 = {_memRequest_bits_data_T_3975[7], _memRequest_bits_data_T_3590[7]};
  wire [1:0]        memRequest_bits_data_hi_hi_15 = {_memRequest_bits_data_T_4745[7], _memRequest_bits_data_T_4360[7]};
  wire [3:0]        memRequest_bits_data_hi_15 = {memRequest_bits_data_hi_hi_15, memRequest_bits_data_hi_lo_15};
  wire [1:0]        memRequest_bits_data_lo_lo_16 = {_memRequest_bits_data_T_2435[8], _memRequest_bits_data_T_2050[8]};
  wire [1:0]        memRequest_bits_data_lo_hi_16 = {_memRequest_bits_data_T_3205[8], _memRequest_bits_data_T_2820[8]};
  wire [3:0]        memRequest_bits_data_lo_16 = {memRequest_bits_data_lo_hi_16, memRequest_bits_data_lo_lo_16};
  wire [1:0]        memRequest_bits_data_hi_lo_16 = {_memRequest_bits_data_T_3975[8], _memRequest_bits_data_T_3590[8]};
  wire [1:0]        memRequest_bits_data_hi_hi_16 = {_memRequest_bits_data_T_4745[8], _memRequest_bits_data_T_4360[8]};
  wire [3:0]        memRequest_bits_data_hi_16 = {memRequest_bits_data_hi_hi_16, memRequest_bits_data_hi_lo_16};
  wire [1:0]        memRequest_bits_data_lo_lo_17 = {_memRequest_bits_data_T_2435[9], _memRequest_bits_data_T_2050[9]};
  wire [1:0]        memRequest_bits_data_lo_hi_17 = {_memRequest_bits_data_T_3205[9], _memRequest_bits_data_T_2820[9]};
  wire [3:0]        memRequest_bits_data_lo_17 = {memRequest_bits_data_lo_hi_17, memRequest_bits_data_lo_lo_17};
  wire [1:0]        memRequest_bits_data_hi_lo_17 = {_memRequest_bits_data_T_3975[9], _memRequest_bits_data_T_3590[9]};
  wire [1:0]        memRequest_bits_data_hi_hi_17 = {_memRequest_bits_data_T_4745[9], _memRequest_bits_data_T_4360[9]};
  wire [3:0]        memRequest_bits_data_hi_17 = {memRequest_bits_data_hi_hi_17, memRequest_bits_data_hi_lo_17};
  wire [1:0]        memRequest_bits_data_lo_lo_18 = {_memRequest_bits_data_T_2435[10], _memRequest_bits_data_T_2050[10]};
  wire [1:0]        memRequest_bits_data_lo_hi_18 = {_memRequest_bits_data_T_3205[10], _memRequest_bits_data_T_2820[10]};
  wire [3:0]        memRequest_bits_data_lo_18 = {memRequest_bits_data_lo_hi_18, memRequest_bits_data_lo_lo_18};
  wire [1:0]        memRequest_bits_data_hi_lo_18 = {_memRequest_bits_data_T_3975[10], _memRequest_bits_data_T_3590[10]};
  wire [1:0]        memRequest_bits_data_hi_hi_18 = {_memRequest_bits_data_T_4745[10], _memRequest_bits_data_T_4360[10]};
  wire [3:0]        memRequest_bits_data_hi_18 = {memRequest_bits_data_hi_hi_18, memRequest_bits_data_hi_lo_18};
  wire [1:0]        memRequest_bits_data_lo_lo_19 = {_memRequest_bits_data_T_2435[11], _memRequest_bits_data_T_2050[11]};
  wire [1:0]        memRequest_bits_data_lo_hi_19 = {_memRequest_bits_data_T_3205[11], _memRequest_bits_data_T_2820[11]};
  wire [3:0]        memRequest_bits_data_lo_19 = {memRequest_bits_data_lo_hi_19, memRequest_bits_data_lo_lo_19};
  wire [1:0]        memRequest_bits_data_hi_lo_19 = {_memRequest_bits_data_T_3975[11], _memRequest_bits_data_T_3590[11]};
  wire [1:0]        memRequest_bits_data_hi_hi_19 = {_memRequest_bits_data_T_4745[11], _memRequest_bits_data_T_4360[11]};
  wire [3:0]        memRequest_bits_data_hi_19 = {memRequest_bits_data_hi_hi_19, memRequest_bits_data_hi_lo_19};
  wire [1:0]        memRequest_bits_data_lo_lo_20 = {_memRequest_bits_data_T_2435[12], _memRequest_bits_data_T_2050[12]};
  wire [1:0]        memRequest_bits_data_lo_hi_20 = {_memRequest_bits_data_T_3205[12], _memRequest_bits_data_T_2820[12]};
  wire [3:0]        memRequest_bits_data_lo_20 = {memRequest_bits_data_lo_hi_20, memRequest_bits_data_lo_lo_20};
  wire [1:0]        memRequest_bits_data_hi_lo_20 = {_memRequest_bits_data_T_3975[12], _memRequest_bits_data_T_3590[12]};
  wire [1:0]        memRequest_bits_data_hi_hi_20 = {_memRequest_bits_data_T_4745[12], _memRequest_bits_data_T_4360[12]};
  wire [3:0]        memRequest_bits_data_hi_20 = {memRequest_bits_data_hi_hi_20, memRequest_bits_data_hi_lo_20};
  wire [1:0]        memRequest_bits_data_lo_lo_21 = {_memRequest_bits_data_T_2435[13], _memRequest_bits_data_T_2050[13]};
  wire [1:0]        memRequest_bits_data_lo_hi_21 = {_memRequest_bits_data_T_3205[13], _memRequest_bits_data_T_2820[13]};
  wire [3:0]        memRequest_bits_data_lo_21 = {memRequest_bits_data_lo_hi_21, memRequest_bits_data_lo_lo_21};
  wire [1:0]        memRequest_bits_data_hi_lo_21 = {_memRequest_bits_data_T_3975[13], _memRequest_bits_data_T_3590[13]};
  wire [1:0]        memRequest_bits_data_hi_hi_21 = {_memRequest_bits_data_T_4745[13], _memRequest_bits_data_T_4360[13]};
  wire [3:0]        memRequest_bits_data_hi_21 = {memRequest_bits_data_hi_hi_21, memRequest_bits_data_hi_lo_21};
  wire [1:0]        memRequest_bits_data_lo_lo_22 = {_memRequest_bits_data_T_2435[14], _memRequest_bits_data_T_2050[14]};
  wire [1:0]        memRequest_bits_data_lo_hi_22 = {_memRequest_bits_data_T_3205[14], _memRequest_bits_data_T_2820[14]};
  wire [3:0]        memRequest_bits_data_lo_22 = {memRequest_bits_data_lo_hi_22, memRequest_bits_data_lo_lo_22};
  wire [1:0]        memRequest_bits_data_hi_lo_22 = {_memRequest_bits_data_T_3975[14], _memRequest_bits_data_T_3590[14]};
  wire [1:0]        memRequest_bits_data_hi_hi_22 = {_memRequest_bits_data_T_4745[14], _memRequest_bits_data_T_4360[14]};
  wire [3:0]        memRequest_bits_data_hi_22 = {memRequest_bits_data_hi_hi_22, memRequest_bits_data_hi_lo_22};
  wire [1:0]        memRequest_bits_data_lo_lo_23 = {_memRequest_bits_data_T_2435[15], _memRequest_bits_data_T_2050[15]};
  wire [1:0]        memRequest_bits_data_lo_hi_23 = {_memRequest_bits_data_T_3205[15], _memRequest_bits_data_T_2820[15]};
  wire [3:0]        memRequest_bits_data_lo_23 = {memRequest_bits_data_lo_hi_23, memRequest_bits_data_lo_lo_23};
  wire [1:0]        memRequest_bits_data_hi_lo_23 = {_memRequest_bits_data_T_3975[15], _memRequest_bits_data_T_3590[15]};
  wire [1:0]        memRequest_bits_data_hi_hi_23 = {_memRequest_bits_data_T_4745[15], _memRequest_bits_data_T_4360[15]};
  wire [3:0]        memRequest_bits_data_hi_23 = {memRequest_bits_data_hi_hi_23, memRequest_bits_data_hi_lo_23};
  wire [1:0]        memRequest_bits_data_lo_lo_24 = {_memRequest_bits_data_T_2435[16], _memRequest_bits_data_T_2050[16]};
  wire [1:0]        memRequest_bits_data_lo_hi_24 = {_memRequest_bits_data_T_3205[16], _memRequest_bits_data_T_2820[16]};
  wire [3:0]        memRequest_bits_data_lo_24 = {memRequest_bits_data_lo_hi_24, memRequest_bits_data_lo_lo_24};
  wire [1:0]        memRequest_bits_data_hi_lo_24 = {_memRequest_bits_data_T_3975[16], _memRequest_bits_data_T_3590[16]};
  wire [1:0]        memRequest_bits_data_hi_hi_24 = {_memRequest_bits_data_T_4745[16], _memRequest_bits_data_T_4360[16]};
  wire [3:0]        memRequest_bits_data_hi_24 = {memRequest_bits_data_hi_hi_24, memRequest_bits_data_hi_lo_24};
  wire [1:0]        memRequest_bits_data_lo_lo_25 = {_memRequest_bits_data_T_2435[17], _memRequest_bits_data_T_2050[17]};
  wire [1:0]        memRequest_bits_data_lo_hi_25 = {_memRequest_bits_data_T_3205[17], _memRequest_bits_data_T_2820[17]};
  wire [3:0]        memRequest_bits_data_lo_25 = {memRequest_bits_data_lo_hi_25, memRequest_bits_data_lo_lo_25};
  wire [1:0]        memRequest_bits_data_hi_lo_25 = {_memRequest_bits_data_T_3975[17], _memRequest_bits_data_T_3590[17]};
  wire [1:0]        memRequest_bits_data_hi_hi_25 = {_memRequest_bits_data_T_4745[17], _memRequest_bits_data_T_4360[17]};
  wire [3:0]        memRequest_bits_data_hi_25 = {memRequest_bits_data_hi_hi_25, memRequest_bits_data_hi_lo_25};
  wire [1:0]        memRequest_bits_data_lo_lo_26 = {_memRequest_bits_data_T_2435[18], _memRequest_bits_data_T_2050[18]};
  wire [1:0]        memRequest_bits_data_lo_hi_26 = {_memRequest_bits_data_T_3205[18], _memRequest_bits_data_T_2820[18]};
  wire [3:0]        memRequest_bits_data_lo_26 = {memRequest_bits_data_lo_hi_26, memRequest_bits_data_lo_lo_26};
  wire [1:0]        memRequest_bits_data_hi_lo_26 = {_memRequest_bits_data_T_3975[18], _memRequest_bits_data_T_3590[18]};
  wire [1:0]        memRequest_bits_data_hi_hi_26 = {_memRequest_bits_data_T_4745[18], _memRequest_bits_data_T_4360[18]};
  wire [3:0]        memRequest_bits_data_hi_26 = {memRequest_bits_data_hi_hi_26, memRequest_bits_data_hi_lo_26};
  wire [1:0]        memRequest_bits_data_lo_lo_27 = {_memRequest_bits_data_T_2435[19], _memRequest_bits_data_T_2050[19]};
  wire [1:0]        memRequest_bits_data_lo_hi_27 = {_memRequest_bits_data_T_3205[19], _memRequest_bits_data_T_2820[19]};
  wire [3:0]        memRequest_bits_data_lo_27 = {memRequest_bits_data_lo_hi_27, memRequest_bits_data_lo_lo_27};
  wire [1:0]        memRequest_bits_data_hi_lo_27 = {_memRequest_bits_data_T_3975[19], _memRequest_bits_data_T_3590[19]};
  wire [1:0]        memRequest_bits_data_hi_hi_27 = {_memRequest_bits_data_T_4745[19], _memRequest_bits_data_T_4360[19]};
  wire [3:0]        memRequest_bits_data_hi_27 = {memRequest_bits_data_hi_hi_27, memRequest_bits_data_hi_lo_27};
  wire [1:0]        memRequest_bits_data_lo_lo_28 = {_memRequest_bits_data_T_2435[20], _memRequest_bits_data_T_2050[20]};
  wire [1:0]        memRequest_bits_data_lo_hi_28 = {_memRequest_bits_data_T_3205[20], _memRequest_bits_data_T_2820[20]};
  wire [3:0]        memRequest_bits_data_lo_28 = {memRequest_bits_data_lo_hi_28, memRequest_bits_data_lo_lo_28};
  wire [1:0]        memRequest_bits_data_hi_lo_28 = {_memRequest_bits_data_T_3975[20], _memRequest_bits_data_T_3590[20]};
  wire [1:0]        memRequest_bits_data_hi_hi_28 = {_memRequest_bits_data_T_4745[20], _memRequest_bits_data_T_4360[20]};
  wire [3:0]        memRequest_bits_data_hi_28 = {memRequest_bits_data_hi_hi_28, memRequest_bits_data_hi_lo_28};
  wire [1:0]        memRequest_bits_data_lo_lo_29 = {_memRequest_bits_data_T_2435[21], _memRequest_bits_data_T_2050[21]};
  wire [1:0]        memRequest_bits_data_lo_hi_29 = {_memRequest_bits_data_T_3205[21], _memRequest_bits_data_T_2820[21]};
  wire [3:0]        memRequest_bits_data_lo_29 = {memRequest_bits_data_lo_hi_29, memRequest_bits_data_lo_lo_29};
  wire [1:0]        memRequest_bits_data_hi_lo_29 = {_memRequest_bits_data_T_3975[21], _memRequest_bits_data_T_3590[21]};
  wire [1:0]        memRequest_bits_data_hi_hi_29 = {_memRequest_bits_data_T_4745[21], _memRequest_bits_data_T_4360[21]};
  wire [3:0]        memRequest_bits_data_hi_29 = {memRequest_bits_data_hi_hi_29, memRequest_bits_data_hi_lo_29};
  wire [1:0]        memRequest_bits_data_lo_lo_30 = {_memRequest_bits_data_T_2435[22], _memRequest_bits_data_T_2050[22]};
  wire [1:0]        memRequest_bits_data_lo_hi_30 = {_memRequest_bits_data_T_3205[22], _memRequest_bits_data_T_2820[22]};
  wire [3:0]        memRequest_bits_data_lo_30 = {memRequest_bits_data_lo_hi_30, memRequest_bits_data_lo_lo_30};
  wire [1:0]        memRequest_bits_data_hi_lo_30 = {_memRequest_bits_data_T_3975[22], _memRequest_bits_data_T_3590[22]};
  wire [1:0]        memRequest_bits_data_hi_hi_30 = {_memRequest_bits_data_T_4745[22], _memRequest_bits_data_T_4360[22]};
  wire [3:0]        memRequest_bits_data_hi_30 = {memRequest_bits_data_hi_hi_30, memRequest_bits_data_hi_lo_30};
  wire [1:0]        memRequest_bits_data_lo_lo_31 = {_memRequest_bits_data_T_2435[23], _memRequest_bits_data_T_2050[23]};
  wire [1:0]        memRequest_bits_data_lo_hi_31 = {_memRequest_bits_data_T_3205[23], _memRequest_bits_data_T_2820[23]};
  wire [3:0]        memRequest_bits_data_lo_31 = {memRequest_bits_data_lo_hi_31, memRequest_bits_data_lo_lo_31};
  wire [1:0]        memRequest_bits_data_hi_lo_31 = {_memRequest_bits_data_T_3975[23], _memRequest_bits_data_T_3590[23]};
  wire [1:0]        memRequest_bits_data_hi_hi_31 = {_memRequest_bits_data_T_4745[23], _memRequest_bits_data_T_4360[23]};
  wire [3:0]        memRequest_bits_data_hi_31 = {memRequest_bits_data_hi_hi_31, memRequest_bits_data_hi_lo_31};
  wire [1:0]        memRequest_bits_data_lo_lo_32 = {_memRequest_bits_data_T_2435[24], _memRequest_bits_data_T_2050[24]};
  wire [1:0]        memRequest_bits_data_lo_hi_32 = {_memRequest_bits_data_T_3205[24], _memRequest_bits_data_T_2820[24]};
  wire [3:0]        memRequest_bits_data_lo_32 = {memRequest_bits_data_lo_hi_32, memRequest_bits_data_lo_lo_32};
  wire [1:0]        memRequest_bits_data_hi_lo_32 = {_memRequest_bits_data_T_3975[24], _memRequest_bits_data_T_3590[24]};
  wire [1:0]        memRequest_bits_data_hi_hi_32 = {_memRequest_bits_data_T_4745[24], _memRequest_bits_data_T_4360[24]};
  wire [3:0]        memRequest_bits_data_hi_32 = {memRequest_bits_data_hi_hi_32, memRequest_bits_data_hi_lo_32};
  wire [1:0]        memRequest_bits_data_lo_lo_33 = {_memRequest_bits_data_T_2435[25], _memRequest_bits_data_T_2050[25]};
  wire [1:0]        memRequest_bits_data_lo_hi_33 = {_memRequest_bits_data_T_3205[25], _memRequest_bits_data_T_2820[25]};
  wire [3:0]        memRequest_bits_data_lo_33 = {memRequest_bits_data_lo_hi_33, memRequest_bits_data_lo_lo_33};
  wire [1:0]        memRequest_bits_data_hi_lo_33 = {_memRequest_bits_data_T_3975[25], _memRequest_bits_data_T_3590[25]};
  wire [1:0]        memRequest_bits_data_hi_hi_33 = {_memRequest_bits_data_T_4745[25], _memRequest_bits_data_T_4360[25]};
  wire [3:0]        memRequest_bits_data_hi_33 = {memRequest_bits_data_hi_hi_33, memRequest_bits_data_hi_lo_33};
  wire [1:0]        memRequest_bits_data_lo_lo_34 = {_memRequest_bits_data_T_2435[26], _memRequest_bits_data_T_2050[26]};
  wire [1:0]        memRequest_bits_data_lo_hi_34 = {_memRequest_bits_data_T_3205[26], _memRequest_bits_data_T_2820[26]};
  wire [3:0]        memRequest_bits_data_lo_34 = {memRequest_bits_data_lo_hi_34, memRequest_bits_data_lo_lo_34};
  wire [1:0]        memRequest_bits_data_hi_lo_34 = {_memRequest_bits_data_T_3975[26], _memRequest_bits_data_T_3590[26]};
  wire [1:0]        memRequest_bits_data_hi_hi_34 = {_memRequest_bits_data_T_4745[26], _memRequest_bits_data_T_4360[26]};
  wire [3:0]        memRequest_bits_data_hi_34 = {memRequest_bits_data_hi_hi_34, memRequest_bits_data_hi_lo_34};
  wire [1:0]        memRequest_bits_data_lo_lo_35 = {_memRequest_bits_data_T_2435[27], _memRequest_bits_data_T_2050[27]};
  wire [1:0]        memRequest_bits_data_lo_hi_35 = {_memRequest_bits_data_T_3205[27], _memRequest_bits_data_T_2820[27]};
  wire [3:0]        memRequest_bits_data_lo_35 = {memRequest_bits_data_lo_hi_35, memRequest_bits_data_lo_lo_35};
  wire [1:0]        memRequest_bits_data_hi_lo_35 = {_memRequest_bits_data_T_3975[27], _memRequest_bits_data_T_3590[27]};
  wire [1:0]        memRequest_bits_data_hi_hi_35 = {_memRequest_bits_data_T_4745[27], _memRequest_bits_data_T_4360[27]};
  wire [3:0]        memRequest_bits_data_hi_35 = {memRequest_bits_data_hi_hi_35, memRequest_bits_data_hi_lo_35};
  wire [1:0]        memRequest_bits_data_lo_lo_36 = {_memRequest_bits_data_T_2435[28], _memRequest_bits_data_T_2050[28]};
  wire [1:0]        memRequest_bits_data_lo_hi_36 = {_memRequest_bits_data_T_3205[28], _memRequest_bits_data_T_2820[28]};
  wire [3:0]        memRequest_bits_data_lo_36 = {memRequest_bits_data_lo_hi_36, memRequest_bits_data_lo_lo_36};
  wire [1:0]        memRequest_bits_data_hi_lo_36 = {_memRequest_bits_data_T_3975[28], _memRequest_bits_data_T_3590[28]};
  wire [1:0]        memRequest_bits_data_hi_hi_36 = {_memRequest_bits_data_T_4745[28], _memRequest_bits_data_T_4360[28]};
  wire [3:0]        memRequest_bits_data_hi_36 = {memRequest_bits_data_hi_hi_36, memRequest_bits_data_hi_lo_36};
  wire [1:0]        memRequest_bits_data_lo_lo_37 = {_memRequest_bits_data_T_2435[29], _memRequest_bits_data_T_2050[29]};
  wire [1:0]        memRequest_bits_data_lo_hi_37 = {_memRequest_bits_data_T_3205[29], _memRequest_bits_data_T_2820[29]};
  wire [3:0]        memRequest_bits_data_lo_37 = {memRequest_bits_data_lo_hi_37, memRequest_bits_data_lo_lo_37};
  wire [1:0]        memRequest_bits_data_hi_lo_37 = {_memRequest_bits_data_T_3975[29], _memRequest_bits_data_T_3590[29]};
  wire [1:0]        memRequest_bits_data_hi_hi_37 = {_memRequest_bits_data_T_4745[29], _memRequest_bits_data_T_4360[29]};
  wire [3:0]        memRequest_bits_data_hi_37 = {memRequest_bits_data_hi_hi_37, memRequest_bits_data_hi_lo_37};
  wire [1:0]        memRequest_bits_data_lo_lo_38 = {_memRequest_bits_data_T_2435[30], _memRequest_bits_data_T_2050[30]};
  wire [1:0]        memRequest_bits_data_lo_hi_38 = {_memRequest_bits_data_T_3205[30], _memRequest_bits_data_T_2820[30]};
  wire [3:0]        memRequest_bits_data_lo_38 = {memRequest_bits_data_lo_hi_38, memRequest_bits_data_lo_lo_38};
  wire [1:0]        memRequest_bits_data_hi_lo_38 = {_memRequest_bits_data_T_3975[30], _memRequest_bits_data_T_3590[30]};
  wire [1:0]        memRequest_bits_data_hi_hi_38 = {_memRequest_bits_data_T_4745[30], _memRequest_bits_data_T_4360[30]};
  wire [3:0]        memRequest_bits_data_hi_38 = {memRequest_bits_data_hi_hi_38, memRequest_bits_data_hi_lo_38};
  wire [1:0]        memRequest_bits_data_lo_lo_39 = {_memRequest_bits_data_T_2435[31], _memRequest_bits_data_T_2050[31]};
  wire [1:0]        memRequest_bits_data_lo_hi_39 = {_memRequest_bits_data_T_3205[31], _memRequest_bits_data_T_2820[31]};
  wire [3:0]        memRequest_bits_data_lo_39 = {memRequest_bits_data_lo_hi_39, memRequest_bits_data_lo_lo_39};
  wire [1:0]        memRequest_bits_data_hi_lo_39 = {_memRequest_bits_data_T_3975[31], _memRequest_bits_data_T_3590[31]};
  wire [1:0]        memRequest_bits_data_hi_hi_39 = {_memRequest_bits_data_T_4745[31], _memRequest_bits_data_T_4360[31]};
  wire [3:0]        memRequest_bits_data_hi_39 = {memRequest_bits_data_hi_hi_39, memRequest_bits_data_hi_lo_39};
  wire [1:0]        memRequest_bits_data_lo_lo_40 = {_memRequest_bits_data_T_2435[32], _memRequest_bits_data_T_2050[32]};
  wire [1:0]        memRequest_bits_data_lo_hi_40 = {_memRequest_bits_data_T_3205[32], _memRequest_bits_data_T_2820[32]};
  wire [3:0]        memRequest_bits_data_lo_40 = {memRequest_bits_data_lo_hi_40, memRequest_bits_data_lo_lo_40};
  wire [1:0]        memRequest_bits_data_hi_lo_40 = {_memRequest_bits_data_T_3975[32], _memRequest_bits_data_T_3590[32]};
  wire [1:0]        memRequest_bits_data_hi_hi_40 = {_memRequest_bits_data_T_4745[32], _memRequest_bits_data_T_4360[32]};
  wire [3:0]        memRequest_bits_data_hi_40 = {memRequest_bits_data_hi_hi_40, memRequest_bits_data_hi_lo_40};
  wire [1:0]        memRequest_bits_data_lo_lo_41 = {_memRequest_bits_data_T_2435[33], _memRequest_bits_data_T_2050[33]};
  wire [1:0]        memRequest_bits_data_lo_hi_41 = {_memRequest_bits_data_T_3205[33], _memRequest_bits_data_T_2820[33]};
  wire [3:0]        memRequest_bits_data_lo_41 = {memRequest_bits_data_lo_hi_41, memRequest_bits_data_lo_lo_41};
  wire [1:0]        memRequest_bits_data_hi_lo_41 = {_memRequest_bits_data_T_3975[33], _memRequest_bits_data_T_3590[33]};
  wire [1:0]        memRequest_bits_data_hi_hi_41 = {_memRequest_bits_data_T_4745[33], _memRequest_bits_data_T_4360[33]};
  wire [3:0]        memRequest_bits_data_hi_41 = {memRequest_bits_data_hi_hi_41, memRequest_bits_data_hi_lo_41};
  wire [1:0]        memRequest_bits_data_lo_lo_42 = {_memRequest_bits_data_T_2435[34], _memRequest_bits_data_T_2050[34]};
  wire [1:0]        memRequest_bits_data_lo_hi_42 = {_memRequest_bits_data_T_3205[34], _memRequest_bits_data_T_2820[34]};
  wire [3:0]        memRequest_bits_data_lo_42 = {memRequest_bits_data_lo_hi_42, memRequest_bits_data_lo_lo_42};
  wire [1:0]        memRequest_bits_data_hi_lo_42 = {_memRequest_bits_data_T_3975[34], _memRequest_bits_data_T_3590[34]};
  wire [1:0]        memRequest_bits_data_hi_hi_42 = {_memRequest_bits_data_T_4745[34], _memRequest_bits_data_T_4360[34]};
  wire [3:0]        memRequest_bits_data_hi_42 = {memRequest_bits_data_hi_hi_42, memRequest_bits_data_hi_lo_42};
  wire [1:0]        memRequest_bits_data_lo_lo_43 = {_memRequest_bits_data_T_2435[35], _memRequest_bits_data_T_2050[35]};
  wire [1:0]        memRequest_bits_data_lo_hi_43 = {_memRequest_bits_data_T_3205[35], _memRequest_bits_data_T_2820[35]};
  wire [3:0]        memRequest_bits_data_lo_43 = {memRequest_bits_data_lo_hi_43, memRequest_bits_data_lo_lo_43};
  wire [1:0]        memRequest_bits_data_hi_lo_43 = {_memRequest_bits_data_T_3975[35], _memRequest_bits_data_T_3590[35]};
  wire [1:0]        memRequest_bits_data_hi_hi_43 = {_memRequest_bits_data_T_4745[35], _memRequest_bits_data_T_4360[35]};
  wire [3:0]        memRequest_bits_data_hi_43 = {memRequest_bits_data_hi_hi_43, memRequest_bits_data_hi_lo_43};
  wire [1:0]        memRequest_bits_data_lo_lo_44 = {_memRequest_bits_data_T_2435[36], _memRequest_bits_data_T_2050[36]};
  wire [1:0]        memRequest_bits_data_lo_hi_44 = {_memRequest_bits_data_T_3205[36], _memRequest_bits_data_T_2820[36]};
  wire [3:0]        memRequest_bits_data_lo_44 = {memRequest_bits_data_lo_hi_44, memRequest_bits_data_lo_lo_44};
  wire [1:0]        memRequest_bits_data_hi_lo_44 = {_memRequest_bits_data_T_3975[36], _memRequest_bits_data_T_3590[36]};
  wire [1:0]        memRequest_bits_data_hi_hi_44 = {_memRequest_bits_data_T_4745[36], _memRequest_bits_data_T_4360[36]};
  wire [3:0]        memRequest_bits_data_hi_44 = {memRequest_bits_data_hi_hi_44, memRequest_bits_data_hi_lo_44};
  wire [1:0]        memRequest_bits_data_lo_lo_45 = {_memRequest_bits_data_T_2435[37], _memRequest_bits_data_T_2050[37]};
  wire [1:0]        memRequest_bits_data_lo_hi_45 = {_memRequest_bits_data_T_3205[37], _memRequest_bits_data_T_2820[37]};
  wire [3:0]        memRequest_bits_data_lo_45 = {memRequest_bits_data_lo_hi_45, memRequest_bits_data_lo_lo_45};
  wire [1:0]        memRequest_bits_data_hi_lo_45 = {_memRequest_bits_data_T_3975[37], _memRequest_bits_data_T_3590[37]};
  wire [1:0]        memRequest_bits_data_hi_hi_45 = {_memRequest_bits_data_T_4745[37], _memRequest_bits_data_T_4360[37]};
  wire [3:0]        memRequest_bits_data_hi_45 = {memRequest_bits_data_hi_hi_45, memRequest_bits_data_hi_lo_45};
  wire [1:0]        memRequest_bits_data_lo_lo_46 = {_memRequest_bits_data_T_2435[38], _memRequest_bits_data_T_2050[38]};
  wire [1:0]        memRequest_bits_data_lo_hi_46 = {_memRequest_bits_data_T_3205[38], _memRequest_bits_data_T_2820[38]};
  wire [3:0]        memRequest_bits_data_lo_46 = {memRequest_bits_data_lo_hi_46, memRequest_bits_data_lo_lo_46};
  wire [1:0]        memRequest_bits_data_hi_lo_46 = {_memRequest_bits_data_T_3975[38], _memRequest_bits_data_T_3590[38]};
  wire [1:0]        memRequest_bits_data_hi_hi_46 = {_memRequest_bits_data_T_4745[38], _memRequest_bits_data_T_4360[38]};
  wire [3:0]        memRequest_bits_data_hi_46 = {memRequest_bits_data_hi_hi_46, memRequest_bits_data_hi_lo_46};
  wire [1:0]        memRequest_bits_data_lo_lo_47 = {_memRequest_bits_data_T_2435[39], _memRequest_bits_data_T_2050[39]};
  wire [1:0]        memRequest_bits_data_lo_hi_47 = {_memRequest_bits_data_T_3205[39], _memRequest_bits_data_T_2820[39]};
  wire [3:0]        memRequest_bits_data_lo_47 = {memRequest_bits_data_lo_hi_47, memRequest_bits_data_lo_lo_47};
  wire [1:0]        memRequest_bits_data_hi_lo_47 = {_memRequest_bits_data_T_3975[39], _memRequest_bits_data_T_3590[39]};
  wire [1:0]        memRequest_bits_data_hi_hi_47 = {_memRequest_bits_data_T_4745[39], _memRequest_bits_data_T_4360[39]};
  wire [3:0]        memRequest_bits_data_hi_47 = {memRequest_bits_data_hi_hi_47, memRequest_bits_data_hi_lo_47};
  wire [1:0]        memRequest_bits_data_lo_lo_48 = {_memRequest_bits_data_T_2435[40], _memRequest_bits_data_T_2050[40]};
  wire [1:0]        memRequest_bits_data_lo_hi_48 = {_memRequest_bits_data_T_3205[40], _memRequest_bits_data_T_2820[40]};
  wire [3:0]        memRequest_bits_data_lo_48 = {memRequest_bits_data_lo_hi_48, memRequest_bits_data_lo_lo_48};
  wire [1:0]        memRequest_bits_data_hi_lo_48 = {_memRequest_bits_data_T_3975[40], _memRequest_bits_data_T_3590[40]};
  wire [1:0]        memRequest_bits_data_hi_hi_48 = {_memRequest_bits_data_T_4745[40], _memRequest_bits_data_T_4360[40]};
  wire [3:0]        memRequest_bits_data_hi_48 = {memRequest_bits_data_hi_hi_48, memRequest_bits_data_hi_lo_48};
  wire [1:0]        memRequest_bits_data_lo_lo_49 = {_memRequest_bits_data_T_2435[41], _memRequest_bits_data_T_2050[41]};
  wire [1:0]        memRequest_bits_data_lo_hi_49 = {_memRequest_bits_data_T_3205[41], _memRequest_bits_data_T_2820[41]};
  wire [3:0]        memRequest_bits_data_lo_49 = {memRequest_bits_data_lo_hi_49, memRequest_bits_data_lo_lo_49};
  wire [1:0]        memRequest_bits_data_hi_lo_49 = {_memRequest_bits_data_T_3975[41], _memRequest_bits_data_T_3590[41]};
  wire [1:0]        memRequest_bits_data_hi_hi_49 = {_memRequest_bits_data_T_4745[41], _memRequest_bits_data_T_4360[41]};
  wire [3:0]        memRequest_bits_data_hi_49 = {memRequest_bits_data_hi_hi_49, memRequest_bits_data_hi_lo_49};
  wire [1:0]        memRequest_bits_data_lo_lo_50 = {_memRequest_bits_data_T_2435[42], _memRequest_bits_data_T_2050[42]};
  wire [1:0]        memRequest_bits_data_lo_hi_50 = {_memRequest_bits_data_T_3205[42], _memRequest_bits_data_T_2820[42]};
  wire [3:0]        memRequest_bits_data_lo_50 = {memRequest_bits_data_lo_hi_50, memRequest_bits_data_lo_lo_50};
  wire [1:0]        memRequest_bits_data_hi_lo_50 = {_memRequest_bits_data_T_3975[42], _memRequest_bits_data_T_3590[42]};
  wire [1:0]        memRequest_bits_data_hi_hi_50 = {_memRequest_bits_data_T_4745[42], _memRequest_bits_data_T_4360[42]};
  wire [3:0]        memRequest_bits_data_hi_50 = {memRequest_bits_data_hi_hi_50, memRequest_bits_data_hi_lo_50};
  wire [1:0]        memRequest_bits_data_lo_lo_51 = {_memRequest_bits_data_T_2435[43], _memRequest_bits_data_T_2050[43]};
  wire [1:0]        memRequest_bits_data_lo_hi_51 = {_memRequest_bits_data_T_3205[43], _memRequest_bits_data_T_2820[43]};
  wire [3:0]        memRequest_bits_data_lo_51 = {memRequest_bits_data_lo_hi_51, memRequest_bits_data_lo_lo_51};
  wire [1:0]        memRequest_bits_data_hi_lo_51 = {_memRequest_bits_data_T_3975[43], _memRequest_bits_data_T_3590[43]};
  wire [1:0]        memRequest_bits_data_hi_hi_51 = {_memRequest_bits_data_T_4745[43], _memRequest_bits_data_T_4360[43]};
  wire [3:0]        memRequest_bits_data_hi_51 = {memRequest_bits_data_hi_hi_51, memRequest_bits_data_hi_lo_51};
  wire [1:0]        memRequest_bits_data_lo_lo_52 = {_memRequest_bits_data_T_2435[44], _memRequest_bits_data_T_2050[44]};
  wire [1:0]        memRequest_bits_data_lo_hi_52 = {_memRequest_bits_data_T_3205[44], _memRequest_bits_data_T_2820[44]};
  wire [3:0]        memRequest_bits_data_lo_52 = {memRequest_bits_data_lo_hi_52, memRequest_bits_data_lo_lo_52};
  wire [1:0]        memRequest_bits_data_hi_lo_52 = {_memRequest_bits_data_T_3975[44], _memRequest_bits_data_T_3590[44]};
  wire [1:0]        memRequest_bits_data_hi_hi_52 = {_memRequest_bits_data_T_4745[44], _memRequest_bits_data_T_4360[44]};
  wire [3:0]        memRequest_bits_data_hi_52 = {memRequest_bits_data_hi_hi_52, memRequest_bits_data_hi_lo_52};
  wire [1:0]        memRequest_bits_data_lo_lo_53 = {_memRequest_bits_data_T_2435[45], _memRequest_bits_data_T_2050[45]};
  wire [1:0]        memRequest_bits_data_lo_hi_53 = {_memRequest_bits_data_T_3205[45], _memRequest_bits_data_T_2820[45]};
  wire [3:0]        memRequest_bits_data_lo_53 = {memRequest_bits_data_lo_hi_53, memRequest_bits_data_lo_lo_53};
  wire [1:0]        memRequest_bits_data_hi_lo_53 = {_memRequest_bits_data_T_3975[45], _memRequest_bits_data_T_3590[45]};
  wire [1:0]        memRequest_bits_data_hi_hi_53 = {_memRequest_bits_data_T_4745[45], _memRequest_bits_data_T_4360[45]};
  wire [3:0]        memRequest_bits_data_hi_53 = {memRequest_bits_data_hi_hi_53, memRequest_bits_data_hi_lo_53};
  wire [1:0]        memRequest_bits_data_lo_lo_54 = {_memRequest_bits_data_T_2435[46], _memRequest_bits_data_T_2050[46]};
  wire [1:0]        memRequest_bits_data_lo_hi_54 = {_memRequest_bits_data_T_3205[46], _memRequest_bits_data_T_2820[46]};
  wire [3:0]        memRequest_bits_data_lo_54 = {memRequest_bits_data_lo_hi_54, memRequest_bits_data_lo_lo_54};
  wire [1:0]        memRequest_bits_data_hi_lo_54 = {_memRequest_bits_data_T_3975[46], _memRequest_bits_data_T_3590[46]};
  wire [1:0]        memRequest_bits_data_hi_hi_54 = {_memRequest_bits_data_T_4745[46], _memRequest_bits_data_T_4360[46]};
  wire [3:0]        memRequest_bits_data_hi_54 = {memRequest_bits_data_hi_hi_54, memRequest_bits_data_hi_lo_54};
  wire [1:0]        memRequest_bits_data_lo_lo_55 = {_memRequest_bits_data_T_2435[47], _memRequest_bits_data_T_2050[47]};
  wire [1:0]        memRequest_bits_data_lo_hi_55 = {_memRequest_bits_data_T_3205[47], _memRequest_bits_data_T_2820[47]};
  wire [3:0]        memRequest_bits_data_lo_55 = {memRequest_bits_data_lo_hi_55, memRequest_bits_data_lo_lo_55};
  wire [1:0]        memRequest_bits_data_hi_lo_55 = {_memRequest_bits_data_T_3975[47], _memRequest_bits_data_T_3590[47]};
  wire [1:0]        memRequest_bits_data_hi_hi_55 = {_memRequest_bits_data_T_4745[47], _memRequest_bits_data_T_4360[47]};
  wire [3:0]        memRequest_bits_data_hi_55 = {memRequest_bits_data_hi_hi_55, memRequest_bits_data_hi_lo_55};
  wire [1:0]        memRequest_bits_data_lo_lo_56 = {_memRequest_bits_data_T_2435[48], _memRequest_bits_data_T_2050[48]};
  wire [1:0]        memRequest_bits_data_lo_hi_56 = {_memRequest_bits_data_T_3205[48], _memRequest_bits_data_T_2820[48]};
  wire [3:0]        memRequest_bits_data_lo_56 = {memRequest_bits_data_lo_hi_56, memRequest_bits_data_lo_lo_56};
  wire [1:0]        memRequest_bits_data_hi_lo_56 = {_memRequest_bits_data_T_3975[48], _memRequest_bits_data_T_3590[48]};
  wire [1:0]        memRequest_bits_data_hi_hi_56 = {_memRequest_bits_data_T_4745[48], _memRequest_bits_data_T_4360[48]};
  wire [3:0]        memRequest_bits_data_hi_56 = {memRequest_bits_data_hi_hi_56, memRequest_bits_data_hi_lo_56};
  wire [1:0]        memRequest_bits_data_lo_lo_57 = {_memRequest_bits_data_T_2435[49], _memRequest_bits_data_T_2050[49]};
  wire [1:0]        memRequest_bits_data_lo_hi_57 = {_memRequest_bits_data_T_3205[49], _memRequest_bits_data_T_2820[49]};
  wire [3:0]        memRequest_bits_data_lo_57 = {memRequest_bits_data_lo_hi_57, memRequest_bits_data_lo_lo_57};
  wire [1:0]        memRequest_bits_data_hi_lo_57 = {_memRequest_bits_data_T_3975[49], _memRequest_bits_data_T_3590[49]};
  wire [1:0]        memRequest_bits_data_hi_hi_57 = {_memRequest_bits_data_T_4745[49], _memRequest_bits_data_T_4360[49]};
  wire [3:0]        memRequest_bits_data_hi_57 = {memRequest_bits_data_hi_hi_57, memRequest_bits_data_hi_lo_57};
  wire [1:0]        memRequest_bits_data_lo_lo_58 = {_memRequest_bits_data_T_2435[50], _memRequest_bits_data_T_2050[50]};
  wire [1:0]        memRequest_bits_data_lo_hi_58 = {_memRequest_bits_data_T_3205[50], _memRequest_bits_data_T_2820[50]};
  wire [3:0]        memRequest_bits_data_lo_58 = {memRequest_bits_data_lo_hi_58, memRequest_bits_data_lo_lo_58};
  wire [1:0]        memRequest_bits_data_hi_lo_58 = {_memRequest_bits_data_T_3975[50], _memRequest_bits_data_T_3590[50]};
  wire [1:0]        memRequest_bits_data_hi_hi_58 = {_memRequest_bits_data_T_4745[50], _memRequest_bits_data_T_4360[50]};
  wire [3:0]        memRequest_bits_data_hi_58 = {memRequest_bits_data_hi_hi_58, memRequest_bits_data_hi_lo_58};
  wire [1:0]        memRequest_bits_data_lo_lo_59 = {_memRequest_bits_data_T_2435[51], _memRequest_bits_data_T_2050[51]};
  wire [1:0]        memRequest_bits_data_lo_hi_59 = {_memRequest_bits_data_T_3205[51], _memRequest_bits_data_T_2820[51]};
  wire [3:0]        memRequest_bits_data_lo_59 = {memRequest_bits_data_lo_hi_59, memRequest_bits_data_lo_lo_59};
  wire [1:0]        memRequest_bits_data_hi_lo_59 = {_memRequest_bits_data_T_3975[51], _memRequest_bits_data_T_3590[51]};
  wire [1:0]        memRequest_bits_data_hi_hi_59 = {_memRequest_bits_data_T_4745[51], _memRequest_bits_data_T_4360[51]};
  wire [3:0]        memRequest_bits_data_hi_59 = {memRequest_bits_data_hi_hi_59, memRequest_bits_data_hi_lo_59};
  wire [1:0]        memRequest_bits_data_lo_lo_60 = {_memRequest_bits_data_T_2435[52], _memRequest_bits_data_T_2050[52]};
  wire [1:0]        memRequest_bits_data_lo_hi_60 = {_memRequest_bits_data_T_3205[52], _memRequest_bits_data_T_2820[52]};
  wire [3:0]        memRequest_bits_data_lo_60 = {memRequest_bits_data_lo_hi_60, memRequest_bits_data_lo_lo_60};
  wire [1:0]        memRequest_bits_data_hi_lo_60 = {_memRequest_bits_data_T_3975[52], _memRequest_bits_data_T_3590[52]};
  wire [1:0]        memRequest_bits_data_hi_hi_60 = {_memRequest_bits_data_T_4745[52], _memRequest_bits_data_T_4360[52]};
  wire [3:0]        memRequest_bits_data_hi_60 = {memRequest_bits_data_hi_hi_60, memRequest_bits_data_hi_lo_60};
  wire [1:0]        memRequest_bits_data_lo_lo_61 = {_memRequest_bits_data_T_2435[53], _memRequest_bits_data_T_2050[53]};
  wire [1:0]        memRequest_bits_data_lo_hi_61 = {_memRequest_bits_data_T_3205[53], _memRequest_bits_data_T_2820[53]};
  wire [3:0]        memRequest_bits_data_lo_61 = {memRequest_bits_data_lo_hi_61, memRequest_bits_data_lo_lo_61};
  wire [1:0]        memRequest_bits_data_hi_lo_61 = {_memRequest_bits_data_T_3975[53], _memRequest_bits_data_T_3590[53]};
  wire [1:0]        memRequest_bits_data_hi_hi_61 = {_memRequest_bits_data_T_4745[53], _memRequest_bits_data_T_4360[53]};
  wire [3:0]        memRequest_bits_data_hi_61 = {memRequest_bits_data_hi_hi_61, memRequest_bits_data_hi_lo_61};
  wire [1:0]        memRequest_bits_data_lo_lo_62 = {_memRequest_bits_data_T_2435[54], _memRequest_bits_data_T_2050[54]};
  wire [1:0]        memRequest_bits_data_lo_hi_62 = {_memRequest_bits_data_T_3205[54], _memRequest_bits_data_T_2820[54]};
  wire [3:0]        memRequest_bits_data_lo_62 = {memRequest_bits_data_lo_hi_62, memRequest_bits_data_lo_lo_62};
  wire [1:0]        memRequest_bits_data_hi_lo_62 = {_memRequest_bits_data_T_3975[54], _memRequest_bits_data_T_3590[54]};
  wire [1:0]        memRequest_bits_data_hi_hi_62 = {_memRequest_bits_data_T_4745[54], _memRequest_bits_data_T_4360[54]};
  wire [3:0]        memRequest_bits_data_hi_62 = {memRequest_bits_data_hi_hi_62, memRequest_bits_data_hi_lo_62};
  wire [1:0]        memRequest_bits_data_lo_lo_63 = {_memRequest_bits_data_T_2435[55], _memRequest_bits_data_T_2050[55]};
  wire [1:0]        memRequest_bits_data_lo_hi_63 = {_memRequest_bits_data_T_3205[55], _memRequest_bits_data_T_2820[55]};
  wire [3:0]        memRequest_bits_data_lo_63 = {memRequest_bits_data_lo_hi_63, memRequest_bits_data_lo_lo_63};
  wire [1:0]        memRequest_bits_data_hi_lo_63 = {_memRequest_bits_data_T_3975[55], _memRequest_bits_data_T_3590[55]};
  wire [1:0]        memRequest_bits_data_hi_hi_63 = {_memRequest_bits_data_T_4745[55], _memRequest_bits_data_T_4360[55]};
  wire [3:0]        memRequest_bits_data_hi_63 = {memRequest_bits_data_hi_hi_63, memRequest_bits_data_hi_lo_63};
  wire [1:0]        memRequest_bits_data_lo_lo_64 = {_memRequest_bits_data_T_2435[56], _memRequest_bits_data_T_2050[56]};
  wire [1:0]        memRequest_bits_data_lo_hi_64 = {_memRequest_bits_data_T_3205[56], _memRequest_bits_data_T_2820[56]};
  wire [3:0]        memRequest_bits_data_lo_64 = {memRequest_bits_data_lo_hi_64, memRequest_bits_data_lo_lo_64};
  wire [1:0]        memRequest_bits_data_hi_lo_64 = {_memRequest_bits_data_T_3975[56], _memRequest_bits_data_T_3590[56]};
  wire [1:0]        memRequest_bits_data_hi_hi_64 = {_memRequest_bits_data_T_4745[56], _memRequest_bits_data_T_4360[56]};
  wire [3:0]        memRequest_bits_data_hi_64 = {memRequest_bits_data_hi_hi_64, memRequest_bits_data_hi_lo_64};
  wire [1:0]        memRequest_bits_data_lo_lo_65 = {_memRequest_bits_data_T_2435[57], _memRequest_bits_data_T_2050[57]};
  wire [1:0]        memRequest_bits_data_lo_hi_65 = {_memRequest_bits_data_T_3205[57], _memRequest_bits_data_T_2820[57]};
  wire [3:0]        memRequest_bits_data_lo_65 = {memRequest_bits_data_lo_hi_65, memRequest_bits_data_lo_lo_65};
  wire [1:0]        memRequest_bits_data_hi_lo_65 = {_memRequest_bits_data_T_3975[57], _memRequest_bits_data_T_3590[57]};
  wire [1:0]        memRequest_bits_data_hi_hi_65 = {_memRequest_bits_data_T_4745[57], _memRequest_bits_data_T_4360[57]};
  wire [3:0]        memRequest_bits_data_hi_65 = {memRequest_bits_data_hi_hi_65, memRequest_bits_data_hi_lo_65};
  wire [1:0]        memRequest_bits_data_lo_lo_66 = {_memRequest_bits_data_T_2435[58], _memRequest_bits_data_T_2050[58]};
  wire [1:0]        memRequest_bits_data_lo_hi_66 = {_memRequest_bits_data_T_3205[58], _memRequest_bits_data_T_2820[58]};
  wire [3:0]        memRequest_bits_data_lo_66 = {memRequest_bits_data_lo_hi_66, memRequest_bits_data_lo_lo_66};
  wire [1:0]        memRequest_bits_data_hi_lo_66 = {_memRequest_bits_data_T_3975[58], _memRequest_bits_data_T_3590[58]};
  wire [1:0]        memRequest_bits_data_hi_hi_66 = {_memRequest_bits_data_T_4745[58], _memRequest_bits_data_T_4360[58]};
  wire [3:0]        memRequest_bits_data_hi_66 = {memRequest_bits_data_hi_hi_66, memRequest_bits_data_hi_lo_66};
  wire [1:0]        memRequest_bits_data_lo_lo_67 = {_memRequest_bits_data_T_2435[59], _memRequest_bits_data_T_2050[59]};
  wire [1:0]        memRequest_bits_data_lo_hi_67 = {_memRequest_bits_data_T_3205[59], _memRequest_bits_data_T_2820[59]};
  wire [3:0]        memRequest_bits_data_lo_67 = {memRequest_bits_data_lo_hi_67, memRequest_bits_data_lo_lo_67};
  wire [1:0]        memRequest_bits_data_hi_lo_67 = {_memRequest_bits_data_T_3975[59], _memRequest_bits_data_T_3590[59]};
  wire [1:0]        memRequest_bits_data_hi_hi_67 = {_memRequest_bits_data_T_4745[59], _memRequest_bits_data_T_4360[59]};
  wire [3:0]        memRequest_bits_data_hi_67 = {memRequest_bits_data_hi_hi_67, memRequest_bits_data_hi_lo_67};
  wire [1:0]        memRequest_bits_data_lo_lo_68 = {_memRequest_bits_data_T_2435[60], _memRequest_bits_data_T_2050[60]};
  wire [1:0]        memRequest_bits_data_lo_hi_68 = {_memRequest_bits_data_T_3205[60], _memRequest_bits_data_T_2820[60]};
  wire [3:0]        memRequest_bits_data_lo_68 = {memRequest_bits_data_lo_hi_68, memRequest_bits_data_lo_lo_68};
  wire [1:0]        memRequest_bits_data_hi_lo_68 = {_memRequest_bits_data_T_3975[60], _memRequest_bits_data_T_3590[60]};
  wire [1:0]        memRequest_bits_data_hi_hi_68 = {_memRequest_bits_data_T_4745[60], _memRequest_bits_data_T_4360[60]};
  wire [3:0]        memRequest_bits_data_hi_68 = {memRequest_bits_data_hi_hi_68, memRequest_bits_data_hi_lo_68};
  wire [1:0]        memRequest_bits_data_lo_lo_69 = {_memRequest_bits_data_T_2435[61], _memRequest_bits_data_T_2050[61]};
  wire [1:0]        memRequest_bits_data_lo_hi_69 = {_memRequest_bits_data_T_3205[61], _memRequest_bits_data_T_2820[61]};
  wire [3:0]        memRequest_bits_data_lo_69 = {memRequest_bits_data_lo_hi_69, memRequest_bits_data_lo_lo_69};
  wire [1:0]        memRequest_bits_data_hi_lo_69 = {_memRequest_bits_data_T_3975[61], _memRequest_bits_data_T_3590[61]};
  wire [1:0]        memRequest_bits_data_hi_hi_69 = {_memRequest_bits_data_T_4745[61], _memRequest_bits_data_T_4360[61]};
  wire [3:0]        memRequest_bits_data_hi_69 = {memRequest_bits_data_hi_hi_69, memRequest_bits_data_hi_lo_69};
  wire [1:0]        memRequest_bits_data_lo_lo_70 = {_memRequest_bits_data_T_2435[62], _memRequest_bits_data_T_2050[62]};
  wire [1:0]        memRequest_bits_data_lo_hi_70 = {_memRequest_bits_data_T_3205[62], _memRequest_bits_data_T_2820[62]};
  wire [3:0]        memRequest_bits_data_lo_70 = {memRequest_bits_data_lo_hi_70, memRequest_bits_data_lo_lo_70};
  wire [1:0]        memRequest_bits_data_hi_lo_70 = {_memRequest_bits_data_T_3975[62], _memRequest_bits_data_T_3590[62]};
  wire [1:0]        memRequest_bits_data_hi_hi_70 = {_memRequest_bits_data_T_4745[62], _memRequest_bits_data_T_4360[62]};
  wire [3:0]        memRequest_bits_data_hi_70 = {memRequest_bits_data_hi_hi_70, memRequest_bits_data_hi_lo_70};
  wire [1:0]        memRequest_bits_data_lo_lo_71 = {_memRequest_bits_data_T_2435[63], _memRequest_bits_data_T_2050[63]};
  wire [1:0]        memRequest_bits_data_lo_hi_71 = {_memRequest_bits_data_T_3205[63], _memRequest_bits_data_T_2820[63]};
  wire [3:0]        memRequest_bits_data_lo_71 = {memRequest_bits_data_lo_hi_71, memRequest_bits_data_lo_lo_71};
  wire [1:0]        memRequest_bits_data_hi_lo_71 = {_memRequest_bits_data_T_3975[63], _memRequest_bits_data_T_3590[63]};
  wire [1:0]        memRequest_bits_data_hi_hi_71 = {_memRequest_bits_data_T_4745[63], _memRequest_bits_data_T_4360[63]};
  wire [3:0]        memRequest_bits_data_hi_71 = {memRequest_bits_data_hi_hi_71, memRequest_bits_data_hi_lo_71};
  wire [1:0]        memRequest_bits_data_lo_lo_72 = {_memRequest_bits_data_T_2435[64], _memRequest_bits_data_T_2050[64]};
  wire [1:0]        memRequest_bits_data_lo_hi_72 = {_memRequest_bits_data_T_3205[64], _memRequest_bits_data_T_2820[64]};
  wire [3:0]        memRequest_bits_data_lo_72 = {memRequest_bits_data_lo_hi_72, memRequest_bits_data_lo_lo_72};
  wire [1:0]        memRequest_bits_data_hi_lo_72 = {_memRequest_bits_data_T_3975[64], _memRequest_bits_data_T_3590[64]};
  wire [1:0]        memRequest_bits_data_hi_hi_72 = {_memRequest_bits_data_T_4745[64], _memRequest_bits_data_T_4360[64]};
  wire [3:0]        memRequest_bits_data_hi_72 = {memRequest_bits_data_hi_hi_72, memRequest_bits_data_hi_lo_72};
  wire [1:0]        memRequest_bits_data_lo_lo_73 = {_memRequest_bits_data_T_2435[65], _memRequest_bits_data_T_2050[65]};
  wire [1:0]        memRequest_bits_data_lo_hi_73 = {_memRequest_bits_data_T_3205[65], _memRequest_bits_data_T_2820[65]};
  wire [3:0]        memRequest_bits_data_lo_73 = {memRequest_bits_data_lo_hi_73, memRequest_bits_data_lo_lo_73};
  wire [1:0]        memRequest_bits_data_hi_lo_73 = {_memRequest_bits_data_T_3975[65], _memRequest_bits_data_T_3590[65]};
  wire [1:0]        memRequest_bits_data_hi_hi_73 = {_memRequest_bits_data_T_4745[65], _memRequest_bits_data_T_4360[65]};
  wire [3:0]        memRequest_bits_data_hi_73 = {memRequest_bits_data_hi_hi_73, memRequest_bits_data_hi_lo_73};
  wire [1:0]        memRequest_bits_data_lo_lo_74 = {_memRequest_bits_data_T_2435[66], _memRequest_bits_data_T_2050[66]};
  wire [1:0]        memRequest_bits_data_lo_hi_74 = {_memRequest_bits_data_T_3205[66], _memRequest_bits_data_T_2820[66]};
  wire [3:0]        memRequest_bits_data_lo_74 = {memRequest_bits_data_lo_hi_74, memRequest_bits_data_lo_lo_74};
  wire [1:0]        memRequest_bits_data_hi_lo_74 = {_memRequest_bits_data_T_3975[66], _memRequest_bits_data_T_3590[66]};
  wire [1:0]        memRequest_bits_data_hi_hi_74 = {_memRequest_bits_data_T_4745[66], _memRequest_bits_data_T_4360[66]};
  wire [3:0]        memRequest_bits_data_hi_74 = {memRequest_bits_data_hi_hi_74, memRequest_bits_data_hi_lo_74};
  wire [1:0]        memRequest_bits_data_lo_lo_75 = {_memRequest_bits_data_T_2435[67], _memRequest_bits_data_T_2050[67]};
  wire [1:0]        memRequest_bits_data_lo_hi_75 = {_memRequest_bits_data_T_3205[67], _memRequest_bits_data_T_2820[67]};
  wire [3:0]        memRequest_bits_data_lo_75 = {memRequest_bits_data_lo_hi_75, memRequest_bits_data_lo_lo_75};
  wire [1:0]        memRequest_bits_data_hi_lo_75 = {_memRequest_bits_data_T_3975[67], _memRequest_bits_data_T_3590[67]};
  wire [1:0]        memRequest_bits_data_hi_hi_75 = {_memRequest_bits_data_T_4745[67], _memRequest_bits_data_T_4360[67]};
  wire [3:0]        memRequest_bits_data_hi_75 = {memRequest_bits_data_hi_hi_75, memRequest_bits_data_hi_lo_75};
  wire [1:0]        memRequest_bits_data_lo_lo_76 = {_memRequest_bits_data_T_2435[68], _memRequest_bits_data_T_2050[68]};
  wire [1:0]        memRequest_bits_data_lo_hi_76 = {_memRequest_bits_data_T_3205[68], _memRequest_bits_data_T_2820[68]};
  wire [3:0]        memRequest_bits_data_lo_76 = {memRequest_bits_data_lo_hi_76, memRequest_bits_data_lo_lo_76};
  wire [1:0]        memRequest_bits_data_hi_lo_76 = {_memRequest_bits_data_T_3975[68], _memRequest_bits_data_T_3590[68]};
  wire [1:0]        memRequest_bits_data_hi_hi_76 = {_memRequest_bits_data_T_4745[68], _memRequest_bits_data_T_4360[68]};
  wire [3:0]        memRequest_bits_data_hi_76 = {memRequest_bits_data_hi_hi_76, memRequest_bits_data_hi_lo_76};
  wire [1:0]        memRequest_bits_data_lo_lo_77 = {_memRequest_bits_data_T_2435[69], _memRequest_bits_data_T_2050[69]};
  wire [1:0]        memRequest_bits_data_lo_hi_77 = {_memRequest_bits_data_T_3205[69], _memRequest_bits_data_T_2820[69]};
  wire [3:0]        memRequest_bits_data_lo_77 = {memRequest_bits_data_lo_hi_77, memRequest_bits_data_lo_lo_77};
  wire [1:0]        memRequest_bits_data_hi_lo_77 = {_memRequest_bits_data_T_3975[69], _memRequest_bits_data_T_3590[69]};
  wire [1:0]        memRequest_bits_data_hi_hi_77 = {_memRequest_bits_data_T_4745[69], _memRequest_bits_data_T_4360[69]};
  wire [3:0]        memRequest_bits_data_hi_77 = {memRequest_bits_data_hi_hi_77, memRequest_bits_data_hi_lo_77};
  wire [1:0]        memRequest_bits_data_lo_lo_78 = {_memRequest_bits_data_T_2435[70], _memRequest_bits_data_T_2050[70]};
  wire [1:0]        memRequest_bits_data_lo_hi_78 = {_memRequest_bits_data_T_3205[70], _memRequest_bits_data_T_2820[70]};
  wire [3:0]        memRequest_bits_data_lo_78 = {memRequest_bits_data_lo_hi_78, memRequest_bits_data_lo_lo_78};
  wire [1:0]        memRequest_bits_data_hi_lo_78 = {_memRequest_bits_data_T_3975[70], _memRequest_bits_data_T_3590[70]};
  wire [1:0]        memRequest_bits_data_hi_hi_78 = {_memRequest_bits_data_T_4745[70], _memRequest_bits_data_T_4360[70]};
  wire [3:0]        memRequest_bits_data_hi_78 = {memRequest_bits_data_hi_hi_78, memRequest_bits_data_hi_lo_78};
  wire [1:0]        memRequest_bits_data_lo_lo_79 = {_memRequest_bits_data_T_2435[71], _memRequest_bits_data_T_2050[71]};
  wire [1:0]        memRequest_bits_data_lo_hi_79 = {_memRequest_bits_data_T_3205[71], _memRequest_bits_data_T_2820[71]};
  wire [3:0]        memRequest_bits_data_lo_79 = {memRequest_bits_data_lo_hi_79, memRequest_bits_data_lo_lo_79};
  wire [1:0]        memRequest_bits_data_hi_lo_79 = {_memRequest_bits_data_T_3975[71], _memRequest_bits_data_T_3590[71]};
  wire [1:0]        memRequest_bits_data_hi_hi_79 = {_memRequest_bits_data_T_4745[71], _memRequest_bits_data_T_4360[71]};
  wire [3:0]        memRequest_bits_data_hi_79 = {memRequest_bits_data_hi_hi_79, memRequest_bits_data_hi_lo_79};
  wire [1:0]        memRequest_bits_data_lo_lo_80 = {_memRequest_bits_data_T_2435[72], _memRequest_bits_data_T_2050[72]};
  wire [1:0]        memRequest_bits_data_lo_hi_80 = {_memRequest_bits_data_T_3205[72], _memRequest_bits_data_T_2820[72]};
  wire [3:0]        memRequest_bits_data_lo_80 = {memRequest_bits_data_lo_hi_80, memRequest_bits_data_lo_lo_80};
  wire [1:0]        memRequest_bits_data_hi_lo_80 = {_memRequest_bits_data_T_3975[72], _memRequest_bits_data_T_3590[72]};
  wire [1:0]        memRequest_bits_data_hi_hi_80 = {_memRequest_bits_data_T_4745[72], _memRequest_bits_data_T_4360[72]};
  wire [3:0]        memRequest_bits_data_hi_80 = {memRequest_bits_data_hi_hi_80, memRequest_bits_data_hi_lo_80};
  wire [1:0]        memRequest_bits_data_lo_lo_81 = {_memRequest_bits_data_T_2435[73], _memRequest_bits_data_T_2050[73]};
  wire [1:0]        memRequest_bits_data_lo_hi_81 = {_memRequest_bits_data_T_3205[73], _memRequest_bits_data_T_2820[73]};
  wire [3:0]        memRequest_bits_data_lo_81 = {memRequest_bits_data_lo_hi_81, memRequest_bits_data_lo_lo_81};
  wire [1:0]        memRequest_bits_data_hi_lo_81 = {_memRequest_bits_data_T_3975[73], _memRequest_bits_data_T_3590[73]};
  wire [1:0]        memRequest_bits_data_hi_hi_81 = {_memRequest_bits_data_T_4745[73], _memRequest_bits_data_T_4360[73]};
  wire [3:0]        memRequest_bits_data_hi_81 = {memRequest_bits_data_hi_hi_81, memRequest_bits_data_hi_lo_81};
  wire [1:0]        memRequest_bits_data_lo_lo_82 = {_memRequest_bits_data_T_2435[74], _memRequest_bits_data_T_2050[74]};
  wire [1:0]        memRequest_bits_data_lo_hi_82 = {_memRequest_bits_data_T_3205[74], _memRequest_bits_data_T_2820[74]};
  wire [3:0]        memRequest_bits_data_lo_82 = {memRequest_bits_data_lo_hi_82, memRequest_bits_data_lo_lo_82};
  wire [1:0]        memRequest_bits_data_hi_lo_82 = {_memRequest_bits_data_T_3975[74], _memRequest_bits_data_T_3590[74]};
  wire [1:0]        memRequest_bits_data_hi_hi_82 = {_memRequest_bits_data_T_4745[74], _memRequest_bits_data_T_4360[74]};
  wire [3:0]        memRequest_bits_data_hi_82 = {memRequest_bits_data_hi_hi_82, memRequest_bits_data_hi_lo_82};
  wire [1:0]        memRequest_bits_data_lo_lo_83 = {_memRequest_bits_data_T_2435[75], _memRequest_bits_data_T_2050[75]};
  wire [1:0]        memRequest_bits_data_lo_hi_83 = {_memRequest_bits_data_T_3205[75], _memRequest_bits_data_T_2820[75]};
  wire [3:0]        memRequest_bits_data_lo_83 = {memRequest_bits_data_lo_hi_83, memRequest_bits_data_lo_lo_83};
  wire [1:0]        memRequest_bits_data_hi_lo_83 = {_memRequest_bits_data_T_3975[75], _memRequest_bits_data_T_3590[75]};
  wire [1:0]        memRequest_bits_data_hi_hi_83 = {_memRequest_bits_data_T_4745[75], _memRequest_bits_data_T_4360[75]};
  wire [3:0]        memRequest_bits_data_hi_83 = {memRequest_bits_data_hi_hi_83, memRequest_bits_data_hi_lo_83};
  wire [1:0]        memRequest_bits_data_lo_lo_84 = {_memRequest_bits_data_T_2435[76], _memRequest_bits_data_T_2050[76]};
  wire [1:0]        memRequest_bits_data_lo_hi_84 = {_memRequest_bits_data_T_3205[76], _memRequest_bits_data_T_2820[76]};
  wire [3:0]        memRequest_bits_data_lo_84 = {memRequest_bits_data_lo_hi_84, memRequest_bits_data_lo_lo_84};
  wire [1:0]        memRequest_bits_data_hi_lo_84 = {_memRequest_bits_data_T_3975[76], _memRequest_bits_data_T_3590[76]};
  wire [1:0]        memRequest_bits_data_hi_hi_84 = {_memRequest_bits_data_T_4745[76], _memRequest_bits_data_T_4360[76]};
  wire [3:0]        memRequest_bits_data_hi_84 = {memRequest_bits_data_hi_hi_84, memRequest_bits_data_hi_lo_84};
  wire [1:0]        memRequest_bits_data_lo_lo_85 = {_memRequest_bits_data_T_2435[77], _memRequest_bits_data_T_2050[77]};
  wire [1:0]        memRequest_bits_data_lo_hi_85 = {_memRequest_bits_data_T_3205[77], _memRequest_bits_data_T_2820[77]};
  wire [3:0]        memRequest_bits_data_lo_85 = {memRequest_bits_data_lo_hi_85, memRequest_bits_data_lo_lo_85};
  wire [1:0]        memRequest_bits_data_hi_lo_85 = {_memRequest_bits_data_T_3975[77], _memRequest_bits_data_T_3590[77]};
  wire [1:0]        memRequest_bits_data_hi_hi_85 = {_memRequest_bits_data_T_4745[77], _memRequest_bits_data_T_4360[77]};
  wire [3:0]        memRequest_bits_data_hi_85 = {memRequest_bits_data_hi_hi_85, memRequest_bits_data_hi_lo_85};
  wire [1:0]        memRequest_bits_data_lo_lo_86 = {_memRequest_bits_data_T_2435[78], _memRequest_bits_data_T_2050[78]};
  wire [1:0]        memRequest_bits_data_lo_hi_86 = {_memRequest_bits_data_T_3205[78], _memRequest_bits_data_T_2820[78]};
  wire [3:0]        memRequest_bits_data_lo_86 = {memRequest_bits_data_lo_hi_86, memRequest_bits_data_lo_lo_86};
  wire [1:0]        memRequest_bits_data_hi_lo_86 = {_memRequest_bits_data_T_3975[78], _memRequest_bits_data_T_3590[78]};
  wire [1:0]        memRequest_bits_data_hi_hi_86 = {_memRequest_bits_data_T_4745[78], _memRequest_bits_data_T_4360[78]};
  wire [3:0]        memRequest_bits_data_hi_86 = {memRequest_bits_data_hi_hi_86, memRequest_bits_data_hi_lo_86};
  wire [1:0]        memRequest_bits_data_lo_lo_87 = {_memRequest_bits_data_T_2435[79], _memRequest_bits_data_T_2050[79]};
  wire [1:0]        memRequest_bits_data_lo_hi_87 = {_memRequest_bits_data_T_3205[79], _memRequest_bits_data_T_2820[79]};
  wire [3:0]        memRequest_bits_data_lo_87 = {memRequest_bits_data_lo_hi_87, memRequest_bits_data_lo_lo_87};
  wire [1:0]        memRequest_bits_data_hi_lo_87 = {_memRequest_bits_data_T_3975[79], _memRequest_bits_data_T_3590[79]};
  wire [1:0]        memRequest_bits_data_hi_hi_87 = {_memRequest_bits_data_T_4745[79], _memRequest_bits_data_T_4360[79]};
  wire [3:0]        memRequest_bits_data_hi_87 = {memRequest_bits_data_hi_hi_87, memRequest_bits_data_hi_lo_87};
  wire [1:0]        memRequest_bits_data_lo_lo_88 = {_memRequest_bits_data_T_2435[80], _memRequest_bits_data_T_2050[80]};
  wire [1:0]        memRequest_bits_data_lo_hi_88 = {_memRequest_bits_data_T_3205[80], _memRequest_bits_data_T_2820[80]};
  wire [3:0]        memRequest_bits_data_lo_88 = {memRequest_bits_data_lo_hi_88, memRequest_bits_data_lo_lo_88};
  wire [1:0]        memRequest_bits_data_hi_lo_88 = {_memRequest_bits_data_T_3975[80], _memRequest_bits_data_T_3590[80]};
  wire [1:0]        memRequest_bits_data_hi_hi_88 = {_memRequest_bits_data_T_4745[80], _memRequest_bits_data_T_4360[80]};
  wire [3:0]        memRequest_bits_data_hi_88 = {memRequest_bits_data_hi_hi_88, memRequest_bits_data_hi_lo_88};
  wire [1:0]        memRequest_bits_data_lo_lo_89 = {_memRequest_bits_data_T_2435[81], _memRequest_bits_data_T_2050[81]};
  wire [1:0]        memRequest_bits_data_lo_hi_89 = {_memRequest_bits_data_T_3205[81], _memRequest_bits_data_T_2820[81]};
  wire [3:0]        memRequest_bits_data_lo_89 = {memRequest_bits_data_lo_hi_89, memRequest_bits_data_lo_lo_89};
  wire [1:0]        memRequest_bits_data_hi_lo_89 = {_memRequest_bits_data_T_3975[81], _memRequest_bits_data_T_3590[81]};
  wire [1:0]        memRequest_bits_data_hi_hi_89 = {_memRequest_bits_data_T_4745[81], _memRequest_bits_data_T_4360[81]};
  wire [3:0]        memRequest_bits_data_hi_89 = {memRequest_bits_data_hi_hi_89, memRequest_bits_data_hi_lo_89};
  wire [1:0]        memRequest_bits_data_lo_lo_90 = {_memRequest_bits_data_T_2435[82], _memRequest_bits_data_T_2050[82]};
  wire [1:0]        memRequest_bits_data_lo_hi_90 = {_memRequest_bits_data_T_3205[82], _memRequest_bits_data_T_2820[82]};
  wire [3:0]        memRequest_bits_data_lo_90 = {memRequest_bits_data_lo_hi_90, memRequest_bits_data_lo_lo_90};
  wire [1:0]        memRequest_bits_data_hi_lo_90 = {_memRequest_bits_data_T_3975[82], _memRequest_bits_data_T_3590[82]};
  wire [1:0]        memRequest_bits_data_hi_hi_90 = {_memRequest_bits_data_T_4745[82], _memRequest_bits_data_T_4360[82]};
  wire [3:0]        memRequest_bits_data_hi_90 = {memRequest_bits_data_hi_hi_90, memRequest_bits_data_hi_lo_90};
  wire [1:0]        memRequest_bits_data_lo_lo_91 = {_memRequest_bits_data_T_2435[83], _memRequest_bits_data_T_2050[83]};
  wire [1:0]        memRequest_bits_data_lo_hi_91 = {_memRequest_bits_data_T_3205[83], _memRequest_bits_data_T_2820[83]};
  wire [3:0]        memRequest_bits_data_lo_91 = {memRequest_bits_data_lo_hi_91, memRequest_bits_data_lo_lo_91};
  wire [1:0]        memRequest_bits_data_hi_lo_91 = {_memRequest_bits_data_T_3975[83], _memRequest_bits_data_T_3590[83]};
  wire [1:0]        memRequest_bits_data_hi_hi_91 = {_memRequest_bits_data_T_4745[83], _memRequest_bits_data_T_4360[83]};
  wire [3:0]        memRequest_bits_data_hi_91 = {memRequest_bits_data_hi_hi_91, memRequest_bits_data_hi_lo_91};
  wire [1:0]        memRequest_bits_data_lo_lo_92 = {_memRequest_bits_data_T_2435[84], _memRequest_bits_data_T_2050[84]};
  wire [1:0]        memRequest_bits_data_lo_hi_92 = {_memRequest_bits_data_T_3205[84], _memRequest_bits_data_T_2820[84]};
  wire [3:0]        memRequest_bits_data_lo_92 = {memRequest_bits_data_lo_hi_92, memRequest_bits_data_lo_lo_92};
  wire [1:0]        memRequest_bits_data_hi_lo_92 = {_memRequest_bits_data_T_3975[84], _memRequest_bits_data_T_3590[84]};
  wire [1:0]        memRequest_bits_data_hi_hi_92 = {_memRequest_bits_data_T_4745[84], _memRequest_bits_data_T_4360[84]};
  wire [3:0]        memRequest_bits_data_hi_92 = {memRequest_bits_data_hi_hi_92, memRequest_bits_data_hi_lo_92};
  wire [1:0]        memRequest_bits_data_lo_lo_93 = {_memRequest_bits_data_T_2435[85], _memRequest_bits_data_T_2050[85]};
  wire [1:0]        memRequest_bits_data_lo_hi_93 = {_memRequest_bits_data_T_3205[85], _memRequest_bits_data_T_2820[85]};
  wire [3:0]        memRequest_bits_data_lo_93 = {memRequest_bits_data_lo_hi_93, memRequest_bits_data_lo_lo_93};
  wire [1:0]        memRequest_bits_data_hi_lo_93 = {_memRequest_bits_data_T_3975[85], _memRequest_bits_data_T_3590[85]};
  wire [1:0]        memRequest_bits_data_hi_hi_93 = {_memRequest_bits_data_T_4745[85], _memRequest_bits_data_T_4360[85]};
  wire [3:0]        memRequest_bits_data_hi_93 = {memRequest_bits_data_hi_hi_93, memRequest_bits_data_hi_lo_93};
  wire [1:0]        memRequest_bits_data_lo_lo_94 = {_memRequest_bits_data_T_2435[86], _memRequest_bits_data_T_2050[86]};
  wire [1:0]        memRequest_bits_data_lo_hi_94 = {_memRequest_bits_data_T_3205[86], _memRequest_bits_data_T_2820[86]};
  wire [3:0]        memRequest_bits_data_lo_94 = {memRequest_bits_data_lo_hi_94, memRequest_bits_data_lo_lo_94};
  wire [1:0]        memRequest_bits_data_hi_lo_94 = {_memRequest_bits_data_T_3975[86], _memRequest_bits_data_T_3590[86]};
  wire [1:0]        memRequest_bits_data_hi_hi_94 = {_memRequest_bits_data_T_4745[86], _memRequest_bits_data_T_4360[86]};
  wire [3:0]        memRequest_bits_data_hi_94 = {memRequest_bits_data_hi_hi_94, memRequest_bits_data_hi_lo_94};
  wire [1:0]        memRequest_bits_data_lo_lo_95 = {_memRequest_bits_data_T_2435[87], _memRequest_bits_data_T_2050[87]};
  wire [1:0]        memRequest_bits_data_lo_hi_95 = {_memRequest_bits_data_T_3205[87], _memRequest_bits_data_T_2820[87]};
  wire [3:0]        memRequest_bits_data_lo_95 = {memRequest_bits_data_lo_hi_95, memRequest_bits_data_lo_lo_95};
  wire [1:0]        memRequest_bits_data_hi_lo_95 = {_memRequest_bits_data_T_3975[87], _memRequest_bits_data_T_3590[87]};
  wire [1:0]        memRequest_bits_data_hi_hi_95 = {_memRequest_bits_data_T_4745[87], _memRequest_bits_data_T_4360[87]};
  wire [3:0]        memRequest_bits_data_hi_95 = {memRequest_bits_data_hi_hi_95, memRequest_bits_data_hi_lo_95};
  wire [1:0]        memRequest_bits_data_lo_lo_96 = {_memRequest_bits_data_T_2435[88], _memRequest_bits_data_T_2050[88]};
  wire [1:0]        memRequest_bits_data_lo_hi_96 = {_memRequest_bits_data_T_3205[88], _memRequest_bits_data_T_2820[88]};
  wire [3:0]        memRequest_bits_data_lo_96 = {memRequest_bits_data_lo_hi_96, memRequest_bits_data_lo_lo_96};
  wire [1:0]        memRequest_bits_data_hi_lo_96 = {_memRequest_bits_data_T_3975[88], _memRequest_bits_data_T_3590[88]};
  wire [1:0]        memRequest_bits_data_hi_hi_96 = {_memRequest_bits_data_T_4745[88], _memRequest_bits_data_T_4360[88]};
  wire [3:0]        memRequest_bits_data_hi_96 = {memRequest_bits_data_hi_hi_96, memRequest_bits_data_hi_lo_96};
  wire [1:0]        memRequest_bits_data_lo_lo_97 = {_memRequest_bits_data_T_2435[89], _memRequest_bits_data_T_2050[89]};
  wire [1:0]        memRequest_bits_data_lo_hi_97 = {_memRequest_bits_data_T_3205[89], _memRequest_bits_data_T_2820[89]};
  wire [3:0]        memRequest_bits_data_lo_97 = {memRequest_bits_data_lo_hi_97, memRequest_bits_data_lo_lo_97};
  wire [1:0]        memRequest_bits_data_hi_lo_97 = {_memRequest_bits_data_T_3975[89], _memRequest_bits_data_T_3590[89]};
  wire [1:0]        memRequest_bits_data_hi_hi_97 = {_memRequest_bits_data_T_4745[89], _memRequest_bits_data_T_4360[89]};
  wire [3:0]        memRequest_bits_data_hi_97 = {memRequest_bits_data_hi_hi_97, memRequest_bits_data_hi_lo_97};
  wire [1:0]        memRequest_bits_data_lo_lo_98 = {_memRequest_bits_data_T_2435[90], _memRequest_bits_data_T_2050[90]};
  wire [1:0]        memRequest_bits_data_lo_hi_98 = {_memRequest_bits_data_T_3205[90], _memRequest_bits_data_T_2820[90]};
  wire [3:0]        memRequest_bits_data_lo_98 = {memRequest_bits_data_lo_hi_98, memRequest_bits_data_lo_lo_98};
  wire [1:0]        memRequest_bits_data_hi_lo_98 = {_memRequest_bits_data_T_3975[90], _memRequest_bits_data_T_3590[90]};
  wire [1:0]        memRequest_bits_data_hi_hi_98 = {_memRequest_bits_data_T_4745[90], _memRequest_bits_data_T_4360[90]};
  wire [3:0]        memRequest_bits_data_hi_98 = {memRequest_bits_data_hi_hi_98, memRequest_bits_data_hi_lo_98};
  wire [1:0]        memRequest_bits_data_lo_lo_99 = {_memRequest_bits_data_T_2435[91], _memRequest_bits_data_T_2050[91]};
  wire [1:0]        memRequest_bits_data_lo_hi_99 = {_memRequest_bits_data_T_3205[91], _memRequest_bits_data_T_2820[91]};
  wire [3:0]        memRequest_bits_data_lo_99 = {memRequest_bits_data_lo_hi_99, memRequest_bits_data_lo_lo_99};
  wire [1:0]        memRequest_bits_data_hi_lo_99 = {_memRequest_bits_data_T_3975[91], _memRequest_bits_data_T_3590[91]};
  wire [1:0]        memRequest_bits_data_hi_hi_99 = {_memRequest_bits_data_T_4745[91], _memRequest_bits_data_T_4360[91]};
  wire [3:0]        memRequest_bits_data_hi_99 = {memRequest_bits_data_hi_hi_99, memRequest_bits_data_hi_lo_99};
  wire [1:0]        memRequest_bits_data_lo_lo_100 = {_memRequest_bits_data_T_2435[92], _memRequest_bits_data_T_2050[92]};
  wire [1:0]        memRequest_bits_data_lo_hi_100 = {_memRequest_bits_data_T_3205[92], _memRequest_bits_data_T_2820[92]};
  wire [3:0]        memRequest_bits_data_lo_100 = {memRequest_bits_data_lo_hi_100, memRequest_bits_data_lo_lo_100};
  wire [1:0]        memRequest_bits_data_hi_lo_100 = {_memRequest_bits_data_T_3975[92], _memRequest_bits_data_T_3590[92]};
  wire [1:0]        memRequest_bits_data_hi_hi_100 = {_memRequest_bits_data_T_4745[92], _memRequest_bits_data_T_4360[92]};
  wire [3:0]        memRequest_bits_data_hi_100 = {memRequest_bits_data_hi_hi_100, memRequest_bits_data_hi_lo_100};
  wire [1:0]        memRequest_bits_data_lo_lo_101 = {_memRequest_bits_data_T_2435[93], _memRequest_bits_data_T_2050[93]};
  wire [1:0]        memRequest_bits_data_lo_hi_101 = {_memRequest_bits_data_T_3205[93], _memRequest_bits_data_T_2820[93]};
  wire [3:0]        memRequest_bits_data_lo_101 = {memRequest_bits_data_lo_hi_101, memRequest_bits_data_lo_lo_101};
  wire [1:0]        memRequest_bits_data_hi_lo_101 = {_memRequest_bits_data_T_3975[93], _memRequest_bits_data_T_3590[93]};
  wire [1:0]        memRequest_bits_data_hi_hi_101 = {_memRequest_bits_data_T_4745[93], _memRequest_bits_data_T_4360[93]};
  wire [3:0]        memRequest_bits_data_hi_101 = {memRequest_bits_data_hi_hi_101, memRequest_bits_data_hi_lo_101};
  wire [1:0]        memRequest_bits_data_lo_lo_102 = {_memRequest_bits_data_T_2435[94], _memRequest_bits_data_T_2050[94]};
  wire [1:0]        memRequest_bits_data_lo_hi_102 = {_memRequest_bits_data_T_3205[94], _memRequest_bits_data_T_2820[94]};
  wire [3:0]        memRequest_bits_data_lo_102 = {memRequest_bits_data_lo_hi_102, memRequest_bits_data_lo_lo_102};
  wire [1:0]        memRequest_bits_data_hi_lo_102 = {_memRequest_bits_data_T_3975[94], _memRequest_bits_data_T_3590[94]};
  wire [1:0]        memRequest_bits_data_hi_hi_102 = {_memRequest_bits_data_T_4745[94], _memRequest_bits_data_T_4360[94]};
  wire [3:0]        memRequest_bits_data_hi_102 = {memRequest_bits_data_hi_hi_102, memRequest_bits_data_hi_lo_102};
  wire [1:0]        memRequest_bits_data_lo_lo_103 = {_memRequest_bits_data_T_2435[95], _memRequest_bits_data_T_2050[95]};
  wire [1:0]        memRequest_bits_data_lo_hi_103 = {_memRequest_bits_data_T_3205[95], _memRequest_bits_data_T_2820[95]};
  wire [3:0]        memRequest_bits_data_lo_103 = {memRequest_bits_data_lo_hi_103, memRequest_bits_data_lo_lo_103};
  wire [1:0]        memRequest_bits_data_hi_lo_103 = {_memRequest_bits_data_T_3975[95], _memRequest_bits_data_T_3590[95]};
  wire [1:0]        memRequest_bits_data_hi_hi_103 = {_memRequest_bits_data_T_4745[95], _memRequest_bits_data_T_4360[95]};
  wire [3:0]        memRequest_bits_data_hi_103 = {memRequest_bits_data_hi_hi_103, memRequest_bits_data_hi_lo_103};
  wire [1:0]        memRequest_bits_data_lo_lo_104 = {_memRequest_bits_data_T_2435[96], _memRequest_bits_data_T_2050[96]};
  wire [1:0]        memRequest_bits_data_lo_hi_104 = {_memRequest_bits_data_T_3205[96], _memRequest_bits_data_T_2820[96]};
  wire [3:0]        memRequest_bits_data_lo_104 = {memRequest_bits_data_lo_hi_104, memRequest_bits_data_lo_lo_104};
  wire [1:0]        memRequest_bits_data_hi_lo_104 = {_memRequest_bits_data_T_3975[96], _memRequest_bits_data_T_3590[96]};
  wire [1:0]        memRequest_bits_data_hi_hi_104 = {_memRequest_bits_data_T_4745[96], _memRequest_bits_data_T_4360[96]};
  wire [3:0]        memRequest_bits_data_hi_104 = {memRequest_bits_data_hi_hi_104, memRequest_bits_data_hi_lo_104};
  wire [1:0]        memRequest_bits_data_lo_lo_105 = {_memRequest_bits_data_T_2435[97], _memRequest_bits_data_T_2050[97]};
  wire [1:0]        memRequest_bits_data_lo_hi_105 = {_memRequest_bits_data_T_3205[97], _memRequest_bits_data_T_2820[97]};
  wire [3:0]        memRequest_bits_data_lo_105 = {memRequest_bits_data_lo_hi_105, memRequest_bits_data_lo_lo_105};
  wire [1:0]        memRequest_bits_data_hi_lo_105 = {_memRequest_bits_data_T_3975[97], _memRequest_bits_data_T_3590[97]};
  wire [1:0]        memRequest_bits_data_hi_hi_105 = {_memRequest_bits_data_T_4745[97], _memRequest_bits_data_T_4360[97]};
  wire [3:0]        memRequest_bits_data_hi_105 = {memRequest_bits_data_hi_hi_105, memRequest_bits_data_hi_lo_105};
  wire [1:0]        memRequest_bits_data_lo_lo_106 = {_memRequest_bits_data_T_2435[98], _memRequest_bits_data_T_2050[98]};
  wire [1:0]        memRequest_bits_data_lo_hi_106 = {_memRequest_bits_data_T_3205[98], _memRequest_bits_data_T_2820[98]};
  wire [3:0]        memRequest_bits_data_lo_106 = {memRequest_bits_data_lo_hi_106, memRequest_bits_data_lo_lo_106};
  wire [1:0]        memRequest_bits_data_hi_lo_106 = {_memRequest_bits_data_T_3975[98], _memRequest_bits_data_T_3590[98]};
  wire [1:0]        memRequest_bits_data_hi_hi_106 = {_memRequest_bits_data_T_4745[98], _memRequest_bits_data_T_4360[98]};
  wire [3:0]        memRequest_bits_data_hi_106 = {memRequest_bits_data_hi_hi_106, memRequest_bits_data_hi_lo_106};
  wire [1:0]        memRequest_bits_data_lo_lo_107 = {_memRequest_bits_data_T_2435[99], _memRequest_bits_data_T_2050[99]};
  wire [1:0]        memRequest_bits_data_lo_hi_107 = {_memRequest_bits_data_T_3205[99], _memRequest_bits_data_T_2820[99]};
  wire [3:0]        memRequest_bits_data_lo_107 = {memRequest_bits_data_lo_hi_107, memRequest_bits_data_lo_lo_107};
  wire [1:0]        memRequest_bits_data_hi_lo_107 = {_memRequest_bits_data_T_3975[99], _memRequest_bits_data_T_3590[99]};
  wire [1:0]        memRequest_bits_data_hi_hi_107 = {_memRequest_bits_data_T_4745[99], _memRequest_bits_data_T_4360[99]};
  wire [3:0]        memRequest_bits_data_hi_107 = {memRequest_bits_data_hi_hi_107, memRequest_bits_data_hi_lo_107};
  wire [1:0]        memRequest_bits_data_lo_lo_108 = {_memRequest_bits_data_T_2435[100], _memRequest_bits_data_T_2050[100]};
  wire [1:0]        memRequest_bits_data_lo_hi_108 = {_memRequest_bits_data_T_3205[100], _memRequest_bits_data_T_2820[100]};
  wire [3:0]        memRequest_bits_data_lo_108 = {memRequest_bits_data_lo_hi_108, memRequest_bits_data_lo_lo_108};
  wire [1:0]        memRequest_bits_data_hi_lo_108 = {_memRequest_bits_data_T_3975[100], _memRequest_bits_data_T_3590[100]};
  wire [1:0]        memRequest_bits_data_hi_hi_108 = {_memRequest_bits_data_T_4745[100], _memRequest_bits_data_T_4360[100]};
  wire [3:0]        memRequest_bits_data_hi_108 = {memRequest_bits_data_hi_hi_108, memRequest_bits_data_hi_lo_108};
  wire [1:0]        memRequest_bits_data_lo_lo_109 = {_memRequest_bits_data_T_2435[101], _memRequest_bits_data_T_2050[101]};
  wire [1:0]        memRequest_bits_data_lo_hi_109 = {_memRequest_bits_data_T_3205[101], _memRequest_bits_data_T_2820[101]};
  wire [3:0]        memRequest_bits_data_lo_109 = {memRequest_bits_data_lo_hi_109, memRequest_bits_data_lo_lo_109};
  wire [1:0]        memRequest_bits_data_hi_lo_109 = {_memRequest_bits_data_T_3975[101], _memRequest_bits_data_T_3590[101]};
  wire [1:0]        memRequest_bits_data_hi_hi_109 = {_memRequest_bits_data_T_4745[101], _memRequest_bits_data_T_4360[101]};
  wire [3:0]        memRequest_bits_data_hi_109 = {memRequest_bits_data_hi_hi_109, memRequest_bits_data_hi_lo_109};
  wire [1:0]        memRequest_bits_data_lo_lo_110 = {_memRequest_bits_data_T_2435[102], _memRequest_bits_data_T_2050[102]};
  wire [1:0]        memRequest_bits_data_lo_hi_110 = {_memRequest_bits_data_T_3205[102], _memRequest_bits_data_T_2820[102]};
  wire [3:0]        memRequest_bits_data_lo_110 = {memRequest_bits_data_lo_hi_110, memRequest_bits_data_lo_lo_110};
  wire [1:0]        memRequest_bits_data_hi_lo_110 = {_memRequest_bits_data_T_3975[102], _memRequest_bits_data_T_3590[102]};
  wire [1:0]        memRequest_bits_data_hi_hi_110 = {_memRequest_bits_data_T_4745[102], _memRequest_bits_data_T_4360[102]};
  wire [3:0]        memRequest_bits_data_hi_110 = {memRequest_bits_data_hi_hi_110, memRequest_bits_data_hi_lo_110};
  wire [1:0]        memRequest_bits_data_lo_lo_111 = {_memRequest_bits_data_T_2435[103], _memRequest_bits_data_T_2050[103]};
  wire [1:0]        memRequest_bits_data_lo_hi_111 = {_memRequest_bits_data_T_3205[103], _memRequest_bits_data_T_2820[103]};
  wire [3:0]        memRequest_bits_data_lo_111 = {memRequest_bits_data_lo_hi_111, memRequest_bits_data_lo_lo_111};
  wire [1:0]        memRequest_bits_data_hi_lo_111 = {_memRequest_bits_data_T_3975[103], _memRequest_bits_data_T_3590[103]};
  wire [1:0]        memRequest_bits_data_hi_hi_111 = {_memRequest_bits_data_T_4745[103], _memRequest_bits_data_T_4360[103]};
  wire [3:0]        memRequest_bits_data_hi_111 = {memRequest_bits_data_hi_hi_111, memRequest_bits_data_hi_lo_111};
  wire [1:0]        memRequest_bits_data_lo_lo_112 = {_memRequest_bits_data_T_2435[104], _memRequest_bits_data_T_2050[104]};
  wire [1:0]        memRequest_bits_data_lo_hi_112 = {_memRequest_bits_data_T_3205[104], _memRequest_bits_data_T_2820[104]};
  wire [3:0]        memRequest_bits_data_lo_112 = {memRequest_bits_data_lo_hi_112, memRequest_bits_data_lo_lo_112};
  wire [1:0]        memRequest_bits_data_hi_lo_112 = {_memRequest_bits_data_T_3975[104], _memRequest_bits_data_T_3590[104]};
  wire [1:0]        memRequest_bits_data_hi_hi_112 = {_memRequest_bits_data_T_4745[104], _memRequest_bits_data_T_4360[104]};
  wire [3:0]        memRequest_bits_data_hi_112 = {memRequest_bits_data_hi_hi_112, memRequest_bits_data_hi_lo_112};
  wire [1:0]        memRequest_bits_data_lo_lo_113 = {_memRequest_bits_data_T_2435[105], _memRequest_bits_data_T_2050[105]};
  wire [1:0]        memRequest_bits_data_lo_hi_113 = {_memRequest_bits_data_T_3205[105], _memRequest_bits_data_T_2820[105]};
  wire [3:0]        memRequest_bits_data_lo_113 = {memRequest_bits_data_lo_hi_113, memRequest_bits_data_lo_lo_113};
  wire [1:0]        memRequest_bits_data_hi_lo_113 = {_memRequest_bits_data_T_3975[105], _memRequest_bits_data_T_3590[105]};
  wire [1:0]        memRequest_bits_data_hi_hi_113 = {_memRequest_bits_data_T_4745[105], _memRequest_bits_data_T_4360[105]};
  wire [3:0]        memRequest_bits_data_hi_113 = {memRequest_bits_data_hi_hi_113, memRequest_bits_data_hi_lo_113};
  wire [1:0]        memRequest_bits_data_lo_lo_114 = {_memRequest_bits_data_T_2435[106], _memRequest_bits_data_T_2050[106]};
  wire [1:0]        memRequest_bits_data_lo_hi_114 = {_memRequest_bits_data_T_3205[106], _memRequest_bits_data_T_2820[106]};
  wire [3:0]        memRequest_bits_data_lo_114 = {memRequest_bits_data_lo_hi_114, memRequest_bits_data_lo_lo_114};
  wire [1:0]        memRequest_bits_data_hi_lo_114 = {_memRequest_bits_data_T_3975[106], _memRequest_bits_data_T_3590[106]};
  wire [1:0]        memRequest_bits_data_hi_hi_114 = {_memRequest_bits_data_T_4745[106], _memRequest_bits_data_T_4360[106]};
  wire [3:0]        memRequest_bits_data_hi_114 = {memRequest_bits_data_hi_hi_114, memRequest_bits_data_hi_lo_114};
  wire [1:0]        memRequest_bits_data_lo_lo_115 = {_memRequest_bits_data_T_2435[107], _memRequest_bits_data_T_2050[107]};
  wire [1:0]        memRequest_bits_data_lo_hi_115 = {_memRequest_bits_data_T_3205[107], _memRequest_bits_data_T_2820[107]};
  wire [3:0]        memRequest_bits_data_lo_115 = {memRequest_bits_data_lo_hi_115, memRequest_bits_data_lo_lo_115};
  wire [1:0]        memRequest_bits_data_hi_lo_115 = {_memRequest_bits_data_T_3975[107], _memRequest_bits_data_T_3590[107]};
  wire [1:0]        memRequest_bits_data_hi_hi_115 = {_memRequest_bits_data_T_4745[107], _memRequest_bits_data_T_4360[107]};
  wire [3:0]        memRequest_bits_data_hi_115 = {memRequest_bits_data_hi_hi_115, memRequest_bits_data_hi_lo_115};
  wire [1:0]        memRequest_bits_data_lo_lo_116 = {_memRequest_bits_data_T_2435[108], _memRequest_bits_data_T_2050[108]};
  wire [1:0]        memRequest_bits_data_lo_hi_116 = {_memRequest_bits_data_T_3205[108], _memRequest_bits_data_T_2820[108]};
  wire [3:0]        memRequest_bits_data_lo_116 = {memRequest_bits_data_lo_hi_116, memRequest_bits_data_lo_lo_116};
  wire [1:0]        memRequest_bits_data_hi_lo_116 = {_memRequest_bits_data_T_3975[108], _memRequest_bits_data_T_3590[108]};
  wire [1:0]        memRequest_bits_data_hi_hi_116 = {_memRequest_bits_data_T_4745[108], _memRequest_bits_data_T_4360[108]};
  wire [3:0]        memRequest_bits_data_hi_116 = {memRequest_bits_data_hi_hi_116, memRequest_bits_data_hi_lo_116};
  wire [1:0]        memRequest_bits_data_lo_lo_117 = {_memRequest_bits_data_T_2435[109], _memRequest_bits_data_T_2050[109]};
  wire [1:0]        memRequest_bits_data_lo_hi_117 = {_memRequest_bits_data_T_3205[109], _memRequest_bits_data_T_2820[109]};
  wire [3:0]        memRequest_bits_data_lo_117 = {memRequest_bits_data_lo_hi_117, memRequest_bits_data_lo_lo_117};
  wire [1:0]        memRequest_bits_data_hi_lo_117 = {_memRequest_bits_data_T_3975[109], _memRequest_bits_data_T_3590[109]};
  wire [1:0]        memRequest_bits_data_hi_hi_117 = {_memRequest_bits_data_T_4745[109], _memRequest_bits_data_T_4360[109]};
  wire [3:0]        memRequest_bits_data_hi_117 = {memRequest_bits_data_hi_hi_117, memRequest_bits_data_hi_lo_117};
  wire [1:0]        memRequest_bits_data_lo_lo_118 = {_memRequest_bits_data_T_2435[110], _memRequest_bits_data_T_2050[110]};
  wire [1:0]        memRequest_bits_data_lo_hi_118 = {_memRequest_bits_data_T_3205[110], _memRequest_bits_data_T_2820[110]};
  wire [3:0]        memRequest_bits_data_lo_118 = {memRequest_bits_data_lo_hi_118, memRequest_bits_data_lo_lo_118};
  wire [1:0]        memRequest_bits_data_hi_lo_118 = {_memRequest_bits_data_T_3975[110], _memRequest_bits_data_T_3590[110]};
  wire [1:0]        memRequest_bits_data_hi_hi_118 = {_memRequest_bits_data_T_4745[110], _memRequest_bits_data_T_4360[110]};
  wire [3:0]        memRequest_bits_data_hi_118 = {memRequest_bits_data_hi_hi_118, memRequest_bits_data_hi_lo_118};
  wire [1:0]        memRequest_bits_data_lo_lo_119 = {_memRequest_bits_data_T_2435[111], _memRequest_bits_data_T_2050[111]};
  wire [1:0]        memRequest_bits_data_lo_hi_119 = {_memRequest_bits_data_T_3205[111], _memRequest_bits_data_T_2820[111]};
  wire [3:0]        memRequest_bits_data_lo_119 = {memRequest_bits_data_lo_hi_119, memRequest_bits_data_lo_lo_119};
  wire [1:0]        memRequest_bits_data_hi_lo_119 = {_memRequest_bits_data_T_3975[111], _memRequest_bits_data_T_3590[111]};
  wire [1:0]        memRequest_bits_data_hi_hi_119 = {_memRequest_bits_data_T_4745[111], _memRequest_bits_data_T_4360[111]};
  wire [3:0]        memRequest_bits_data_hi_119 = {memRequest_bits_data_hi_hi_119, memRequest_bits_data_hi_lo_119};
  wire [1:0]        memRequest_bits_data_lo_lo_120 = {_memRequest_bits_data_T_2435[112], _memRequest_bits_data_T_2050[112]};
  wire [1:0]        memRequest_bits_data_lo_hi_120 = {_memRequest_bits_data_T_3205[112], _memRequest_bits_data_T_2820[112]};
  wire [3:0]        memRequest_bits_data_lo_120 = {memRequest_bits_data_lo_hi_120, memRequest_bits_data_lo_lo_120};
  wire [1:0]        memRequest_bits_data_hi_lo_120 = {_memRequest_bits_data_T_3975[112], _memRequest_bits_data_T_3590[112]};
  wire [1:0]        memRequest_bits_data_hi_hi_120 = {_memRequest_bits_data_T_4745[112], _memRequest_bits_data_T_4360[112]};
  wire [3:0]        memRequest_bits_data_hi_120 = {memRequest_bits_data_hi_hi_120, memRequest_bits_data_hi_lo_120};
  wire [1:0]        memRequest_bits_data_lo_lo_121 = {_memRequest_bits_data_T_2435[113], _memRequest_bits_data_T_2050[113]};
  wire [1:0]        memRequest_bits_data_lo_hi_121 = {_memRequest_bits_data_T_3205[113], _memRequest_bits_data_T_2820[113]};
  wire [3:0]        memRequest_bits_data_lo_121 = {memRequest_bits_data_lo_hi_121, memRequest_bits_data_lo_lo_121};
  wire [1:0]        memRequest_bits_data_hi_lo_121 = {_memRequest_bits_data_T_3975[113], _memRequest_bits_data_T_3590[113]};
  wire [1:0]        memRequest_bits_data_hi_hi_121 = {_memRequest_bits_data_T_4745[113], _memRequest_bits_data_T_4360[113]};
  wire [3:0]        memRequest_bits_data_hi_121 = {memRequest_bits_data_hi_hi_121, memRequest_bits_data_hi_lo_121};
  wire [1:0]        memRequest_bits_data_lo_lo_122 = {_memRequest_bits_data_T_2435[114], _memRequest_bits_data_T_2050[114]};
  wire [1:0]        memRequest_bits_data_lo_hi_122 = {_memRequest_bits_data_T_3205[114], _memRequest_bits_data_T_2820[114]};
  wire [3:0]        memRequest_bits_data_lo_122 = {memRequest_bits_data_lo_hi_122, memRequest_bits_data_lo_lo_122};
  wire [1:0]        memRequest_bits_data_hi_lo_122 = {_memRequest_bits_data_T_3975[114], _memRequest_bits_data_T_3590[114]};
  wire [1:0]        memRequest_bits_data_hi_hi_122 = {_memRequest_bits_data_T_4745[114], _memRequest_bits_data_T_4360[114]};
  wire [3:0]        memRequest_bits_data_hi_122 = {memRequest_bits_data_hi_hi_122, memRequest_bits_data_hi_lo_122};
  wire [1:0]        memRequest_bits_data_lo_lo_123 = {_memRequest_bits_data_T_2435[115], _memRequest_bits_data_T_2050[115]};
  wire [1:0]        memRequest_bits_data_lo_hi_123 = {_memRequest_bits_data_T_3205[115], _memRequest_bits_data_T_2820[115]};
  wire [3:0]        memRequest_bits_data_lo_123 = {memRequest_bits_data_lo_hi_123, memRequest_bits_data_lo_lo_123};
  wire [1:0]        memRequest_bits_data_hi_lo_123 = {_memRequest_bits_data_T_3975[115], _memRequest_bits_data_T_3590[115]};
  wire [1:0]        memRequest_bits_data_hi_hi_123 = {_memRequest_bits_data_T_4745[115], _memRequest_bits_data_T_4360[115]};
  wire [3:0]        memRequest_bits_data_hi_123 = {memRequest_bits_data_hi_hi_123, memRequest_bits_data_hi_lo_123};
  wire [1:0]        memRequest_bits_data_lo_lo_124 = {_memRequest_bits_data_T_2435[116], _memRequest_bits_data_T_2050[116]};
  wire [1:0]        memRequest_bits_data_lo_hi_124 = {_memRequest_bits_data_T_3205[116], _memRequest_bits_data_T_2820[116]};
  wire [3:0]        memRequest_bits_data_lo_124 = {memRequest_bits_data_lo_hi_124, memRequest_bits_data_lo_lo_124};
  wire [1:0]        memRequest_bits_data_hi_lo_124 = {_memRequest_bits_data_T_3975[116], _memRequest_bits_data_T_3590[116]};
  wire [1:0]        memRequest_bits_data_hi_hi_124 = {_memRequest_bits_data_T_4745[116], _memRequest_bits_data_T_4360[116]};
  wire [3:0]        memRequest_bits_data_hi_124 = {memRequest_bits_data_hi_hi_124, memRequest_bits_data_hi_lo_124};
  wire [1:0]        memRequest_bits_data_lo_lo_125 = {_memRequest_bits_data_T_2435[117], _memRequest_bits_data_T_2050[117]};
  wire [1:0]        memRequest_bits_data_lo_hi_125 = {_memRequest_bits_data_T_3205[117], _memRequest_bits_data_T_2820[117]};
  wire [3:0]        memRequest_bits_data_lo_125 = {memRequest_bits_data_lo_hi_125, memRequest_bits_data_lo_lo_125};
  wire [1:0]        memRequest_bits_data_hi_lo_125 = {_memRequest_bits_data_T_3975[117], _memRequest_bits_data_T_3590[117]};
  wire [1:0]        memRequest_bits_data_hi_hi_125 = {_memRequest_bits_data_T_4745[117], _memRequest_bits_data_T_4360[117]};
  wire [3:0]        memRequest_bits_data_hi_125 = {memRequest_bits_data_hi_hi_125, memRequest_bits_data_hi_lo_125};
  wire [1:0]        memRequest_bits_data_lo_lo_126 = {_memRequest_bits_data_T_2435[118], _memRequest_bits_data_T_2050[118]};
  wire [1:0]        memRequest_bits_data_lo_hi_126 = {_memRequest_bits_data_T_3205[118], _memRequest_bits_data_T_2820[118]};
  wire [3:0]        memRequest_bits_data_lo_126 = {memRequest_bits_data_lo_hi_126, memRequest_bits_data_lo_lo_126};
  wire [1:0]        memRequest_bits_data_hi_lo_126 = {_memRequest_bits_data_T_3975[118], _memRequest_bits_data_T_3590[118]};
  wire [1:0]        memRequest_bits_data_hi_hi_126 = {_memRequest_bits_data_T_4745[118], _memRequest_bits_data_T_4360[118]};
  wire [3:0]        memRequest_bits_data_hi_126 = {memRequest_bits_data_hi_hi_126, memRequest_bits_data_hi_lo_126};
  wire [1:0]        memRequest_bits_data_lo_lo_127 = {_memRequest_bits_data_T_2435[119], _memRequest_bits_data_T_2050[119]};
  wire [1:0]        memRequest_bits_data_lo_hi_127 = {_memRequest_bits_data_T_3205[119], _memRequest_bits_data_T_2820[119]};
  wire [3:0]        memRequest_bits_data_lo_127 = {memRequest_bits_data_lo_hi_127, memRequest_bits_data_lo_lo_127};
  wire [1:0]        memRequest_bits_data_hi_lo_127 = {_memRequest_bits_data_T_3975[119], _memRequest_bits_data_T_3590[119]};
  wire [1:0]        memRequest_bits_data_hi_hi_127 = {_memRequest_bits_data_T_4745[119], _memRequest_bits_data_T_4360[119]};
  wire [3:0]        memRequest_bits_data_hi_127 = {memRequest_bits_data_hi_hi_127, memRequest_bits_data_hi_lo_127};
  wire [1:0]        memRequest_bits_data_lo_lo_128 = {_memRequest_bits_data_T_2435[120], _memRequest_bits_data_T_2050[120]};
  wire [1:0]        memRequest_bits_data_lo_hi_128 = {_memRequest_bits_data_T_3205[120], _memRequest_bits_data_T_2820[120]};
  wire [3:0]        memRequest_bits_data_lo_128 = {memRequest_bits_data_lo_hi_128, memRequest_bits_data_lo_lo_128};
  wire [1:0]        memRequest_bits_data_hi_lo_128 = {_memRequest_bits_data_T_3975[120], _memRequest_bits_data_T_3590[120]};
  wire [1:0]        memRequest_bits_data_hi_hi_128 = {_memRequest_bits_data_T_4745[120], _memRequest_bits_data_T_4360[120]};
  wire [3:0]        memRequest_bits_data_hi_128 = {memRequest_bits_data_hi_hi_128, memRequest_bits_data_hi_lo_128};
  wire [1:0]        memRequest_bits_data_lo_lo_129 = {_memRequest_bits_data_T_2435[121], _memRequest_bits_data_T_2050[121]};
  wire [1:0]        memRequest_bits_data_lo_hi_129 = {_memRequest_bits_data_T_3205[121], _memRequest_bits_data_T_2820[121]};
  wire [3:0]        memRequest_bits_data_lo_129 = {memRequest_bits_data_lo_hi_129, memRequest_bits_data_lo_lo_129};
  wire [1:0]        memRequest_bits_data_hi_lo_129 = {_memRequest_bits_data_T_3975[121], _memRequest_bits_data_T_3590[121]};
  wire [1:0]        memRequest_bits_data_hi_hi_129 = {_memRequest_bits_data_T_4745[121], _memRequest_bits_data_T_4360[121]};
  wire [3:0]        memRequest_bits_data_hi_129 = {memRequest_bits_data_hi_hi_129, memRequest_bits_data_hi_lo_129};
  wire [1:0]        memRequest_bits_data_lo_lo_130 = {_memRequest_bits_data_T_2435[122], _memRequest_bits_data_T_2050[122]};
  wire [1:0]        memRequest_bits_data_lo_hi_130 = {_memRequest_bits_data_T_3205[122], _memRequest_bits_data_T_2820[122]};
  wire [3:0]        memRequest_bits_data_lo_130 = {memRequest_bits_data_lo_hi_130, memRequest_bits_data_lo_lo_130};
  wire [1:0]        memRequest_bits_data_hi_lo_130 = {_memRequest_bits_data_T_3975[122], _memRequest_bits_data_T_3590[122]};
  wire [1:0]        memRequest_bits_data_hi_hi_130 = {_memRequest_bits_data_T_4745[122], _memRequest_bits_data_T_4360[122]};
  wire [3:0]        memRequest_bits_data_hi_130 = {memRequest_bits_data_hi_hi_130, memRequest_bits_data_hi_lo_130};
  wire [1:0]        memRequest_bits_data_lo_lo_131 = {_memRequest_bits_data_T_2435[123], _memRequest_bits_data_T_2050[123]};
  wire [1:0]        memRequest_bits_data_lo_hi_131 = {_memRequest_bits_data_T_3205[123], _memRequest_bits_data_T_2820[123]};
  wire [3:0]        memRequest_bits_data_lo_131 = {memRequest_bits_data_lo_hi_131, memRequest_bits_data_lo_lo_131};
  wire [1:0]        memRequest_bits_data_hi_lo_131 = {_memRequest_bits_data_T_3975[123], _memRequest_bits_data_T_3590[123]};
  wire [1:0]        memRequest_bits_data_hi_hi_131 = {_memRequest_bits_data_T_4745[123], _memRequest_bits_data_T_4360[123]};
  wire [3:0]        memRequest_bits_data_hi_131 = {memRequest_bits_data_hi_hi_131, memRequest_bits_data_hi_lo_131};
  wire [1:0]        memRequest_bits_data_lo_lo_132 = {_memRequest_bits_data_T_2435[124], _memRequest_bits_data_T_2050[124]};
  wire [1:0]        memRequest_bits_data_lo_hi_132 = {_memRequest_bits_data_T_3205[124], _memRequest_bits_data_T_2820[124]};
  wire [3:0]        memRequest_bits_data_lo_132 = {memRequest_bits_data_lo_hi_132, memRequest_bits_data_lo_lo_132};
  wire [1:0]        memRequest_bits_data_hi_lo_132 = {_memRequest_bits_data_T_3975[124], _memRequest_bits_data_T_3590[124]};
  wire [1:0]        memRequest_bits_data_hi_hi_132 = {_memRequest_bits_data_T_4745[124], _memRequest_bits_data_T_4360[124]};
  wire [3:0]        memRequest_bits_data_hi_132 = {memRequest_bits_data_hi_hi_132, memRequest_bits_data_hi_lo_132};
  wire [1:0]        memRequest_bits_data_lo_lo_133 = {_memRequest_bits_data_T_2435[125], _memRequest_bits_data_T_2050[125]};
  wire [1:0]        memRequest_bits_data_lo_hi_133 = {_memRequest_bits_data_T_3205[125], _memRequest_bits_data_T_2820[125]};
  wire [3:0]        memRequest_bits_data_lo_133 = {memRequest_bits_data_lo_hi_133, memRequest_bits_data_lo_lo_133};
  wire [1:0]        memRequest_bits_data_hi_lo_133 = {_memRequest_bits_data_T_3975[125], _memRequest_bits_data_T_3590[125]};
  wire [1:0]        memRequest_bits_data_hi_hi_133 = {_memRequest_bits_data_T_4745[125], _memRequest_bits_data_T_4360[125]};
  wire [3:0]        memRequest_bits_data_hi_133 = {memRequest_bits_data_hi_hi_133, memRequest_bits_data_hi_lo_133};
  wire [1:0]        memRequest_bits_data_lo_lo_134 = {_memRequest_bits_data_T_2435[126], _memRequest_bits_data_T_2050[126]};
  wire [1:0]        memRequest_bits_data_lo_hi_134 = {_memRequest_bits_data_T_3205[126], _memRequest_bits_data_T_2820[126]};
  wire [3:0]        memRequest_bits_data_lo_134 = {memRequest_bits_data_lo_hi_134, memRequest_bits_data_lo_lo_134};
  wire [1:0]        memRequest_bits_data_hi_lo_134 = {_memRequest_bits_data_T_3975[126], _memRequest_bits_data_T_3590[126]};
  wire [1:0]        memRequest_bits_data_hi_hi_134 = {_memRequest_bits_data_T_4745[126], _memRequest_bits_data_T_4360[126]};
  wire [3:0]        memRequest_bits_data_hi_134 = {memRequest_bits_data_hi_hi_134, memRequest_bits_data_hi_lo_134};
  wire [1:0]        memRequest_bits_data_lo_lo_135 = {_memRequest_bits_data_T_2435[127], _memRequest_bits_data_T_2050[127]};
  wire [1:0]        memRequest_bits_data_lo_hi_135 = {_memRequest_bits_data_T_3205[127], _memRequest_bits_data_T_2820[127]};
  wire [3:0]        memRequest_bits_data_lo_135 = {memRequest_bits_data_lo_hi_135, memRequest_bits_data_lo_lo_135};
  wire [1:0]        memRequest_bits_data_hi_lo_135 = {_memRequest_bits_data_T_3975[127], _memRequest_bits_data_T_3590[127]};
  wire [1:0]        memRequest_bits_data_hi_hi_135 = {_memRequest_bits_data_T_4745[127], _memRequest_bits_data_T_4360[127]};
  wire [3:0]        memRequest_bits_data_hi_135 = {memRequest_bits_data_hi_hi_135, memRequest_bits_data_hi_lo_135};
  wire [1:0]        memRequest_bits_data_lo_lo_136 = {_memRequest_bits_data_T_2435[128], _memRequest_bits_data_T_2050[128]};
  wire [1:0]        memRequest_bits_data_lo_hi_136 = {_memRequest_bits_data_T_3205[128], _memRequest_bits_data_T_2820[128]};
  wire [3:0]        memRequest_bits_data_lo_136 = {memRequest_bits_data_lo_hi_136, memRequest_bits_data_lo_lo_136};
  wire [1:0]        memRequest_bits_data_hi_lo_136 = {_memRequest_bits_data_T_3975[128], _memRequest_bits_data_T_3590[128]};
  wire [1:0]        memRequest_bits_data_hi_hi_136 = {_memRequest_bits_data_T_4745[128], _memRequest_bits_data_T_4360[128]};
  wire [3:0]        memRequest_bits_data_hi_136 = {memRequest_bits_data_hi_hi_136, memRequest_bits_data_hi_lo_136};
  wire [1:0]        memRequest_bits_data_lo_lo_137 = {_memRequest_bits_data_T_2435[129], _memRequest_bits_data_T_2050[129]};
  wire [1:0]        memRequest_bits_data_lo_hi_137 = {_memRequest_bits_data_T_3205[129], _memRequest_bits_data_T_2820[129]};
  wire [3:0]        memRequest_bits_data_lo_137 = {memRequest_bits_data_lo_hi_137, memRequest_bits_data_lo_lo_137};
  wire [1:0]        memRequest_bits_data_hi_lo_137 = {_memRequest_bits_data_T_3975[129], _memRequest_bits_data_T_3590[129]};
  wire [1:0]        memRequest_bits_data_hi_hi_137 = {_memRequest_bits_data_T_4745[129], _memRequest_bits_data_T_4360[129]};
  wire [3:0]        memRequest_bits_data_hi_137 = {memRequest_bits_data_hi_hi_137, memRequest_bits_data_hi_lo_137};
  wire [1:0]        memRequest_bits_data_lo_lo_138 = {_memRequest_bits_data_T_2435[130], _memRequest_bits_data_T_2050[130]};
  wire [1:0]        memRequest_bits_data_lo_hi_138 = {_memRequest_bits_data_T_3205[130], _memRequest_bits_data_T_2820[130]};
  wire [3:0]        memRequest_bits_data_lo_138 = {memRequest_bits_data_lo_hi_138, memRequest_bits_data_lo_lo_138};
  wire [1:0]        memRequest_bits_data_hi_lo_138 = {_memRequest_bits_data_T_3975[130], _memRequest_bits_data_T_3590[130]};
  wire [1:0]        memRequest_bits_data_hi_hi_138 = {_memRequest_bits_data_T_4745[130], _memRequest_bits_data_T_4360[130]};
  wire [3:0]        memRequest_bits_data_hi_138 = {memRequest_bits_data_hi_hi_138, memRequest_bits_data_hi_lo_138};
  wire [1:0]        memRequest_bits_data_lo_lo_139 = {_memRequest_bits_data_T_2435[131], _memRequest_bits_data_T_2050[131]};
  wire [1:0]        memRequest_bits_data_lo_hi_139 = {_memRequest_bits_data_T_3205[131], _memRequest_bits_data_T_2820[131]};
  wire [3:0]        memRequest_bits_data_lo_139 = {memRequest_bits_data_lo_hi_139, memRequest_bits_data_lo_lo_139};
  wire [1:0]        memRequest_bits_data_hi_lo_139 = {_memRequest_bits_data_T_3975[131], _memRequest_bits_data_T_3590[131]};
  wire [1:0]        memRequest_bits_data_hi_hi_139 = {_memRequest_bits_data_T_4745[131], _memRequest_bits_data_T_4360[131]};
  wire [3:0]        memRequest_bits_data_hi_139 = {memRequest_bits_data_hi_hi_139, memRequest_bits_data_hi_lo_139};
  wire [1:0]        memRequest_bits_data_lo_lo_140 = {_memRequest_bits_data_T_2435[132], _memRequest_bits_data_T_2050[132]};
  wire [1:0]        memRequest_bits_data_lo_hi_140 = {_memRequest_bits_data_T_3205[132], _memRequest_bits_data_T_2820[132]};
  wire [3:0]        memRequest_bits_data_lo_140 = {memRequest_bits_data_lo_hi_140, memRequest_bits_data_lo_lo_140};
  wire [1:0]        memRequest_bits_data_hi_lo_140 = {_memRequest_bits_data_T_3975[132], _memRequest_bits_data_T_3590[132]};
  wire [1:0]        memRequest_bits_data_hi_hi_140 = {_memRequest_bits_data_T_4745[132], _memRequest_bits_data_T_4360[132]};
  wire [3:0]        memRequest_bits_data_hi_140 = {memRequest_bits_data_hi_hi_140, memRequest_bits_data_hi_lo_140};
  wire [1:0]        memRequest_bits_data_lo_lo_141 = {_memRequest_bits_data_T_2435[133], _memRequest_bits_data_T_2050[133]};
  wire [1:0]        memRequest_bits_data_lo_hi_141 = {_memRequest_bits_data_T_3205[133], _memRequest_bits_data_T_2820[133]};
  wire [3:0]        memRequest_bits_data_lo_141 = {memRequest_bits_data_lo_hi_141, memRequest_bits_data_lo_lo_141};
  wire [1:0]        memRequest_bits_data_hi_lo_141 = {_memRequest_bits_data_T_3975[133], _memRequest_bits_data_T_3590[133]};
  wire [1:0]        memRequest_bits_data_hi_hi_141 = {_memRequest_bits_data_T_4745[133], _memRequest_bits_data_T_4360[133]};
  wire [3:0]        memRequest_bits_data_hi_141 = {memRequest_bits_data_hi_hi_141, memRequest_bits_data_hi_lo_141};
  wire [1:0]        memRequest_bits_data_lo_lo_142 = {_memRequest_bits_data_T_2435[134], _memRequest_bits_data_T_2050[134]};
  wire [1:0]        memRequest_bits_data_lo_hi_142 = {_memRequest_bits_data_T_3205[134], _memRequest_bits_data_T_2820[134]};
  wire [3:0]        memRequest_bits_data_lo_142 = {memRequest_bits_data_lo_hi_142, memRequest_bits_data_lo_lo_142};
  wire [1:0]        memRequest_bits_data_hi_lo_142 = {_memRequest_bits_data_T_3975[134], _memRequest_bits_data_T_3590[134]};
  wire [1:0]        memRequest_bits_data_hi_hi_142 = {_memRequest_bits_data_T_4745[134], _memRequest_bits_data_T_4360[134]};
  wire [3:0]        memRequest_bits_data_hi_142 = {memRequest_bits_data_hi_hi_142, memRequest_bits_data_hi_lo_142};
  wire [1:0]        memRequest_bits_data_lo_lo_143 = {_memRequest_bits_data_T_2435[135], _memRequest_bits_data_T_2050[135]};
  wire [1:0]        memRequest_bits_data_lo_hi_143 = {_memRequest_bits_data_T_3205[135], _memRequest_bits_data_T_2820[135]};
  wire [3:0]        memRequest_bits_data_lo_143 = {memRequest_bits_data_lo_hi_143, memRequest_bits_data_lo_lo_143};
  wire [1:0]        memRequest_bits_data_hi_lo_143 = {_memRequest_bits_data_T_3975[135], _memRequest_bits_data_T_3590[135]};
  wire [1:0]        memRequest_bits_data_hi_hi_143 = {_memRequest_bits_data_T_4745[135], _memRequest_bits_data_T_4360[135]};
  wire [3:0]        memRequest_bits_data_hi_143 = {memRequest_bits_data_hi_hi_143, memRequest_bits_data_hi_lo_143};
  wire [1:0]        memRequest_bits_data_lo_lo_144 = {_memRequest_bits_data_T_2435[136], _memRequest_bits_data_T_2050[136]};
  wire [1:0]        memRequest_bits_data_lo_hi_144 = {_memRequest_bits_data_T_3205[136], _memRequest_bits_data_T_2820[136]};
  wire [3:0]        memRequest_bits_data_lo_144 = {memRequest_bits_data_lo_hi_144, memRequest_bits_data_lo_lo_144};
  wire [1:0]        memRequest_bits_data_hi_lo_144 = {_memRequest_bits_data_T_3975[136], _memRequest_bits_data_T_3590[136]};
  wire [1:0]        memRequest_bits_data_hi_hi_144 = {_memRequest_bits_data_T_4745[136], _memRequest_bits_data_T_4360[136]};
  wire [3:0]        memRequest_bits_data_hi_144 = {memRequest_bits_data_hi_hi_144, memRequest_bits_data_hi_lo_144};
  wire [1:0]        memRequest_bits_data_lo_lo_145 = {_memRequest_bits_data_T_2435[137], _memRequest_bits_data_T_2050[137]};
  wire [1:0]        memRequest_bits_data_lo_hi_145 = {_memRequest_bits_data_T_3205[137], _memRequest_bits_data_T_2820[137]};
  wire [3:0]        memRequest_bits_data_lo_145 = {memRequest_bits_data_lo_hi_145, memRequest_bits_data_lo_lo_145};
  wire [1:0]        memRequest_bits_data_hi_lo_145 = {_memRequest_bits_data_T_3975[137], _memRequest_bits_data_T_3590[137]};
  wire [1:0]        memRequest_bits_data_hi_hi_145 = {_memRequest_bits_data_T_4745[137], _memRequest_bits_data_T_4360[137]};
  wire [3:0]        memRequest_bits_data_hi_145 = {memRequest_bits_data_hi_hi_145, memRequest_bits_data_hi_lo_145};
  wire [1:0]        memRequest_bits_data_lo_lo_146 = {_memRequest_bits_data_T_2435[138], _memRequest_bits_data_T_2050[138]};
  wire [1:0]        memRequest_bits_data_lo_hi_146 = {_memRequest_bits_data_T_3205[138], _memRequest_bits_data_T_2820[138]};
  wire [3:0]        memRequest_bits_data_lo_146 = {memRequest_bits_data_lo_hi_146, memRequest_bits_data_lo_lo_146};
  wire [1:0]        memRequest_bits_data_hi_lo_146 = {_memRequest_bits_data_T_3975[138], _memRequest_bits_data_T_3590[138]};
  wire [1:0]        memRequest_bits_data_hi_hi_146 = {_memRequest_bits_data_T_4745[138], _memRequest_bits_data_T_4360[138]};
  wire [3:0]        memRequest_bits_data_hi_146 = {memRequest_bits_data_hi_hi_146, memRequest_bits_data_hi_lo_146};
  wire [1:0]        memRequest_bits_data_lo_lo_147 = {_memRequest_bits_data_T_2435[139], _memRequest_bits_data_T_2050[139]};
  wire [1:0]        memRequest_bits_data_lo_hi_147 = {_memRequest_bits_data_T_3205[139], _memRequest_bits_data_T_2820[139]};
  wire [3:0]        memRequest_bits_data_lo_147 = {memRequest_bits_data_lo_hi_147, memRequest_bits_data_lo_lo_147};
  wire [1:0]        memRequest_bits_data_hi_lo_147 = {_memRequest_bits_data_T_3975[139], _memRequest_bits_data_T_3590[139]};
  wire [1:0]        memRequest_bits_data_hi_hi_147 = {_memRequest_bits_data_T_4745[139], _memRequest_bits_data_T_4360[139]};
  wire [3:0]        memRequest_bits_data_hi_147 = {memRequest_bits_data_hi_hi_147, memRequest_bits_data_hi_lo_147};
  wire [1:0]        memRequest_bits_data_lo_lo_148 = {_memRequest_bits_data_T_2435[140], _memRequest_bits_data_T_2050[140]};
  wire [1:0]        memRequest_bits_data_lo_hi_148 = {_memRequest_bits_data_T_3205[140], _memRequest_bits_data_T_2820[140]};
  wire [3:0]        memRequest_bits_data_lo_148 = {memRequest_bits_data_lo_hi_148, memRequest_bits_data_lo_lo_148};
  wire [1:0]        memRequest_bits_data_hi_lo_148 = {_memRequest_bits_data_T_3975[140], _memRequest_bits_data_T_3590[140]};
  wire [1:0]        memRequest_bits_data_hi_hi_148 = {_memRequest_bits_data_T_4745[140], _memRequest_bits_data_T_4360[140]};
  wire [3:0]        memRequest_bits_data_hi_148 = {memRequest_bits_data_hi_hi_148, memRequest_bits_data_hi_lo_148};
  wire [1:0]        memRequest_bits_data_lo_lo_149 = {_memRequest_bits_data_T_2435[141], _memRequest_bits_data_T_2050[141]};
  wire [1:0]        memRequest_bits_data_lo_hi_149 = {_memRequest_bits_data_T_3205[141], _memRequest_bits_data_T_2820[141]};
  wire [3:0]        memRequest_bits_data_lo_149 = {memRequest_bits_data_lo_hi_149, memRequest_bits_data_lo_lo_149};
  wire [1:0]        memRequest_bits_data_hi_lo_149 = {_memRequest_bits_data_T_3975[141], _memRequest_bits_data_T_3590[141]};
  wire [1:0]        memRequest_bits_data_hi_hi_149 = {_memRequest_bits_data_T_4745[141], _memRequest_bits_data_T_4360[141]};
  wire [3:0]        memRequest_bits_data_hi_149 = {memRequest_bits_data_hi_hi_149, memRequest_bits_data_hi_lo_149};
  wire [1:0]        memRequest_bits_data_lo_lo_150 = {_memRequest_bits_data_T_2435[142], _memRequest_bits_data_T_2050[142]};
  wire [1:0]        memRequest_bits_data_lo_hi_150 = {_memRequest_bits_data_T_3205[142], _memRequest_bits_data_T_2820[142]};
  wire [3:0]        memRequest_bits_data_lo_150 = {memRequest_bits_data_lo_hi_150, memRequest_bits_data_lo_lo_150};
  wire [1:0]        memRequest_bits_data_hi_lo_150 = {_memRequest_bits_data_T_3975[142], _memRequest_bits_data_T_3590[142]};
  wire [1:0]        memRequest_bits_data_hi_hi_150 = {_memRequest_bits_data_T_4745[142], _memRequest_bits_data_T_4360[142]};
  wire [3:0]        memRequest_bits_data_hi_150 = {memRequest_bits_data_hi_hi_150, memRequest_bits_data_hi_lo_150};
  wire [1:0]        memRequest_bits_data_lo_lo_151 = {_memRequest_bits_data_T_2435[143], _memRequest_bits_data_T_2050[143]};
  wire [1:0]        memRequest_bits_data_lo_hi_151 = {_memRequest_bits_data_T_3205[143], _memRequest_bits_data_T_2820[143]};
  wire [3:0]        memRequest_bits_data_lo_151 = {memRequest_bits_data_lo_hi_151, memRequest_bits_data_lo_lo_151};
  wire [1:0]        memRequest_bits_data_hi_lo_151 = {_memRequest_bits_data_T_3975[143], _memRequest_bits_data_T_3590[143]};
  wire [1:0]        memRequest_bits_data_hi_hi_151 = {_memRequest_bits_data_T_4745[143], _memRequest_bits_data_T_4360[143]};
  wire [3:0]        memRequest_bits_data_hi_151 = {memRequest_bits_data_hi_hi_151, memRequest_bits_data_hi_lo_151};
  wire [1:0]        memRequest_bits_data_lo_lo_152 = {_memRequest_bits_data_T_2435[144], _memRequest_bits_data_T_2050[144]};
  wire [1:0]        memRequest_bits_data_lo_hi_152 = {_memRequest_bits_data_T_3205[144], _memRequest_bits_data_T_2820[144]};
  wire [3:0]        memRequest_bits_data_lo_152 = {memRequest_bits_data_lo_hi_152, memRequest_bits_data_lo_lo_152};
  wire [1:0]        memRequest_bits_data_hi_lo_152 = {_memRequest_bits_data_T_3975[144], _memRequest_bits_data_T_3590[144]};
  wire [1:0]        memRequest_bits_data_hi_hi_152 = {_memRequest_bits_data_T_4745[144], _memRequest_bits_data_T_4360[144]};
  wire [3:0]        memRequest_bits_data_hi_152 = {memRequest_bits_data_hi_hi_152, memRequest_bits_data_hi_lo_152};
  wire [1:0]        memRequest_bits_data_lo_lo_153 = {_memRequest_bits_data_T_2435[145], _memRequest_bits_data_T_2050[145]};
  wire [1:0]        memRequest_bits_data_lo_hi_153 = {_memRequest_bits_data_T_3205[145], _memRequest_bits_data_T_2820[145]};
  wire [3:0]        memRequest_bits_data_lo_153 = {memRequest_bits_data_lo_hi_153, memRequest_bits_data_lo_lo_153};
  wire [1:0]        memRequest_bits_data_hi_lo_153 = {_memRequest_bits_data_T_3975[145], _memRequest_bits_data_T_3590[145]};
  wire [1:0]        memRequest_bits_data_hi_hi_153 = {_memRequest_bits_data_T_4745[145], _memRequest_bits_data_T_4360[145]};
  wire [3:0]        memRequest_bits_data_hi_153 = {memRequest_bits_data_hi_hi_153, memRequest_bits_data_hi_lo_153};
  wire [1:0]        memRequest_bits_data_lo_lo_154 = {_memRequest_bits_data_T_2435[146], _memRequest_bits_data_T_2050[146]};
  wire [1:0]        memRequest_bits_data_lo_hi_154 = {_memRequest_bits_data_T_3205[146], _memRequest_bits_data_T_2820[146]};
  wire [3:0]        memRequest_bits_data_lo_154 = {memRequest_bits_data_lo_hi_154, memRequest_bits_data_lo_lo_154};
  wire [1:0]        memRequest_bits_data_hi_lo_154 = {_memRequest_bits_data_T_3975[146], _memRequest_bits_data_T_3590[146]};
  wire [1:0]        memRequest_bits_data_hi_hi_154 = {_memRequest_bits_data_T_4745[146], _memRequest_bits_data_T_4360[146]};
  wire [3:0]        memRequest_bits_data_hi_154 = {memRequest_bits_data_hi_hi_154, memRequest_bits_data_hi_lo_154};
  wire [1:0]        memRequest_bits_data_lo_lo_155 = {_memRequest_bits_data_T_2435[147], _memRequest_bits_data_T_2050[147]};
  wire [1:0]        memRequest_bits_data_lo_hi_155 = {_memRequest_bits_data_T_3205[147], _memRequest_bits_data_T_2820[147]};
  wire [3:0]        memRequest_bits_data_lo_155 = {memRequest_bits_data_lo_hi_155, memRequest_bits_data_lo_lo_155};
  wire [1:0]        memRequest_bits_data_hi_lo_155 = {_memRequest_bits_data_T_3975[147], _memRequest_bits_data_T_3590[147]};
  wire [1:0]        memRequest_bits_data_hi_hi_155 = {_memRequest_bits_data_T_4745[147], _memRequest_bits_data_T_4360[147]};
  wire [3:0]        memRequest_bits_data_hi_155 = {memRequest_bits_data_hi_hi_155, memRequest_bits_data_hi_lo_155};
  wire [1:0]        memRequest_bits_data_lo_lo_156 = {_memRequest_bits_data_T_2435[148], _memRequest_bits_data_T_2050[148]};
  wire [1:0]        memRequest_bits_data_lo_hi_156 = {_memRequest_bits_data_T_3205[148], _memRequest_bits_data_T_2820[148]};
  wire [3:0]        memRequest_bits_data_lo_156 = {memRequest_bits_data_lo_hi_156, memRequest_bits_data_lo_lo_156};
  wire [1:0]        memRequest_bits_data_hi_lo_156 = {_memRequest_bits_data_T_3975[148], _memRequest_bits_data_T_3590[148]};
  wire [1:0]        memRequest_bits_data_hi_hi_156 = {_memRequest_bits_data_T_4745[148], _memRequest_bits_data_T_4360[148]};
  wire [3:0]        memRequest_bits_data_hi_156 = {memRequest_bits_data_hi_hi_156, memRequest_bits_data_hi_lo_156};
  wire [1:0]        memRequest_bits_data_lo_lo_157 = {_memRequest_bits_data_T_2435[149], _memRequest_bits_data_T_2050[149]};
  wire [1:0]        memRequest_bits_data_lo_hi_157 = {_memRequest_bits_data_T_3205[149], _memRequest_bits_data_T_2820[149]};
  wire [3:0]        memRequest_bits_data_lo_157 = {memRequest_bits_data_lo_hi_157, memRequest_bits_data_lo_lo_157};
  wire [1:0]        memRequest_bits_data_hi_lo_157 = {_memRequest_bits_data_T_3975[149], _memRequest_bits_data_T_3590[149]};
  wire [1:0]        memRequest_bits_data_hi_hi_157 = {_memRequest_bits_data_T_4745[149], _memRequest_bits_data_T_4360[149]};
  wire [3:0]        memRequest_bits_data_hi_157 = {memRequest_bits_data_hi_hi_157, memRequest_bits_data_hi_lo_157};
  wire [1:0]        memRequest_bits_data_lo_lo_158 = {_memRequest_bits_data_T_2435[150], _memRequest_bits_data_T_2050[150]};
  wire [1:0]        memRequest_bits_data_lo_hi_158 = {_memRequest_bits_data_T_3205[150], _memRequest_bits_data_T_2820[150]};
  wire [3:0]        memRequest_bits_data_lo_158 = {memRequest_bits_data_lo_hi_158, memRequest_bits_data_lo_lo_158};
  wire [1:0]        memRequest_bits_data_hi_lo_158 = {_memRequest_bits_data_T_3975[150], _memRequest_bits_data_T_3590[150]};
  wire [1:0]        memRequest_bits_data_hi_hi_158 = {_memRequest_bits_data_T_4745[150], _memRequest_bits_data_T_4360[150]};
  wire [3:0]        memRequest_bits_data_hi_158 = {memRequest_bits_data_hi_hi_158, memRequest_bits_data_hi_lo_158};
  wire [1:0]        memRequest_bits_data_lo_lo_159 = {_memRequest_bits_data_T_2435[151], _memRequest_bits_data_T_2050[151]};
  wire [1:0]        memRequest_bits_data_lo_hi_159 = {_memRequest_bits_data_T_3205[151], _memRequest_bits_data_T_2820[151]};
  wire [3:0]        memRequest_bits_data_lo_159 = {memRequest_bits_data_lo_hi_159, memRequest_bits_data_lo_lo_159};
  wire [1:0]        memRequest_bits_data_hi_lo_159 = {_memRequest_bits_data_T_3975[151], _memRequest_bits_data_T_3590[151]};
  wire [1:0]        memRequest_bits_data_hi_hi_159 = {_memRequest_bits_data_T_4745[151], _memRequest_bits_data_T_4360[151]};
  wire [3:0]        memRequest_bits_data_hi_159 = {memRequest_bits_data_hi_hi_159, memRequest_bits_data_hi_lo_159};
  wire [1:0]        memRequest_bits_data_lo_lo_160 = {_memRequest_bits_data_T_2435[152], _memRequest_bits_data_T_2050[152]};
  wire [1:0]        memRequest_bits_data_lo_hi_160 = {_memRequest_bits_data_T_3205[152], _memRequest_bits_data_T_2820[152]};
  wire [3:0]        memRequest_bits_data_lo_160 = {memRequest_bits_data_lo_hi_160, memRequest_bits_data_lo_lo_160};
  wire [1:0]        memRequest_bits_data_hi_lo_160 = {_memRequest_bits_data_T_3975[152], _memRequest_bits_data_T_3590[152]};
  wire [1:0]        memRequest_bits_data_hi_hi_160 = {_memRequest_bits_data_T_4745[152], _memRequest_bits_data_T_4360[152]};
  wire [3:0]        memRequest_bits_data_hi_160 = {memRequest_bits_data_hi_hi_160, memRequest_bits_data_hi_lo_160};
  wire [1:0]        memRequest_bits_data_lo_lo_161 = {_memRequest_bits_data_T_2435[153], _memRequest_bits_data_T_2050[153]};
  wire [1:0]        memRequest_bits_data_lo_hi_161 = {_memRequest_bits_data_T_3205[153], _memRequest_bits_data_T_2820[153]};
  wire [3:0]        memRequest_bits_data_lo_161 = {memRequest_bits_data_lo_hi_161, memRequest_bits_data_lo_lo_161};
  wire [1:0]        memRequest_bits_data_hi_lo_161 = {_memRequest_bits_data_T_3975[153], _memRequest_bits_data_T_3590[153]};
  wire [1:0]        memRequest_bits_data_hi_hi_161 = {_memRequest_bits_data_T_4745[153], _memRequest_bits_data_T_4360[153]};
  wire [3:0]        memRequest_bits_data_hi_161 = {memRequest_bits_data_hi_hi_161, memRequest_bits_data_hi_lo_161};
  wire [1:0]        memRequest_bits_data_lo_lo_162 = {_memRequest_bits_data_T_2435[154], _memRequest_bits_data_T_2050[154]};
  wire [1:0]        memRequest_bits_data_lo_hi_162 = {_memRequest_bits_data_T_3205[154], _memRequest_bits_data_T_2820[154]};
  wire [3:0]        memRequest_bits_data_lo_162 = {memRequest_bits_data_lo_hi_162, memRequest_bits_data_lo_lo_162};
  wire [1:0]        memRequest_bits_data_hi_lo_162 = {_memRequest_bits_data_T_3975[154], _memRequest_bits_data_T_3590[154]};
  wire [1:0]        memRequest_bits_data_hi_hi_162 = {_memRequest_bits_data_T_4745[154], _memRequest_bits_data_T_4360[154]};
  wire [3:0]        memRequest_bits_data_hi_162 = {memRequest_bits_data_hi_hi_162, memRequest_bits_data_hi_lo_162};
  wire [1:0]        memRequest_bits_data_lo_lo_163 = {_memRequest_bits_data_T_2435[155], _memRequest_bits_data_T_2050[155]};
  wire [1:0]        memRequest_bits_data_lo_hi_163 = {_memRequest_bits_data_T_3205[155], _memRequest_bits_data_T_2820[155]};
  wire [3:0]        memRequest_bits_data_lo_163 = {memRequest_bits_data_lo_hi_163, memRequest_bits_data_lo_lo_163};
  wire [1:0]        memRequest_bits_data_hi_lo_163 = {_memRequest_bits_data_T_3975[155], _memRequest_bits_data_T_3590[155]};
  wire [1:0]        memRequest_bits_data_hi_hi_163 = {_memRequest_bits_data_T_4745[155], _memRequest_bits_data_T_4360[155]};
  wire [3:0]        memRequest_bits_data_hi_163 = {memRequest_bits_data_hi_hi_163, memRequest_bits_data_hi_lo_163};
  wire [1:0]        memRequest_bits_data_lo_lo_164 = {_memRequest_bits_data_T_2435[156], _memRequest_bits_data_T_2050[156]};
  wire [1:0]        memRequest_bits_data_lo_hi_164 = {_memRequest_bits_data_T_3205[156], _memRequest_bits_data_T_2820[156]};
  wire [3:0]        memRequest_bits_data_lo_164 = {memRequest_bits_data_lo_hi_164, memRequest_bits_data_lo_lo_164};
  wire [1:0]        memRequest_bits_data_hi_lo_164 = {_memRequest_bits_data_T_3975[156], _memRequest_bits_data_T_3590[156]};
  wire [1:0]        memRequest_bits_data_hi_hi_164 = {_memRequest_bits_data_T_4745[156], _memRequest_bits_data_T_4360[156]};
  wire [3:0]        memRequest_bits_data_hi_164 = {memRequest_bits_data_hi_hi_164, memRequest_bits_data_hi_lo_164};
  wire [1:0]        memRequest_bits_data_lo_lo_165 = {_memRequest_bits_data_T_2435[157], _memRequest_bits_data_T_2050[157]};
  wire [1:0]        memRequest_bits_data_lo_hi_165 = {_memRequest_bits_data_T_3205[157], _memRequest_bits_data_T_2820[157]};
  wire [3:0]        memRequest_bits_data_lo_165 = {memRequest_bits_data_lo_hi_165, memRequest_bits_data_lo_lo_165};
  wire [1:0]        memRequest_bits_data_hi_lo_165 = {_memRequest_bits_data_T_3975[157], _memRequest_bits_data_T_3590[157]};
  wire [1:0]        memRequest_bits_data_hi_hi_165 = {_memRequest_bits_data_T_4745[157], _memRequest_bits_data_T_4360[157]};
  wire [3:0]        memRequest_bits_data_hi_165 = {memRequest_bits_data_hi_hi_165, memRequest_bits_data_hi_lo_165};
  wire [1:0]        memRequest_bits_data_lo_lo_166 = {_memRequest_bits_data_T_2435[158], _memRequest_bits_data_T_2050[158]};
  wire [1:0]        memRequest_bits_data_lo_hi_166 = {_memRequest_bits_data_T_3205[158], _memRequest_bits_data_T_2820[158]};
  wire [3:0]        memRequest_bits_data_lo_166 = {memRequest_bits_data_lo_hi_166, memRequest_bits_data_lo_lo_166};
  wire [1:0]        memRequest_bits_data_hi_lo_166 = {_memRequest_bits_data_T_3975[158], _memRequest_bits_data_T_3590[158]};
  wire [1:0]        memRequest_bits_data_hi_hi_166 = {_memRequest_bits_data_T_4745[158], _memRequest_bits_data_T_4360[158]};
  wire [3:0]        memRequest_bits_data_hi_166 = {memRequest_bits_data_hi_hi_166, memRequest_bits_data_hi_lo_166};
  wire [1:0]        memRequest_bits_data_lo_lo_167 = {_memRequest_bits_data_T_2435[159], _memRequest_bits_data_T_2050[159]};
  wire [1:0]        memRequest_bits_data_lo_hi_167 = {_memRequest_bits_data_T_3205[159], _memRequest_bits_data_T_2820[159]};
  wire [3:0]        memRequest_bits_data_lo_167 = {memRequest_bits_data_lo_hi_167, memRequest_bits_data_lo_lo_167};
  wire [1:0]        memRequest_bits_data_hi_lo_167 = {_memRequest_bits_data_T_3975[159], _memRequest_bits_data_T_3590[159]};
  wire [1:0]        memRequest_bits_data_hi_hi_167 = {_memRequest_bits_data_T_4745[159], _memRequest_bits_data_T_4360[159]};
  wire [3:0]        memRequest_bits_data_hi_167 = {memRequest_bits_data_hi_hi_167, memRequest_bits_data_hi_lo_167};
  wire [1:0]        memRequest_bits_data_lo_lo_168 = {_memRequest_bits_data_T_2435[160], _memRequest_bits_data_T_2050[160]};
  wire [1:0]        memRequest_bits_data_lo_hi_168 = {_memRequest_bits_data_T_3205[160], _memRequest_bits_data_T_2820[160]};
  wire [3:0]        memRequest_bits_data_lo_168 = {memRequest_bits_data_lo_hi_168, memRequest_bits_data_lo_lo_168};
  wire [1:0]        memRequest_bits_data_hi_lo_168 = {_memRequest_bits_data_T_3975[160], _memRequest_bits_data_T_3590[160]};
  wire [1:0]        memRequest_bits_data_hi_hi_168 = {_memRequest_bits_data_T_4745[160], _memRequest_bits_data_T_4360[160]};
  wire [3:0]        memRequest_bits_data_hi_168 = {memRequest_bits_data_hi_hi_168, memRequest_bits_data_hi_lo_168};
  wire [1:0]        memRequest_bits_data_lo_lo_169 = {_memRequest_bits_data_T_2435[161], _memRequest_bits_data_T_2050[161]};
  wire [1:0]        memRequest_bits_data_lo_hi_169 = {_memRequest_bits_data_T_3205[161], _memRequest_bits_data_T_2820[161]};
  wire [3:0]        memRequest_bits_data_lo_169 = {memRequest_bits_data_lo_hi_169, memRequest_bits_data_lo_lo_169};
  wire [1:0]        memRequest_bits_data_hi_lo_169 = {_memRequest_bits_data_T_3975[161], _memRequest_bits_data_T_3590[161]};
  wire [1:0]        memRequest_bits_data_hi_hi_169 = {_memRequest_bits_data_T_4745[161], _memRequest_bits_data_T_4360[161]};
  wire [3:0]        memRequest_bits_data_hi_169 = {memRequest_bits_data_hi_hi_169, memRequest_bits_data_hi_lo_169};
  wire [1:0]        memRequest_bits_data_lo_lo_170 = {_memRequest_bits_data_T_2435[162], _memRequest_bits_data_T_2050[162]};
  wire [1:0]        memRequest_bits_data_lo_hi_170 = {_memRequest_bits_data_T_3205[162], _memRequest_bits_data_T_2820[162]};
  wire [3:0]        memRequest_bits_data_lo_170 = {memRequest_bits_data_lo_hi_170, memRequest_bits_data_lo_lo_170};
  wire [1:0]        memRequest_bits_data_hi_lo_170 = {_memRequest_bits_data_T_3975[162], _memRequest_bits_data_T_3590[162]};
  wire [1:0]        memRequest_bits_data_hi_hi_170 = {_memRequest_bits_data_T_4745[162], _memRequest_bits_data_T_4360[162]};
  wire [3:0]        memRequest_bits_data_hi_170 = {memRequest_bits_data_hi_hi_170, memRequest_bits_data_hi_lo_170};
  wire [1:0]        memRequest_bits_data_lo_lo_171 = {_memRequest_bits_data_T_2435[163], _memRequest_bits_data_T_2050[163]};
  wire [1:0]        memRequest_bits_data_lo_hi_171 = {_memRequest_bits_data_T_3205[163], _memRequest_bits_data_T_2820[163]};
  wire [3:0]        memRequest_bits_data_lo_171 = {memRequest_bits_data_lo_hi_171, memRequest_bits_data_lo_lo_171};
  wire [1:0]        memRequest_bits_data_hi_lo_171 = {_memRequest_bits_data_T_3975[163], _memRequest_bits_data_T_3590[163]};
  wire [1:0]        memRequest_bits_data_hi_hi_171 = {_memRequest_bits_data_T_4745[163], _memRequest_bits_data_T_4360[163]};
  wire [3:0]        memRequest_bits_data_hi_171 = {memRequest_bits_data_hi_hi_171, memRequest_bits_data_hi_lo_171};
  wire [1:0]        memRequest_bits_data_lo_lo_172 = {_memRequest_bits_data_T_2435[164], _memRequest_bits_data_T_2050[164]};
  wire [1:0]        memRequest_bits_data_lo_hi_172 = {_memRequest_bits_data_T_3205[164], _memRequest_bits_data_T_2820[164]};
  wire [3:0]        memRequest_bits_data_lo_172 = {memRequest_bits_data_lo_hi_172, memRequest_bits_data_lo_lo_172};
  wire [1:0]        memRequest_bits_data_hi_lo_172 = {_memRequest_bits_data_T_3975[164], _memRequest_bits_data_T_3590[164]};
  wire [1:0]        memRequest_bits_data_hi_hi_172 = {_memRequest_bits_data_T_4745[164], _memRequest_bits_data_T_4360[164]};
  wire [3:0]        memRequest_bits_data_hi_172 = {memRequest_bits_data_hi_hi_172, memRequest_bits_data_hi_lo_172};
  wire [1:0]        memRequest_bits_data_lo_lo_173 = {_memRequest_bits_data_T_2435[165], _memRequest_bits_data_T_2050[165]};
  wire [1:0]        memRequest_bits_data_lo_hi_173 = {_memRequest_bits_data_T_3205[165], _memRequest_bits_data_T_2820[165]};
  wire [3:0]        memRequest_bits_data_lo_173 = {memRequest_bits_data_lo_hi_173, memRequest_bits_data_lo_lo_173};
  wire [1:0]        memRequest_bits_data_hi_lo_173 = {_memRequest_bits_data_T_3975[165], _memRequest_bits_data_T_3590[165]};
  wire [1:0]        memRequest_bits_data_hi_hi_173 = {_memRequest_bits_data_T_4745[165], _memRequest_bits_data_T_4360[165]};
  wire [3:0]        memRequest_bits_data_hi_173 = {memRequest_bits_data_hi_hi_173, memRequest_bits_data_hi_lo_173};
  wire [1:0]        memRequest_bits_data_lo_lo_174 = {_memRequest_bits_data_T_2435[166], _memRequest_bits_data_T_2050[166]};
  wire [1:0]        memRequest_bits_data_lo_hi_174 = {_memRequest_bits_data_T_3205[166], _memRequest_bits_data_T_2820[166]};
  wire [3:0]        memRequest_bits_data_lo_174 = {memRequest_bits_data_lo_hi_174, memRequest_bits_data_lo_lo_174};
  wire [1:0]        memRequest_bits_data_hi_lo_174 = {_memRequest_bits_data_T_3975[166], _memRequest_bits_data_T_3590[166]};
  wire [1:0]        memRequest_bits_data_hi_hi_174 = {_memRequest_bits_data_T_4745[166], _memRequest_bits_data_T_4360[166]};
  wire [3:0]        memRequest_bits_data_hi_174 = {memRequest_bits_data_hi_hi_174, memRequest_bits_data_hi_lo_174};
  wire [1:0]        memRequest_bits_data_lo_lo_175 = {_memRequest_bits_data_T_2435[167], _memRequest_bits_data_T_2050[167]};
  wire [1:0]        memRequest_bits_data_lo_hi_175 = {_memRequest_bits_data_T_3205[167], _memRequest_bits_data_T_2820[167]};
  wire [3:0]        memRequest_bits_data_lo_175 = {memRequest_bits_data_lo_hi_175, memRequest_bits_data_lo_lo_175};
  wire [1:0]        memRequest_bits_data_hi_lo_175 = {_memRequest_bits_data_T_3975[167], _memRequest_bits_data_T_3590[167]};
  wire [1:0]        memRequest_bits_data_hi_hi_175 = {_memRequest_bits_data_T_4745[167], _memRequest_bits_data_T_4360[167]};
  wire [3:0]        memRequest_bits_data_hi_175 = {memRequest_bits_data_hi_hi_175, memRequest_bits_data_hi_lo_175};
  wire [1:0]        memRequest_bits_data_lo_lo_176 = {_memRequest_bits_data_T_2435[168], _memRequest_bits_data_T_2050[168]};
  wire [1:0]        memRequest_bits_data_lo_hi_176 = {_memRequest_bits_data_T_3205[168], _memRequest_bits_data_T_2820[168]};
  wire [3:0]        memRequest_bits_data_lo_176 = {memRequest_bits_data_lo_hi_176, memRequest_bits_data_lo_lo_176};
  wire [1:0]        memRequest_bits_data_hi_lo_176 = {_memRequest_bits_data_T_3975[168], _memRequest_bits_data_T_3590[168]};
  wire [1:0]        memRequest_bits_data_hi_hi_176 = {_memRequest_bits_data_T_4745[168], _memRequest_bits_data_T_4360[168]};
  wire [3:0]        memRequest_bits_data_hi_176 = {memRequest_bits_data_hi_hi_176, memRequest_bits_data_hi_lo_176};
  wire [1:0]        memRequest_bits_data_lo_lo_177 = {_memRequest_bits_data_T_2435[169], _memRequest_bits_data_T_2050[169]};
  wire [1:0]        memRequest_bits_data_lo_hi_177 = {_memRequest_bits_data_T_3205[169], _memRequest_bits_data_T_2820[169]};
  wire [3:0]        memRequest_bits_data_lo_177 = {memRequest_bits_data_lo_hi_177, memRequest_bits_data_lo_lo_177};
  wire [1:0]        memRequest_bits_data_hi_lo_177 = {_memRequest_bits_data_T_3975[169], _memRequest_bits_data_T_3590[169]};
  wire [1:0]        memRequest_bits_data_hi_hi_177 = {_memRequest_bits_data_T_4745[169], _memRequest_bits_data_T_4360[169]};
  wire [3:0]        memRequest_bits_data_hi_177 = {memRequest_bits_data_hi_hi_177, memRequest_bits_data_hi_lo_177};
  wire [1:0]        memRequest_bits_data_lo_lo_178 = {_memRequest_bits_data_T_2435[170], _memRequest_bits_data_T_2050[170]};
  wire [1:0]        memRequest_bits_data_lo_hi_178 = {_memRequest_bits_data_T_3205[170], _memRequest_bits_data_T_2820[170]};
  wire [3:0]        memRequest_bits_data_lo_178 = {memRequest_bits_data_lo_hi_178, memRequest_bits_data_lo_lo_178};
  wire [1:0]        memRequest_bits_data_hi_lo_178 = {_memRequest_bits_data_T_3975[170], _memRequest_bits_data_T_3590[170]};
  wire [1:0]        memRequest_bits_data_hi_hi_178 = {_memRequest_bits_data_T_4745[170], _memRequest_bits_data_T_4360[170]};
  wire [3:0]        memRequest_bits_data_hi_178 = {memRequest_bits_data_hi_hi_178, memRequest_bits_data_hi_lo_178};
  wire [1:0]        memRequest_bits_data_lo_lo_179 = {_memRequest_bits_data_T_2435[171], _memRequest_bits_data_T_2050[171]};
  wire [1:0]        memRequest_bits_data_lo_hi_179 = {_memRequest_bits_data_T_3205[171], _memRequest_bits_data_T_2820[171]};
  wire [3:0]        memRequest_bits_data_lo_179 = {memRequest_bits_data_lo_hi_179, memRequest_bits_data_lo_lo_179};
  wire [1:0]        memRequest_bits_data_hi_lo_179 = {_memRequest_bits_data_T_3975[171], _memRequest_bits_data_T_3590[171]};
  wire [1:0]        memRequest_bits_data_hi_hi_179 = {_memRequest_bits_data_T_4745[171], _memRequest_bits_data_T_4360[171]};
  wire [3:0]        memRequest_bits_data_hi_179 = {memRequest_bits_data_hi_hi_179, memRequest_bits_data_hi_lo_179};
  wire [1:0]        memRequest_bits_data_lo_lo_180 = {_memRequest_bits_data_T_2435[172], _memRequest_bits_data_T_2050[172]};
  wire [1:0]        memRequest_bits_data_lo_hi_180 = {_memRequest_bits_data_T_3205[172], _memRequest_bits_data_T_2820[172]};
  wire [3:0]        memRequest_bits_data_lo_180 = {memRequest_bits_data_lo_hi_180, memRequest_bits_data_lo_lo_180};
  wire [1:0]        memRequest_bits_data_hi_lo_180 = {_memRequest_bits_data_T_3975[172], _memRequest_bits_data_T_3590[172]};
  wire [1:0]        memRequest_bits_data_hi_hi_180 = {_memRequest_bits_data_T_4745[172], _memRequest_bits_data_T_4360[172]};
  wire [3:0]        memRequest_bits_data_hi_180 = {memRequest_bits_data_hi_hi_180, memRequest_bits_data_hi_lo_180};
  wire [1:0]        memRequest_bits_data_lo_lo_181 = {_memRequest_bits_data_T_2435[173], _memRequest_bits_data_T_2050[173]};
  wire [1:0]        memRequest_bits_data_lo_hi_181 = {_memRequest_bits_data_T_3205[173], _memRequest_bits_data_T_2820[173]};
  wire [3:0]        memRequest_bits_data_lo_181 = {memRequest_bits_data_lo_hi_181, memRequest_bits_data_lo_lo_181};
  wire [1:0]        memRequest_bits_data_hi_lo_181 = {_memRequest_bits_data_T_3975[173], _memRequest_bits_data_T_3590[173]};
  wire [1:0]        memRequest_bits_data_hi_hi_181 = {_memRequest_bits_data_T_4745[173], _memRequest_bits_data_T_4360[173]};
  wire [3:0]        memRequest_bits_data_hi_181 = {memRequest_bits_data_hi_hi_181, memRequest_bits_data_hi_lo_181};
  wire [1:0]        memRequest_bits_data_lo_lo_182 = {_memRequest_bits_data_T_2435[174], _memRequest_bits_data_T_2050[174]};
  wire [1:0]        memRequest_bits_data_lo_hi_182 = {_memRequest_bits_data_T_3205[174], _memRequest_bits_data_T_2820[174]};
  wire [3:0]        memRequest_bits_data_lo_182 = {memRequest_bits_data_lo_hi_182, memRequest_bits_data_lo_lo_182};
  wire [1:0]        memRequest_bits_data_hi_lo_182 = {_memRequest_bits_data_T_3975[174], _memRequest_bits_data_T_3590[174]};
  wire [1:0]        memRequest_bits_data_hi_hi_182 = {_memRequest_bits_data_T_4745[174], _memRequest_bits_data_T_4360[174]};
  wire [3:0]        memRequest_bits_data_hi_182 = {memRequest_bits_data_hi_hi_182, memRequest_bits_data_hi_lo_182};
  wire [1:0]        memRequest_bits_data_lo_lo_183 = {_memRequest_bits_data_T_2435[175], _memRequest_bits_data_T_2050[175]};
  wire [1:0]        memRequest_bits_data_lo_hi_183 = {_memRequest_bits_data_T_3205[175], _memRequest_bits_data_T_2820[175]};
  wire [3:0]        memRequest_bits_data_lo_183 = {memRequest_bits_data_lo_hi_183, memRequest_bits_data_lo_lo_183};
  wire [1:0]        memRequest_bits_data_hi_lo_183 = {_memRequest_bits_data_T_3975[175], _memRequest_bits_data_T_3590[175]};
  wire [1:0]        memRequest_bits_data_hi_hi_183 = {_memRequest_bits_data_T_4745[175], _memRequest_bits_data_T_4360[175]};
  wire [3:0]        memRequest_bits_data_hi_183 = {memRequest_bits_data_hi_hi_183, memRequest_bits_data_hi_lo_183};
  wire [1:0]        memRequest_bits_data_lo_lo_184 = {_memRequest_bits_data_T_2435[176], _memRequest_bits_data_T_2050[176]};
  wire [1:0]        memRequest_bits_data_lo_hi_184 = {_memRequest_bits_data_T_3205[176], _memRequest_bits_data_T_2820[176]};
  wire [3:0]        memRequest_bits_data_lo_184 = {memRequest_bits_data_lo_hi_184, memRequest_bits_data_lo_lo_184};
  wire [1:0]        memRequest_bits_data_hi_lo_184 = {_memRequest_bits_data_T_3975[176], _memRequest_bits_data_T_3590[176]};
  wire [1:0]        memRequest_bits_data_hi_hi_184 = {_memRequest_bits_data_T_4745[176], _memRequest_bits_data_T_4360[176]};
  wire [3:0]        memRequest_bits_data_hi_184 = {memRequest_bits_data_hi_hi_184, memRequest_bits_data_hi_lo_184};
  wire [1:0]        memRequest_bits_data_lo_lo_185 = {_memRequest_bits_data_T_2435[177], _memRequest_bits_data_T_2050[177]};
  wire [1:0]        memRequest_bits_data_lo_hi_185 = {_memRequest_bits_data_T_3205[177], _memRequest_bits_data_T_2820[177]};
  wire [3:0]        memRequest_bits_data_lo_185 = {memRequest_bits_data_lo_hi_185, memRequest_bits_data_lo_lo_185};
  wire [1:0]        memRequest_bits_data_hi_lo_185 = {_memRequest_bits_data_T_3975[177], _memRequest_bits_data_T_3590[177]};
  wire [1:0]        memRequest_bits_data_hi_hi_185 = {_memRequest_bits_data_T_4745[177], _memRequest_bits_data_T_4360[177]};
  wire [3:0]        memRequest_bits_data_hi_185 = {memRequest_bits_data_hi_hi_185, memRequest_bits_data_hi_lo_185};
  wire [1:0]        memRequest_bits_data_lo_lo_186 = {_memRequest_bits_data_T_2435[178], _memRequest_bits_data_T_2050[178]};
  wire [1:0]        memRequest_bits_data_lo_hi_186 = {_memRequest_bits_data_T_3205[178], _memRequest_bits_data_T_2820[178]};
  wire [3:0]        memRequest_bits_data_lo_186 = {memRequest_bits_data_lo_hi_186, memRequest_bits_data_lo_lo_186};
  wire [1:0]        memRequest_bits_data_hi_lo_186 = {_memRequest_bits_data_T_3975[178], _memRequest_bits_data_T_3590[178]};
  wire [1:0]        memRequest_bits_data_hi_hi_186 = {_memRequest_bits_data_T_4745[178], _memRequest_bits_data_T_4360[178]};
  wire [3:0]        memRequest_bits_data_hi_186 = {memRequest_bits_data_hi_hi_186, memRequest_bits_data_hi_lo_186};
  wire [1:0]        memRequest_bits_data_lo_lo_187 = {_memRequest_bits_data_T_2435[179], _memRequest_bits_data_T_2050[179]};
  wire [1:0]        memRequest_bits_data_lo_hi_187 = {_memRequest_bits_data_T_3205[179], _memRequest_bits_data_T_2820[179]};
  wire [3:0]        memRequest_bits_data_lo_187 = {memRequest_bits_data_lo_hi_187, memRequest_bits_data_lo_lo_187};
  wire [1:0]        memRequest_bits_data_hi_lo_187 = {_memRequest_bits_data_T_3975[179], _memRequest_bits_data_T_3590[179]};
  wire [1:0]        memRequest_bits_data_hi_hi_187 = {_memRequest_bits_data_T_4745[179], _memRequest_bits_data_T_4360[179]};
  wire [3:0]        memRequest_bits_data_hi_187 = {memRequest_bits_data_hi_hi_187, memRequest_bits_data_hi_lo_187};
  wire [1:0]        memRequest_bits_data_lo_lo_188 = {_memRequest_bits_data_T_2435[180], _memRequest_bits_data_T_2050[180]};
  wire [1:0]        memRequest_bits_data_lo_hi_188 = {_memRequest_bits_data_T_3205[180], _memRequest_bits_data_T_2820[180]};
  wire [3:0]        memRequest_bits_data_lo_188 = {memRequest_bits_data_lo_hi_188, memRequest_bits_data_lo_lo_188};
  wire [1:0]        memRequest_bits_data_hi_lo_188 = {_memRequest_bits_data_T_3975[180], _memRequest_bits_data_T_3590[180]};
  wire [1:0]        memRequest_bits_data_hi_hi_188 = {_memRequest_bits_data_T_4745[180], _memRequest_bits_data_T_4360[180]};
  wire [3:0]        memRequest_bits_data_hi_188 = {memRequest_bits_data_hi_hi_188, memRequest_bits_data_hi_lo_188};
  wire [1:0]        memRequest_bits_data_lo_lo_189 = {_memRequest_bits_data_T_2435[181], _memRequest_bits_data_T_2050[181]};
  wire [1:0]        memRequest_bits_data_lo_hi_189 = {_memRequest_bits_data_T_3205[181], _memRequest_bits_data_T_2820[181]};
  wire [3:0]        memRequest_bits_data_lo_189 = {memRequest_bits_data_lo_hi_189, memRequest_bits_data_lo_lo_189};
  wire [1:0]        memRequest_bits_data_hi_lo_189 = {_memRequest_bits_data_T_3975[181], _memRequest_bits_data_T_3590[181]};
  wire [1:0]        memRequest_bits_data_hi_hi_189 = {_memRequest_bits_data_T_4745[181], _memRequest_bits_data_T_4360[181]};
  wire [3:0]        memRequest_bits_data_hi_189 = {memRequest_bits_data_hi_hi_189, memRequest_bits_data_hi_lo_189};
  wire [1:0]        memRequest_bits_data_lo_lo_190 = {_memRequest_bits_data_T_2435[182], _memRequest_bits_data_T_2050[182]};
  wire [1:0]        memRequest_bits_data_lo_hi_190 = {_memRequest_bits_data_T_3205[182], _memRequest_bits_data_T_2820[182]};
  wire [3:0]        memRequest_bits_data_lo_190 = {memRequest_bits_data_lo_hi_190, memRequest_bits_data_lo_lo_190};
  wire [1:0]        memRequest_bits_data_hi_lo_190 = {_memRequest_bits_data_T_3975[182], _memRequest_bits_data_T_3590[182]};
  wire [1:0]        memRequest_bits_data_hi_hi_190 = {_memRequest_bits_data_T_4745[182], _memRequest_bits_data_T_4360[182]};
  wire [3:0]        memRequest_bits_data_hi_190 = {memRequest_bits_data_hi_hi_190, memRequest_bits_data_hi_lo_190};
  wire [1:0]        memRequest_bits_data_lo_lo_191 = {_memRequest_bits_data_T_2435[183], _memRequest_bits_data_T_2050[183]};
  wire [1:0]        memRequest_bits_data_lo_hi_191 = {_memRequest_bits_data_T_3205[183], _memRequest_bits_data_T_2820[183]};
  wire [3:0]        memRequest_bits_data_lo_191 = {memRequest_bits_data_lo_hi_191, memRequest_bits_data_lo_lo_191};
  wire [1:0]        memRequest_bits_data_hi_lo_191 = {_memRequest_bits_data_T_3975[183], _memRequest_bits_data_T_3590[183]};
  wire [1:0]        memRequest_bits_data_hi_hi_191 = {_memRequest_bits_data_T_4745[183], _memRequest_bits_data_T_4360[183]};
  wire [3:0]        memRequest_bits_data_hi_191 = {memRequest_bits_data_hi_hi_191, memRequest_bits_data_hi_lo_191};
  wire [1:0]        memRequest_bits_data_lo_lo_192 = {_memRequest_bits_data_T_2435[184], _memRequest_bits_data_T_2050[184]};
  wire [1:0]        memRequest_bits_data_lo_hi_192 = {_memRequest_bits_data_T_3205[184], _memRequest_bits_data_T_2820[184]};
  wire [3:0]        memRequest_bits_data_lo_192 = {memRequest_bits_data_lo_hi_192, memRequest_bits_data_lo_lo_192};
  wire [1:0]        memRequest_bits_data_hi_lo_192 = {_memRequest_bits_data_T_3975[184], _memRequest_bits_data_T_3590[184]};
  wire [1:0]        memRequest_bits_data_hi_hi_192 = {_memRequest_bits_data_T_4745[184], _memRequest_bits_data_T_4360[184]};
  wire [3:0]        memRequest_bits_data_hi_192 = {memRequest_bits_data_hi_hi_192, memRequest_bits_data_hi_lo_192};
  wire [1:0]        memRequest_bits_data_lo_lo_193 = {_memRequest_bits_data_T_2435[185], _memRequest_bits_data_T_2050[185]};
  wire [1:0]        memRequest_bits_data_lo_hi_193 = {_memRequest_bits_data_T_3205[185], _memRequest_bits_data_T_2820[185]};
  wire [3:0]        memRequest_bits_data_lo_193 = {memRequest_bits_data_lo_hi_193, memRequest_bits_data_lo_lo_193};
  wire [1:0]        memRequest_bits_data_hi_lo_193 = {_memRequest_bits_data_T_3975[185], _memRequest_bits_data_T_3590[185]};
  wire [1:0]        memRequest_bits_data_hi_hi_193 = {_memRequest_bits_data_T_4745[185], _memRequest_bits_data_T_4360[185]};
  wire [3:0]        memRequest_bits_data_hi_193 = {memRequest_bits_data_hi_hi_193, memRequest_bits_data_hi_lo_193};
  wire [1:0]        memRequest_bits_data_lo_lo_194 = {_memRequest_bits_data_T_2435[186], _memRequest_bits_data_T_2050[186]};
  wire [1:0]        memRequest_bits_data_lo_hi_194 = {_memRequest_bits_data_T_3205[186], _memRequest_bits_data_T_2820[186]};
  wire [3:0]        memRequest_bits_data_lo_194 = {memRequest_bits_data_lo_hi_194, memRequest_bits_data_lo_lo_194};
  wire [1:0]        memRequest_bits_data_hi_lo_194 = {_memRequest_bits_data_T_3975[186], _memRequest_bits_data_T_3590[186]};
  wire [1:0]        memRequest_bits_data_hi_hi_194 = {_memRequest_bits_data_T_4745[186], _memRequest_bits_data_T_4360[186]};
  wire [3:0]        memRequest_bits_data_hi_194 = {memRequest_bits_data_hi_hi_194, memRequest_bits_data_hi_lo_194};
  wire [1:0]        memRequest_bits_data_lo_lo_195 = {_memRequest_bits_data_T_2435[187], _memRequest_bits_data_T_2050[187]};
  wire [1:0]        memRequest_bits_data_lo_hi_195 = {_memRequest_bits_data_T_3205[187], _memRequest_bits_data_T_2820[187]};
  wire [3:0]        memRequest_bits_data_lo_195 = {memRequest_bits_data_lo_hi_195, memRequest_bits_data_lo_lo_195};
  wire [1:0]        memRequest_bits_data_hi_lo_195 = {_memRequest_bits_data_T_3975[187], _memRequest_bits_data_T_3590[187]};
  wire [1:0]        memRequest_bits_data_hi_hi_195 = {_memRequest_bits_data_T_4745[187], _memRequest_bits_data_T_4360[187]};
  wire [3:0]        memRequest_bits_data_hi_195 = {memRequest_bits_data_hi_hi_195, memRequest_bits_data_hi_lo_195};
  wire [1:0]        memRequest_bits_data_lo_lo_196 = {_memRequest_bits_data_T_2435[188], _memRequest_bits_data_T_2050[188]};
  wire [1:0]        memRequest_bits_data_lo_hi_196 = {_memRequest_bits_data_T_3205[188], _memRequest_bits_data_T_2820[188]};
  wire [3:0]        memRequest_bits_data_lo_196 = {memRequest_bits_data_lo_hi_196, memRequest_bits_data_lo_lo_196};
  wire [1:0]        memRequest_bits_data_hi_lo_196 = {_memRequest_bits_data_T_3975[188], _memRequest_bits_data_T_3590[188]};
  wire [1:0]        memRequest_bits_data_hi_hi_196 = {_memRequest_bits_data_T_4745[188], _memRequest_bits_data_T_4360[188]};
  wire [3:0]        memRequest_bits_data_hi_196 = {memRequest_bits_data_hi_hi_196, memRequest_bits_data_hi_lo_196};
  wire [1:0]        memRequest_bits_data_lo_lo_197 = {_memRequest_bits_data_T_2435[189], _memRequest_bits_data_T_2050[189]};
  wire [1:0]        memRequest_bits_data_lo_hi_197 = {_memRequest_bits_data_T_3205[189], _memRequest_bits_data_T_2820[189]};
  wire [3:0]        memRequest_bits_data_lo_197 = {memRequest_bits_data_lo_hi_197, memRequest_bits_data_lo_lo_197};
  wire [1:0]        memRequest_bits_data_hi_lo_197 = {_memRequest_bits_data_T_3975[189], _memRequest_bits_data_T_3590[189]};
  wire [1:0]        memRequest_bits_data_hi_hi_197 = {_memRequest_bits_data_T_4745[189], _memRequest_bits_data_T_4360[189]};
  wire [3:0]        memRequest_bits_data_hi_197 = {memRequest_bits_data_hi_hi_197, memRequest_bits_data_hi_lo_197};
  wire [1:0]        memRequest_bits_data_lo_lo_198 = {_memRequest_bits_data_T_2435[190], _memRequest_bits_data_T_2050[190]};
  wire [1:0]        memRequest_bits_data_lo_hi_198 = {_memRequest_bits_data_T_3205[190], _memRequest_bits_data_T_2820[190]};
  wire [3:0]        memRequest_bits_data_lo_198 = {memRequest_bits_data_lo_hi_198, memRequest_bits_data_lo_lo_198};
  wire [1:0]        memRequest_bits_data_hi_lo_198 = {_memRequest_bits_data_T_3975[190], _memRequest_bits_data_T_3590[190]};
  wire [1:0]        memRequest_bits_data_hi_hi_198 = {_memRequest_bits_data_T_4745[190], _memRequest_bits_data_T_4360[190]};
  wire [3:0]        memRequest_bits_data_hi_198 = {memRequest_bits_data_hi_hi_198, memRequest_bits_data_hi_lo_198};
  wire [1:0]        memRequest_bits_data_lo_lo_199 = {_memRequest_bits_data_T_2435[191], _memRequest_bits_data_T_2050[191]};
  wire [1:0]        memRequest_bits_data_lo_hi_199 = {_memRequest_bits_data_T_3205[191], _memRequest_bits_data_T_2820[191]};
  wire [3:0]        memRequest_bits_data_lo_199 = {memRequest_bits_data_lo_hi_199, memRequest_bits_data_lo_lo_199};
  wire [1:0]        memRequest_bits_data_hi_lo_199 = {_memRequest_bits_data_T_3975[191], _memRequest_bits_data_T_3590[191]};
  wire [1:0]        memRequest_bits_data_hi_hi_199 = {_memRequest_bits_data_T_4745[191], _memRequest_bits_data_T_4360[191]};
  wire [3:0]        memRequest_bits_data_hi_199 = {memRequest_bits_data_hi_hi_199, memRequest_bits_data_hi_lo_199};
  wire [1:0]        memRequest_bits_data_lo_lo_200 = {_memRequest_bits_data_T_2435[192], _memRequest_bits_data_T_2050[192]};
  wire [1:0]        memRequest_bits_data_lo_hi_200 = {_memRequest_bits_data_T_3205[192], _memRequest_bits_data_T_2820[192]};
  wire [3:0]        memRequest_bits_data_lo_200 = {memRequest_bits_data_lo_hi_200, memRequest_bits_data_lo_lo_200};
  wire [1:0]        memRequest_bits_data_hi_lo_200 = {_memRequest_bits_data_T_3975[192], _memRequest_bits_data_T_3590[192]};
  wire [1:0]        memRequest_bits_data_hi_hi_200 = {_memRequest_bits_data_T_4745[192], _memRequest_bits_data_T_4360[192]};
  wire [3:0]        memRequest_bits_data_hi_200 = {memRequest_bits_data_hi_hi_200, memRequest_bits_data_hi_lo_200};
  wire [1:0]        memRequest_bits_data_lo_lo_201 = {_memRequest_bits_data_T_2435[193], _memRequest_bits_data_T_2050[193]};
  wire [1:0]        memRequest_bits_data_lo_hi_201 = {_memRequest_bits_data_T_3205[193], _memRequest_bits_data_T_2820[193]};
  wire [3:0]        memRequest_bits_data_lo_201 = {memRequest_bits_data_lo_hi_201, memRequest_bits_data_lo_lo_201};
  wire [1:0]        memRequest_bits_data_hi_lo_201 = {_memRequest_bits_data_T_3975[193], _memRequest_bits_data_T_3590[193]};
  wire [1:0]        memRequest_bits_data_hi_hi_201 = {_memRequest_bits_data_T_4745[193], _memRequest_bits_data_T_4360[193]};
  wire [3:0]        memRequest_bits_data_hi_201 = {memRequest_bits_data_hi_hi_201, memRequest_bits_data_hi_lo_201};
  wire [1:0]        memRequest_bits_data_lo_lo_202 = {_memRequest_bits_data_T_2435[194], _memRequest_bits_data_T_2050[194]};
  wire [1:0]        memRequest_bits_data_lo_hi_202 = {_memRequest_bits_data_T_3205[194], _memRequest_bits_data_T_2820[194]};
  wire [3:0]        memRequest_bits_data_lo_202 = {memRequest_bits_data_lo_hi_202, memRequest_bits_data_lo_lo_202};
  wire [1:0]        memRequest_bits_data_hi_lo_202 = {_memRequest_bits_data_T_3975[194], _memRequest_bits_data_T_3590[194]};
  wire [1:0]        memRequest_bits_data_hi_hi_202 = {_memRequest_bits_data_T_4745[194], _memRequest_bits_data_T_4360[194]};
  wire [3:0]        memRequest_bits_data_hi_202 = {memRequest_bits_data_hi_hi_202, memRequest_bits_data_hi_lo_202};
  wire [1:0]        memRequest_bits_data_lo_lo_203 = {_memRequest_bits_data_T_2435[195], _memRequest_bits_data_T_2050[195]};
  wire [1:0]        memRequest_bits_data_lo_hi_203 = {_memRequest_bits_data_T_3205[195], _memRequest_bits_data_T_2820[195]};
  wire [3:0]        memRequest_bits_data_lo_203 = {memRequest_bits_data_lo_hi_203, memRequest_bits_data_lo_lo_203};
  wire [1:0]        memRequest_bits_data_hi_lo_203 = {_memRequest_bits_data_T_3975[195], _memRequest_bits_data_T_3590[195]};
  wire [1:0]        memRequest_bits_data_hi_hi_203 = {_memRequest_bits_data_T_4745[195], _memRequest_bits_data_T_4360[195]};
  wire [3:0]        memRequest_bits_data_hi_203 = {memRequest_bits_data_hi_hi_203, memRequest_bits_data_hi_lo_203};
  wire [1:0]        memRequest_bits_data_lo_lo_204 = {_memRequest_bits_data_T_2435[196], _memRequest_bits_data_T_2050[196]};
  wire [1:0]        memRequest_bits_data_lo_hi_204 = {_memRequest_bits_data_T_3205[196], _memRequest_bits_data_T_2820[196]};
  wire [3:0]        memRequest_bits_data_lo_204 = {memRequest_bits_data_lo_hi_204, memRequest_bits_data_lo_lo_204};
  wire [1:0]        memRequest_bits_data_hi_lo_204 = {_memRequest_bits_data_T_3975[196], _memRequest_bits_data_T_3590[196]};
  wire [1:0]        memRequest_bits_data_hi_hi_204 = {_memRequest_bits_data_T_4745[196], _memRequest_bits_data_T_4360[196]};
  wire [3:0]        memRequest_bits_data_hi_204 = {memRequest_bits_data_hi_hi_204, memRequest_bits_data_hi_lo_204};
  wire [1:0]        memRequest_bits_data_lo_lo_205 = {_memRequest_bits_data_T_2435[197], _memRequest_bits_data_T_2050[197]};
  wire [1:0]        memRequest_bits_data_lo_hi_205 = {_memRequest_bits_data_T_3205[197], _memRequest_bits_data_T_2820[197]};
  wire [3:0]        memRequest_bits_data_lo_205 = {memRequest_bits_data_lo_hi_205, memRequest_bits_data_lo_lo_205};
  wire [1:0]        memRequest_bits_data_hi_lo_205 = {_memRequest_bits_data_T_3975[197], _memRequest_bits_data_T_3590[197]};
  wire [1:0]        memRequest_bits_data_hi_hi_205 = {_memRequest_bits_data_T_4745[197], _memRequest_bits_data_T_4360[197]};
  wire [3:0]        memRequest_bits_data_hi_205 = {memRequest_bits_data_hi_hi_205, memRequest_bits_data_hi_lo_205};
  wire [1:0]        memRequest_bits_data_lo_lo_206 = {_memRequest_bits_data_T_2435[198], _memRequest_bits_data_T_2050[198]};
  wire [1:0]        memRequest_bits_data_lo_hi_206 = {_memRequest_bits_data_T_3205[198], _memRequest_bits_data_T_2820[198]};
  wire [3:0]        memRequest_bits_data_lo_206 = {memRequest_bits_data_lo_hi_206, memRequest_bits_data_lo_lo_206};
  wire [1:0]        memRequest_bits_data_hi_lo_206 = {_memRequest_bits_data_T_3975[198], _memRequest_bits_data_T_3590[198]};
  wire [1:0]        memRequest_bits_data_hi_hi_206 = {_memRequest_bits_data_T_4745[198], _memRequest_bits_data_T_4360[198]};
  wire [3:0]        memRequest_bits_data_hi_206 = {memRequest_bits_data_hi_hi_206, memRequest_bits_data_hi_lo_206};
  wire [1:0]        memRequest_bits_data_lo_lo_207 = {_memRequest_bits_data_T_2435[199], _memRequest_bits_data_T_2050[199]};
  wire [1:0]        memRequest_bits_data_lo_hi_207 = {_memRequest_bits_data_T_3205[199], _memRequest_bits_data_T_2820[199]};
  wire [3:0]        memRequest_bits_data_lo_207 = {memRequest_bits_data_lo_hi_207, memRequest_bits_data_lo_lo_207};
  wire [1:0]        memRequest_bits_data_hi_lo_207 = {_memRequest_bits_data_T_3975[199], _memRequest_bits_data_T_3590[199]};
  wire [1:0]        memRequest_bits_data_hi_hi_207 = {_memRequest_bits_data_T_4745[199], _memRequest_bits_data_T_4360[199]};
  wire [3:0]        memRequest_bits_data_hi_207 = {memRequest_bits_data_hi_hi_207, memRequest_bits_data_hi_lo_207};
  wire [1:0]        memRequest_bits_data_lo_lo_208 = {_memRequest_bits_data_T_2435[200], _memRequest_bits_data_T_2050[200]};
  wire [1:0]        memRequest_bits_data_lo_hi_208 = {_memRequest_bits_data_T_3205[200], _memRequest_bits_data_T_2820[200]};
  wire [3:0]        memRequest_bits_data_lo_208 = {memRequest_bits_data_lo_hi_208, memRequest_bits_data_lo_lo_208};
  wire [1:0]        memRequest_bits_data_hi_lo_208 = {_memRequest_bits_data_T_3975[200], _memRequest_bits_data_T_3590[200]};
  wire [1:0]        memRequest_bits_data_hi_hi_208 = {_memRequest_bits_data_T_4745[200], _memRequest_bits_data_T_4360[200]};
  wire [3:0]        memRequest_bits_data_hi_208 = {memRequest_bits_data_hi_hi_208, memRequest_bits_data_hi_lo_208};
  wire [1:0]        memRequest_bits_data_lo_lo_209 = {_memRequest_bits_data_T_2435[201], _memRequest_bits_data_T_2050[201]};
  wire [1:0]        memRequest_bits_data_lo_hi_209 = {_memRequest_bits_data_T_3205[201], _memRequest_bits_data_T_2820[201]};
  wire [3:0]        memRequest_bits_data_lo_209 = {memRequest_bits_data_lo_hi_209, memRequest_bits_data_lo_lo_209};
  wire [1:0]        memRequest_bits_data_hi_lo_209 = {_memRequest_bits_data_T_3975[201], _memRequest_bits_data_T_3590[201]};
  wire [1:0]        memRequest_bits_data_hi_hi_209 = {_memRequest_bits_data_T_4745[201], _memRequest_bits_data_T_4360[201]};
  wire [3:0]        memRequest_bits_data_hi_209 = {memRequest_bits_data_hi_hi_209, memRequest_bits_data_hi_lo_209};
  wire [1:0]        memRequest_bits_data_lo_lo_210 = {_memRequest_bits_data_T_2435[202], _memRequest_bits_data_T_2050[202]};
  wire [1:0]        memRequest_bits_data_lo_hi_210 = {_memRequest_bits_data_T_3205[202], _memRequest_bits_data_T_2820[202]};
  wire [3:0]        memRequest_bits_data_lo_210 = {memRequest_bits_data_lo_hi_210, memRequest_bits_data_lo_lo_210};
  wire [1:0]        memRequest_bits_data_hi_lo_210 = {_memRequest_bits_data_T_3975[202], _memRequest_bits_data_T_3590[202]};
  wire [1:0]        memRequest_bits_data_hi_hi_210 = {_memRequest_bits_data_T_4745[202], _memRequest_bits_data_T_4360[202]};
  wire [3:0]        memRequest_bits_data_hi_210 = {memRequest_bits_data_hi_hi_210, memRequest_bits_data_hi_lo_210};
  wire [1:0]        memRequest_bits_data_lo_lo_211 = {_memRequest_bits_data_T_2435[203], _memRequest_bits_data_T_2050[203]};
  wire [1:0]        memRequest_bits_data_lo_hi_211 = {_memRequest_bits_data_T_3205[203], _memRequest_bits_data_T_2820[203]};
  wire [3:0]        memRequest_bits_data_lo_211 = {memRequest_bits_data_lo_hi_211, memRequest_bits_data_lo_lo_211};
  wire [1:0]        memRequest_bits_data_hi_lo_211 = {_memRequest_bits_data_T_3975[203], _memRequest_bits_data_T_3590[203]};
  wire [1:0]        memRequest_bits_data_hi_hi_211 = {_memRequest_bits_data_T_4745[203], _memRequest_bits_data_T_4360[203]};
  wire [3:0]        memRequest_bits_data_hi_211 = {memRequest_bits_data_hi_hi_211, memRequest_bits_data_hi_lo_211};
  wire [1:0]        memRequest_bits_data_lo_lo_212 = {_memRequest_bits_data_T_2435[204], _memRequest_bits_data_T_2050[204]};
  wire [1:0]        memRequest_bits_data_lo_hi_212 = {_memRequest_bits_data_T_3205[204], _memRequest_bits_data_T_2820[204]};
  wire [3:0]        memRequest_bits_data_lo_212 = {memRequest_bits_data_lo_hi_212, memRequest_bits_data_lo_lo_212};
  wire [1:0]        memRequest_bits_data_hi_lo_212 = {_memRequest_bits_data_T_3975[204], _memRequest_bits_data_T_3590[204]};
  wire [1:0]        memRequest_bits_data_hi_hi_212 = {_memRequest_bits_data_T_4745[204], _memRequest_bits_data_T_4360[204]};
  wire [3:0]        memRequest_bits_data_hi_212 = {memRequest_bits_data_hi_hi_212, memRequest_bits_data_hi_lo_212};
  wire [1:0]        memRequest_bits_data_lo_lo_213 = {_memRequest_bits_data_T_2435[205], _memRequest_bits_data_T_2050[205]};
  wire [1:0]        memRequest_bits_data_lo_hi_213 = {_memRequest_bits_data_T_3205[205], _memRequest_bits_data_T_2820[205]};
  wire [3:0]        memRequest_bits_data_lo_213 = {memRequest_bits_data_lo_hi_213, memRequest_bits_data_lo_lo_213};
  wire [1:0]        memRequest_bits_data_hi_lo_213 = {_memRequest_bits_data_T_3975[205], _memRequest_bits_data_T_3590[205]};
  wire [1:0]        memRequest_bits_data_hi_hi_213 = {_memRequest_bits_data_T_4745[205], _memRequest_bits_data_T_4360[205]};
  wire [3:0]        memRequest_bits_data_hi_213 = {memRequest_bits_data_hi_hi_213, memRequest_bits_data_hi_lo_213};
  wire [1:0]        memRequest_bits_data_lo_lo_214 = {_memRequest_bits_data_T_2435[206], _memRequest_bits_data_T_2050[206]};
  wire [1:0]        memRequest_bits_data_lo_hi_214 = {_memRequest_bits_data_T_3205[206], _memRequest_bits_data_T_2820[206]};
  wire [3:0]        memRequest_bits_data_lo_214 = {memRequest_bits_data_lo_hi_214, memRequest_bits_data_lo_lo_214};
  wire [1:0]        memRequest_bits_data_hi_lo_214 = {_memRequest_bits_data_T_3975[206], _memRequest_bits_data_T_3590[206]};
  wire [1:0]        memRequest_bits_data_hi_hi_214 = {_memRequest_bits_data_T_4745[206], _memRequest_bits_data_T_4360[206]};
  wire [3:0]        memRequest_bits_data_hi_214 = {memRequest_bits_data_hi_hi_214, memRequest_bits_data_hi_lo_214};
  wire [1:0]        memRequest_bits_data_lo_lo_215 = {_memRequest_bits_data_T_2435[207], _memRequest_bits_data_T_2050[207]};
  wire [1:0]        memRequest_bits_data_lo_hi_215 = {_memRequest_bits_data_T_3205[207], _memRequest_bits_data_T_2820[207]};
  wire [3:0]        memRequest_bits_data_lo_215 = {memRequest_bits_data_lo_hi_215, memRequest_bits_data_lo_lo_215};
  wire [1:0]        memRequest_bits_data_hi_lo_215 = {_memRequest_bits_data_T_3975[207], _memRequest_bits_data_T_3590[207]};
  wire [1:0]        memRequest_bits_data_hi_hi_215 = {_memRequest_bits_data_T_4745[207], _memRequest_bits_data_T_4360[207]};
  wire [3:0]        memRequest_bits_data_hi_215 = {memRequest_bits_data_hi_hi_215, memRequest_bits_data_hi_lo_215};
  wire [1:0]        memRequest_bits_data_lo_lo_216 = {_memRequest_bits_data_T_2435[208], _memRequest_bits_data_T_2050[208]};
  wire [1:0]        memRequest_bits_data_lo_hi_216 = {_memRequest_bits_data_T_3205[208], _memRequest_bits_data_T_2820[208]};
  wire [3:0]        memRequest_bits_data_lo_216 = {memRequest_bits_data_lo_hi_216, memRequest_bits_data_lo_lo_216};
  wire [1:0]        memRequest_bits_data_hi_lo_216 = {_memRequest_bits_data_T_3975[208], _memRequest_bits_data_T_3590[208]};
  wire [1:0]        memRequest_bits_data_hi_hi_216 = {_memRequest_bits_data_T_4745[208], _memRequest_bits_data_T_4360[208]};
  wire [3:0]        memRequest_bits_data_hi_216 = {memRequest_bits_data_hi_hi_216, memRequest_bits_data_hi_lo_216};
  wire [1:0]        memRequest_bits_data_lo_lo_217 = {_memRequest_bits_data_T_2435[209], _memRequest_bits_data_T_2050[209]};
  wire [1:0]        memRequest_bits_data_lo_hi_217 = {_memRequest_bits_data_T_3205[209], _memRequest_bits_data_T_2820[209]};
  wire [3:0]        memRequest_bits_data_lo_217 = {memRequest_bits_data_lo_hi_217, memRequest_bits_data_lo_lo_217};
  wire [1:0]        memRequest_bits_data_hi_lo_217 = {_memRequest_bits_data_T_3975[209], _memRequest_bits_data_T_3590[209]};
  wire [1:0]        memRequest_bits_data_hi_hi_217 = {_memRequest_bits_data_T_4745[209], _memRequest_bits_data_T_4360[209]};
  wire [3:0]        memRequest_bits_data_hi_217 = {memRequest_bits_data_hi_hi_217, memRequest_bits_data_hi_lo_217};
  wire [1:0]        memRequest_bits_data_lo_lo_218 = {_memRequest_bits_data_T_2435[210], _memRequest_bits_data_T_2050[210]};
  wire [1:0]        memRequest_bits_data_lo_hi_218 = {_memRequest_bits_data_T_3205[210], _memRequest_bits_data_T_2820[210]};
  wire [3:0]        memRequest_bits_data_lo_218 = {memRequest_bits_data_lo_hi_218, memRequest_bits_data_lo_lo_218};
  wire [1:0]        memRequest_bits_data_hi_lo_218 = {_memRequest_bits_data_T_3975[210], _memRequest_bits_data_T_3590[210]};
  wire [1:0]        memRequest_bits_data_hi_hi_218 = {_memRequest_bits_data_T_4745[210], _memRequest_bits_data_T_4360[210]};
  wire [3:0]        memRequest_bits_data_hi_218 = {memRequest_bits_data_hi_hi_218, memRequest_bits_data_hi_lo_218};
  wire [1:0]        memRequest_bits_data_lo_lo_219 = {_memRequest_bits_data_T_2435[211], _memRequest_bits_data_T_2050[211]};
  wire [1:0]        memRequest_bits_data_lo_hi_219 = {_memRequest_bits_data_T_3205[211], _memRequest_bits_data_T_2820[211]};
  wire [3:0]        memRequest_bits_data_lo_219 = {memRequest_bits_data_lo_hi_219, memRequest_bits_data_lo_lo_219};
  wire [1:0]        memRequest_bits_data_hi_lo_219 = {_memRequest_bits_data_T_3975[211], _memRequest_bits_data_T_3590[211]};
  wire [1:0]        memRequest_bits_data_hi_hi_219 = {_memRequest_bits_data_T_4745[211], _memRequest_bits_data_T_4360[211]};
  wire [3:0]        memRequest_bits_data_hi_219 = {memRequest_bits_data_hi_hi_219, memRequest_bits_data_hi_lo_219};
  wire [1:0]        memRequest_bits_data_lo_lo_220 = {_memRequest_bits_data_T_2435[212], _memRequest_bits_data_T_2050[212]};
  wire [1:0]        memRequest_bits_data_lo_hi_220 = {_memRequest_bits_data_T_3205[212], _memRequest_bits_data_T_2820[212]};
  wire [3:0]        memRequest_bits_data_lo_220 = {memRequest_bits_data_lo_hi_220, memRequest_bits_data_lo_lo_220};
  wire [1:0]        memRequest_bits_data_hi_lo_220 = {_memRequest_bits_data_T_3975[212], _memRequest_bits_data_T_3590[212]};
  wire [1:0]        memRequest_bits_data_hi_hi_220 = {_memRequest_bits_data_T_4745[212], _memRequest_bits_data_T_4360[212]};
  wire [3:0]        memRequest_bits_data_hi_220 = {memRequest_bits_data_hi_hi_220, memRequest_bits_data_hi_lo_220};
  wire [1:0]        memRequest_bits_data_lo_lo_221 = {_memRequest_bits_data_T_2435[213], _memRequest_bits_data_T_2050[213]};
  wire [1:0]        memRequest_bits_data_lo_hi_221 = {_memRequest_bits_data_T_3205[213], _memRequest_bits_data_T_2820[213]};
  wire [3:0]        memRequest_bits_data_lo_221 = {memRequest_bits_data_lo_hi_221, memRequest_bits_data_lo_lo_221};
  wire [1:0]        memRequest_bits_data_hi_lo_221 = {_memRequest_bits_data_T_3975[213], _memRequest_bits_data_T_3590[213]};
  wire [1:0]        memRequest_bits_data_hi_hi_221 = {_memRequest_bits_data_T_4745[213], _memRequest_bits_data_T_4360[213]};
  wire [3:0]        memRequest_bits_data_hi_221 = {memRequest_bits_data_hi_hi_221, memRequest_bits_data_hi_lo_221};
  wire [1:0]        memRequest_bits_data_lo_lo_222 = {_memRequest_bits_data_T_2435[214], _memRequest_bits_data_T_2050[214]};
  wire [1:0]        memRequest_bits_data_lo_hi_222 = {_memRequest_bits_data_T_3205[214], _memRequest_bits_data_T_2820[214]};
  wire [3:0]        memRequest_bits_data_lo_222 = {memRequest_bits_data_lo_hi_222, memRequest_bits_data_lo_lo_222};
  wire [1:0]        memRequest_bits_data_hi_lo_222 = {_memRequest_bits_data_T_3975[214], _memRequest_bits_data_T_3590[214]};
  wire [1:0]        memRequest_bits_data_hi_hi_222 = {_memRequest_bits_data_T_4745[214], _memRequest_bits_data_T_4360[214]};
  wire [3:0]        memRequest_bits_data_hi_222 = {memRequest_bits_data_hi_hi_222, memRequest_bits_data_hi_lo_222};
  wire [1:0]        memRequest_bits_data_lo_lo_223 = {_memRequest_bits_data_T_2435[215], _memRequest_bits_data_T_2050[215]};
  wire [1:0]        memRequest_bits_data_lo_hi_223 = {_memRequest_bits_data_T_3205[215], _memRequest_bits_data_T_2820[215]};
  wire [3:0]        memRequest_bits_data_lo_223 = {memRequest_bits_data_lo_hi_223, memRequest_bits_data_lo_lo_223};
  wire [1:0]        memRequest_bits_data_hi_lo_223 = {_memRequest_bits_data_T_3975[215], _memRequest_bits_data_T_3590[215]};
  wire [1:0]        memRequest_bits_data_hi_hi_223 = {_memRequest_bits_data_T_4745[215], _memRequest_bits_data_T_4360[215]};
  wire [3:0]        memRequest_bits_data_hi_223 = {memRequest_bits_data_hi_hi_223, memRequest_bits_data_hi_lo_223};
  wire [1:0]        memRequest_bits_data_lo_lo_224 = {_memRequest_bits_data_T_2435[216], _memRequest_bits_data_T_2050[216]};
  wire [1:0]        memRequest_bits_data_lo_hi_224 = {_memRequest_bits_data_T_3205[216], _memRequest_bits_data_T_2820[216]};
  wire [3:0]        memRequest_bits_data_lo_224 = {memRequest_bits_data_lo_hi_224, memRequest_bits_data_lo_lo_224};
  wire [1:0]        memRequest_bits_data_hi_lo_224 = {_memRequest_bits_data_T_3975[216], _memRequest_bits_data_T_3590[216]};
  wire [1:0]        memRequest_bits_data_hi_hi_224 = {_memRequest_bits_data_T_4745[216], _memRequest_bits_data_T_4360[216]};
  wire [3:0]        memRequest_bits_data_hi_224 = {memRequest_bits_data_hi_hi_224, memRequest_bits_data_hi_lo_224};
  wire [1:0]        memRequest_bits_data_lo_lo_225 = {_memRequest_bits_data_T_2435[217], _memRequest_bits_data_T_2050[217]};
  wire [1:0]        memRequest_bits_data_lo_hi_225 = {_memRequest_bits_data_T_3205[217], _memRequest_bits_data_T_2820[217]};
  wire [3:0]        memRequest_bits_data_lo_225 = {memRequest_bits_data_lo_hi_225, memRequest_bits_data_lo_lo_225};
  wire [1:0]        memRequest_bits_data_hi_lo_225 = {_memRequest_bits_data_T_3975[217], _memRequest_bits_data_T_3590[217]};
  wire [1:0]        memRequest_bits_data_hi_hi_225 = {_memRequest_bits_data_T_4745[217], _memRequest_bits_data_T_4360[217]};
  wire [3:0]        memRequest_bits_data_hi_225 = {memRequest_bits_data_hi_hi_225, memRequest_bits_data_hi_lo_225};
  wire [1:0]        memRequest_bits_data_lo_lo_226 = {_memRequest_bits_data_T_2435[218], _memRequest_bits_data_T_2050[218]};
  wire [1:0]        memRequest_bits_data_lo_hi_226 = {_memRequest_bits_data_T_3205[218], _memRequest_bits_data_T_2820[218]};
  wire [3:0]        memRequest_bits_data_lo_226 = {memRequest_bits_data_lo_hi_226, memRequest_bits_data_lo_lo_226};
  wire [1:0]        memRequest_bits_data_hi_lo_226 = {_memRequest_bits_data_T_3975[218], _memRequest_bits_data_T_3590[218]};
  wire [1:0]        memRequest_bits_data_hi_hi_226 = {_memRequest_bits_data_T_4745[218], _memRequest_bits_data_T_4360[218]};
  wire [3:0]        memRequest_bits_data_hi_226 = {memRequest_bits_data_hi_hi_226, memRequest_bits_data_hi_lo_226};
  wire [1:0]        memRequest_bits_data_lo_lo_227 = {_memRequest_bits_data_T_2435[219], _memRequest_bits_data_T_2050[219]};
  wire [1:0]        memRequest_bits_data_lo_hi_227 = {_memRequest_bits_data_T_3205[219], _memRequest_bits_data_T_2820[219]};
  wire [3:0]        memRequest_bits_data_lo_227 = {memRequest_bits_data_lo_hi_227, memRequest_bits_data_lo_lo_227};
  wire [1:0]        memRequest_bits_data_hi_lo_227 = {_memRequest_bits_data_T_3975[219], _memRequest_bits_data_T_3590[219]};
  wire [1:0]        memRequest_bits_data_hi_hi_227 = {_memRequest_bits_data_T_4745[219], _memRequest_bits_data_T_4360[219]};
  wire [3:0]        memRequest_bits_data_hi_227 = {memRequest_bits_data_hi_hi_227, memRequest_bits_data_hi_lo_227};
  wire [1:0]        memRequest_bits_data_lo_lo_228 = {_memRequest_bits_data_T_2435[220], _memRequest_bits_data_T_2050[220]};
  wire [1:0]        memRequest_bits_data_lo_hi_228 = {_memRequest_bits_data_T_3205[220], _memRequest_bits_data_T_2820[220]};
  wire [3:0]        memRequest_bits_data_lo_228 = {memRequest_bits_data_lo_hi_228, memRequest_bits_data_lo_lo_228};
  wire [1:0]        memRequest_bits_data_hi_lo_228 = {_memRequest_bits_data_T_3975[220], _memRequest_bits_data_T_3590[220]};
  wire [1:0]        memRequest_bits_data_hi_hi_228 = {_memRequest_bits_data_T_4745[220], _memRequest_bits_data_T_4360[220]};
  wire [3:0]        memRequest_bits_data_hi_228 = {memRequest_bits_data_hi_hi_228, memRequest_bits_data_hi_lo_228};
  wire [1:0]        memRequest_bits_data_lo_lo_229 = {_memRequest_bits_data_T_2435[221], _memRequest_bits_data_T_2050[221]};
  wire [1:0]        memRequest_bits_data_lo_hi_229 = {_memRequest_bits_data_T_3205[221], _memRequest_bits_data_T_2820[221]};
  wire [3:0]        memRequest_bits_data_lo_229 = {memRequest_bits_data_lo_hi_229, memRequest_bits_data_lo_lo_229};
  wire [1:0]        memRequest_bits_data_hi_lo_229 = {_memRequest_bits_data_T_3975[221], _memRequest_bits_data_T_3590[221]};
  wire [1:0]        memRequest_bits_data_hi_hi_229 = {_memRequest_bits_data_T_4745[221], _memRequest_bits_data_T_4360[221]};
  wire [3:0]        memRequest_bits_data_hi_229 = {memRequest_bits_data_hi_hi_229, memRequest_bits_data_hi_lo_229};
  wire [1:0]        memRequest_bits_data_lo_lo_230 = {_memRequest_bits_data_T_2435[222], _memRequest_bits_data_T_2050[222]};
  wire [1:0]        memRequest_bits_data_lo_hi_230 = {_memRequest_bits_data_T_3205[222], _memRequest_bits_data_T_2820[222]};
  wire [3:0]        memRequest_bits_data_lo_230 = {memRequest_bits_data_lo_hi_230, memRequest_bits_data_lo_lo_230};
  wire [1:0]        memRequest_bits_data_hi_lo_230 = {_memRequest_bits_data_T_3975[222], _memRequest_bits_data_T_3590[222]};
  wire [1:0]        memRequest_bits_data_hi_hi_230 = {_memRequest_bits_data_T_4745[222], _memRequest_bits_data_T_4360[222]};
  wire [3:0]        memRequest_bits_data_hi_230 = {memRequest_bits_data_hi_hi_230, memRequest_bits_data_hi_lo_230};
  wire [1:0]        memRequest_bits_data_lo_lo_231 = {_memRequest_bits_data_T_2435[223], _memRequest_bits_data_T_2050[223]};
  wire [1:0]        memRequest_bits_data_lo_hi_231 = {_memRequest_bits_data_T_3205[223], _memRequest_bits_data_T_2820[223]};
  wire [3:0]        memRequest_bits_data_lo_231 = {memRequest_bits_data_lo_hi_231, memRequest_bits_data_lo_lo_231};
  wire [1:0]        memRequest_bits_data_hi_lo_231 = {_memRequest_bits_data_T_3975[223], _memRequest_bits_data_T_3590[223]};
  wire [1:0]        memRequest_bits_data_hi_hi_231 = {_memRequest_bits_data_T_4745[223], _memRequest_bits_data_T_4360[223]};
  wire [3:0]        memRequest_bits_data_hi_231 = {memRequest_bits_data_hi_hi_231, memRequest_bits_data_hi_lo_231};
  wire [1:0]        memRequest_bits_data_lo_lo_232 = {_memRequest_bits_data_T_2435[224], _memRequest_bits_data_T_2050[224]};
  wire [1:0]        memRequest_bits_data_lo_hi_232 = {_memRequest_bits_data_T_3205[224], _memRequest_bits_data_T_2820[224]};
  wire [3:0]        memRequest_bits_data_lo_232 = {memRequest_bits_data_lo_hi_232, memRequest_bits_data_lo_lo_232};
  wire [1:0]        memRequest_bits_data_hi_lo_232 = {_memRequest_bits_data_T_3975[224], _memRequest_bits_data_T_3590[224]};
  wire [1:0]        memRequest_bits_data_hi_hi_232 = {_memRequest_bits_data_T_4745[224], _memRequest_bits_data_T_4360[224]};
  wire [3:0]        memRequest_bits_data_hi_232 = {memRequest_bits_data_hi_hi_232, memRequest_bits_data_hi_lo_232};
  wire [1:0]        memRequest_bits_data_lo_lo_233 = {_memRequest_bits_data_T_2435[225], _memRequest_bits_data_T_2050[225]};
  wire [1:0]        memRequest_bits_data_lo_hi_233 = {_memRequest_bits_data_T_3205[225], _memRequest_bits_data_T_2820[225]};
  wire [3:0]        memRequest_bits_data_lo_233 = {memRequest_bits_data_lo_hi_233, memRequest_bits_data_lo_lo_233};
  wire [1:0]        memRequest_bits_data_hi_lo_233 = {_memRequest_bits_data_T_3975[225], _memRequest_bits_data_T_3590[225]};
  wire [1:0]        memRequest_bits_data_hi_hi_233 = {_memRequest_bits_data_T_4745[225], _memRequest_bits_data_T_4360[225]};
  wire [3:0]        memRequest_bits_data_hi_233 = {memRequest_bits_data_hi_hi_233, memRequest_bits_data_hi_lo_233};
  wire [1:0]        memRequest_bits_data_lo_lo_234 = {_memRequest_bits_data_T_2435[226], _memRequest_bits_data_T_2050[226]};
  wire [1:0]        memRequest_bits_data_lo_hi_234 = {_memRequest_bits_data_T_3205[226], _memRequest_bits_data_T_2820[226]};
  wire [3:0]        memRequest_bits_data_lo_234 = {memRequest_bits_data_lo_hi_234, memRequest_bits_data_lo_lo_234};
  wire [1:0]        memRequest_bits_data_hi_lo_234 = {_memRequest_bits_data_T_3975[226], _memRequest_bits_data_T_3590[226]};
  wire [1:0]        memRequest_bits_data_hi_hi_234 = {_memRequest_bits_data_T_4745[226], _memRequest_bits_data_T_4360[226]};
  wire [3:0]        memRequest_bits_data_hi_234 = {memRequest_bits_data_hi_hi_234, memRequest_bits_data_hi_lo_234};
  wire [1:0]        memRequest_bits_data_lo_lo_235 = {_memRequest_bits_data_T_2435[227], _memRequest_bits_data_T_2050[227]};
  wire [1:0]        memRequest_bits_data_lo_hi_235 = {_memRequest_bits_data_T_3205[227], _memRequest_bits_data_T_2820[227]};
  wire [3:0]        memRequest_bits_data_lo_235 = {memRequest_bits_data_lo_hi_235, memRequest_bits_data_lo_lo_235};
  wire [1:0]        memRequest_bits_data_hi_lo_235 = {_memRequest_bits_data_T_3975[227], _memRequest_bits_data_T_3590[227]};
  wire [1:0]        memRequest_bits_data_hi_hi_235 = {_memRequest_bits_data_T_4745[227], _memRequest_bits_data_T_4360[227]};
  wire [3:0]        memRequest_bits_data_hi_235 = {memRequest_bits_data_hi_hi_235, memRequest_bits_data_hi_lo_235};
  wire [1:0]        memRequest_bits_data_lo_lo_236 = {_memRequest_bits_data_T_2435[228], _memRequest_bits_data_T_2050[228]};
  wire [1:0]        memRequest_bits_data_lo_hi_236 = {_memRequest_bits_data_T_3205[228], _memRequest_bits_data_T_2820[228]};
  wire [3:0]        memRequest_bits_data_lo_236 = {memRequest_bits_data_lo_hi_236, memRequest_bits_data_lo_lo_236};
  wire [1:0]        memRequest_bits_data_hi_lo_236 = {_memRequest_bits_data_T_3975[228], _memRequest_bits_data_T_3590[228]};
  wire [1:0]        memRequest_bits_data_hi_hi_236 = {_memRequest_bits_data_T_4745[228], _memRequest_bits_data_T_4360[228]};
  wire [3:0]        memRequest_bits_data_hi_236 = {memRequest_bits_data_hi_hi_236, memRequest_bits_data_hi_lo_236};
  wire [1:0]        memRequest_bits_data_lo_lo_237 = {_memRequest_bits_data_T_2435[229], _memRequest_bits_data_T_2050[229]};
  wire [1:0]        memRequest_bits_data_lo_hi_237 = {_memRequest_bits_data_T_3205[229], _memRequest_bits_data_T_2820[229]};
  wire [3:0]        memRequest_bits_data_lo_237 = {memRequest_bits_data_lo_hi_237, memRequest_bits_data_lo_lo_237};
  wire [1:0]        memRequest_bits_data_hi_lo_237 = {_memRequest_bits_data_T_3975[229], _memRequest_bits_data_T_3590[229]};
  wire [1:0]        memRequest_bits_data_hi_hi_237 = {_memRequest_bits_data_T_4745[229], _memRequest_bits_data_T_4360[229]};
  wire [3:0]        memRequest_bits_data_hi_237 = {memRequest_bits_data_hi_hi_237, memRequest_bits_data_hi_lo_237};
  wire [1:0]        memRequest_bits_data_lo_lo_238 = {_memRequest_bits_data_T_2435[230], _memRequest_bits_data_T_2050[230]};
  wire [1:0]        memRequest_bits_data_lo_hi_238 = {_memRequest_bits_data_T_3205[230], _memRequest_bits_data_T_2820[230]};
  wire [3:0]        memRequest_bits_data_lo_238 = {memRequest_bits_data_lo_hi_238, memRequest_bits_data_lo_lo_238};
  wire [1:0]        memRequest_bits_data_hi_lo_238 = {_memRequest_bits_data_T_3975[230], _memRequest_bits_data_T_3590[230]};
  wire [1:0]        memRequest_bits_data_hi_hi_238 = {_memRequest_bits_data_T_4745[230], _memRequest_bits_data_T_4360[230]};
  wire [3:0]        memRequest_bits_data_hi_238 = {memRequest_bits_data_hi_hi_238, memRequest_bits_data_hi_lo_238};
  wire [1:0]        memRequest_bits_data_lo_lo_239 = {_memRequest_bits_data_T_2435[231], _memRequest_bits_data_T_2050[231]};
  wire [1:0]        memRequest_bits_data_lo_hi_239 = {_memRequest_bits_data_T_3205[231], _memRequest_bits_data_T_2820[231]};
  wire [3:0]        memRequest_bits_data_lo_239 = {memRequest_bits_data_lo_hi_239, memRequest_bits_data_lo_lo_239};
  wire [1:0]        memRequest_bits_data_hi_lo_239 = {_memRequest_bits_data_T_3975[231], _memRequest_bits_data_T_3590[231]};
  wire [1:0]        memRequest_bits_data_hi_hi_239 = {_memRequest_bits_data_T_4745[231], _memRequest_bits_data_T_4360[231]};
  wire [3:0]        memRequest_bits_data_hi_239 = {memRequest_bits_data_hi_hi_239, memRequest_bits_data_hi_lo_239};
  wire [1:0]        memRequest_bits_data_lo_lo_240 = {_memRequest_bits_data_T_2435[232], _memRequest_bits_data_T_2050[232]};
  wire [1:0]        memRequest_bits_data_lo_hi_240 = {_memRequest_bits_data_T_3205[232], _memRequest_bits_data_T_2820[232]};
  wire [3:0]        memRequest_bits_data_lo_240 = {memRequest_bits_data_lo_hi_240, memRequest_bits_data_lo_lo_240};
  wire [1:0]        memRequest_bits_data_hi_lo_240 = {_memRequest_bits_data_T_3975[232], _memRequest_bits_data_T_3590[232]};
  wire [1:0]        memRequest_bits_data_hi_hi_240 = {_memRequest_bits_data_T_4745[232], _memRequest_bits_data_T_4360[232]};
  wire [3:0]        memRequest_bits_data_hi_240 = {memRequest_bits_data_hi_hi_240, memRequest_bits_data_hi_lo_240};
  wire [1:0]        memRequest_bits_data_lo_lo_241 = {_memRequest_bits_data_T_2435[233], _memRequest_bits_data_T_2050[233]};
  wire [1:0]        memRequest_bits_data_lo_hi_241 = {_memRequest_bits_data_T_3205[233], _memRequest_bits_data_T_2820[233]};
  wire [3:0]        memRequest_bits_data_lo_241 = {memRequest_bits_data_lo_hi_241, memRequest_bits_data_lo_lo_241};
  wire [1:0]        memRequest_bits_data_hi_lo_241 = {_memRequest_bits_data_T_3975[233], _memRequest_bits_data_T_3590[233]};
  wire [1:0]        memRequest_bits_data_hi_hi_241 = {_memRequest_bits_data_T_4745[233], _memRequest_bits_data_T_4360[233]};
  wire [3:0]        memRequest_bits_data_hi_241 = {memRequest_bits_data_hi_hi_241, memRequest_bits_data_hi_lo_241};
  wire [1:0]        memRequest_bits_data_lo_lo_242 = {_memRequest_bits_data_T_2435[234], _memRequest_bits_data_T_2050[234]};
  wire [1:0]        memRequest_bits_data_lo_hi_242 = {_memRequest_bits_data_T_3205[234], _memRequest_bits_data_T_2820[234]};
  wire [3:0]        memRequest_bits_data_lo_242 = {memRequest_bits_data_lo_hi_242, memRequest_bits_data_lo_lo_242};
  wire [1:0]        memRequest_bits_data_hi_lo_242 = {_memRequest_bits_data_T_3975[234], _memRequest_bits_data_T_3590[234]};
  wire [1:0]        memRequest_bits_data_hi_hi_242 = {_memRequest_bits_data_T_4745[234], _memRequest_bits_data_T_4360[234]};
  wire [3:0]        memRequest_bits_data_hi_242 = {memRequest_bits_data_hi_hi_242, memRequest_bits_data_hi_lo_242};
  wire [1:0]        memRequest_bits_data_lo_lo_243 = {_memRequest_bits_data_T_2435[235], _memRequest_bits_data_T_2050[235]};
  wire [1:0]        memRequest_bits_data_lo_hi_243 = {_memRequest_bits_data_T_3205[235], _memRequest_bits_data_T_2820[235]};
  wire [3:0]        memRequest_bits_data_lo_243 = {memRequest_bits_data_lo_hi_243, memRequest_bits_data_lo_lo_243};
  wire [1:0]        memRequest_bits_data_hi_lo_243 = {_memRequest_bits_data_T_3975[235], _memRequest_bits_data_T_3590[235]};
  wire [1:0]        memRequest_bits_data_hi_hi_243 = {_memRequest_bits_data_T_4745[235], _memRequest_bits_data_T_4360[235]};
  wire [3:0]        memRequest_bits_data_hi_243 = {memRequest_bits_data_hi_hi_243, memRequest_bits_data_hi_lo_243};
  wire [1:0]        memRequest_bits_data_lo_lo_244 = {_memRequest_bits_data_T_2435[236], _memRequest_bits_data_T_2050[236]};
  wire [1:0]        memRequest_bits_data_lo_hi_244 = {_memRequest_bits_data_T_3205[236], _memRequest_bits_data_T_2820[236]};
  wire [3:0]        memRequest_bits_data_lo_244 = {memRequest_bits_data_lo_hi_244, memRequest_bits_data_lo_lo_244};
  wire [1:0]        memRequest_bits_data_hi_lo_244 = {_memRequest_bits_data_T_3975[236], _memRequest_bits_data_T_3590[236]};
  wire [1:0]        memRequest_bits_data_hi_hi_244 = {_memRequest_bits_data_T_4745[236], _memRequest_bits_data_T_4360[236]};
  wire [3:0]        memRequest_bits_data_hi_244 = {memRequest_bits_data_hi_hi_244, memRequest_bits_data_hi_lo_244};
  wire [1:0]        memRequest_bits_data_lo_lo_245 = {_memRequest_bits_data_T_2435[237], _memRequest_bits_data_T_2050[237]};
  wire [1:0]        memRequest_bits_data_lo_hi_245 = {_memRequest_bits_data_T_3205[237], _memRequest_bits_data_T_2820[237]};
  wire [3:0]        memRequest_bits_data_lo_245 = {memRequest_bits_data_lo_hi_245, memRequest_bits_data_lo_lo_245};
  wire [1:0]        memRequest_bits_data_hi_lo_245 = {_memRequest_bits_data_T_3975[237], _memRequest_bits_data_T_3590[237]};
  wire [1:0]        memRequest_bits_data_hi_hi_245 = {_memRequest_bits_data_T_4745[237], _memRequest_bits_data_T_4360[237]};
  wire [3:0]        memRequest_bits_data_hi_245 = {memRequest_bits_data_hi_hi_245, memRequest_bits_data_hi_lo_245};
  wire [1:0]        memRequest_bits_data_lo_lo_246 = {_memRequest_bits_data_T_2435[238], _memRequest_bits_data_T_2050[238]};
  wire [1:0]        memRequest_bits_data_lo_hi_246 = {_memRequest_bits_data_T_3205[238], _memRequest_bits_data_T_2820[238]};
  wire [3:0]        memRequest_bits_data_lo_246 = {memRequest_bits_data_lo_hi_246, memRequest_bits_data_lo_lo_246};
  wire [1:0]        memRequest_bits_data_hi_lo_246 = {_memRequest_bits_data_T_3975[238], _memRequest_bits_data_T_3590[238]};
  wire [1:0]        memRequest_bits_data_hi_hi_246 = {_memRequest_bits_data_T_4745[238], _memRequest_bits_data_T_4360[238]};
  wire [3:0]        memRequest_bits_data_hi_246 = {memRequest_bits_data_hi_hi_246, memRequest_bits_data_hi_lo_246};
  wire [1:0]        memRequest_bits_data_lo_lo_247 = {_memRequest_bits_data_T_2435[239], _memRequest_bits_data_T_2050[239]};
  wire [1:0]        memRequest_bits_data_lo_hi_247 = {_memRequest_bits_data_T_3205[239], _memRequest_bits_data_T_2820[239]};
  wire [3:0]        memRequest_bits_data_lo_247 = {memRequest_bits_data_lo_hi_247, memRequest_bits_data_lo_lo_247};
  wire [1:0]        memRequest_bits_data_hi_lo_247 = {_memRequest_bits_data_T_3975[239], _memRequest_bits_data_T_3590[239]};
  wire [1:0]        memRequest_bits_data_hi_hi_247 = {_memRequest_bits_data_T_4745[239], _memRequest_bits_data_T_4360[239]};
  wire [3:0]        memRequest_bits_data_hi_247 = {memRequest_bits_data_hi_hi_247, memRequest_bits_data_hi_lo_247};
  wire [1:0]        memRequest_bits_data_lo_lo_248 = {_memRequest_bits_data_T_2435[240], _memRequest_bits_data_T_2050[240]};
  wire [1:0]        memRequest_bits_data_lo_hi_248 = {_memRequest_bits_data_T_3205[240], _memRequest_bits_data_T_2820[240]};
  wire [3:0]        memRequest_bits_data_lo_248 = {memRequest_bits_data_lo_hi_248, memRequest_bits_data_lo_lo_248};
  wire [1:0]        memRequest_bits_data_hi_lo_248 = {_memRequest_bits_data_T_3975[240], _memRequest_bits_data_T_3590[240]};
  wire [1:0]        memRequest_bits_data_hi_hi_248 = {_memRequest_bits_data_T_4745[240], _memRequest_bits_data_T_4360[240]};
  wire [3:0]        memRequest_bits_data_hi_248 = {memRequest_bits_data_hi_hi_248, memRequest_bits_data_hi_lo_248};
  wire [1:0]        memRequest_bits_data_lo_lo_249 = {_memRequest_bits_data_T_2435[241], _memRequest_bits_data_T_2050[241]};
  wire [1:0]        memRequest_bits_data_lo_hi_249 = {_memRequest_bits_data_T_3205[241], _memRequest_bits_data_T_2820[241]};
  wire [3:0]        memRequest_bits_data_lo_249 = {memRequest_bits_data_lo_hi_249, memRequest_bits_data_lo_lo_249};
  wire [1:0]        memRequest_bits_data_hi_lo_249 = {_memRequest_bits_data_T_3975[241], _memRequest_bits_data_T_3590[241]};
  wire [1:0]        memRequest_bits_data_hi_hi_249 = {_memRequest_bits_data_T_4745[241], _memRequest_bits_data_T_4360[241]};
  wire [3:0]        memRequest_bits_data_hi_249 = {memRequest_bits_data_hi_hi_249, memRequest_bits_data_hi_lo_249};
  wire [1:0]        memRequest_bits_data_lo_lo_250 = {_memRequest_bits_data_T_2435[242], _memRequest_bits_data_T_2050[242]};
  wire [1:0]        memRequest_bits_data_lo_hi_250 = {_memRequest_bits_data_T_3205[242], _memRequest_bits_data_T_2820[242]};
  wire [3:0]        memRequest_bits_data_lo_250 = {memRequest_bits_data_lo_hi_250, memRequest_bits_data_lo_lo_250};
  wire [1:0]        memRequest_bits_data_hi_lo_250 = {_memRequest_bits_data_T_3975[242], _memRequest_bits_data_T_3590[242]};
  wire [1:0]        memRequest_bits_data_hi_hi_250 = {_memRequest_bits_data_T_4745[242], _memRequest_bits_data_T_4360[242]};
  wire [3:0]        memRequest_bits_data_hi_250 = {memRequest_bits_data_hi_hi_250, memRequest_bits_data_hi_lo_250};
  wire [1:0]        memRequest_bits_data_lo_lo_251 = {_memRequest_bits_data_T_2435[243], _memRequest_bits_data_T_2050[243]};
  wire [1:0]        memRequest_bits_data_lo_hi_251 = {_memRequest_bits_data_T_3205[243], _memRequest_bits_data_T_2820[243]};
  wire [3:0]        memRequest_bits_data_lo_251 = {memRequest_bits_data_lo_hi_251, memRequest_bits_data_lo_lo_251};
  wire [1:0]        memRequest_bits_data_hi_lo_251 = {_memRequest_bits_data_T_3975[243], _memRequest_bits_data_T_3590[243]};
  wire [1:0]        memRequest_bits_data_hi_hi_251 = {_memRequest_bits_data_T_4745[243], _memRequest_bits_data_T_4360[243]};
  wire [3:0]        memRequest_bits_data_hi_251 = {memRequest_bits_data_hi_hi_251, memRequest_bits_data_hi_lo_251};
  wire [1:0]        memRequest_bits_data_lo_lo_252 = {_memRequest_bits_data_T_2435[244], _memRequest_bits_data_T_2050[244]};
  wire [1:0]        memRequest_bits_data_lo_hi_252 = {_memRequest_bits_data_T_3205[244], _memRequest_bits_data_T_2820[244]};
  wire [3:0]        memRequest_bits_data_lo_252 = {memRequest_bits_data_lo_hi_252, memRequest_bits_data_lo_lo_252};
  wire [1:0]        memRequest_bits_data_hi_lo_252 = {_memRequest_bits_data_T_3975[244], _memRequest_bits_data_T_3590[244]};
  wire [1:0]        memRequest_bits_data_hi_hi_252 = {_memRequest_bits_data_T_4745[244], _memRequest_bits_data_T_4360[244]};
  wire [3:0]        memRequest_bits_data_hi_252 = {memRequest_bits_data_hi_hi_252, memRequest_bits_data_hi_lo_252};
  wire [1:0]        memRequest_bits_data_lo_lo_253 = {_memRequest_bits_data_T_2435[245], _memRequest_bits_data_T_2050[245]};
  wire [1:0]        memRequest_bits_data_lo_hi_253 = {_memRequest_bits_data_T_3205[245], _memRequest_bits_data_T_2820[245]};
  wire [3:0]        memRequest_bits_data_lo_253 = {memRequest_bits_data_lo_hi_253, memRequest_bits_data_lo_lo_253};
  wire [1:0]        memRequest_bits_data_hi_lo_253 = {_memRequest_bits_data_T_3975[245], _memRequest_bits_data_T_3590[245]};
  wire [1:0]        memRequest_bits_data_hi_hi_253 = {_memRequest_bits_data_T_4745[245], _memRequest_bits_data_T_4360[245]};
  wire [3:0]        memRequest_bits_data_hi_253 = {memRequest_bits_data_hi_hi_253, memRequest_bits_data_hi_lo_253};
  wire [1:0]        memRequest_bits_data_lo_lo_254 = {_memRequest_bits_data_T_2435[246], _memRequest_bits_data_T_2050[246]};
  wire [1:0]        memRequest_bits_data_lo_hi_254 = {_memRequest_bits_data_T_3205[246], _memRequest_bits_data_T_2820[246]};
  wire [3:0]        memRequest_bits_data_lo_254 = {memRequest_bits_data_lo_hi_254, memRequest_bits_data_lo_lo_254};
  wire [1:0]        memRequest_bits_data_hi_lo_254 = {_memRequest_bits_data_T_3975[246], _memRequest_bits_data_T_3590[246]};
  wire [1:0]        memRequest_bits_data_hi_hi_254 = {_memRequest_bits_data_T_4745[246], _memRequest_bits_data_T_4360[246]};
  wire [3:0]        memRequest_bits_data_hi_254 = {memRequest_bits_data_hi_hi_254, memRequest_bits_data_hi_lo_254};
  wire [1:0]        memRequest_bits_data_lo_lo_255 = {_memRequest_bits_data_T_2435[247], _memRequest_bits_data_T_2050[247]};
  wire [1:0]        memRequest_bits_data_lo_hi_255 = {_memRequest_bits_data_T_3205[247], _memRequest_bits_data_T_2820[247]};
  wire [3:0]        memRequest_bits_data_lo_255 = {memRequest_bits_data_lo_hi_255, memRequest_bits_data_lo_lo_255};
  wire [1:0]        memRequest_bits_data_hi_lo_255 = {_memRequest_bits_data_T_3975[247], _memRequest_bits_data_T_3590[247]};
  wire [1:0]        memRequest_bits_data_hi_hi_255 = {_memRequest_bits_data_T_4745[247], _memRequest_bits_data_T_4360[247]};
  wire [3:0]        memRequest_bits_data_hi_255 = {memRequest_bits_data_hi_hi_255, memRequest_bits_data_hi_lo_255};
  wire [1:0]        memRequest_bits_data_lo_lo_256 = {_memRequest_bits_data_T_2435[248], _memRequest_bits_data_T_2050[248]};
  wire [1:0]        memRequest_bits_data_lo_hi_256 = {_memRequest_bits_data_T_3205[248], _memRequest_bits_data_T_2820[248]};
  wire [3:0]        memRequest_bits_data_lo_256 = {memRequest_bits_data_lo_hi_256, memRequest_bits_data_lo_lo_256};
  wire [1:0]        memRequest_bits_data_hi_lo_256 = {_memRequest_bits_data_T_3975[248], _memRequest_bits_data_T_3590[248]};
  wire [1:0]        memRequest_bits_data_hi_hi_256 = {_memRequest_bits_data_T_4745[248], _memRequest_bits_data_T_4360[248]};
  wire [3:0]        memRequest_bits_data_hi_256 = {memRequest_bits_data_hi_hi_256, memRequest_bits_data_hi_lo_256};
  wire [1:0]        memRequest_bits_data_lo_lo_257 = {_memRequest_bits_data_T_2435[249], _memRequest_bits_data_T_2050[249]};
  wire [1:0]        memRequest_bits_data_lo_hi_257 = {_memRequest_bits_data_T_3205[249], _memRequest_bits_data_T_2820[249]};
  wire [3:0]        memRequest_bits_data_lo_257 = {memRequest_bits_data_lo_hi_257, memRequest_bits_data_lo_lo_257};
  wire [1:0]        memRequest_bits_data_hi_lo_257 = {_memRequest_bits_data_T_3975[249], _memRequest_bits_data_T_3590[249]};
  wire [1:0]        memRequest_bits_data_hi_hi_257 = {_memRequest_bits_data_T_4745[249], _memRequest_bits_data_T_4360[249]};
  wire [3:0]        memRequest_bits_data_hi_257 = {memRequest_bits_data_hi_hi_257, memRequest_bits_data_hi_lo_257};
  wire [1:0]        memRequest_bits_data_lo_lo_258 = {_memRequest_bits_data_T_2435[250], _memRequest_bits_data_T_2050[250]};
  wire [1:0]        memRequest_bits_data_lo_hi_258 = {_memRequest_bits_data_T_3205[250], _memRequest_bits_data_T_2820[250]};
  wire [3:0]        memRequest_bits_data_lo_258 = {memRequest_bits_data_lo_hi_258, memRequest_bits_data_lo_lo_258};
  wire [1:0]        memRequest_bits_data_hi_lo_258 = {_memRequest_bits_data_T_3975[250], _memRequest_bits_data_T_3590[250]};
  wire [1:0]        memRequest_bits_data_hi_hi_258 = {_memRequest_bits_data_T_4745[250], _memRequest_bits_data_T_4360[250]};
  wire [3:0]        memRequest_bits_data_hi_258 = {memRequest_bits_data_hi_hi_258, memRequest_bits_data_hi_lo_258};
  wire [1:0]        memRequest_bits_data_lo_lo_259 = {_memRequest_bits_data_T_2435[251], _memRequest_bits_data_T_2050[251]};
  wire [1:0]        memRequest_bits_data_lo_hi_259 = {_memRequest_bits_data_T_3205[251], _memRequest_bits_data_T_2820[251]};
  wire [3:0]        memRequest_bits_data_lo_259 = {memRequest_bits_data_lo_hi_259, memRequest_bits_data_lo_lo_259};
  wire [1:0]        memRequest_bits_data_hi_lo_259 = {_memRequest_bits_data_T_3975[251], _memRequest_bits_data_T_3590[251]};
  wire [1:0]        memRequest_bits_data_hi_hi_259 = {_memRequest_bits_data_T_4745[251], _memRequest_bits_data_T_4360[251]};
  wire [3:0]        memRequest_bits_data_hi_259 = {memRequest_bits_data_hi_hi_259, memRequest_bits_data_hi_lo_259};
  wire [1:0]        memRequest_bits_data_lo_lo_260 = {_memRequest_bits_data_T_2435[252], _memRequest_bits_data_T_2050[252]};
  wire [1:0]        memRequest_bits_data_lo_hi_260 = {_memRequest_bits_data_T_3205[252], _memRequest_bits_data_T_2820[252]};
  wire [3:0]        memRequest_bits_data_lo_260 = {memRequest_bits_data_lo_hi_260, memRequest_bits_data_lo_lo_260};
  wire [1:0]        memRequest_bits_data_hi_lo_260 = {_memRequest_bits_data_T_3975[252], _memRequest_bits_data_T_3590[252]};
  wire [1:0]        memRequest_bits_data_hi_hi_260 = {_memRequest_bits_data_T_4745[252], _memRequest_bits_data_T_4360[252]};
  wire [3:0]        memRequest_bits_data_hi_260 = {memRequest_bits_data_hi_hi_260, memRequest_bits_data_hi_lo_260};
  wire [1:0]        memRequest_bits_data_lo_lo_261 = {_memRequest_bits_data_T_2435[253], _memRequest_bits_data_T_2050[253]};
  wire [1:0]        memRequest_bits_data_lo_hi_261 = {_memRequest_bits_data_T_3205[253], _memRequest_bits_data_T_2820[253]};
  wire [3:0]        memRequest_bits_data_lo_261 = {memRequest_bits_data_lo_hi_261, memRequest_bits_data_lo_lo_261};
  wire [1:0]        memRequest_bits_data_hi_lo_261 = {_memRequest_bits_data_T_3975[253], _memRequest_bits_data_T_3590[253]};
  wire [1:0]        memRequest_bits_data_hi_hi_261 = {_memRequest_bits_data_T_4745[253], _memRequest_bits_data_T_4360[253]};
  wire [3:0]        memRequest_bits_data_hi_261 = {memRequest_bits_data_hi_hi_261, memRequest_bits_data_hi_lo_261};
  wire [1:0]        memRequest_bits_data_lo_lo_262 = {_memRequest_bits_data_T_2435[254], _memRequest_bits_data_T_2050[254]};
  wire [1:0]        memRequest_bits_data_lo_hi_262 = {_memRequest_bits_data_T_3205[254], _memRequest_bits_data_T_2820[254]};
  wire [3:0]        memRequest_bits_data_lo_262 = {memRequest_bits_data_lo_hi_262, memRequest_bits_data_lo_lo_262};
  wire [1:0]        memRequest_bits_data_hi_lo_262 = {_memRequest_bits_data_T_3975[254], _memRequest_bits_data_T_3590[254]};
  wire [1:0]        memRequest_bits_data_hi_hi_262 = {_memRequest_bits_data_T_4745[254], _memRequest_bits_data_T_4360[254]};
  wire [3:0]        memRequest_bits_data_hi_262 = {memRequest_bits_data_hi_hi_262, memRequest_bits_data_hi_lo_262};
  wire [1:0]        memRequest_bits_data_lo_lo_263 = {_memRequest_bits_data_T_2435[255], _memRequest_bits_data_T_2050[255]};
  wire [1:0]        memRequest_bits_data_lo_hi_263 = {_memRequest_bits_data_T_3205[255], _memRequest_bits_data_T_2820[255]};
  wire [3:0]        memRequest_bits_data_lo_263 = {memRequest_bits_data_lo_hi_263, memRequest_bits_data_lo_lo_263};
  wire [1:0]        memRequest_bits_data_hi_lo_263 = {_memRequest_bits_data_T_3975[255], _memRequest_bits_data_T_3590[255]};
  wire [1:0]        memRequest_bits_data_hi_hi_263 = {_memRequest_bits_data_T_4745[255], _memRequest_bits_data_T_4360[255]};
  wire [3:0]        memRequest_bits_data_hi_263 = {memRequest_bits_data_hi_hi_263, memRequest_bits_data_hi_lo_263};
  wire [1:0]        memRequest_bits_data_lo_lo_264 = {_memRequest_bits_data_T_2435[256], _memRequest_bits_data_T_2050[256]};
  wire [1:0]        memRequest_bits_data_lo_hi_264 = {_memRequest_bits_data_T_3205[256], _memRequest_bits_data_T_2820[256]};
  wire [3:0]        memRequest_bits_data_lo_264 = {memRequest_bits_data_lo_hi_264, memRequest_bits_data_lo_lo_264};
  wire [1:0]        memRequest_bits_data_hi_lo_264 = {_memRequest_bits_data_T_3975[256], _memRequest_bits_data_T_3590[256]};
  wire [1:0]        memRequest_bits_data_hi_hi_264 = {_memRequest_bits_data_T_4745[256], _memRequest_bits_data_T_4360[256]};
  wire [3:0]        memRequest_bits_data_hi_264 = {memRequest_bits_data_hi_hi_264, memRequest_bits_data_hi_lo_264};
  wire [1:0]        memRequest_bits_data_lo_lo_265 = {_memRequest_bits_data_T_2435[257], _memRequest_bits_data_T_2050[257]};
  wire [1:0]        memRequest_bits_data_lo_hi_265 = {_memRequest_bits_data_T_3205[257], _memRequest_bits_data_T_2820[257]};
  wire [3:0]        memRequest_bits_data_lo_265 = {memRequest_bits_data_lo_hi_265, memRequest_bits_data_lo_lo_265};
  wire [1:0]        memRequest_bits_data_hi_lo_265 = {_memRequest_bits_data_T_3975[257], _memRequest_bits_data_T_3590[257]};
  wire [1:0]        memRequest_bits_data_hi_hi_265 = {_memRequest_bits_data_T_4745[257], _memRequest_bits_data_T_4360[257]};
  wire [3:0]        memRequest_bits_data_hi_265 = {memRequest_bits_data_hi_hi_265, memRequest_bits_data_hi_lo_265};
  wire [1:0]        memRequest_bits_data_lo_lo_266 = {_memRequest_bits_data_T_2435[258], _memRequest_bits_data_T_2050[258]};
  wire [1:0]        memRequest_bits_data_lo_hi_266 = {_memRequest_bits_data_T_3205[258], _memRequest_bits_data_T_2820[258]};
  wire [3:0]        memRequest_bits_data_lo_266 = {memRequest_bits_data_lo_hi_266, memRequest_bits_data_lo_lo_266};
  wire [1:0]        memRequest_bits_data_hi_lo_266 = {_memRequest_bits_data_T_3975[258], _memRequest_bits_data_T_3590[258]};
  wire [1:0]        memRequest_bits_data_hi_hi_266 = {_memRequest_bits_data_T_4745[258], _memRequest_bits_data_T_4360[258]};
  wire [3:0]        memRequest_bits_data_hi_266 = {memRequest_bits_data_hi_hi_266, memRequest_bits_data_hi_lo_266};
  wire [1:0]        memRequest_bits_data_lo_lo_267 = {_memRequest_bits_data_T_2435[259], _memRequest_bits_data_T_2050[259]};
  wire [1:0]        memRequest_bits_data_lo_hi_267 = {_memRequest_bits_data_T_3205[259], _memRequest_bits_data_T_2820[259]};
  wire [3:0]        memRequest_bits_data_lo_267 = {memRequest_bits_data_lo_hi_267, memRequest_bits_data_lo_lo_267};
  wire [1:0]        memRequest_bits_data_hi_lo_267 = {_memRequest_bits_data_T_3975[259], _memRequest_bits_data_T_3590[259]};
  wire [1:0]        memRequest_bits_data_hi_hi_267 = {_memRequest_bits_data_T_4745[259], _memRequest_bits_data_T_4360[259]};
  wire [3:0]        memRequest_bits_data_hi_267 = {memRequest_bits_data_hi_hi_267, memRequest_bits_data_hi_lo_267};
  wire [1:0]        memRequest_bits_data_lo_lo_268 = {_memRequest_bits_data_T_2435[260], _memRequest_bits_data_T_2050[260]};
  wire [1:0]        memRequest_bits_data_lo_hi_268 = {_memRequest_bits_data_T_3205[260], _memRequest_bits_data_T_2820[260]};
  wire [3:0]        memRequest_bits_data_lo_268 = {memRequest_bits_data_lo_hi_268, memRequest_bits_data_lo_lo_268};
  wire [1:0]        memRequest_bits_data_hi_lo_268 = {_memRequest_bits_data_T_3975[260], _memRequest_bits_data_T_3590[260]};
  wire [1:0]        memRequest_bits_data_hi_hi_268 = {_memRequest_bits_data_T_4745[260], _memRequest_bits_data_T_4360[260]};
  wire [3:0]        memRequest_bits_data_hi_268 = {memRequest_bits_data_hi_hi_268, memRequest_bits_data_hi_lo_268};
  wire [1:0]        memRequest_bits_data_lo_lo_269 = {_memRequest_bits_data_T_2435[261], _memRequest_bits_data_T_2050[261]};
  wire [1:0]        memRequest_bits_data_lo_hi_269 = {_memRequest_bits_data_T_3205[261], _memRequest_bits_data_T_2820[261]};
  wire [3:0]        memRequest_bits_data_lo_269 = {memRequest_bits_data_lo_hi_269, memRequest_bits_data_lo_lo_269};
  wire [1:0]        memRequest_bits_data_hi_lo_269 = {_memRequest_bits_data_T_3975[261], _memRequest_bits_data_T_3590[261]};
  wire [1:0]        memRequest_bits_data_hi_hi_269 = {_memRequest_bits_data_T_4745[261], _memRequest_bits_data_T_4360[261]};
  wire [3:0]        memRequest_bits_data_hi_269 = {memRequest_bits_data_hi_hi_269, memRequest_bits_data_hi_lo_269};
  wire [1:0]        memRequest_bits_data_lo_lo_270 = {_memRequest_bits_data_T_2435[262], _memRequest_bits_data_T_2050[262]};
  wire [1:0]        memRequest_bits_data_lo_hi_270 = {_memRequest_bits_data_T_3205[262], _memRequest_bits_data_T_2820[262]};
  wire [3:0]        memRequest_bits_data_lo_270 = {memRequest_bits_data_lo_hi_270, memRequest_bits_data_lo_lo_270};
  wire [1:0]        memRequest_bits_data_hi_lo_270 = {_memRequest_bits_data_T_3975[262], _memRequest_bits_data_T_3590[262]};
  wire [1:0]        memRequest_bits_data_hi_hi_270 = {_memRequest_bits_data_T_4745[262], _memRequest_bits_data_T_4360[262]};
  wire [3:0]        memRequest_bits_data_hi_270 = {memRequest_bits_data_hi_hi_270, memRequest_bits_data_hi_lo_270};
  wire [1:0]        memRequest_bits_data_lo_lo_271 = {_memRequest_bits_data_T_2435[263], _memRequest_bits_data_T_2050[263]};
  wire [1:0]        memRequest_bits_data_lo_hi_271 = {_memRequest_bits_data_T_3205[263], _memRequest_bits_data_T_2820[263]};
  wire [3:0]        memRequest_bits_data_lo_271 = {memRequest_bits_data_lo_hi_271, memRequest_bits_data_lo_lo_271};
  wire [1:0]        memRequest_bits_data_hi_lo_271 = {_memRequest_bits_data_T_3975[263], _memRequest_bits_data_T_3590[263]};
  wire [1:0]        memRequest_bits_data_hi_hi_271 = {_memRequest_bits_data_T_4745[263], _memRequest_bits_data_T_4360[263]};
  wire [3:0]        memRequest_bits_data_hi_271 = {memRequest_bits_data_hi_hi_271, memRequest_bits_data_hi_lo_271};
  wire [1:0]        memRequest_bits_data_lo_lo_272 = {_memRequest_bits_data_T_2435[264], _memRequest_bits_data_T_2050[264]};
  wire [1:0]        memRequest_bits_data_lo_hi_272 = {_memRequest_bits_data_T_3205[264], _memRequest_bits_data_T_2820[264]};
  wire [3:0]        memRequest_bits_data_lo_272 = {memRequest_bits_data_lo_hi_272, memRequest_bits_data_lo_lo_272};
  wire [1:0]        memRequest_bits_data_hi_lo_272 = {_memRequest_bits_data_T_3975[264], _memRequest_bits_data_T_3590[264]};
  wire [1:0]        memRequest_bits_data_hi_hi_272 = {_memRequest_bits_data_T_4745[264], _memRequest_bits_data_T_4360[264]};
  wire [3:0]        memRequest_bits_data_hi_272 = {memRequest_bits_data_hi_hi_272, memRequest_bits_data_hi_lo_272};
  wire [1:0]        memRequest_bits_data_lo_lo_273 = {_memRequest_bits_data_T_2435[265], _memRequest_bits_data_T_2050[265]};
  wire [1:0]        memRequest_bits_data_lo_hi_273 = {_memRequest_bits_data_T_3205[265], _memRequest_bits_data_T_2820[265]};
  wire [3:0]        memRequest_bits_data_lo_273 = {memRequest_bits_data_lo_hi_273, memRequest_bits_data_lo_lo_273};
  wire [1:0]        memRequest_bits_data_hi_lo_273 = {_memRequest_bits_data_T_3975[265], _memRequest_bits_data_T_3590[265]};
  wire [1:0]        memRequest_bits_data_hi_hi_273 = {_memRequest_bits_data_T_4745[265], _memRequest_bits_data_T_4360[265]};
  wire [3:0]        memRequest_bits_data_hi_273 = {memRequest_bits_data_hi_hi_273, memRequest_bits_data_hi_lo_273};
  wire [1:0]        memRequest_bits_data_lo_lo_274 = {_memRequest_bits_data_T_2435[266], _memRequest_bits_data_T_2050[266]};
  wire [1:0]        memRequest_bits_data_lo_hi_274 = {_memRequest_bits_data_T_3205[266], _memRequest_bits_data_T_2820[266]};
  wire [3:0]        memRequest_bits_data_lo_274 = {memRequest_bits_data_lo_hi_274, memRequest_bits_data_lo_lo_274};
  wire [1:0]        memRequest_bits_data_hi_lo_274 = {_memRequest_bits_data_T_3975[266], _memRequest_bits_data_T_3590[266]};
  wire [1:0]        memRequest_bits_data_hi_hi_274 = {_memRequest_bits_data_T_4745[266], _memRequest_bits_data_T_4360[266]};
  wire [3:0]        memRequest_bits_data_hi_274 = {memRequest_bits_data_hi_hi_274, memRequest_bits_data_hi_lo_274};
  wire [1:0]        memRequest_bits_data_lo_lo_275 = {_memRequest_bits_data_T_2435[267], _memRequest_bits_data_T_2050[267]};
  wire [1:0]        memRequest_bits_data_lo_hi_275 = {_memRequest_bits_data_T_3205[267], _memRequest_bits_data_T_2820[267]};
  wire [3:0]        memRequest_bits_data_lo_275 = {memRequest_bits_data_lo_hi_275, memRequest_bits_data_lo_lo_275};
  wire [1:0]        memRequest_bits_data_hi_lo_275 = {_memRequest_bits_data_T_3975[267], _memRequest_bits_data_T_3590[267]};
  wire [1:0]        memRequest_bits_data_hi_hi_275 = {_memRequest_bits_data_T_4745[267], _memRequest_bits_data_T_4360[267]};
  wire [3:0]        memRequest_bits_data_hi_275 = {memRequest_bits_data_hi_hi_275, memRequest_bits_data_hi_lo_275};
  wire [1:0]        memRequest_bits_data_lo_lo_276 = {_memRequest_bits_data_T_2435[268], _memRequest_bits_data_T_2050[268]};
  wire [1:0]        memRequest_bits_data_lo_hi_276 = {_memRequest_bits_data_T_3205[268], _memRequest_bits_data_T_2820[268]};
  wire [3:0]        memRequest_bits_data_lo_276 = {memRequest_bits_data_lo_hi_276, memRequest_bits_data_lo_lo_276};
  wire [1:0]        memRequest_bits_data_hi_lo_276 = {_memRequest_bits_data_T_3975[268], _memRequest_bits_data_T_3590[268]};
  wire [1:0]        memRequest_bits_data_hi_hi_276 = {_memRequest_bits_data_T_4745[268], _memRequest_bits_data_T_4360[268]};
  wire [3:0]        memRequest_bits_data_hi_276 = {memRequest_bits_data_hi_hi_276, memRequest_bits_data_hi_lo_276};
  wire [1:0]        memRequest_bits_data_lo_lo_277 = {_memRequest_bits_data_T_2435[269], _memRequest_bits_data_T_2050[269]};
  wire [1:0]        memRequest_bits_data_lo_hi_277 = {_memRequest_bits_data_T_3205[269], _memRequest_bits_data_T_2820[269]};
  wire [3:0]        memRequest_bits_data_lo_277 = {memRequest_bits_data_lo_hi_277, memRequest_bits_data_lo_lo_277};
  wire [1:0]        memRequest_bits_data_hi_lo_277 = {_memRequest_bits_data_T_3975[269], _memRequest_bits_data_T_3590[269]};
  wire [1:0]        memRequest_bits_data_hi_hi_277 = {_memRequest_bits_data_T_4745[269], _memRequest_bits_data_T_4360[269]};
  wire [3:0]        memRequest_bits_data_hi_277 = {memRequest_bits_data_hi_hi_277, memRequest_bits_data_hi_lo_277};
  wire [1:0]        memRequest_bits_data_lo_lo_278 = {_memRequest_bits_data_T_2435[270], _memRequest_bits_data_T_2050[270]};
  wire [1:0]        memRequest_bits_data_lo_hi_278 = {_memRequest_bits_data_T_3205[270], _memRequest_bits_data_T_2820[270]};
  wire [3:0]        memRequest_bits_data_lo_278 = {memRequest_bits_data_lo_hi_278, memRequest_bits_data_lo_lo_278};
  wire [1:0]        memRequest_bits_data_hi_lo_278 = {_memRequest_bits_data_T_3975[270], _memRequest_bits_data_T_3590[270]};
  wire [1:0]        memRequest_bits_data_hi_hi_278 = {_memRequest_bits_data_T_4745[270], _memRequest_bits_data_T_4360[270]};
  wire [3:0]        memRequest_bits_data_hi_278 = {memRequest_bits_data_hi_hi_278, memRequest_bits_data_hi_lo_278};
  wire [1:0]        memRequest_bits_data_lo_lo_279 = {_memRequest_bits_data_T_2435[271], _memRequest_bits_data_T_2050[271]};
  wire [1:0]        memRequest_bits_data_lo_hi_279 = {_memRequest_bits_data_T_3205[271], _memRequest_bits_data_T_2820[271]};
  wire [3:0]        memRequest_bits_data_lo_279 = {memRequest_bits_data_lo_hi_279, memRequest_bits_data_lo_lo_279};
  wire [1:0]        memRequest_bits_data_hi_lo_279 = {_memRequest_bits_data_T_3975[271], _memRequest_bits_data_T_3590[271]};
  wire [1:0]        memRequest_bits_data_hi_hi_279 = {_memRequest_bits_data_T_4745[271], _memRequest_bits_data_T_4360[271]};
  wire [3:0]        memRequest_bits_data_hi_279 = {memRequest_bits_data_hi_hi_279, memRequest_bits_data_hi_lo_279};
  wire [1:0]        memRequest_bits_data_lo_lo_280 = {_memRequest_bits_data_T_2435[272], _memRequest_bits_data_T_2050[272]};
  wire [1:0]        memRequest_bits_data_lo_hi_280 = {_memRequest_bits_data_T_3205[272], _memRequest_bits_data_T_2820[272]};
  wire [3:0]        memRequest_bits_data_lo_280 = {memRequest_bits_data_lo_hi_280, memRequest_bits_data_lo_lo_280};
  wire [1:0]        memRequest_bits_data_hi_lo_280 = {_memRequest_bits_data_T_3975[272], _memRequest_bits_data_T_3590[272]};
  wire [1:0]        memRequest_bits_data_hi_hi_280 = {_memRequest_bits_data_T_4745[272], _memRequest_bits_data_T_4360[272]};
  wire [3:0]        memRequest_bits_data_hi_280 = {memRequest_bits_data_hi_hi_280, memRequest_bits_data_hi_lo_280};
  wire [1:0]        memRequest_bits_data_lo_lo_281 = {_memRequest_bits_data_T_2435[273], _memRequest_bits_data_T_2050[273]};
  wire [1:0]        memRequest_bits_data_lo_hi_281 = {_memRequest_bits_data_T_3205[273], _memRequest_bits_data_T_2820[273]};
  wire [3:0]        memRequest_bits_data_lo_281 = {memRequest_bits_data_lo_hi_281, memRequest_bits_data_lo_lo_281};
  wire [1:0]        memRequest_bits_data_hi_lo_281 = {_memRequest_bits_data_T_3975[273], _memRequest_bits_data_T_3590[273]};
  wire [1:0]        memRequest_bits_data_hi_hi_281 = {_memRequest_bits_data_T_4745[273], _memRequest_bits_data_T_4360[273]};
  wire [3:0]        memRequest_bits_data_hi_281 = {memRequest_bits_data_hi_hi_281, memRequest_bits_data_hi_lo_281};
  wire [1:0]        memRequest_bits_data_lo_lo_282 = {_memRequest_bits_data_T_2435[274], _memRequest_bits_data_T_2050[274]};
  wire [1:0]        memRequest_bits_data_lo_hi_282 = {_memRequest_bits_data_T_3205[274], _memRequest_bits_data_T_2820[274]};
  wire [3:0]        memRequest_bits_data_lo_282 = {memRequest_bits_data_lo_hi_282, memRequest_bits_data_lo_lo_282};
  wire [1:0]        memRequest_bits_data_hi_lo_282 = {_memRequest_bits_data_T_3975[274], _memRequest_bits_data_T_3590[274]};
  wire [1:0]        memRequest_bits_data_hi_hi_282 = {_memRequest_bits_data_T_4745[274], _memRequest_bits_data_T_4360[274]};
  wire [3:0]        memRequest_bits_data_hi_282 = {memRequest_bits_data_hi_hi_282, memRequest_bits_data_hi_lo_282};
  wire [1:0]        memRequest_bits_data_lo_lo_283 = {_memRequest_bits_data_T_2435[275], _memRequest_bits_data_T_2050[275]};
  wire [1:0]        memRequest_bits_data_lo_hi_283 = {_memRequest_bits_data_T_3205[275], _memRequest_bits_data_T_2820[275]};
  wire [3:0]        memRequest_bits_data_lo_283 = {memRequest_bits_data_lo_hi_283, memRequest_bits_data_lo_lo_283};
  wire [1:0]        memRequest_bits_data_hi_lo_283 = {_memRequest_bits_data_T_3975[275], _memRequest_bits_data_T_3590[275]};
  wire [1:0]        memRequest_bits_data_hi_hi_283 = {_memRequest_bits_data_T_4745[275], _memRequest_bits_data_T_4360[275]};
  wire [3:0]        memRequest_bits_data_hi_283 = {memRequest_bits_data_hi_hi_283, memRequest_bits_data_hi_lo_283};
  wire [1:0]        memRequest_bits_data_lo_lo_284 = {_memRequest_bits_data_T_2435[276], _memRequest_bits_data_T_2050[276]};
  wire [1:0]        memRequest_bits_data_lo_hi_284 = {_memRequest_bits_data_T_3205[276], _memRequest_bits_data_T_2820[276]};
  wire [3:0]        memRequest_bits_data_lo_284 = {memRequest_bits_data_lo_hi_284, memRequest_bits_data_lo_lo_284};
  wire [1:0]        memRequest_bits_data_hi_lo_284 = {_memRequest_bits_data_T_3975[276], _memRequest_bits_data_T_3590[276]};
  wire [1:0]        memRequest_bits_data_hi_hi_284 = {_memRequest_bits_data_T_4745[276], _memRequest_bits_data_T_4360[276]};
  wire [3:0]        memRequest_bits_data_hi_284 = {memRequest_bits_data_hi_hi_284, memRequest_bits_data_hi_lo_284};
  wire [1:0]        memRequest_bits_data_lo_lo_285 = {_memRequest_bits_data_T_2435[277], _memRequest_bits_data_T_2050[277]};
  wire [1:0]        memRequest_bits_data_lo_hi_285 = {_memRequest_bits_data_T_3205[277], _memRequest_bits_data_T_2820[277]};
  wire [3:0]        memRequest_bits_data_lo_285 = {memRequest_bits_data_lo_hi_285, memRequest_bits_data_lo_lo_285};
  wire [1:0]        memRequest_bits_data_hi_lo_285 = {_memRequest_bits_data_T_3975[277], _memRequest_bits_data_T_3590[277]};
  wire [1:0]        memRequest_bits_data_hi_hi_285 = {_memRequest_bits_data_T_4745[277], _memRequest_bits_data_T_4360[277]};
  wire [3:0]        memRequest_bits_data_hi_285 = {memRequest_bits_data_hi_hi_285, memRequest_bits_data_hi_lo_285};
  wire [1:0]        memRequest_bits_data_lo_lo_286 = {_memRequest_bits_data_T_2435[278], _memRequest_bits_data_T_2050[278]};
  wire [1:0]        memRequest_bits_data_lo_hi_286 = {_memRequest_bits_data_T_3205[278], _memRequest_bits_data_T_2820[278]};
  wire [3:0]        memRequest_bits_data_lo_286 = {memRequest_bits_data_lo_hi_286, memRequest_bits_data_lo_lo_286};
  wire [1:0]        memRequest_bits_data_hi_lo_286 = {_memRequest_bits_data_T_3975[278], _memRequest_bits_data_T_3590[278]};
  wire [1:0]        memRequest_bits_data_hi_hi_286 = {_memRequest_bits_data_T_4745[278], _memRequest_bits_data_T_4360[278]};
  wire [3:0]        memRequest_bits_data_hi_286 = {memRequest_bits_data_hi_hi_286, memRequest_bits_data_hi_lo_286};
  wire [1:0]        memRequest_bits_data_lo_lo_287 = {_memRequest_bits_data_T_2435[279], _memRequest_bits_data_T_2050[279]};
  wire [1:0]        memRequest_bits_data_lo_hi_287 = {_memRequest_bits_data_T_3205[279], _memRequest_bits_data_T_2820[279]};
  wire [3:0]        memRequest_bits_data_lo_287 = {memRequest_bits_data_lo_hi_287, memRequest_bits_data_lo_lo_287};
  wire [1:0]        memRequest_bits_data_hi_lo_287 = {_memRequest_bits_data_T_3975[279], _memRequest_bits_data_T_3590[279]};
  wire [1:0]        memRequest_bits_data_hi_hi_287 = {_memRequest_bits_data_T_4745[279], _memRequest_bits_data_T_4360[279]};
  wire [3:0]        memRequest_bits_data_hi_287 = {memRequest_bits_data_hi_hi_287, memRequest_bits_data_hi_lo_287};
  wire [1:0]        memRequest_bits_data_lo_lo_288 = {_memRequest_bits_data_T_2435[280], _memRequest_bits_data_T_2050[280]};
  wire [1:0]        memRequest_bits_data_lo_hi_288 = {_memRequest_bits_data_T_3205[280], _memRequest_bits_data_T_2820[280]};
  wire [3:0]        memRequest_bits_data_lo_288 = {memRequest_bits_data_lo_hi_288, memRequest_bits_data_lo_lo_288};
  wire [1:0]        memRequest_bits_data_hi_lo_288 = {_memRequest_bits_data_T_3975[280], _memRequest_bits_data_T_3590[280]};
  wire [1:0]        memRequest_bits_data_hi_hi_288 = {_memRequest_bits_data_T_4745[280], _memRequest_bits_data_T_4360[280]};
  wire [3:0]        memRequest_bits_data_hi_288 = {memRequest_bits_data_hi_hi_288, memRequest_bits_data_hi_lo_288};
  wire [1:0]        memRequest_bits_data_lo_lo_289 = {_memRequest_bits_data_T_2435[281], _memRequest_bits_data_T_2050[281]};
  wire [1:0]        memRequest_bits_data_lo_hi_289 = {_memRequest_bits_data_T_3205[281], _memRequest_bits_data_T_2820[281]};
  wire [3:0]        memRequest_bits_data_lo_289 = {memRequest_bits_data_lo_hi_289, memRequest_bits_data_lo_lo_289};
  wire [1:0]        memRequest_bits_data_hi_lo_289 = {_memRequest_bits_data_T_3975[281], _memRequest_bits_data_T_3590[281]};
  wire [1:0]        memRequest_bits_data_hi_hi_289 = {_memRequest_bits_data_T_4745[281], _memRequest_bits_data_T_4360[281]};
  wire [3:0]        memRequest_bits_data_hi_289 = {memRequest_bits_data_hi_hi_289, memRequest_bits_data_hi_lo_289};
  wire [1:0]        memRequest_bits_data_lo_lo_290 = {_memRequest_bits_data_T_2435[282], _memRequest_bits_data_T_2050[282]};
  wire [1:0]        memRequest_bits_data_lo_hi_290 = {_memRequest_bits_data_T_3205[282], _memRequest_bits_data_T_2820[282]};
  wire [3:0]        memRequest_bits_data_lo_290 = {memRequest_bits_data_lo_hi_290, memRequest_bits_data_lo_lo_290};
  wire [1:0]        memRequest_bits_data_hi_lo_290 = {_memRequest_bits_data_T_3975[282], _memRequest_bits_data_T_3590[282]};
  wire [1:0]        memRequest_bits_data_hi_hi_290 = {_memRequest_bits_data_T_4745[282], _memRequest_bits_data_T_4360[282]};
  wire [3:0]        memRequest_bits_data_hi_290 = {memRequest_bits_data_hi_hi_290, memRequest_bits_data_hi_lo_290};
  wire [1:0]        memRequest_bits_data_lo_lo_291 = {_memRequest_bits_data_T_2435[283], _memRequest_bits_data_T_2050[283]};
  wire [1:0]        memRequest_bits_data_lo_hi_291 = {_memRequest_bits_data_T_3205[283], _memRequest_bits_data_T_2820[283]};
  wire [3:0]        memRequest_bits_data_lo_291 = {memRequest_bits_data_lo_hi_291, memRequest_bits_data_lo_lo_291};
  wire [1:0]        memRequest_bits_data_hi_lo_291 = {_memRequest_bits_data_T_3975[283], _memRequest_bits_data_T_3590[283]};
  wire [1:0]        memRequest_bits_data_hi_hi_291 = {_memRequest_bits_data_T_4745[283], _memRequest_bits_data_T_4360[283]};
  wire [3:0]        memRequest_bits_data_hi_291 = {memRequest_bits_data_hi_hi_291, memRequest_bits_data_hi_lo_291};
  wire [1:0]        memRequest_bits_data_lo_lo_292 = {_memRequest_bits_data_T_2435[284], _memRequest_bits_data_T_2050[284]};
  wire [1:0]        memRequest_bits_data_lo_hi_292 = {_memRequest_bits_data_T_3205[284], _memRequest_bits_data_T_2820[284]};
  wire [3:0]        memRequest_bits_data_lo_292 = {memRequest_bits_data_lo_hi_292, memRequest_bits_data_lo_lo_292};
  wire [1:0]        memRequest_bits_data_hi_lo_292 = {_memRequest_bits_data_T_3975[284], _memRequest_bits_data_T_3590[284]};
  wire [1:0]        memRequest_bits_data_hi_hi_292 = {_memRequest_bits_data_T_4745[284], _memRequest_bits_data_T_4360[284]};
  wire [3:0]        memRequest_bits_data_hi_292 = {memRequest_bits_data_hi_hi_292, memRequest_bits_data_hi_lo_292};
  wire [1:0]        memRequest_bits_data_lo_lo_293 = {_memRequest_bits_data_T_2435[285], _memRequest_bits_data_T_2050[285]};
  wire [1:0]        memRequest_bits_data_lo_hi_293 = {_memRequest_bits_data_T_3205[285], _memRequest_bits_data_T_2820[285]};
  wire [3:0]        memRequest_bits_data_lo_293 = {memRequest_bits_data_lo_hi_293, memRequest_bits_data_lo_lo_293};
  wire [1:0]        memRequest_bits_data_hi_lo_293 = {_memRequest_bits_data_T_3975[285], _memRequest_bits_data_T_3590[285]};
  wire [1:0]        memRequest_bits_data_hi_hi_293 = {_memRequest_bits_data_T_4745[285], _memRequest_bits_data_T_4360[285]};
  wire [3:0]        memRequest_bits_data_hi_293 = {memRequest_bits_data_hi_hi_293, memRequest_bits_data_hi_lo_293};
  wire [1:0]        memRequest_bits_data_lo_lo_294 = {_memRequest_bits_data_T_2435[286], _memRequest_bits_data_T_2050[286]};
  wire [1:0]        memRequest_bits_data_lo_hi_294 = {_memRequest_bits_data_T_3205[286], _memRequest_bits_data_T_2820[286]};
  wire [3:0]        memRequest_bits_data_lo_294 = {memRequest_bits_data_lo_hi_294, memRequest_bits_data_lo_lo_294};
  wire [1:0]        memRequest_bits_data_hi_lo_294 = {_memRequest_bits_data_T_3975[286], _memRequest_bits_data_T_3590[286]};
  wire [1:0]        memRequest_bits_data_hi_hi_294 = {_memRequest_bits_data_T_4745[286], _memRequest_bits_data_T_4360[286]};
  wire [3:0]        memRequest_bits_data_hi_294 = {memRequest_bits_data_hi_hi_294, memRequest_bits_data_hi_lo_294};
  wire [1:0]        memRequest_bits_data_lo_lo_295 = {_memRequest_bits_data_T_2435[287], _memRequest_bits_data_T_2050[287]};
  wire [1:0]        memRequest_bits_data_lo_hi_295 = {_memRequest_bits_data_T_3205[287], _memRequest_bits_data_T_2820[287]};
  wire [3:0]        memRequest_bits_data_lo_295 = {memRequest_bits_data_lo_hi_295, memRequest_bits_data_lo_lo_295};
  wire [1:0]        memRequest_bits_data_hi_lo_295 = {_memRequest_bits_data_T_3975[287], _memRequest_bits_data_T_3590[287]};
  wire [1:0]        memRequest_bits_data_hi_hi_295 = {_memRequest_bits_data_T_4745[287], _memRequest_bits_data_T_4360[287]};
  wire [3:0]        memRequest_bits_data_hi_295 = {memRequest_bits_data_hi_hi_295, memRequest_bits_data_hi_lo_295};
  wire [1:0]        memRequest_bits_data_lo_lo_296 = {_memRequest_bits_data_T_2435[288], _memRequest_bits_data_T_2050[288]};
  wire [1:0]        memRequest_bits_data_lo_hi_296 = {_memRequest_bits_data_T_3205[288], _memRequest_bits_data_T_2820[288]};
  wire [3:0]        memRequest_bits_data_lo_296 = {memRequest_bits_data_lo_hi_296, memRequest_bits_data_lo_lo_296};
  wire [1:0]        memRequest_bits_data_hi_lo_296 = {_memRequest_bits_data_T_3975[288], _memRequest_bits_data_T_3590[288]};
  wire [1:0]        memRequest_bits_data_hi_hi_296 = {_memRequest_bits_data_T_4745[288], _memRequest_bits_data_T_4360[288]};
  wire [3:0]        memRequest_bits_data_hi_296 = {memRequest_bits_data_hi_hi_296, memRequest_bits_data_hi_lo_296};
  wire [1:0]        memRequest_bits_data_lo_lo_297 = {_memRequest_bits_data_T_2435[289], _memRequest_bits_data_T_2050[289]};
  wire [1:0]        memRequest_bits_data_lo_hi_297 = {_memRequest_bits_data_T_3205[289], _memRequest_bits_data_T_2820[289]};
  wire [3:0]        memRequest_bits_data_lo_297 = {memRequest_bits_data_lo_hi_297, memRequest_bits_data_lo_lo_297};
  wire [1:0]        memRequest_bits_data_hi_lo_297 = {_memRequest_bits_data_T_3975[289], _memRequest_bits_data_T_3590[289]};
  wire [1:0]        memRequest_bits_data_hi_hi_297 = {_memRequest_bits_data_T_4745[289], _memRequest_bits_data_T_4360[289]};
  wire [3:0]        memRequest_bits_data_hi_297 = {memRequest_bits_data_hi_hi_297, memRequest_bits_data_hi_lo_297};
  wire [1:0]        memRequest_bits_data_lo_lo_298 = {_memRequest_bits_data_T_2435[290], _memRequest_bits_data_T_2050[290]};
  wire [1:0]        memRequest_bits_data_lo_hi_298 = {_memRequest_bits_data_T_3205[290], _memRequest_bits_data_T_2820[290]};
  wire [3:0]        memRequest_bits_data_lo_298 = {memRequest_bits_data_lo_hi_298, memRequest_bits_data_lo_lo_298};
  wire [1:0]        memRequest_bits_data_hi_lo_298 = {_memRequest_bits_data_T_3975[290], _memRequest_bits_data_T_3590[290]};
  wire [1:0]        memRequest_bits_data_hi_hi_298 = {_memRequest_bits_data_T_4745[290], _memRequest_bits_data_T_4360[290]};
  wire [3:0]        memRequest_bits_data_hi_298 = {memRequest_bits_data_hi_hi_298, memRequest_bits_data_hi_lo_298};
  wire [1:0]        memRequest_bits_data_lo_lo_299 = {_memRequest_bits_data_T_2435[291], _memRequest_bits_data_T_2050[291]};
  wire [1:0]        memRequest_bits_data_lo_hi_299 = {_memRequest_bits_data_T_3205[291], _memRequest_bits_data_T_2820[291]};
  wire [3:0]        memRequest_bits_data_lo_299 = {memRequest_bits_data_lo_hi_299, memRequest_bits_data_lo_lo_299};
  wire [1:0]        memRequest_bits_data_hi_lo_299 = {_memRequest_bits_data_T_3975[291], _memRequest_bits_data_T_3590[291]};
  wire [1:0]        memRequest_bits_data_hi_hi_299 = {_memRequest_bits_data_T_4745[291], _memRequest_bits_data_T_4360[291]};
  wire [3:0]        memRequest_bits_data_hi_299 = {memRequest_bits_data_hi_hi_299, memRequest_bits_data_hi_lo_299};
  wire [1:0]        memRequest_bits_data_lo_lo_300 = {_memRequest_bits_data_T_2435[292], _memRequest_bits_data_T_2050[292]};
  wire [1:0]        memRequest_bits_data_lo_hi_300 = {_memRequest_bits_data_T_3205[292], _memRequest_bits_data_T_2820[292]};
  wire [3:0]        memRequest_bits_data_lo_300 = {memRequest_bits_data_lo_hi_300, memRequest_bits_data_lo_lo_300};
  wire [1:0]        memRequest_bits_data_hi_lo_300 = {_memRequest_bits_data_T_3975[292], _memRequest_bits_data_T_3590[292]};
  wire [1:0]        memRequest_bits_data_hi_hi_300 = {_memRequest_bits_data_T_4745[292], _memRequest_bits_data_T_4360[292]};
  wire [3:0]        memRequest_bits_data_hi_300 = {memRequest_bits_data_hi_hi_300, memRequest_bits_data_hi_lo_300};
  wire [1:0]        memRequest_bits_data_lo_lo_301 = {_memRequest_bits_data_T_2435[293], _memRequest_bits_data_T_2050[293]};
  wire [1:0]        memRequest_bits_data_lo_hi_301 = {_memRequest_bits_data_T_3205[293], _memRequest_bits_data_T_2820[293]};
  wire [3:0]        memRequest_bits_data_lo_301 = {memRequest_bits_data_lo_hi_301, memRequest_bits_data_lo_lo_301};
  wire [1:0]        memRequest_bits_data_hi_lo_301 = {_memRequest_bits_data_T_3975[293], _memRequest_bits_data_T_3590[293]};
  wire [1:0]        memRequest_bits_data_hi_hi_301 = {_memRequest_bits_data_T_4745[293], _memRequest_bits_data_T_4360[293]};
  wire [3:0]        memRequest_bits_data_hi_301 = {memRequest_bits_data_hi_hi_301, memRequest_bits_data_hi_lo_301};
  wire [1:0]        memRequest_bits_data_lo_lo_302 = {_memRequest_bits_data_T_2435[294], _memRequest_bits_data_T_2050[294]};
  wire [1:0]        memRequest_bits_data_lo_hi_302 = {_memRequest_bits_data_T_3205[294], _memRequest_bits_data_T_2820[294]};
  wire [3:0]        memRequest_bits_data_lo_302 = {memRequest_bits_data_lo_hi_302, memRequest_bits_data_lo_lo_302};
  wire [1:0]        memRequest_bits_data_hi_lo_302 = {_memRequest_bits_data_T_3975[294], _memRequest_bits_data_T_3590[294]};
  wire [1:0]        memRequest_bits_data_hi_hi_302 = {_memRequest_bits_data_T_4745[294], _memRequest_bits_data_T_4360[294]};
  wire [3:0]        memRequest_bits_data_hi_302 = {memRequest_bits_data_hi_hi_302, memRequest_bits_data_hi_lo_302};
  wire [1:0]        memRequest_bits_data_lo_lo_303 = {_memRequest_bits_data_T_2435[295], _memRequest_bits_data_T_2050[295]};
  wire [1:0]        memRequest_bits_data_lo_hi_303 = {_memRequest_bits_data_T_3205[295], _memRequest_bits_data_T_2820[295]};
  wire [3:0]        memRequest_bits_data_lo_303 = {memRequest_bits_data_lo_hi_303, memRequest_bits_data_lo_lo_303};
  wire [1:0]        memRequest_bits_data_hi_lo_303 = {_memRequest_bits_data_T_3975[295], _memRequest_bits_data_T_3590[295]};
  wire [1:0]        memRequest_bits_data_hi_hi_303 = {_memRequest_bits_data_T_4745[295], _memRequest_bits_data_T_4360[295]};
  wire [3:0]        memRequest_bits_data_hi_303 = {memRequest_bits_data_hi_hi_303, memRequest_bits_data_hi_lo_303};
  wire [1:0]        memRequest_bits_data_lo_lo_304 = {_memRequest_bits_data_T_2435[296], _memRequest_bits_data_T_2050[296]};
  wire [1:0]        memRequest_bits_data_lo_hi_304 = {_memRequest_bits_data_T_3205[296], _memRequest_bits_data_T_2820[296]};
  wire [3:0]        memRequest_bits_data_lo_304 = {memRequest_bits_data_lo_hi_304, memRequest_bits_data_lo_lo_304};
  wire [1:0]        memRequest_bits_data_hi_lo_304 = {_memRequest_bits_data_T_3975[296], _memRequest_bits_data_T_3590[296]};
  wire [1:0]        memRequest_bits_data_hi_hi_304 = {_memRequest_bits_data_T_4745[296], _memRequest_bits_data_T_4360[296]};
  wire [3:0]        memRequest_bits_data_hi_304 = {memRequest_bits_data_hi_hi_304, memRequest_bits_data_hi_lo_304};
  wire [1:0]        memRequest_bits_data_lo_lo_305 = {_memRequest_bits_data_T_2435[297], _memRequest_bits_data_T_2050[297]};
  wire [1:0]        memRequest_bits_data_lo_hi_305 = {_memRequest_bits_data_T_3205[297], _memRequest_bits_data_T_2820[297]};
  wire [3:0]        memRequest_bits_data_lo_305 = {memRequest_bits_data_lo_hi_305, memRequest_bits_data_lo_lo_305};
  wire [1:0]        memRequest_bits_data_hi_lo_305 = {_memRequest_bits_data_T_3975[297], _memRequest_bits_data_T_3590[297]};
  wire [1:0]        memRequest_bits_data_hi_hi_305 = {_memRequest_bits_data_T_4745[297], _memRequest_bits_data_T_4360[297]};
  wire [3:0]        memRequest_bits_data_hi_305 = {memRequest_bits_data_hi_hi_305, memRequest_bits_data_hi_lo_305};
  wire [1:0]        memRequest_bits_data_lo_lo_306 = {_memRequest_bits_data_T_2435[298], _memRequest_bits_data_T_2050[298]};
  wire [1:0]        memRequest_bits_data_lo_hi_306 = {_memRequest_bits_data_T_3205[298], _memRequest_bits_data_T_2820[298]};
  wire [3:0]        memRequest_bits_data_lo_306 = {memRequest_bits_data_lo_hi_306, memRequest_bits_data_lo_lo_306};
  wire [1:0]        memRequest_bits_data_hi_lo_306 = {_memRequest_bits_data_T_3975[298], _memRequest_bits_data_T_3590[298]};
  wire [1:0]        memRequest_bits_data_hi_hi_306 = {_memRequest_bits_data_T_4745[298], _memRequest_bits_data_T_4360[298]};
  wire [3:0]        memRequest_bits_data_hi_306 = {memRequest_bits_data_hi_hi_306, memRequest_bits_data_hi_lo_306};
  wire [1:0]        memRequest_bits_data_lo_lo_307 = {_memRequest_bits_data_T_2435[299], _memRequest_bits_data_T_2050[299]};
  wire [1:0]        memRequest_bits_data_lo_hi_307 = {_memRequest_bits_data_T_3205[299], _memRequest_bits_data_T_2820[299]};
  wire [3:0]        memRequest_bits_data_lo_307 = {memRequest_bits_data_lo_hi_307, memRequest_bits_data_lo_lo_307};
  wire [1:0]        memRequest_bits_data_hi_lo_307 = {_memRequest_bits_data_T_3975[299], _memRequest_bits_data_T_3590[299]};
  wire [1:0]        memRequest_bits_data_hi_hi_307 = {_memRequest_bits_data_T_4745[299], _memRequest_bits_data_T_4360[299]};
  wire [3:0]        memRequest_bits_data_hi_307 = {memRequest_bits_data_hi_hi_307, memRequest_bits_data_hi_lo_307};
  wire [1:0]        memRequest_bits_data_lo_lo_308 = {_memRequest_bits_data_T_2435[300], _memRequest_bits_data_T_2050[300]};
  wire [1:0]        memRequest_bits_data_lo_hi_308 = {_memRequest_bits_data_T_3205[300], _memRequest_bits_data_T_2820[300]};
  wire [3:0]        memRequest_bits_data_lo_308 = {memRequest_bits_data_lo_hi_308, memRequest_bits_data_lo_lo_308};
  wire [1:0]        memRequest_bits_data_hi_lo_308 = {_memRequest_bits_data_T_3975[300], _memRequest_bits_data_T_3590[300]};
  wire [1:0]        memRequest_bits_data_hi_hi_308 = {_memRequest_bits_data_T_4745[300], _memRequest_bits_data_T_4360[300]};
  wire [3:0]        memRequest_bits_data_hi_308 = {memRequest_bits_data_hi_hi_308, memRequest_bits_data_hi_lo_308};
  wire [1:0]        memRequest_bits_data_lo_lo_309 = {_memRequest_bits_data_T_2435[301], _memRequest_bits_data_T_2050[301]};
  wire [1:0]        memRequest_bits_data_lo_hi_309 = {_memRequest_bits_data_T_3205[301], _memRequest_bits_data_T_2820[301]};
  wire [3:0]        memRequest_bits_data_lo_309 = {memRequest_bits_data_lo_hi_309, memRequest_bits_data_lo_lo_309};
  wire [1:0]        memRequest_bits_data_hi_lo_309 = {_memRequest_bits_data_T_3975[301], _memRequest_bits_data_T_3590[301]};
  wire [1:0]        memRequest_bits_data_hi_hi_309 = {_memRequest_bits_data_T_4745[301], _memRequest_bits_data_T_4360[301]};
  wire [3:0]        memRequest_bits_data_hi_309 = {memRequest_bits_data_hi_hi_309, memRequest_bits_data_hi_lo_309};
  wire [1:0]        memRequest_bits_data_lo_lo_310 = {_memRequest_bits_data_T_2435[302], _memRequest_bits_data_T_2050[302]};
  wire [1:0]        memRequest_bits_data_lo_hi_310 = {_memRequest_bits_data_T_3205[302], _memRequest_bits_data_T_2820[302]};
  wire [3:0]        memRequest_bits_data_lo_310 = {memRequest_bits_data_lo_hi_310, memRequest_bits_data_lo_lo_310};
  wire [1:0]        memRequest_bits_data_hi_lo_310 = {_memRequest_bits_data_T_3975[302], _memRequest_bits_data_T_3590[302]};
  wire [1:0]        memRequest_bits_data_hi_hi_310 = {_memRequest_bits_data_T_4745[302], _memRequest_bits_data_T_4360[302]};
  wire [3:0]        memRequest_bits_data_hi_310 = {memRequest_bits_data_hi_hi_310, memRequest_bits_data_hi_lo_310};
  wire [1:0]        memRequest_bits_data_lo_lo_311 = {_memRequest_bits_data_T_2435[303], _memRequest_bits_data_T_2050[303]};
  wire [1:0]        memRequest_bits_data_lo_hi_311 = {_memRequest_bits_data_T_3205[303], _memRequest_bits_data_T_2820[303]};
  wire [3:0]        memRequest_bits_data_lo_311 = {memRequest_bits_data_lo_hi_311, memRequest_bits_data_lo_lo_311};
  wire [1:0]        memRequest_bits_data_hi_lo_311 = {_memRequest_bits_data_T_3975[303], _memRequest_bits_data_T_3590[303]};
  wire [1:0]        memRequest_bits_data_hi_hi_311 = {_memRequest_bits_data_T_4745[303], _memRequest_bits_data_T_4360[303]};
  wire [3:0]        memRequest_bits_data_hi_311 = {memRequest_bits_data_hi_hi_311, memRequest_bits_data_hi_lo_311};
  wire [1:0]        memRequest_bits_data_lo_lo_312 = {_memRequest_bits_data_T_2435[304], _memRequest_bits_data_T_2050[304]};
  wire [1:0]        memRequest_bits_data_lo_hi_312 = {_memRequest_bits_data_T_3205[304], _memRequest_bits_data_T_2820[304]};
  wire [3:0]        memRequest_bits_data_lo_312 = {memRequest_bits_data_lo_hi_312, memRequest_bits_data_lo_lo_312};
  wire [1:0]        memRequest_bits_data_hi_lo_312 = {_memRequest_bits_data_T_3975[304], _memRequest_bits_data_T_3590[304]};
  wire [1:0]        memRequest_bits_data_hi_hi_312 = {_memRequest_bits_data_T_4745[304], _memRequest_bits_data_T_4360[304]};
  wire [3:0]        memRequest_bits_data_hi_312 = {memRequest_bits_data_hi_hi_312, memRequest_bits_data_hi_lo_312};
  wire [1:0]        memRequest_bits_data_lo_lo_313 = {_memRequest_bits_data_T_2435[305], _memRequest_bits_data_T_2050[305]};
  wire [1:0]        memRequest_bits_data_lo_hi_313 = {_memRequest_bits_data_T_3205[305], _memRequest_bits_data_T_2820[305]};
  wire [3:0]        memRequest_bits_data_lo_313 = {memRequest_bits_data_lo_hi_313, memRequest_bits_data_lo_lo_313};
  wire [1:0]        memRequest_bits_data_hi_lo_313 = {_memRequest_bits_data_T_3975[305], _memRequest_bits_data_T_3590[305]};
  wire [1:0]        memRequest_bits_data_hi_hi_313 = {_memRequest_bits_data_T_4745[305], _memRequest_bits_data_T_4360[305]};
  wire [3:0]        memRequest_bits_data_hi_313 = {memRequest_bits_data_hi_hi_313, memRequest_bits_data_hi_lo_313};
  wire [1:0]        memRequest_bits_data_lo_lo_314 = {_memRequest_bits_data_T_2435[306], _memRequest_bits_data_T_2050[306]};
  wire [1:0]        memRequest_bits_data_lo_hi_314 = {_memRequest_bits_data_T_3205[306], _memRequest_bits_data_T_2820[306]};
  wire [3:0]        memRequest_bits_data_lo_314 = {memRequest_bits_data_lo_hi_314, memRequest_bits_data_lo_lo_314};
  wire [1:0]        memRequest_bits_data_hi_lo_314 = {_memRequest_bits_data_T_3975[306], _memRequest_bits_data_T_3590[306]};
  wire [1:0]        memRequest_bits_data_hi_hi_314 = {_memRequest_bits_data_T_4745[306], _memRequest_bits_data_T_4360[306]};
  wire [3:0]        memRequest_bits_data_hi_314 = {memRequest_bits_data_hi_hi_314, memRequest_bits_data_hi_lo_314};
  wire [1:0]        memRequest_bits_data_lo_lo_315 = {_memRequest_bits_data_T_2435[307], _memRequest_bits_data_T_2050[307]};
  wire [1:0]        memRequest_bits_data_lo_hi_315 = {_memRequest_bits_data_T_3205[307], _memRequest_bits_data_T_2820[307]};
  wire [3:0]        memRequest_bits_data_lo_315 = {memRequest_bits_data_lo_hi_315, memRequest_bits_data_lo_lo_315};
  wire [1:0]        memRequest_bits_data_hi_lo_315 = {_memRequest_bits_data_T_3975[307], _memRequest_bits_data_T_3590[307]};
  wire [1:0]        memRequest_bits_data_hi_hi_315 = {_memRequest_bits_data_T_4745[307], _memRequest_bits_data_T_4360[307]};
  wire [3:0]        memRequest_bits_data_hi_315 = {memRequest_bits_data_hi_hi_315, memRequest_bits_data_hi_lo_315};
  wire [1:0]        memRequest_bits_data_lo_lo_316 = {_memRequest_bits_data_T_2435[308], _memRequest_bits_data_T_2050[308]};
  wire [1:0]        memRequest_bits_data_lo_hi_316 = {_memRequest_bits_data_T_3205[308], _memRequest_bits_data_T_2820[308]};
  wire [3:0]        memRequest_bits_data_lo_316 = {memRequest_bits_data_lo_hi_316, memRequest_bits_data_lo_lo_316};
  wire [1:0]        memRequest_bits_data_hi_lo_316 = {_memRequest_bits_data_T_3975[308], _memRequest_bits_data_T_3590[308]};
  wire [1:0]        memRequest_bits_data_hi_hi_316 = {_memRequest_bits_data_T_4745[308], _memRequest_bits_data_T_4360[308]};
  wire [3:0]        memRequest_bits_data_hi_316 = {memRequest_bits_data_hi_hi_316, memRequest_bits_data_hi_lo_316};
  wire [1:0]        memRequest_bits_data_lo_lo_317 = {_memRequest_bits_data_T_2435[309], _memRequest_bits_data_T_2050[309]};
  wire [1:0]        memRequest_bits_data_lo_hi_317 = {_memRequest_bits_data_T_3205[309], _memRequest_bits_data_T_2820[309]};
  wire [3:0]        memRequest_bits_data_lo_317 = {memRequest_bits_data_lo_hi_317, memRequest_bits_data_lo_lo_317};
  wire [1:0]        memRequest_bits_data_hi_lo_317 = {_memRequest_bits_data_T_3975[309], _memRequest_bits_data_T_3590[309]};
  wire [1:0]        memRequest_bits_data_hi_hi_317 = {_memRequest_bits_data_T_4745[309], _memRequest_bits_data_T_4360[309]};
  wire [3:0]        memRequest_bits_data_hi_317 = {memRequest_bits_data_hi_hi_317, memRequest_bits_data_hi_lo_317};
  wire [1:0]        memRequest_bits_data_lo_lo_318 = {_memRequest_bits_data_T_2435[310], _memRequest_bits_data_T_2050[310]};
  wire [1:0]        memRequest_bits_data_lo_hi_318 = {_memRequest_bits_data_T_3205[310], _memRequest_bits_data_T_2820[310]};
  wire [3:0]        memRequest_bits_data_lo_318 = {memRequest_bits_data_lo_hi_318, memRequest_bits_data_lo_lo_318};
  wire [1:0]        memRequest_bits_data_hi_lo_318 = {_memRequest_bits_data_T_3975[310], _memRequest_bits_data_T_3590[310]};
  wire [1:0]        memRequest_bits_data_hi_hi_318 = {_memRequest_bits_data_T_4745[310], _memRequest_bits_data_T_4360[310]};
  wire [3:0]        memRequest_bits_data_hi_318 = {memRequest_bits_data_hi_hi_318, memRequest_bits_data_hi_lo_318};
  wire [1:0]        memRequest_bits_data_lo_lo_319 = {_memRequest_bits_data_T_2435[311], _memRequest_bits_data_T_2050[311]};
  wire [1:0]        memRequest_bits_data_lo_hi_319 = {_memRequest_bits_data_T_3205[311], _memRequest_bits_data_T_2820[311]};
  wire [3:0]        memRequest_bits_data_lo_319 = {memRequest_bits_data_lo_hi_319, memRequest_bits_data_lo_lo_319};
  wire [1:0]        memRequest_bits_data_hi_lo_319 = {_memRequest_bits_data_T_3975[311], _memRequest_bits_data_T_3590[311]};
  wire [1:0]        memRequest_bits_data_hi_hi_319 = {_memRequest_bits_data_T_4745[311], _memRequest_bits_data_T_4360[311]};
  wire [3:0]        memRequest_bits_data_hi_319 = {memRequest_bits_data_hi_hi_319, memRequest_bits_data_hi_lo_319};
  wire [1:0]        memRequest_bits_data_lo_lo_320 = {_memRequest_bits_data_T_2435[312], _memRequest_bits_data_T_2050[312]};
  wire [1:0]        memRequest_bits_data_lo_hi_320 = {_memRequest_bits_data_T_3205[312], _memRequest_bits_data_T_2820[312]};
  wire [3:0]        memRequest_bits_data_lo_320 = {memRequest_bits_data_lo_hi_320, memRequest_bits_data_lo_lo_320};
  wire [1:0]        memRequest_bits_data_hi_lo_320 = {_memRequest_bits_data_T_3975[312], _memRequest_bits_data_T_3590[312]};
  wire [1:0]        memRequest_bits_data_hi_hi_320 = {_memRequest_bits_data_T_4745[312], _memRequest_bits_data_T_4360[312]};
  wire [3:0]        memRequest_bits_data_hi_320 = {memRequest_bits_data_hi_hi_320, memRequest_bits_data_hi_lo_320};
  wire [1:0]        memRequest_bits_data_lo_lo_321 = {_memRequest_bits_data_T_2435[313], _memRequest_bits_data_T_2050[313]};
  wire [1:0]        memRequest_bits_data_lo_hi_321 = {_memRequest_bits_data_T_3205[313], _memRequest_bits_data_T_2820[313]};
  wire [3:0]        memRequest_bits_data_lo_321 = {memRequest_bits_data_lo_hi_321, memRequest_bits_data_lo_lo_321};
  wire [1:0]        memRequest_bits_data_hi_lo_321 = {_memRequest_bits_data_T_3975[313], _memRequest_bits_data_T_3590[313]};
  wire [1:0]        memRequest_bits_data_hi_hi_321 = {_memRequest_bits_data_T_4745[313], _memRequest_bits_data_T_4360[313]};
  wire [3:0]        memRequest_bits_data_hi_321 = {memRequest_bits_data_hi_hi_321, memRequest_bits_data_hi_lo_321};
  wire [1:0]        memRequest_bits_data_lo_lo_322 = {_memRequest_bits_data_T_2435[314], _memRequest_bits_data_T_2050[314]};
  wire [1:0]        memRequest_bits_data_lo_hi_322 = {_memRequest_bits_data_T_3205[314], _memRequest_bits_data_T_2820[314]};
  wire [3:0]        memRequest_bits_data_lo_322 = {memRequest_bits_data_lo_hi_322, memRequest_bits_data_lo_lo_322};
  wire [1:0]        memRequest_bits_data_hi_lo_322 = {_memRequest_bits_data_T_3975[314], _memRequest_bits_data_T_3590[314]};
  wire [1:0]        memRequest_bits_data_hi_hi_322 = {_memRequest_bits_data_T_4745[314], _memRequest_bits_data_T_4360[314]};
  wire [3:0]        memRequest_bits_data_hi_322 = {memRequest_bits_data_hi_hi_322, memRequest_bits_data_hi_lo_322};
  wire [1:0]        memRequest_bits_data_lo_lo_323 = {_memRequest_bits_data_T_2435[315], _memRequest_bits_data_T_2050[315]};
  wire [1:0]        memRequest_bits_data_lo_hi_323 = {_memRequest_bits_data_T_3205[315], _memRequest_bits_data_T_2820[315]};
  wire [3:0]        memRequest_bits_data_lo_323 = {memRequest_bits_data_lo_hi_323, memRequest_bits_data_lo_lo_323};
  wire [1:0]        memRequest_bits_data_hi_lo_323 = {_memRequest_bits_data_T_3975[315], _memRequest_bits_data_T_3590[315]};
  wire [1:0]        memRequest_bits_data_hi_hi_323 = {_memRequest_bits_data_T_4745[315], _memRequest_bits_data_T_4360[315]};
  wire [3:0]        memRequest_bits_data_hi_323 = {memRequest_bits_data_hi_hi_323, memRequest_bits_data_hi_lo_323};
  wire [1:0]        memRequest_bits_data_lo_lo_324 = {_memRequest_bits_data_T_2435[316], _memRequest_bits_data_T_2050[316]};
  wire [1:0]        memRequest_bits_data_lo_hi_324 = {_memRequest_bits_data_T_3205[316], _memRequest_bits_data_T_2820[316]};
  wire [3:0]        memRequest_bits_data_lo_324 = {memRequest_bits_data_lo_hi_324, memRequest_bits_data_lo_lo_324};
  wire [1:0]        memRequest_bits_data_hi_lo_324 = {_memRequest_bits_data_T_3975[316], _memRequest_bits_data_T_3590[316]};
  wire [1:0]        memRequest_bits_data_hi_hi_324 = {_memRequest_bits_data_T_4745[316], _memRequest_bits_data_T_4360[316]};
  wire [3:0]        memRequest_bits_data_hi_324 = {memRequest_bits_data_hi_hi_324, memRequest_bits_data_hi_lo_324};
  wire [1:0]        memRequest_bits_data_lo_lo_325 = {_memRequest_bits_data_T_2435[317], _memRequest_bits_data_T_2050[317]};
  wire [1:0]        memRequest_bits_data_lo_hi_325 = {_memRequest_bits_data_T_3205[317], _memRequest_bits_data_T_2820[317]};
  wire [3:0]        memRequest_bits_data_lo_325 = {memRequest_bits_data_lo_hi_325, memRequest_bits_data_lo_lo_325};
  wire [1:0]        memRequest_bits_data_hi_lo_325 = {_memRequest_bits_data_T_3975[317], _memRequest_bits_data_T_3590[317]};
  wire [1:0]        memRequest_bits_data_hi_hi_325 = {_memRequest_bits_data_T_4745[317], _memRequest_bits_data_T_4360[317]};
  wire [3:0]        memRequest_bits_data_hi_325 = {memRequest_bits_data_hi_hi_325, memRequest_bits_data_hi_lo_325};
  wire [1:0]        memRequest_bits_data_lo_lo_326 = {_memRequest_bits_data_T_2435[318], _memRequest_bits_data_T_2050[318]};
  wire [1:0]        memRequest_bits_data_lo_hi_326 = {_memRequest_bits_data_T_3205[318], _memRequest_bits_data_T_2820[318]};
  wire [3:0]        memRequest_bits_data_lo_326 = {memRequest_bits_data_lo_hi_326, memRequest_bits_data_lo_lo_326};
  wire [1:0]        memRequest_bits_data_hi_lo_326 = {_memRequest_bits_data_T_3975[318], _memRequest_bits_data_T_3590[318]};
  wire [1:0]        memRequest_bits_data_hi_hi_326 = {_memRequest_bits_data_T_4745[318], _memRequest_bits_data_T_4360[318]};
  wire [3:0]        memRequest_bits_data_hi_326 = {memRequest_bits_data_hi_hi_326, memRequest_bits_data_hi_lo_326};
  wire [1:0]        memRequest_bits_data_lo_lo_327 = {_memRequest_bits_data_T_2435[319], _memRequest_bits_data_T_2050[319]};
  wire [1:0]        memRequest_bits_data_lo_hi_327 = {_memRequest_bits_data_T_3205[319], _memRequest_bits_data_T_2820[319]};
  wire [3:0]        memRequest_bits_data_lo_327 = {memRequest_bits_data_lo_hi_327, memRequest_bits_data_lo_lo_327};
  wire [1:0]        memRequest_bits_data_hi_lo_327 = {_memRequest_bits_data_T_3975[319], _memRequest_bits_data_T_3590[319]};
  wire [1:0]        memRequest_bits_data_hi_hi_327 = {_memRequest_bits_data_T_4745[319], _memRequest_bits_data_T_4360[319]};
  wire [3:0]        memRequest_bits_data_hi_327 = {memRequest_bits_data_hi_hi_327, memRequest_bits_data_hi_lo_327};
  wire [1:0]        memRequest_bits_data_lo_lo_328 = {_memRequest_bits_data_T_2435[320], _memRequest_bits_data_T_2050[320]};
  wire [1:0]        memRequest_bits_data_lo_hi_328 = {_memRequest_bits_data_T_3205[320], _memRequest_bits_data_T_2820[320]};
  wire [3:0]        memRequest_bits_data_lo_328 = {memRequest_bits_data_lo_hi_328, memRequest_bits_data_lo_lo_328};
  wire [1:0]        memRequest_bits_data_hi_lo_328 = {_memRequest_bits_data_T_3975[320], _memRequest_bits_data_T_3590[320]};
  wire [1:0]        memRequest_bits_data_hi_hi_328 = {_memRequest_bits_data_T_4745[320], _memRequest_bits_data_T_4360[320]};
  wire [3:0]        memRequest_bits_data_hi_328 = {memRequest_bits_data_hi_hi_328, memRequest_bits_data_hi_lo_328};
  wire [1:0]        memRequest_bits_data_lo_lo_329 = {_memRequest_bits_data_T_2435[321], _memRequest_bits_data_T_2050[321]};
  wire [1:0]        memRequest_bits_data_lo_hi_329 = {_memRequest_bits_data_T_3205[321], _memRequest_bits_data_T_2820[321]};
  wire [3:0]        memRequest_bits_data_lo_329 = {memRequest_bits_data_lo_hi_329, memRequest_bits_data_lo_lo_329};
  wire [1:0]        memRequest_bits_data_hi_lo_329 = {_memRequest_bits_data_T_3975[321], _memRequest_bits_data_T_3590[321]};
  wire [1:0]        memRequest_bits_data_hi_hi_329 = {_memRequest_bits_data_T_4745[321], _memRequest_bits_data_T_4360[321]};
  wire [3:0]        memRequest_bits_data_hi_329 = {memRequest_bits_data_hi_hi_329, memRequest_bits_data_hi_lo_329};
  wire [1:0]        memRequest_bits_data_lo_lo_330 = {_memRequest_bits_data_T_2435[322], _memRequest_bits_data_T_2050[322]};
  wire [1:0]        memRequest_bits_data_lo_hi_330 = {_memRequest_bits_data_T_3205[322], _memRequest_bits_data_T_2820[322]};
  wire [3:0]        memRequest_bits_data_lo_330 = {memRequest_bits_data_lo_hi_330, memRequest_bits_data_lo_lo_330};
  wire [1:0]        memRequest_bits_data_hi_lo_330 = {_memRequest_bits_data_T_3975[322], _memRequest_bits_data_T_3590[322]};
  wire [1:0]        memRequest_bits_data_hi_hi_330 = {_memRequest_bits_data_T_4745[322], _memRequest_bits_data_T_4360[322]};
  wire [3:0]        memRequest_bits_data_hi_330 = {memRequest_bits_data_hi_hi_330, memRequest_bits_data_hi_lo_330};
  wire [1:0]        memRequest_bits_data_lo_lo_331 = {_memRequest_bits_data_T_2435[323], _memRequest_bits_data_T_2050[323]};
  wire [1:0]        memRequest_bits_data_lo_hi_331 = {_memRequest_bits_data_T_3205[323], _memRequest_bits_data_T_2820[323]};
  wire [3:0]        memRequest_bits_data_lo_331 = {memRequest_bits_data_lo_hi_331, memRequest_bits_data_lo_lo_331};
  wire [1:0]        memRequest_bits_data_hi_lo_331 = {_memRequest_bits_data_T_3975[323], _memRequest_bits_data_T_3590[323]};
  wire [1:0]        memRequest_bits_data_hi_hi_331 = {_memRequest_bits_data_T_4745[323], _memRequest_bits_data_T_4360[323]};
  wire [3:0]        memRequest_bits_data_hi_331 = {memRequest_bits_data_hi_hi_331, memRequest_bits_data_hi_lo_331};
  wire [1:0]        memRequest_bits_data_lo_lo_332 = {_memRequest_bits_data_T_2435[324], _memRequest_bits_data_T_2050[324]};
  wire [1:0]        memRequest_bits_data_lo_hi_332 = {_memRequest_bits_data_T_3205[324], _memRequest_bits_data_T_2820[324]};
  wire [3:0]        memRequest_bits_data_lo_332 = {memRequest_bits_data_lo_hi_332, memRequest_bits_data_lo_lo_332};
  wire [1:0]        memRequest_bits_data_hi_lo_332 = {_memRequest_bits_data_T_3975[324], _memRequest_bits_data_T_3590[324]};
  wire [1:0]        memRequest_bits_data_hi_hi_332 = {_memRequest_bits_data_T_4745[324], _memRequest_bits_data_T_4360[324]};
  wire [3:0]        memRequest_bits_data_hi_332 = {memRequest_bits_data_hi_hi_332, memRequest_bits_data_hi_lo_332};
  wire [1:0]        memRequest_bits_data_lo_lo_333 = {_memRequest_bits_data_T_2435[325], _memRequest_bits_data_T_2050[325]};
  wire [1:0]        memRequest_bits_data_lo_hi_333 = {_memRequest_bits_data_T_3205[325], _memRequest_bits_data_T_2820[325]};
  wire [3:0]        memRequest_bits_data_lo_333 = {memRequest_bits_data_lo_hi_333, memRequest_bits_data_lo_lo_333};
  wire [1:0]        memRequest_bits_data_hi_lo_333 = {_memRequest_bits_data_T_3975[325], _memRequest_bits_data_T_3590[325]};
  wire [1:0]        memRequest_bits_data_hi_hi_333 = {_memRequest_bits_data_T_4745[325], _memRequest_bits_data_T_4360[325]};
  wire [3:0]        memRequest_bits_data_hi_333 = {memRequest_bits_data_hi_hi_333, memRequest_bits_data_hi_lo_333};
  wire [1:0]        memRequest_bits_data_lo_lo_334 = {_memRequest_bits_data_T_2435[326], _memRequest_bits_data_T_2050[326]};
  wire [1:0]        memRequest_bits_data_lo_hi_334 = {_memRequest_bits_data_T_3205[326], _memRequest_bits_data_T_2820[326]};
  wire [3:0]        memRequest_bits_data_lo_334 = {memRequest_bits_data_lo_hi_334, memRequest_bits_data_lo_lo_334};
  wire [1:0]        memRequest_bits_data_hi_lo_334 = {_memRequest_bits_data_T_3975[326], _memRequest_bits_data_T_3590[326]};
  wire [1:0]        memRequest_bits_data_hi_hi_334 = {_memRequest_bits_data_T_4745[326], _memRequest_bits_data_T_4360[326]};
  wire [3:0]        memRequest_bits_data_hi_334 = {memRequest_bits_data_hi_hi_334, memRequest_bits_data_hi_lo_334};
  wire [1:0]        memRequest_bits_data_lo_lo_335 = {_memRequest_bits_data_T_2435[327], _memRequest_bits_data_T_2050[327]};
  wire [1:0]        memRequest_bits_data_lo_hi_335 = {_memRequest_bits_data_T_3205[327], _memRequest_bits_data_T_2820[327]};
  wire [3:0]        memRequest_bits_data_lo_335 = {memRequest_bits_data_lo_hi_335, memRequest_bits_data_lo_lo_335};
  wire [1:0]        memRequest_bits_data_hi_lo_335 = {_memRequest_bits_data_T_3975[327], _memRequest_bits_data_T_3590[327]};
  wire [1:0]        memRequest_bits_data_hi_hi_335 = {_memRequest_bits_data_T_4745[327], _memRequest_bits_data_T_4360[327]};
  wire [3:0]        memRequest_bits_data_hi_335 = {memRequest_bits_data_hi_hi_335, memRequest_bits_data_hi_lo_335};
  wire [1:0]        memRequest_bits_data_lo_lo_336 = {_memRequest_bits_data_T_2435[328], _memRequest_bits_data_T_2050[328]};
  wire [1:0]        memRequest_bits_data_lo_hi_336 = {_memRequest_bits_data_T_3205[328], _memRequest_bits_data_T_2820[328]};
  wire [3:0]        memRequest_bits_data_lo_336 = {memRequest_bits_data_lo_hi_336, memRequest_bits_data_lo_lo_336};
  wire [1:0]        memRequest_bits_data_hi_lo_336 = {_memRequest_bits_data_T_3975[328], _memRequest_bits_data_T_3590[328]};
  wire [1:0]        memRequest_bits_data_hi_hi_336 = {_memRequest_bits_data_T_4745[328], _memRequest_bits_data_T_4360[328]};
  wire [3:0]        memRequest_bits_data_hi_336 = {memRequest_bits_data_hi_hi_336, memRequest_bits_data_hi_lo_336};
  wire [1:0]        memRequest_bits_data_lo_lo_337 = {_memRequest_bits_data_T_2435[329], _memRequest_bits_data_T_2050[329]};
  wire [1:0]        memRequest_bits_data_lo_hi_337 = {_memRequest_bits_data_T_3205[329], _memRequest_bits_data_T_2820[329]};
  wire [3:0]        memRequest_bits_data_lo_337 = {memRequest_bits_data_lo_hi_337, memRequest_bits_data_lo_lo_337};
  wire [1:0]        memRequest_bits_data_hi_lo_337 = {_memRequest_bits_data_T_3975[329], _memRequest_bits_data_T_3590[329]};
  wire [1:0]        memRequest_bits_data_hi_hi_337 = {_memRequest_bits_data_T_4745[329], _memRequest_bits_data_T_4360[329]};
  wire [3:0]        memRequest_bits_data_hi_337 = {memRequest_bits_data_hi_hi_337, memRequest_bits_data_hi_lo_337};
  wire [1:0]        memRequest_bits_data_lo_lo_338 = {_memRequest_bits_data_T_2435[330], _memRequest_bits_data_T_2050[330]};
  wire [1:0]        memRequest_bits_data_lo_hi_338 = {_memRequest_bits_data_T_3205[330], _memRequest_bits_data_T_2820[330]};
  wire [3:0]        memRequest_bits_data_lo_338 = {memRequest_bits_data_lo_hi_338, memRequest_bits_data_lo_lo_338};
  wire [1:0]        memRequest_bits_data_hi_lo_338 = {_memRequest_bits_data_T_3975[330], _memRequest_bits_data_T_3590[330]};
  wire [1:0]        memRequest_bits_data_hi_hi_338 = {_memRequest_bits_data_T_4745[330], _memRequest_bits_data_T_4360[330]};
  wire [3:0]        memRequest_bits_data_hi_338 = {memRequest_bits_data_hi_hi_338, memRequest_bits_data_hi_lo_338};
  wire [1:0]        memRequest_bits_data_lo_lo_339 = {_memRequest_bits_data_T_2435[331], _memRequest_bits_data_T_2050[331]};
  wire [1:0]        memRequest_bits_data_lo_hi_339 = {_memRequest_bits_data_T_3205[331], _memRequest_bits_data_T_2820[331]};
  wire [3:0]        memRequest_bits_data_lo_339 = {memRequest_bits_data_lo_hi_339, memRequest_bits_data_lo_lo_339};
  wire [1:0]        memRequest_bits_data_hi_lo_339 = {_memRequest_bits_data_T_3975[331], _memRequest_bits_data_T_3590[331]};
  wire [1:0]        memRequest_bits_data_hi_hi_339 = {_memRequest_bits_data_T_4745[331], _memRequest_bits_data_T_4360[331]};
  wire [3:0]        memRequest_bits_data_hi_339 = {memRequest_bits_data_hi_hi_339, memRequest_bits_data_hi_lo_339};
  wire [1:0]        memRequest_bits_data_lo_lo_340 = {_memRequest_bits_data_T_2435[332], _memRequest_bits_data_T_2050[332]};
  wire [1:0]        memRequest_bits_data_lo_hi_340 = {_memRequest_bits_data_T_3205[332], _memRequest_bits_data_T_2820[332]};
  wire [3:0]        memRequest_bits_data_lo_340 = {memRequest_bits_data_lo_hi_340, memRequest_bits_data_lo_lo_340};
  wire [1:0]        memRequest_bits_data_hi_lo_340 = {_memRequest_bits_data_T_3975[332], _memRequest_bits_data_T_3590[332]};
  wire [1:0]        memRequest_bits_data_hi_hi_340 = {_memRequest_bits_data_T_4745[332], _memRequest_bits_data_T_4360[332]};
  wire [3:0]        memRequest_bits_data_hi_340 = {memRequest_bits_data_hi_hi_340, memRequest_bits_data_hi_lo_340};
  wire [1:0]        memRequest_bits_data_lo_lo_341 = {_memRequest_bits_data_T_2435[333], _memRequest_bits_data_T_2050[333]};
  wire [1:0]        memRequest_bits_data_lo_hi_341 = {_memRequest_bits_data_T_3205[333], _memRequest_bits_data_T_2820[333]};
  wire [3:0]        memRequest_bits_data_lo_341 = {memRequest_bits_data_lo_hi_341, memRequest_bits_data_lo_lo_341};
  wire [1:0]        memRequest_bits_data_hi_lo_341 = {_memRequest_bits_data_T_3975[333], _memRequest_bits_data_T_3590[333]};
  wire [1:0]        memRequest_bits_data_hi_hi_341 = {_memRequest_bits_data_T_4745[333], _memRequest_bits_data_T_4360[333]};
  wire [3:0]        memRequest_bits_data_hi_341 = {memRequest_bits_data_hi_hi_341, memRequest_bits_data_hi_lo_341};
  wire [1:0]        memRequest_bits_data_lo_lo_342 = {_memRequest_bits_data_T_2435[334], _memRequest_bits_data_T_2050[334]};
  wire [1:0]        memRequest_bits_data_lo_hi_342 = {_memRequest_bits_data_T_3205[334], _memRequest_bits_data_T_2820[334]};
  wire [3:0]        memRequest_bits_data_lo_342 = {memRequest_bits_data_lo_hi_342, memRequest_bits_data_lo_lo_342};
  wire [1:0]        memRequest_bits_data_hi_lo_342 = {_memRequest_bits_data_T_3975[334], _memRequest_bits_data_T_3590[334]};
  wire [1:0]        memRequest_bits_data_hi_hi_342 = {_memRequest_bits_data_T_4745[334], _memRequest_bits_data_T_4360[334]};
  wire [3:0]        memRequest_bits_data_hi_342 = {memRequest_bits_data_hi_hi_342, memRequest_bits_data_hi_lo_342};
  wire [1:0]        memRequest_bits_data_lo_lo_343 = {_memRequest_bits_data_T_2435[335], _memRequest_bits_data_T_2050[335]};
  wire [1:0]        memRequest_bits_data_lo_hi_343 = {_memRequest_bits_data_T_3205[335], _memRequest_bits_data_T_2820[335]};
  wire [3:0]        memRequest_bits_data_lo_343 = {memRequest_bits_data_lo_hi_343, memRequest_bits_data_lo_lo_343};
  wire [1:0]        memRequest_bits_data_hi_lo_343 = {_memRequest_bits_data_T_3975[335], _memRequest_bits_data_T_3590[335]};
  wire [1:0]        memRequest_bits_data_hi_hi_343 = {_memRequest_bits_data_T_4745[335], _memRequest_bits_data_T_4360[335]};
  wire [3:0]        memRequest_bits_data_hi_343 = {memRequest_bits_data_hi_hi_343, memRequest_bits_data_hi_lo_343};
  wire [1:0]        memRequest_bits_data_lo_lo_344 = {_memRequest_bits_data_T_2435[336], _memRequest_bits_data_T_2050[336]};
  wire [1:0]        memRequest_bits_data_lo_hi_344 = {_memRequest_bits_data_T_3205[336], _memRequest_bits_data_T_2820[336]};
  wire [3:0]        memRequest_bits_data_lo_344 = {memRequest_bits_data_lo_hi_344, memRequest_bits_data_lo_lo_344};
  wire [1:0]        memRequest_bits_data_hi_lo_344 = {_memRequest_bits_data_T_3975[336], _memRequest_bits_data_T_3590[336]};
  wire [1:0]        memRequest_bits_data_hi_hi_344 = {_memRequest_bits_data_T_4745[336], _memRequest_bits_data_T_4360[336]};
  wire [3:0]        memRequest_bits_data_hi_344 = {memRequest_bits_data_hi_hi_344, memRequest_bits_data_hi_lo_344};
  wire [1:0]        memRequest_bits_data_lo_lo_345 = {_memRequest_bits_data_T_2435[337], _memRequest_bits_data_T_2050[337]};
  wire [1:0]        memRequest_bits_data_lo_hi_345 = {_memRequest_bits_data_T_3205[337], _memRequest_bits_data_T_2820[337]};
  wire [3:0]        memRequest_bits_data_lo_345 = {memRequest_bits_data_lo_hi_345, memRequest_bits_data_lo_lo_345};
  wire [1:0]        memRequest_bits_data_hi_lo_345 = {_memRequest_bits_data_T_3975[337], _memRequest_bits_data_T_3590[337]};
  wire [1:0]        memRequest_bits_data_hi_hi_345 = {_memRequest_bits_data_T_4745[337], _memRequest_bits_data_T_4360[337]};
  wire [3:0]        memRequest_bits_data_hi_345 = {memRequest_bits_data_hi_hi_345, memRequest_bits_data_hi_lo_345};
  wire [1:0]        memRequest_bits_data_lo_lo_346 = {_memRequest_bits_data_T_2435[338], _memRequest_bits_data_T_2050[338]};
  wire [1:0]        memRequest_bits_data_lo_hi_346 = {_memRequest_bits_data_T_3205[338], _memRequest_bits_data_T_2820[338]};
  wire [3:0]        memRequest_bits_data_lo_346 = {memRequest_bits_data_lo_hi_346, memRequest_bits_data_lo_lo_346};
  wire [1:0]        memRequest_bits_data_hi_lo_346 = {_memRequest_bits_data_T_3975[338], _memRequest_bits_data_T_3590[338]};
  wire [1:0]        memRequest_bits_data_hi_hi_346 = {_memRequest_bits_data_T_4745[338], _memRequest_bits_data_T_4360[338]};
  wire [3:0]        memRequest_bits_data_hi_346 = {memRequest_bits_data_hi_hi_346, memRequest_bits_data_hi_lo_346};
  wire [1:0]        memRequest_bits_data_lo_lo_347 = {_memRequest_bits_data_T_2435[339], _memRequest_bits_data_T_2050[339]};
  wire [1:0]        memRequest_bits_data_lo_hi_347 = {_memRequest_bits_data_T_3205[339], _memRequest_bits_data_T_2820[339]};
  wire [3:0]        memRequest_bits_data_lo_347 = {memRequest_bits_data_lo_hi_347, memRequest_bits_data_lo_lo_347};
  wire [1:0]        memRequest_bits_data_hi_lo_347 = {_memRequest_bits_data_T_3975[339], _memRequest_bits_data_T_3590[339]};
  wire [1:0]        memRequest_bits_data_hi_hi_347 = {_memRequest_bits_data_T_4745[339], _memRequest_bits_data_T_4360[339]};
  wire [3:0]        memRequest_bits_data_hi_347 = {memRequest_bits_data_hi_hi_347, memRequest_bits_data_hi_lo_347};
  wire [1:0]        memRequest_bits_data_lo_lo_348 = {_memRequest_bits_data_T_2435[340], _memRequest_bits_data_T_2050[340]};
  wire [1:0]        memRequest_bits_data_lo_hi_348 = {_memRequest_bits_data_T_3205[340], _memRequest_bits_data_T_2820[340]};
  wire [3:0]        memRequest_bits_data_lo_348 = {memRequest_bits_data_lo_hi_348, memRequest_bits_data_lo_lo_348};
  wire [1:0]        memRequest_bits_data_hi_lo_348 = {_memRequest_bits_data_T_3975[340], _memRequest_bits_data_T_3590[340]};
  wire [1:0]        memRequest_bits_data_hi_hi_348 = {_memRequest_bits_data_T_4745[340], _memRequest_bits_data_T_4360[340]};
  wire [3:0]        memRequest_bits_data_hi_348 = {memRequest_bits_data_hi_hi_348, memRequest_bits_data_hi_lo_348};
  wire [1:0]        memRequest_bits_data_lo_lo_349 = {_memRequest_bits_data_T_2435[341], _memRequest_bits_data_T_2050[341]};
  wire [1:0]        memRequest_bits_data_lo_hi_349 = {_memRequest_bits_data_T_3205[341], _memRequest_bits_data_T_2820[341]};
  wire [3:0]        memRequest_bits_data_lo_349 = {memRequest_bits_data_lo_hi_349, memRequest_bits_data_lo_lo_349};
  wire [1:0]        memRequest_bits_data_hi_lo_349 = {_memRequest_bits_data_T_3975[341], _memRequest_bits_data_T_3590[341]};
  wire [1:0]        memRequest_bits_data_hi_hi_349 = {_memRequest_bits_data_T_4745[341], _memRequest_bits_data_T_4360[341]};
  wire [3:0]        memRequest_bits_data_hi_349 = {memRequest_bits_data_hi_hi_349, memRequest_bits_data_hi_lo_349};
  wire [1:0]        memRequest_bits_data_lo_lo_350 = {_memRequest_bits_data_T_2435[342], _memRequest_bits_data_T_2050[342]};
  wire [1:0]        memRequest_bits_data_lo_hi_350 = {_memRequest_bits_data_T_3205[342], _memRequest_bits_data_T_2820[342]};
  wire [3:0]        memRequest_bits_data_lo_350 = {memRequest_bits_data_lo_hi_350, memRequest_bits_data_lo_lo_350};
  wire [1:0]        memRequest_bits_data_hi_lo_350 = {_memRequest_bits_data_T_3975[342], _memRequest_bits_data_T_3590[342]};
  wire [1:0]        memRequest_bits_data_hi_hi_350 = {_memRequest_bits_data_T_4745[342], _memRequest_bits_data_T_4360[342]};
  wire [3:0]        memRequest_bits_data_hi_350 = {memRequest_bits_data_hi_hi_350, memRequest_bits_data_hi_lo_350};
  wire [1:0]        memRequest_bits_data_lo_lo_351 = {_memRequest_bits_data_T_2435[343], _memRequest_bits_data_T_2050[343]};
  wire [1:0]        memRequest_bits_data_lo_hi_351 = {_memRequest_bits_data_T_3205[343], _memRequest_bits_data_T_2820[343]};
  wire [3:0]        memRequest_bits_data_lo_351 = {memRequest_bits_data_lo_hi_351, memRequest_bits_data_lo_lo_351};
  wire [1:0]        memRequest_bits_data_hi_lo_351 = {_memRequest_bits_data_T_3975[343], _memRequest_bits_data_T_3590[343]};
  wire [1:0]        memRequest_bits_data_hi_hi_351 = {_memRequest_bits_data_T_4745[343], _memRequest_bits_data_T_4360[343]};
  wire [3:0]        memRequest_bits_data_hi_351 = {memRequest_bits_data_hi_hi_351, memRequest_bits_data_hi_lo_351};
  wire [1:0]        memRequest_bits_data_lo_lo_352 = {_memRequest_bits_data_T_2435[344], _memRequest_bits_data_T_2050[344]};
  wire [1:0]        memRequest_bits_data_lo_hi_352 = {_memRequest_bits_data_T_3205[344], _memRequest_bits_data_T_2820[344]};
  wire [3:0]        memRequest_bits_data_lo_352 = {memRequest_bits_data_lo_hi_352, memRequest_bits_data_lo_lo_352};
  wire [1:0]        memRequest_bits_data_hi_lo_352 = {_memRequest_bits_data_T_3975[344], _memRequest_bits_data_T_3590[344]};
  wire [1:0]        memRequest_bits_data_hi_hi_352 = {_memRequest_bits_data_T_4745[344], _memRequest_bits_data_T_4360[344]};
  wire [3:0]        memRequest_bits_data_hi_352 = {memRequest_bits_data_hi_hi_352, memRequest_bits_data_hi_lo_352};
  wire [1:0]        memRequest_bits_data_lo_lo_353 = {_memRequest_bits_data_T_2435[345], _memRequest_bits_data_T_2050[345]};
  wire [1:0]        memRequest_bits_data_lo_hi_353 = {_memRequest_bits_data_T_3205[345], _memRequest_bits_data_T_2820[345]};
  wire [3:0]        memRequest_bits_data_lo_353 = {memRequest_bits_data_lo_hi_353, memRequest_bits_data_lo_lo_353};
  wire [1:0]        memRequest_bits_data_hi_lo_353 = {_memRequest_bits_data_T_3975[345], _memRequest_bits_data_T_3590[345]};
  wire [1:0]        memRequest_bits_data_hi_hi_353 = {_memRequest_bits_data_T_4745[345], _memRequest_bits_data_T_4360[345]};
  wire [3:0]        memRequest_bits_data_hi_353 = {memRequest_bits_data_hi_hi_353, memRequest_bits_data_hi_lo_353};
  wire [1:0]        memRequest_bits_data_lo_lo_354 = {_memRequest_bits_data_T_2435[346], _memRequest_bits_data_T_2050[346]};
  wire [1:0]        memRequest_bits_data_lo_hi_354 = {_memRequest_bits_data_T_3205[346], _memRequest_bits_data_T_2820[346]};
  wire [3:0]        memRequest_bits_data_lo_354 = {memRequest_bits_data_lo_hi_354, memRequest_bits_data_lo_lo_354};
  wire [1:0]        memRequest_bits_data_hi_lo_354 = {_memRequest_bits_data_T_3975[346], _memRequest_bits_data_T_3590[346]};
  wire [1:0]        memRequest_bits_data_hi_hi_354 = {_memRequest_bits_data_T_4745[346], _memRequest_bits_data_T_4360[346]};
  wire [3:0]        memRequest_bits_data_hi_354 = {memRequest_bits_data_hi_hi_354, memRequest_bits_data_hi_lo_354};
  wire [1:0]        memRequest_bits_data_lo_lo_355 = {_memRequest_bits_data_T_2435[347], _memRequest_bits_data_T_2050[347]};
  wire [1:0]        memRequest_bits_data_lo_hi_355 = {_memRequest_bits_data_T_3205[347], _memRequest_bits_data_T_2820[347]};
  wire [3:0]        memRequest_bits_data_lo_355 = {memRequest_bits_data_lo_hi_355, memRequest_bits_data_lo_lo_355};
  wire [1:0]        memRequest_bits_data_hi_lo_355 = {_memRequest_bits_data_T_3975[347], _memRequest_bits_data_T_3590[347]};
  wire [1:0]        memRequest_bits_data_hi_hi_355 = {_memRequest_bits_data_T_4745[347], _memRequest_bits_data_T_4360[347]};
  wire [3:0]        memRequest_bits_data_hi_355 = {memRequest_bits_data_hi_hi_355, memRequest_bits_data_hi_lo_355};
  wire [1:0]        memRequest_bits_data_lo_lo_356 = {_memRequest_bits_data_T_2435[348], _memRequest_bits_data_T_2050[348]};
  wire [1:0]        memRequest_bits_data_lo_hi_356 = {_memRequest_bits_data_T_3205[348], _memRequest_bits_data_T_2820[348]};
  wire [3:0]        memRequest_bits_data_lo_356 = {memRequest_bits_data_lo_hi_356, memRequest_bits_data_lo_lo_356};
  wire [1:0]        memRequest_bits_data_hi_lo_356 = {_memRequest_bits_data_T_3975[348], _memRequest_bits_data_T_3590[348]};
  wire [1:0]        memRequest_bits_data_hi_hi_356 = {_memRequest_bits_data_T_4745[348], _memRequest_bits_data_T_4360[348]};
  wire [3:0]        memRequest_bits_data_hi_356 = {memRequest_bits_data_hi_hi_356, memRequest_bits_data_hi_lo_356};
  wire [1:0]        memRequest_bits_data_lo_lo_357 = {_memRequest_bits_data_T_2435[349], _memRequest_bits_data_T_2050[349]};
  wire [1:0]        memRequest_bits_data_lo_hi_357 = {_memRequest_bits_data_T_3205[349], _memRequest_bits_data_T_2820[349]};
  wire [3:0]        memRequest_bits_data_lo_357 = {memRequest_bits_data_lo_hi_357, memRequest_bits_data_lo_lo_357};
  wire [1:0]        memRequest_bits_data_hi_lo_357 = {_memRequest_bits_data_T_3975[349], _memRequest_bits_data_T_3590[349]};
  wire [1:0]        memRequest_bits_data_hi_hi_357 = {_memRequest_bits_data_T_4745[349], _memRequest_bits_data_T_4360[349]};
  wire [3:0]        memRequest_bits_data_hi_357 = {memRequest_bits_data_hi_hi_357, memRequest_bits_data_hi_lo_357};
  wire [1:0]        memRequest_bits_data_lo_lo_358 = {_memRequest_bits_data_T_2435[350], _memRequest_bits_data_T_2050[350]};
  wire [1:0]        memRequest_bits_data_lo_hi_358 = {_memRequest_bits_data_T_3205[350], _memRequest_bits_data_T_2820[350]};
  wire [3:0]        memRequest_bits_data_lo_358 = {memRequest_bits_data_lo_hi_358, memRequest_bits_data_lo_lo_358};
  wire [1:0]        memRequest_bits_data_hi_lo_358 = {_memRequest_bits_data_T_3975[350], _memRequest_bits_data_T_3590[350]};
  wire [1:0]        memRequest_bits_data_hi_hi_358 = {_memRequest_bits_data_T_4745[350], _memRequest_bits_data_T_4360[350]};
  wire [3:0]        memRequest_bits_data_hi_358 = {memRequest_bits_data_hi_hi_358, memRequest_bits_data_hi_lo_358};
  wire [1:0]        memRequest_bits_data_lo_lo_359 = {_memRequest_bits_data_T_2435[351], _memRequest_bits_data_T_2050[351]};
  wire [1:0]        memRequest_bits_data_lo_hi_359 = {_memRequest_bits_data_T_3205[351], _memRequest_bits_data_T_2820[351]};
  wire [3:0]        memRequest_bits_data_lo_359 = {memRequest_bits_data_lo_hi_359, memRequest_bits_data_lo_lo_359};
  wire [1:0]        memRequest_bits_data_hi_lo_359 = {_memRequest_bits_data_T_3975[351], _memRequest_bits_data_T_3590[351]};
  wire [1:0]        memRequest_bits_data_hi_hi_359 = {_memRequest_bits_data_T_4745[351], _memRequest_bits_data_T_4360[351]};
  wire [3:0]        memRequest_bits_data_hi_359 = {memRequest_bits_data_hi_hi_359, memRequest_bits_data_hi_lo_359};
  wire [1:0]        memRequest_bits_data_lo_lo_360 = {_memRequest_bits_data_T_2435[352], _memRequest_bits_data_T_2050[352]};
  wire [1:0]        memRequest_bits_data_lo_hi_360 = {_memRequest_bits_data_T_3205[352], _memRequest_bits_data_T_2820[352]};
  wire [3:0]        memRequest_bits_data_lo_360 = {memRequest_bits_data_lo_hi_360, memRequest_bits_data_lo_lo_360};
  wire [1:0]        memRequest_bits_data_hi_lo_360 = {_memRequest_bits_data_T_3975[352], _memRequest_bits_data_T_3590[352]};
  wire [1:0]        memRequest_bits_data_hi_hi_360 = {_memRequest_bits_data_T_4745[352], _memRequest_bits_data_T_4360[352]};
  wire [3:0]        memRequest_bits_data_hi_360 = {memRequest_bits_data_hi_hi_360, memRequest_bits_data_hi_lo_360};
  wire [1:0]        memRequest_bits_data_lo_lo_361 = {_memRequest_bits_data_T_2435[353], _memRequest_bits_data_T_2050[353]};
  wire [1:0]        memRequest_bits_data_lo_hi_361 = {_memRequest_bits_data_T_3205[353], _memRequest_bits_data_T_2820[353]};
  wire [3:0]        memRequest_bits_data_lo_361 = {memRequest_bits_data_lo_hi_361, memRequest_bits_data_lo_lo_361};
  wire [1:0]        memRequest_bits_data_hi_lo_361 = {_memRequest_bits_data_T_3975[353], _memRequest_bits_data_T_3590[353]};
  wire [1:0]        memRequest_bits_data_hi_hi_361 = {_memRequest_bits_data_T_4745[353], _memRequest_bits_data_T_4360[353]};
  wire [3:0]        memRequest_bits_data_hi_361 = {memRequest_bits_data_hi_hi_361, memRequest_bits_data_hi_lo_361};
  wire [1:0]        memRequest_bits_data_lo_lo_362 = {_memRequest_bits_data_T_2435[354], _memRequest_bits_data_T_2050[354]};
  wire [1:0]        memRequest_bits_data_lo_hi_362 = {_memRequest_bits_data_T_3205[354], _memRequest_bits_data_T_2820[354]};
  wire [3:0]        memRequest_bits_data_lo_362 = {memRequest_bits_data_lo_hi_362, memRequest_bits_data_lo_lo_362};
  wire [1:0]        memRequest_bits_data_hi_lo_362 = {_memRequest_bits_data_T_3975[354], _memRequest_bits_data_T_3590[354]};
  wire [1:0]        memRequest_bits_data_hi_hi_362 = {_memRequest_bits_data_T_4745[354], _memRequest_bits_data_T_4360[354]};
  wire [3:0]        memRequest_bits_data_hi_362 = {memRequest_bits_data_hi_hi_362, memRequest_bits_data_hi_lo_362};
  wire [1:0]        memRequest_bits_data_lo_lo_363 = {_memRequest_bits_data_T_2435[355], _memRequest_bits_data_T_2050[355]};
  wire [1:0]        memRequest_bits_data_lo_hi_363 = {_memRequest_bits_data_T_3205[355], _memRequest_bits_data_T_2820[355]};
  wire [3:0]        memRequest_bits_data_lo_363 = {memRequest_bits_data_lo_hi_363, memRequest_bits_data_lo_lo_363};
  wire [1:0]        memRequest_bits_data_hi_lo_363 = {_memRequest_bits_data_T_3975[355], _memRequest_bits_data_T_3590[355]};
  wire [1:0]        memRequest_bits_data_hi_hi_363 = {_memRequest_bits_data_T_4745[355], _memRequest_bits_data_T_4360[355]};
  wire [3:0]        memRequest_bits_data_hi_363 = {memRequest_bits_data_hi_hi_363, memRequest_bits_data_hi_lo_363};
  wire [1:0]        memRequest_bits_data_lo_lo_364 = {_memRequest_bits_data_T_2435[356], _memRequest_bits_data_T_2050[356]};
  wire [1:0]        memRequest_bits_data_lo_hi_364 = {_memRequest_bits_data_T_3205[356], _memRequest_bits_data_T_2820[356]};
  wire [3:0]        memRequest_bits_data_lo_364 = {memRequest_bits_data_lo_hi_364, memRequest_bits_data_lo_lo_364};
  wire [1:0]        memRequest_bits_data_hi_lo_364 = {_memRequest_bits_data_T_3975[356], _memRequest_bits_data_T_3590[356]};
  wire [1:0]        memRequest_bits_data_hi_hi_364 = {_memRequest_bits_data_T_4745[356], _memRequest_bits_data_T_4360[356]};
  wire [3:0]        memRequest_bits_data_hi_364 = {memRequest_bits_data_hi_hi_364, memRequest_bits_data_hi_lo_364};
  wire [1:0]        memRequest_bits_data_lo_lo_365 = {_memRequest_bits_data_T_2435[357], _memRequest_bits_data_T_2050[357]};
  wire [1:0]        memRequest_bits_data_lo_hi_365 = {_memRequest_bits_data_T_3205[357], _memRequest_bits_data_T_2820[357]};
  wire [3:0]        memRequest_bits_data_lo_365 = {memRequest_bits_data_lo_hi_365, memRequest_bits_data_lo_lo_365};
  wire [1:0]        memRequest_bits_data_hi_lo_365 = {_memRequest_bits_data_T_3975[357], _memRequest_bits_data_T_3590[357]};
  wire [1:0]        memRequest_bits_data_hi_hi_365 = {_memRequest_bits_data_T_4745[357], _memRequest_bits_data_T_4360[357]};
  wire [3:0]        memRequest_bits_data_hi_365 = {memRequest_bits_data_hi_hi_365, memRequest_bits_data_hi_lo_365};
  wire [1:0]        memRequest_bits_data_lo_lo_366 = {_memRequest_bits_data_T_2435[358], _memRequest_bits_data_T_2050[358]};
  wire [1:0]        memRequest_bits_data_lo_hi_366 = {_memRequest_bits_data_T_3205[358], _memRequest_bits_data_T_2820[358]};
  wire [3:0]        memRequest_bits_data_lo_366 = {memRequest_bits_data_lo_hi_366, memRequest_bits_data_lo_lo_366};
  wire [1:0]        memRequest_bits_data_hi_lo_366 = {_memRequest_bits_data_T_3975[358], _memRequest_bits_data_T_3590[358]};
  wire [1:0]        memRequest_bits_data_hi_hi_366 = {_memRequest_bits_data_T_4745[358], _memRequest_bits_data_T_4360[358]};
  wire [3:0]        memRequest_bits_data_hi_366 = {memRequest_bits_data_hi_hi_366, memRequest_bits_data_hi_lo_366};
  wire [1:0]        memRequest_bits_data_lo_lo_367 = {_memRequest_bits_data_T_2435[359], _memRequest_bits_data_T_2050[359]};
  wire [1:0]        memRequest_bits_data_lo_hi_367 = {_memRequest_bits_data_T_3205[359], _memRequest_bits_data_T_2820[359]};
  wire [3:0]        memRequest_bits_data_lo_367 = {memRequest_bits_data_lo_hi_367, memRequest_bits_data_lo_lo_367};
  wire [1:0]        memRequest_bits_data_hi_lo_367 = {_memRequest_bits_data_T_3975[359], _memRequest_bits_data_T_3590[359]};
  wire [1:0]        memRequest_bits_data_hi_hi_367 = {_memRequest_bits_data_T_4745[359], _memRequest_bits_data_T_4360[359]};
  wire [3:0]        memRequest_bits_data_hi_367 = {memRequest_bits_data_hi_hi_367, memRequest_bits_data_hi_lo_367};
  wire [1:0]        memRequest_bits_data_lo_lo_368 = {_memRequest_bits_data_T_2435[360], _memRequest_bits_data_T_2050[360]};
  wire [1:0]        memRequest_bits_data_lo_hi_368 = {_memRequest_bits_data_T_3205[360], _memRequest_bits_data_T_2820[360]};
  wire [3:0]        memRequest_bits_data_lo_368 = {memRequest_bits_data_lo_hi_368, memRequest_bits_data_lo_lo_368};
  wire [1:0]        memRequest_bits_data_hi_lo_368 = {_memRequest_bits_data_T_3975[360], _memRequest_bits_data_T_3590[360]};
  wire [1:0]        memRequest_bits_data_hi_hi_368 = {_memRequest_bits_data_T_4745[360], _memRequest_bits_data_T_4360[360]};
  wire [3:0]        memRequest_bits_data_hi_368 = {memRequest_bits_data_hi_hi_368, memRequest_bits_data_hi_lo_368};
  wire [1:0]        memRequest_bits_data_lo_lo_369 = {_memRequest_bits_data_T_2435[361], _memRequest_bits_data_T_2050[361]};
  wire [1:0]        memRequest_bits_data_lo_hi_369 = {_memRequest_bits_data_T_3205[361], _memRequest_bits_data_T_2820[361]};
  wire [3:0]        memRequest_bits_data_lo_369 = {memRequest_bits_data_lo_hi_369, memRequest_bits_data_lo_lo_369};
  wire [1:0]        memRequest_bits_data_hi_lo_369 = {_memRequest_bits_data_T_3975[361], _memRequest_bits_data_T_3590[361]};
  wire [1:0]        memRequest_bits_data_hi_hi_369 = {_memRequest_bits_data_T_4745[361], _memRequest_bits_data_T_4360[361]};
  wire [3:0]        memRequest_bits_data_hi_369 = {memRequest_bits_data_hi_hi_369, memRequest_bits_data_hi_lo_369};
  wire [1:0]        memRequest_bits_data_lo_lo_370 = {_memRequest_bits_data_T_2435[362], _memRequest_bits_data_T_2050[362]};
  wire [1:0]        memRequest_bits_data_lo_hi_370 = {_memRequest_bits_data_T_3205[362], _memRequest_bits_data_T_2820[362]};
  wire [3:0]        memRequest_bits_data_lo_370 = {memRequest_bits_data_lo_hi_370, memRequest_bits_data_lo_lo_370};
  wire [1:0]        memRequest_bits_data_hi_lo_370 = {_memRequest_bits_data_T_3975[362], _memRequest_bits_data_T_3590[362]};
  wire [1:0]        memRequest_bits_data_hi_hi_370 = {_memRequest_bits_data_T_4745[362], _memRequest_bits_data_T_4360[362]};
  wire [3:0]        memRequest_bits_data_hi_370 = {memRequest_bits_data_hi_hi_370, memRequest_bits_data_hi_lo_370};
  wire [1:0]        memRequest_bits_data_lo_lo_371 = {_memRequest_bits_data_T_2435[363], _memRequest_bits_data_T_2050[363]};
  wire [1:0]        memRequest_bits_data_lo_hi_371 = {_memRequest_bits_data_T_3205[363], _memRequest_bits_data_T_2820[363]};
  wire [3:0]        memRequest_bits_data_lo_371 = {memRequest_bits_data_lo_hi_371, memRequest_bits_data_lo_lo_371};
  wire [1:0]        memRequest_bits_data_hi_lo_371 = {_memRequest_bits_data_T_3975[363], _memRequest_bits_data_T_3590[363]};
  wire [1:0]        memRequest_bits_data_hi_hi_371 = {_memRequest_bits_data_T_4745[363], _memRequest_bits_data_T_4360[363]};
  wire [3:0]        memRequest_bits_data_hi_371 = {memRequest_bits_data_hi_hi_371, memRequest_bits_data_hi_lo_371};
  wire [1:0]        memRequest_bits_data_lo_lo_372 = {_memRequest_bits_data_T_2435[364], _memRequest_bits_data_T_2050[364]};
  wire [1:0]        memRequest_bits_data_lo_hi_372 = {_memRequest_bits_data_T_3205[364], _memRequest_bits_data_T_2820[364]};
  wire [3:0]        memRequest_bits_data_lo_372 = {memRequest_bits_data_lo_hi_372, memRequest_bits_data_lo_lo_372};
  wire [1:0]        memRequest_bits_data_hi_lo_372 = {_memRequest_bits_data_T_3975[364], _memRequest_bits_data_T_3590[364]};
  wire [1:0]        memRequest_bits_data_hi_hi_372 = {_memRequest_bits_data_T_4745[364], _memRequest_bits_data_T_4360[364]};
  wire [3:0]        memRequest_bits_data_hi_372 = {memRequest_bits_data_hi_hi_372, memRequest_bits_data_hi_lo_372};
  wire [1:0]        memRequest_bits_data_lo_lo_373 = {_memRequest_bits_data_T_2435[365], _memRequest_bits_data_T_2050[365]};
  wire [1:0]        memRequest_bits_data_lo_hi_373 = {_memRequest_bits_data_T_3205[365], _memRequest_bits_data_T_2820[365]};
  wire [3:0]        memRequest_bits_data_lo_373 = {memRequest_bits_data_lo_hi_373, memRequest_bits_data_lo_lo_373};
  wire [1:0]        memRequest_bits_data_hi_lo_373 = {_memRequest_bits_data_T_3975[365], _memRequest_bits_data_T_3590[365]};
  wire [1:0]        memRequest_bits_data_hi_hi_373 = {_memRequest_bits_data_T_4745[365], _memRequest_bits_data_T_4360[365]};
  wire [3:0]        memRequest_bits_data_hi_373 = {memRequest_bits_data_hi_hi_373, memRequest_bits_data_hi_lo_373};
  wire [1:0]        memRequest_bits_data_lo_lo_374 = {_memRequest_bits_data_T_2435[366], _memRequest_bits_data_T_2050[366]};
  wire [1:0]        memRequest_bits_data_lo_hi_374 = {_memRequest_bits_data_T_3205[366], _memRequest_bits_data_T_2820[366]};
  wire [3:0]        memRequest_bits_data_lo_374 = {memRequest_bits_data_lo_hi_374, memRequest_bits_data_lo_lo_374};
  wire [1:0]        memRequest_bits_data_hi_lo_374 = {_memRequest_bits_data_T_3975[366], _memRequest_bits_data_T_3590[366]};
  wire [1:0]        memRequest_bits_data_hi_hi_374 = {_memRequest_bits_data_T_4745[366], _memRequest_bits_data_T_4360[366]};
  wire [3:0]        memRequest_bits_data_hi_374 = {memRequest_bits_data_hi_hi_374, memRequest_bits_data_hi_lo_374};
  wire [1:0]        memRequest_bits_data_lo_lo_375 = {_memRequest_bits_data_T_2435[367], _memRequest_bits_data_T_2050[367]};
  wire [1:0]        memRequest_bits_data_lo_hi_375 = {_memRequest_bits_data_T_3205[367], _memRequest_bits_data_T_2820[367]};
  wire [3:0]        memRequest_bits_data_lo_375 = {memRequest_bits_data_lo_hi_375, memRequest_bits_data_lo_lo_375};
  wire [1:0]        memRequest_bits_data_hi_lo_375 = {_memRequest_bits_data_T_3975[367], _memRequest_bits_data_T_3590[367]};
  wire [1:0]        memRequest_bits_data_hi_hi_375 = {_memRequest_bits_data_T_4745[367], _memRequest_bits_data_T_4360[367]};
  wire [3:0]        memRequest_bits_data_hi_375 = {memRequest_bits_data_hi_hi_375, memRequest_bits_data_hi_lo_375};
  wire [1:0]        memRequest_bits_data_lo_lo_376 = {_memRequest_bits_data_T_2435[368], _memRequest_bits_data_T_2050[368]};
  wire [1:0]        memRequest_bits_data_lo_hi_376 = {_memRequest_bits_data_T_3205[368], _memRequest_bits_data_T_2820[368]};
  wire [3:0]        memRequest_bits_data_lo_376 = {memRequest_bits_data_lo_hi_376, memRequest_bits_data_lo_lo_376};
  wire [1:0]        memRequest_bits_data_hi_lo_376 = {_memRequest_bits_data_T_3975[368], _memRequest_bits_data_T_3590[368]};
  wire [1:0]        memRequest_bits_data_hi_hi_376 = {_memRequest_bits_data_T_4745[368], _memRequest_bits_data_T_4360[368]};
  wire [3:0]        memRequest_bits_data_hi_376 = {memRequest_bits_data_hi_hi_376, memRequest_bits_data_hi_lo_376};
  wire [1:0]        memRequest_bits_data_lo_lo_377 = {_memRequest_bits_data_T_2435[369], _memRequest_bits_data_T_2050[369]};
  wire [1:0]        memRequest_bits_data_lo_hi_377 = {_memRequest_bits_data_T_3205[369], _memRequest_bits_data_T_2820[369]};
  wire [3:0]        memRequest_bits_data_lo_377 = {memRequest_bits_data_lo_hi_377, memRequest_bits_data_lo_lo_377};
  wire [1:0]        memRequest_bits_data_hi_lo_377 = {_memRequest_bits_data_T_3975[369], _memRequest_bits_data_T_3590[369]};
  wire [1:0]        memRequest_bits_data_hi_hi_377 = {_memRequest_bits_data_T_4745[369], _memRequest_bits_data_T_4360[369]};
  wire [3:0]        memRequest_bits_data_hi_377 = {memRequest_bits_data_hi_hi_377, memRequest_bits_data_hi_lo_377};
  wire [1:0]        memRequest_bits_data_lo_lo_378 = {_memRequest_bits_data_T_2435[370], _memRequest_bits_data_T_2050[370]};
  wire [1:0]        memRequest_bits_data_lo_hi_378 = {_memRequest_bits_data_T_3205[370], _memRequest_bits_data_T_2820[370]};
  wire [3:0]        memRequest_bits_data_lo_378 = {memRequest_bits_data_lo_hi_378, memRequest_bits_data_lo_lo_378};
  wire [1:0]        memRequest_bits_data_hi_lo_378 = {_memRequest_bits_data_T_3975[370], _memRequest_bits_data_T_3590[370]};
  wire [1:0]        memRequest_bits_data_hi_hi_378 = {_memRequest_bits_data_T_4745[370], _memRequest_bits_data_T_4360[370]};
  wire [3:0]        memRequest_bits_data_hi_378 = {memRequest_bits_data_hi_hi_378, memRequest_bits_data_hi_lo_378};
  wire [1:0]        memRequest_bits_data_lo_lo_379 = {_memRequest_bits_data_T_2435[371], _memRequest_bits_data_T_2050[371]};
  wire [1:0]        memRequest_bits_data_lo_hi_379 = {_memRequest_bits_data_T_3205[371], _memRequest_bits_data_T_2820[371]};
  wire [3:0]        memRequest_bits_data_lo_379 = {memRequest_bits_data_lo_hi_379, memRequest_bits_data_lo_lo_379};
  wire [1:0]        memRequest_bits_data_hi_lo_379 = {_memRequest_bits_data_T_3975[371], _memRequest_bits_data_T_3590[371]};
  wire [1:0]        memRequest_bits_data_hi_hi_379 = {_memRequest_bits_data_T_4745[371], _memRequest_bits_data_T_4360[371]};
  wire [3:0]        memRequest_bits_data_hi_379 = {memRequest_bits_data_hi_hi_379, memRequest_bits_data_hi_lo_379};
  wire [1:0]        memRequest_bits_data_lo_lo_380 = {_memRequest_bits_data_T_2435[372], _memRequest_bits_data_T_2050[372]};
  wire [1:0]        memRequest_bits_data_lo_hi_380 = {_memRequest_bits_data_T_3205[372], _memRequest_bits_data_T_2820[372]};
  wire [3:0]        memRequest_bits_data_lo_380 = {memRequest_bits_data_lo_hi_380, memRequest_bits_data_lo_lo_380};
  wire [1:0]        memRequest_bits_data_hi_lo_380 = {_memRequest_bits_data_T_3975[372], _memRequest_bits_data_T_3590[372]};
  wire [1:0]        memRequest_bits_data_hi_hi_380 = {_memRequest_bits_data_T_4745[372], _memRequest_bits_data_T_4360[372]};
  wire [3:0]        memRequest_bits_data_hi_380 = {memRequest_bits_data_hi_hi_380, memRequest_bits_data_hi_lo_380};
  wire [1:0]        memRequest_bits_data_lo_lo_381 = {_memRequest_bits_data_T_2435[373], _memRequest_bits_data_T_2050[373]};
  wire [1:0]        memRequest_bits_data_lo_hi_381 = {_memRequest_bits_data_T_3205[373], _memRequest_bits_data_T_2820[373]};
  wire [3:0]        memRequest_bits_data_lo_381 = {memRequest_bits_data_lo_hi_381, memRequest_bits_data_lo_lo_381};
  wire [1:0]        memRequest_bits_data_hi_lo_381 = {_memRequest_bits_data_T_3975[373], _memRequest_bits_data_T_3590[373]};
  wire [1:0]        memRequest_bits_data_hi_hi_381 = {_memRequest_bits_data_T_4745[373], _memRequest_bits_data_T_4360[373]};
  wire [3:0]        memRequest_bits_data_hi_381 = {memRequest_bits_data_hi_hi_381, memRequest_bits_data_hi_lo_381};
  wire [1:0]        memRequest_bits_data_lo_lo_382 = {_memRequest_bits_data_T_2435[374], _memRequest_bits_data_T_2050[374]};
  wire [1:0]        memRequest_bits_data_lo_hi_382 = {_memRequest_bits_data_T_3205[374], _memRequest_bits_data_T_2820[374]};
  wire [3:0]        memRequest_bits_data_lo_382 = {memRequest_bits_data_lo_hi_382, memRequest_bits_data_lo_lo_382};
  wire [1:0]        memRequest_bits_data_hi_lo_382 = {_memRequest_bits_data_T_3975[374], _memRequest_bits_data_T_3590[374]};
  wire [1:0]        memRequest_bits_data_hi_hi_382 = {_memRequest_bits_data_T_4745[374], _memRequest_bits_data_T_4360[374]};
  wire [3:0]        memRequest_bits_data_hi_382 = {memRequest_bits_data_hi_hi_382, memRequest_bits_data_hi_lo_382};
  wire [1:0]        memRequest_bits_data_lo_lo_383 = {_memRequest_bits_data_T_2435[375], _memRequest_bits_data_T_2050[375]};
  wire [1:0]        memRequest_bits_data_lo_hi_383 = {_memRequest_bits_data_T_3205[375], _memRequest_bits_data_T_2820[375]};
  wire [3:0]        memRequest_bits_data_lo_383 = {memRequest_bits_data_lo_hi_383, memRequest_bits_data_lo_lo_383};
  wire [1:0]        memRequest_bits_data_hi_lo_383 = {_memRequest_bits_data_T_3975[375], _memRequest_bits_data_T_3590[375]};
  wire [1:0]        memRequest_bits_data_hi_hi_383 = {_memRequest_bits_data_T_4745[375], _memRequest_bits_data_T_4360[375]};
  wire [3:0]        memRequest_bits_data_hi_383 = {memRequest_bits_data_hi_hi_383, memRequest_bits_data_hi_lo_383};
  wire [1:0]        memRequest_bits_data_lo_lo_384 = {_memRequest_bits_data_T_2435[376], _memRequest_bits_data_T_2050[376]};
  wire [1:0]        memRequest_bits_data_lo_hi_384 = {_memRequest_bits_data_T_3205[376], _memRequest_bits_data_T_2820[376]};
  wire [3:0]        memRequest_bits_data_lo_384 = {memRequest_bits_data_lo_hi_384, memRequest_bits_data_lo_lo_384};
  wire [1:0]        memRequest_bits_data_hi_lo_384 = {_memRequest_bits_data_T_3975[376], _memRequest_bits_data_T_3590[376]};
  wire [1:0]        memRequest_bits_data_hi_hi_384 = {_memRequest_bits_data_T_4745[376], _memRequest_bits_data_T_4360[376]};
  wire [3:0]        memRequest_bits_data_hi_384 = {memRequest_bits_data_hi_hi_384, memRequest_bits_data_hi_lo_384};
  wire [1:0]        memRequest_bits_data_lo_lo_385 = {_memRequest_bits_data_T_2435[377], _memRequest_bits_data_T_2050[377]};
  wire [1:0]        memRequest_bits_data_lo_hi_385 = {_memRequest_bits_data_T_3205[377], _memRequest_bits_data_T_2820[377]};
  wire [3:0]        memRequest_bits_data_lo_385 = {memRequest_bits_data_lo_hi_385, memRequest_bits_data_lo_lo_385};
  wire [1:0]        memRequest_bits_data_hi_lo_385 = {_memRequest_bits_data_T_3975[377], _memRequest_bits_data_T_3590[377]};
  wire [1:0]        memRequest_bits_data_hi_hi_385 = {_memRequest_bits_data_T_4745[377], _memRequest_bits_data_T_4360[377]};
  wire [3:0]        memRequest_bits_data_hi_385 = {memRequest_bits_data_hi_hi_385, memRequest_bits_data_hi_lo_385};
  wire [1:0]        memRequest_bits_data_lo_lo_386 = {_memRequest_bits_data_T_2435[378], _memRequest_bits_data_T_2050[378]};
  wire [1:0]        memRequest_bits_data_lo_hi_386 = {_memRequest_bits_data_T_3205[378], _memRequest_bits_data_T_2820[378]};
  wire [3:0]        memRequest_bits_data_lo_386 = {memRequest_bits_data_lo_hi_386, memRequest_bits_data_lo_lo_386};
  wire [1:0]        memRequest_bits_data_hi_lo_386 = {_memRequest_bits_data_T_3975[378], _memRequest_bits_data_T_3590[378]};
  wire [1:0]        memRequest_bits_data_hi_hi_386 = {_memRequest_bits_data_T_4745[378], _memRequest_bits_data_T_4360[378]};
  wire [3:0]        memRequest_bits_data_hi_386 = {memRequest_bits_data_hi_hi_386, memRequest_bits_data_hi_lo_386};
  wire [1:0]        memRequest_bits_data_lo_lo_387 = {_memRequest_bits_data_T_2435[379], _memRequest_bits_data_T_2050[379]};
  wire [1:0]        memRequest_bits_data_lo_hi_387 = {_memRequest_bits_data_T_3205[379], _memRequest_bits_data_T_2820[379]};
  wire [3:0]        memRequest_bits_data_lo_387 = {memRequest_bits_data_lo_hi_387, memRequest_bits_data_lo_lo_387};
  wire [1:0]        memRequest_bits_data_hi_lo_387 = {_memRequest_bits_data_T_3975[379], _memRequest_bits_data_T_3590[379]};
  wire [1:0]        memRequest_bits_data_hi_hi_387 = {_memRequest_bits_data_T_4745[379], _memRequest_bits_data_T_4360[379]};
  wire [3:0]        memRequest_bits_data_hi_387 = {memRequest_bits_data_hi_hi_387, memRequest_bits_data_hi_lo_387};
  wire [1:0]        memRequest_bits_data_lo_lo_388 = {_memRequest_bits_data_T_2435[380], _memRequest_bits_data_T_2050[380]};
  wire [1:0]        memRequest_bits_data_lo_hi_388 = {_memRequest_bits_data_T_3205[380], _memRequest_bits_data_T_2820[380]};
  wire [3:0]        memRequest_bits_data_lo_388 = {memRequest_bits_data_lo_hi_388, memRequest_bits_data_lo_lo_388};
  wire [1:0]        memRequest_bits_data_hi_lo_388 = {_memRequest_bits_data_T_3975[380], _memRequest_bits_data_T_3590[380]};
  wire [1:0]        memRequest_bits_data_hi_hi_388 = {_memRequest_bits_data_T_4745[380], _memRequest_bits_data_T_4360[380]};
  wire [3:0]        memRequest_bits_data_hi_388 = {memRequest_bits_data_hi_hi_388, memRequest_bits_data_hi_lo_388};
  wire [1:0]        memRequest_bits_data_lo_lo_389 = {_memRequest_bits_data_T_2435[381], _memRequest_bits_data_T_2050[381]};
  wire [1:0]        memRequest_bits_data_lo_hi_389 = {_memRequest_bits_data_T_3205[381], _memRequest_bits_data_T_2820[381]};
  wire [3:0]        memRequest_bits_data_lo_389 = {memRequest_bits_data_lo_hi_389, memRequest_bits_data_lo_lo_389};
  wire [1:0]        memRequest_bits_data_hi_lo_389 = {_memRequest_bits_data_T_3975[381], _memRequest_bits_data_T_3590[381]};
  wire [1:0]        memRequest_bits_data_hi_hi_389 = {_memRequest_bits_data_T_4745[381], _memRequest_bits_data_T_4360[381]};
  wire [3:0]        memRequest_bits_data_hi_389 = {memRequest_bits_data_hi_hi_389, memRequest_bits_data_hi_lo_389};
  wire [1:0]        memRequest_bits_data_lo_lo_390 = {_memRequest_bits_data_T_2435[382], _memRequest_bits_data_T_2050[382]};
  wire [1:0]        memRequest_bits_data_lo_hi_390 = {_memRequest_bits_data_T_3205[382], _memRequest_bits_data_T_2820[382]};
  wire [3:0]        memRequest_bits_data_lo_390 = {memRequest_bits_data_lo_hi_390, memRequest_bits_data_lo_lo_390};
  wire [1:0]        memRequest_bits_data_hi_lo_390 = {_memRequest_bits_data_T_3975[382], _memRequest_bits_data_T_3590[382]};
  wire [1:0]        memRequest_bits_data_hi_hi_390 = {_memRequest_bits_data_T_4745[382], _memRequest_bits_data_T_4360[382]};
  wire [3:0]        memRequest_bits_data_hi_390 = {memRequest_bits_data_hi_hi_390, memRequest_bits_data_hi_lo_390};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_9, memRequest_bits_data_lo_9, memRequest_bits_data_hi_8, memRequest_bits_data_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_12, memRequest_bits_data_lo_12, memRequest_bits_data_hi_11, memRequest_bits_data_lo_11};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_10, memRequest_bits_data_lo_10};
  wire [39:0]       memRequest_bits_data_lo_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_15, memRequest_bits_data_lo_15, memRequest_bits_data_hi_14, memRequest_bits_data_lo_14};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_13, memRequest_bits_data_lo_13};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_18, memRequest_bits_data_lo_18, memRequest_bits_data_hi_17, memRequest_bits_data_lo_17};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_16, memRequest_bits_data_lo_16};
  wire [47:0]       memRequest_bits_data_lo_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_lo_lo_lo_hi_lo_8};
  wire [87:0]       memRequest_bits_data_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_21, memRequest_bits_data_lo_21, memRequest_bits_data_hi_20, memRequest_bits_data_lo_20};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_19, memRequest_bits_data_lo_19};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_24, memRequest_bits_data_lo_24, memRequest_bits_data_hi_23, memRequest_bits_data_lo_23};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_22, memRequest_bits_data_lo_22};
  wire [47:0]       memRequest_bits_data_lo_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_27, memRequest_bits_data_lo_27, memRequest_bits_data_hi_26, memRequest_bits_data_lo_26};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_25, memRequest_bits_data_lo_25};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_30, memRequest_bits_data_lo_30, memRequest_bits_data_hi_29, memRequest_bits_data_lo_29};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_28, memRequest_bits_data_lo_28};
  wire [47:0]       memRequest_bits_data_lo_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_hi_8, memRequest_bits_data_lo_lo_lo_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_lo_lo_hi_lo_8};
  wire [183:0]      memRequest_bits_data_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_33, memRequest_bits_data_lo_33, memRequest_bits_data_hi_32, memRequest_bits_data_lo_32};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_31, memRequest_bits_data_lo_31};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_36, memRequest_bits_data_lo_36, memRequest_bits_data_hi_35, memRequest_bits_data_lo_35};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_34, memRequest_bits_data_lo_34};
  wire [47:0]       memRequest_bits_data_lo_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_39, memRequest_bits_data_lo_39, memRequest_bits_data_hi_38, memRequest_bits_data_lo_38};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_37, memRequest_bits_data_lo_37};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_42, memRequest_bits_data_lo_42, memRequest_bits_data_hi_41, memRequest_bits_data_lo_41};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_40, memRequest_bits_data_lo_40};
  wire [47:0]       memRequest_bits_data_lo_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_hi_8, memRequest_bits_data_lo_lo_lo_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_lo_hi_8, memRequest_bits_data_lo_lo_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_45, memRequest_bits_data_lo_45, memRequest_bits_data_hi_44, memRequest_bits_data_lo_44};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_43, memRequest_bits_data_lo_43};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_48, memRequest_bits_data_lo_48, memRequest_bits_data_hi_47, memRequest_bits_data_lo_47};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_46, memRequest_bits_data_lo_46};
  wire [47:0]       memRequest_bits_data_lo_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_lo_hi_8, memRequest_bits_data_lo_lo_lo_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_51, memRequest_bits_data_lo_51, memRequest_bits_data_hi_50, memRequest_bits_data_lo_50};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_49, memRequest_bits_data_lo_49};
  wire [15:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_54, memRequest_bits_data_lo_54, memRequest_bits_data_hi_53, memRequest_bits_data_lo_53};
  wire [23:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_52, memRequest_bits_data_lo_52};
  wire [47:0]       memRequest_bits_data_lo_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_hi_8, memRequest_bits_data_lo_lo_lo_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_hi_8, memRequest_bits_data_lo_lo_lo_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_lo_hi_lo_8};
  wire [375:0]      memRequest_bits_data_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_57, memRequest_bits_data_lo_57, memRequest_bits_data_hi_56, memRequest_bits_data_lo_56};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_55, memRequest_bits_data_lo_55};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_60, memRequest_bits_data_lo_60, memRequest_bits_data_hi_59, memRequest_bits_data_lo_59};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_58, memRequest_bits_data_lo_58};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_lo_hi_8, memRequest_bits_data_lo_lo_hi_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_63, memRequest_bits_data_lo_63, memRequest_bits_data_hi_62, memRequest_bits_data_lo_62};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_61, memRequest_bits_data_lo_61};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_66, memRequest_bits_data_lo_66, memRequest_bits_data_hi_65, memRequest_bits_data_lo_65};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_64, memRequest_bits_data_lo_64};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_lo_hi_8, memRequest_bits_data_lo_lo_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_69, memRequest_bits_data_lo_69, memRequest_bits_data_hi_68, memRequest_bits_data_lo_68};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_67, memRequest_bits_data_lo_67};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_72, memRequest_bits_data_lo_72, memRequest_bits_data_hi_71, memRequest_bits_data_lo_71};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_70, memRequest_bits_data_lo_70};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_lo_hi_8, memRequest_bits_data_lo_lo_hi_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_75, memRequest_bits_data_lo_75, memRequest_bits_data_hi_74, memRequest_bits_data_lo_74};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_73, memRequest_bits_data_lo_73};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_78, memRequest_bits_data_lo_78, memRequest_bits_data_hi_77, memRequest_bits_data_lo_77};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_76, memRequest_bits_data_lo_76};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_hi_lo_8};
  wire [191:0]      memRequest_bits_data_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_lo_hi_8, memRequest_bits_data_lo_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_81, memRequest_bits_data_lo_81, memRequest_bits_data_hi_80, memRequest_bits_data_lo_80};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_79, memRequest_bits_data_lo_79};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_84, memRequest_bits_data_lo_84, memRequest_bits_data_hi_83, memRequest_bits_data_lo_83};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_82, memRequest_bits_data_lo_82};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_lo_hi_8, memRequest_bits_data_lo_lo_hi_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_87, memRequest_bits_data_lo_87, memRequest_bits_data_hi_86, memRequest_bits_data_lo_86};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_85, memRequest_bits_data_lo_85};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_90, memRequest_bits_data_lo_90, memRequest_bits_data_hi_89, memRequest_bits_data_lo_89};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_88, memRequest_bits_data_lo_88};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_lo_hi_8, memRequest_bits_data_lo_lo_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_93, memRequest_bits_data_lo_93, memRequest_bits_data_hi_92, memRequest_bits_data_lo_92};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_91, memRequest_bits_data_lo_91};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_96, memRequest_bits_data_lo_96, memRequest_bits_data_hi_95, memRequest_bits_data_lo_95};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_94, memRequest_bits_data_lo_94};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_lo_hi_8, memRequest_bits_data_lo_lo_hi_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_99, memRequest_bits_data_lo_99, memRequest_bits_data_hi_98, memRequest_bits_data_lo_98};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_97, memRequest_bits_data_lo_97};
  wire [15:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_102, memRequest_bits_data_lo_102, memRequest_bits_data_hi_101, memRequest_bits_data_lo_101};
  wire [23:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_100, memRequest_bits_data_lo_100};
  wire [47:0]       memRequest_bits_data_lo_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_hi_8, memRequest_bits_data_lo_lo_hi_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_hi_8, memRequest_bits_data_lo_lo_hi_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_hi_8, memRequest_bits_data_lo_lo_hi_hi_lo_8};
  wire [383:0]      memRequest_bits_data_lo_lo_hi_8 = {memRequest_bits_data_lo_lo_hi_hi_8, memRequest_bits_data_lo_lo_hi_lo_8};
  wire [759:0]      memRequest_bits_data_lo_lo_391 = {memRequest_bits_data_lo_lo_hi_8, memRequest_bits_data_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_105, memRequest_bits_data_lo_105, memRequest_bits_data_hi_104, memRequest_bits_data_lo_104};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_hi, memRequest_bits_data_hi_103, memRequest_bits_data_lo_103};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_108, memRequest_bits_data_lo_108, memRequest_bits_data_hi_107, memRequest_bits_data_lo_107};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_106, memRequest_bits_data_lo_106};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_111, memRequest_bits_data_lo_111, memRequest_bits_data_hi_110, memRequest_bits_data_lo_110};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_109, memRequest_bits_data_lo_109};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_114, memRequest_bits_data_lo_114, memRequest_bits_data_hi_113, memRequest_bits_data_lo_113};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_112, memRequest_bits_data_lo_112};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_lo_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_117, memRequest_bits_data_lo_117, memRequest_bits_data_hi_116, memRequest_bits_data_lo_116};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_115, memRequest_bits_data_lo_115};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_120, memRequest_bits_data_lo_120, memRequest_bits_data_hi_119, memRequest_bits_data_lo_119};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_118, memRequest_bits_data_lo_118};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_123, memRequest_bits_data_lo_123, memRequest_bits_data_hi_122, memRequest_bits_data_lo_122};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_121, memRequest_bits_data_lo_121};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_126, memRequest_bits_data_lo_126, memRequest_bits_data_hi_125, memRequest_bits_data_lo_125};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_124, memRequest_bits_data_lo_124};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_lo_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_lo_hi_lo_8};
  wire [191:0]      memRequest_bits_data_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_129, memRequest_bits_data_lo_129, memRequest_bits_data_hi_128, memRequest_bits_data_lo_128};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_127, memRequest_bits_data_lo_127};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_132, memRequest_bits_data_lo_132, memRequest_bits_data_hi_131, memRequest_bits_data_lo_131};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_130, memRequest_bits_data_lo_130};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_lo_hi_8, memRequest_bits_data_lo_hi_lo_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_135, memRequest_bits_data_lo_135, memRequest_bits_data_hi_134, memRequest_bits_data_lo_134};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_133, memRequest_bits_data_lo_133};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_138, memRequest_bits_data_lo_138, memRequest_bits_data_hi_137, memRequest_bits_data_lo_137};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_136, memRequest_bits_data_lo_136};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_141, memRequest_bits_data_lo_141, memRequest_bits_data_hi_140, memRequest_bits_data_lo_140};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_139, memRequest_bits_data_lo_139};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_144, memRequest_bits_data_lo_144, memRequest_bits_data_hi_143, memRequest_bits_data_lo_143};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_142, memRequest_bits_data_lo_142};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_147, memRequest_bits_data_lo_147, memRequest_bits_data_hi_146, memRequest_bits_data_lo_146};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_145, memRequest_bits_data_lo_145};
  wire [15:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_150, memRequest_bits_data_lo_150, memRequest_bits_data_hi_149, memRequest_bits_data_lo_149};
  wire [23:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_148, memRequest_bits_data_lo_148};
  wire [47:0]       memRequest_bits_data_lo_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_hi_8, memRequest_bits_data_lo_hi_lo_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_lo_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_hi_lo_8};
  wire [383:0]      memRequest_bits_data_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_153, memRequest_bits_data_lo_153, memRequest_bits_data_hi_152, memRequest_bits_data_lo_152};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_151, memRequest_bits_data_lo_151};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_156, memRequest_bits_data_lo_156, memRequest_bits_data_hi_155, memRequest_bits_data_lo_155};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_154, memRequest_bits_data_lo_154};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_lo_hi_8, memRequest_bits_data_lo_hi_hi_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_159, memRequest_bits_data_lo_159, memRequest_bits_data_hi_158, memRequest_bits_data_lo_158};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_157, memRequest_bits_data_lo_157};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_162, memRequest_bits_data_lo_162, memRequest_bits_data_hi_161, memRequest_bits_data_lo_161};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_160, memRequest_bits_data_lo_160};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_lo_hi_8, memRequest_bits_data_lo_hi_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_165, memRequest_bits_data_lo_165, memRequest_bits_data_hi_164, memRequest_bits_data_lo_164};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_163, memRequest_bits_data_lo_163};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_168, memRequest_bits_data_lo_168, memRequest_bits_data_hi_167, memRequest_bits_data_lo_167};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_166, memRequest_bits_data_lo_166};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_lo_hi_8, memRequest_bits_data_lo_hi_hi_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_171, memRequest_bits_data_lo_171, memRequest_bits_data_hi_170, memRequest_bits_data_lo_170};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_169, memRequest_bits_data_lo_169};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_174, memRequest_bits_data_lo_174, memRequest_bits_data_hi_173, memRequest_bits_data_lo_173};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_172, memRequest_bits_data_lo_172};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_hi_lo_8};
  wire [191:0]      memRequest_bits_data_lo_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_lo_hi_8, memRequest_bits_data_lo_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_177, memRequest_bits_data_lo_177, memRequest_bits_data_hi_176, memRequest_bits_data_lo_176};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_175, memRequest_bits_data_lo_175};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_180, memRequest_bits_data_lo_180, memRequest_bits_data_hi_179, memRequest_bits_data_lo_179};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_178, memRequest_bits_data_lo_178};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_lo_hi_8, memRequest_bits_data_lo_hi_hi_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_183, memRequest_bits_data_lo_183, memRequest_bits_data_hi_182, memRequest_bits_data_lo_182};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_181, memRequest_bits_data_lo_181};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_186, memRequest_bits_data_lo_186, memRequest_bits_data_hi_185, memRequest_bits_data_lo_185};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_184, memRequest_bits_data_lo_184};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_hi_8, memRequest_bits_data_lo_hi_hi_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_lo_hi_8, memRequest_bits_data_lo_hi_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_189, memRequest_bits_data_lo_189, memRequest_bits_data_hi_188, memRequest_bits_data_lo_188};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_187, memRequest_bits_data_lo_187};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_192, memRequest_bits_data_lo_192, memRequest_bits_data_hi_191, memRequest_bits_data_lo_191};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_190, memRequest_bits_data_lo_190};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_lo_hi_8, memRequest_bits_data_lo_hi_hi_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_195, memRequest_bits_data_lo_195, memRequest_bits_data_hi_194, memRequest_bits_data_lo_194};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_193, memRequest_bits_data_lo_193};
  wire [15:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_198, memRequest_bits_data_lo_198, memRequest_bits_data_hi_197, memRequest_bits_data_lo_197};
  wire [23:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_196, memRequest_bits_data_lo_196};
  wire [47:0]       memRequest_bits_data_lo_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_lo_hi_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_hi_lo_8};
  wire [383:0]      memRequest_bits_data_lo_hi_hi_8 = {memRequest_bits_data_lo_hi_hi_hi_8, memRequest_bits_data_lo_hi_hi_lo_8};
  wire [767:0]      memRequest_bits_data_lo_hi_391 = {memRequest_bits_data_lo_hi_hi_8, memRequest_bits_data_lo_hi_lo_8};
  wire [1527:0]     memRequest_bits_data_lo_391 = {memRequest_bits_data_lo_hi_391, memRequest_bits_data_lo_lo_391};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_201, memRequest_bits_data_lo_201, memRequest_bits_data_hi_200, memRequest_bits_data_lo_200};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_hi, memRequest_bits_data_hi_199, memRequest_bits_data_lo_199};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_204, memRequest_bits_data_lo_204, memRequest_bits_data_hi_203, memRequest_bits_data_lo_203};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_202, memRequest_bits_data_lo_202};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_207, memRequest_bits_data_lo_207, memRequest_bits_data_hi_206, memRequest_bits_data_lo_206};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_205, memRequest_bits_data_lo_205};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_210, memRequest_bits_data_lo_210, memRequest_bits_data_hi_209, memRequest_bits_data_lo_209};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_208, memRequest_bits_data_lo_208};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_hi_8, memRequest_bits_data_hi_lo_lo_lo_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_213, memRequest_bits_data_lo_213, memRequest_bits_data_hi_212, memRequest_bits_data_lo_212};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_211, memRequest_bits_data_lo_211};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_216, memRequest_bits_data_lo_216, memRequest_bits_data_hi_215, memRequest_bits_data_lo_215};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_214, memRequest_bits_data_lo_214};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_219, memRequest_bits_data_lo_219, memRequest_bits_data_hi_218, memRequest_bits_data_lo_218};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_217, memRequest_bits_data_lo_217};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_222, memRequest_bits_data_lo_222, memRequest_bits_data_hi_221, memRequest_bits_data_lo_221};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_220, memRequest_bits_data_lo_220};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_hi_8, memRequest_bits_data_hi_lo_lo_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_hi_8, memRequest_bits_data_hi_lo_lo_lo_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_225, memRequest_bits_data_lo_225, memRequest_bits_data_hi_224, memRequest_bits_data_lo_224};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_223, memRequest_bits_data_lo_223};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_228, memRequest_bits_data_lo_228, memRequest_bits_data_hi_227, memRequest_bits_data_lo_227};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_226, memRequest_bits_data_lo_226};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_231, memRequest_bits_data_lo_231, memRequest_bits_data_hi_230, memRequest_bits_data_lo_230};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_229, memRequest_bits_data_lo_229};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_234, memRequest_bits_data_lo_234, memRequest_bits_data_hi_233, memRequest_bits_data_lo_233};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_232, memRequest_bits_data_lo_232};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_lo_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_237, memRequest_bits_data_lo_237, memRequest_bits_data_hi_236, memRequest_bits_data_lo_236};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_235, memRequest_bits_data_lo_235};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_240, memRequest_bits_data_lo_240, memRequest_bits_data_hi_239, memRequest_bits_data_lo_239};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_238, memRequest_bits_data_lo_238};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_243, memRequest_bits_data_lo_243, memRequest_bits_data_hi_242, memRequest_bits_data_lo_242};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_241, memRequest_bits_data_lo_241};
  wire [15:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_246, memRequest_bits_data_lo_246, memRequest_bits_data_hi_245, memRequest_bits_data_lo_245};
  wire [23:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_244, memRequest_bits_data_lo_244};
  wire [47:0]       memRequest_bits_data_hi_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_hi_8, memRequest_bits_data_hi_lo_lo_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_hi_8, memRequest_bits_data_hi_lo_lo_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_lo_hi_hi_8, memRequest_bits_data_hi_lo_lo_hi_lo_8};
  wire [383:0]      memRequest_bits_data_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_249, memRequest_bits_data_lo_249, memRequest_bits_data_hi_248, memRequest_bits_data_lo_248};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_247, memRequest_bits_data_lo_247};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_252, memRequest_bits_data_lo_252, memRequest_bits_data_hi_251, memRequest_bits_data_lo_251};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_250, memRequest_bits_data_lo_250};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_lo_hi_8, memRequest_bits_data_hi_lo_hi_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_255, memRequest_bits_data_lo_255, memRequest_bits_data_hi_254, memRequest_bits_data_lo_254};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_253, memRequest_bits_data_lo_253};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_258, memRequest_bits_data_lo_258, memRequest_bits_data_hi_257, memRequest_bits_data_lo_257};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_256, memRequest_bits_data_lo_256};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_261, memRequest_bits_data_lo_261, memRequest_bits_data_hi_260, memRequest_bits_data_lo_260};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_259, memRequest_bits_data_lo_259};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_264, memRequest_bits_data_lo_264, memRequest_bits_data_hi_263, memRequest_bits_data_lo_263};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_262, memRequest_bits_data_lo_262};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_lo_hi_8, memRequest_bits_data_hi_lo_hi_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_267, memRequest_bits_data_lo_267, memRequest_bits_data_hi_266, memRequest_bits_data_lo_266};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_265, memRequest_bits_data_lo_265};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_270, memRequest_bits_data_lo_270, memRequest_bits_data_hi_269, memRequest_bits_data_lo_269};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_268, memRequest_bits_data_lo_268};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_lo_hi_8, memRequest_bits_data_hi_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_273, memRequest_bits_data_lo_273, memRequest_bits_data_hi_272, memRequest_bits_data_lo_272};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_271, memRequest_bits_data_lo_271};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_276, memRequest_bits_data_lo_276, memRequest_bits_data_hi_275, memRequest_bits_data_lo_275};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_274, memRequest_bits_data_lo_274};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_lo_hi_8, memRequest_bits_data_hi_lo_hi_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_279, memRequest_bits_data_lo_279, memRequest_bits_data_hi_278, memRequest_bits_data_lo_278};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_277, memRequest_bits_data_lo_277};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_282, memRequest_bits_data_lo_282, memRequest_bits_data_hi_281, memRequest_bits_data_lo_281};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_280, memRequest_bits_data_lo_280};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_lo_hi_8, memRequest_bits_data_hi_lo_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_285, memRequest_bits_data_lo_285, memRequest_bits_data_hi_284, memRequest_bits_data_lo_284};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_283, memRequest_bits_data_lo_283};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_288, memRequest_bits_data_lo_288, memRequest_bits_data_hi_287, memRequest_bits_data_lo_287};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_286, memRequest_bits_data_lo_286};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_lo_hi_8, memRequest_bits_data_hi_lo_hi_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_291, memRequest_bits_data_lo_291, memRequest_bits_data_hi_290, memRequest_bits_data_lo_290};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_289, memRequest_bits_data_lo_289};
  wire [15:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_294, memRequest_bits_data_lo_294, memRequest_bits_data_hi_293, memRequest_bits_data_lo_293};
  wire [23:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_292, memRequest_bits_data_lo_292};
  wire [47:0]       memRequest_bits_data_hi_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_hi_8, memRequest_bits_data_hi_lo_hi_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_hi_8, memRequest_bits_data_hi_lo_hi_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_hi_8, memRequest_bits_data_hi_lo_hi_hi_lo_8};
  wire [383:0]      memRequest_bits_data_hi_lo_hi_8 = {memRequest_bits_data_hi_lo_hi_hi_8, memRequest_bits_data_hi_lo_hi_lo_8};
  wire [767:0]      memRequest_bits_data_hi_lo_391 = {memRequest_bits_data_hi_lo_hi_8, memRequest_bits_data_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_297, memRequest_bits_data_lo_297, memRequest_bits_data_hi_296, memRequest_bits_data_lo_296};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_hi, memRequest_bits_data_hi_295, memRequest_bits_data_lo_295};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_300, memRequest_bits_data_lo_300, memRequest_bits_data_hi_299, memRequest_bits_data_lo_299};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_hi, memRequest_bits_data_hi_298, memRequest_bits_data_lo_298};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_303, memRequest_bits_data_lo_303, memRequest_bits_data_hi_302, memRequest_bits_data_lo_302};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_hi, memRequest_bits_data_hi_301, memRequest_bits_data_lo_301};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_306, memRequest_bits_data_lo_306, memRequest_bits_data_hi_305, memRequest_bits_data_lo_305};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_hi, memRequest_bits_data_hi_304, memRequest_bits_data_lo_304};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_hi_8, memRequest_bits_data_hi_hi_lo_lo_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_309, memRequest_bits_data_lo_309, memRequest_bits_data_hi_308, memRequest_bits_data_lo_308};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_hi, memRequest_bits_data_hi_307, memRequest_bits_data_lo_307};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_312, memRequest_bits_data_lo_312, memRequest_bits_data_hi_311, memRequest_bits_data_lo_311};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_hi, memRequest_bits_data_hi_310, memRequest_bits_data_lo_310};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_315, memRequest_bits_data_lo_315, memRequest_bits_data_hi_314, memRequest_bits_data_lo_314};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_hi, memRequest_bits_data_hi_313, memRequest_bits_data_lo_313};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_318, memRequest_bits_data_lo_318, memRequest_bits_data_hi_317, memRequest_bits_data_lo_317};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_hi, memRequest_bits_data_hi_316, memRequest_bits_data_lo_316};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_hi_8, memRequest_bits_data_hi_hi_lo_lo_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_321, memRequest_bits_data_lo_321, memRequest_bits_data_hi_320, memRequest_bits_data_lo_320};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_hi, memRequest_bits_data_hi_319, memRequest_bits_data_lo_319};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_324, memRequest_bits_data_lo_324, memRequest_bits_data_hi_323, memRequest_bits_data_lo_323};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_hi, memRequest_bits_data_hi_322, memRequest_bits_data_lo_322};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_lo_hi_8, memRequest_bits_data_hi_hi_lo_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_327, memRequest_bits_data_lo_327, memRequest_bits_data_hi_326, memRequest_bits_data_lo_326};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_hi, memRequest_bits_data_hi_325, memRequest_bits_data_lo_325};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_330, memRequest_bits_data_lo_330, memRequest_bits_data_hi_329, memRequest_bits_data_lo_329};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_hi, memRequest_bits_data_hi_328, memRequest_bits_data_lo_328};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_hi_8, memRequest_bits_data_hi_hi_lo_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_333, memRequest_bits_data_lo_333, memRequest_bits_data_hi_332, memRequest_bits_data_lo_332};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_hi, memRequest_bits_data_hi_331, memRequest_bits_data_lo_331};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_336, memRequest_bits_data_lo_336, memRequest_bits_data_hi_335, memRequest_bits_data_lo_335};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_hi, memRequest_bits_data_hi_334, memRequest_bits_data_lo_334};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_339, memRequest_bits_data_lo_339, memRequest_bits_data_hi_338, memRequest_bits_data_lo_338};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_hi, memRequest_bits_data_hi_337, memRequest_bits_data_lo_337};
  wire [15:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_342, memRequest_bits_data_lo_342, memRequest_bits_data_hi_341, memRequest_bits_data_lo_341};
  wire [23:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_hi, memRequest_bits_data_hi_340, memRequest_bits_data_lo_340};
  wire [47:0]       memRequest_bits_data_hi_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_lo_hi_hi_8, memRequest_bits_data_hi_hi_lo_hi_lo_8};
  wire [383:0]      memRequest_bits_data_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_hi = {memRequest_bits_data_hi_345, memRequest_bits_data_lo_345, memRequest_bits_data_hi_344, memRequest_bits_data_lo_344};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_hi, memRequest_bits_data_hi_343, memRequest_bits_data_lo_343};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_hi = {memRequest_bits_data_hi_348, memRequest_bits_data_lo_348, memRequest_bits_data_hi_347, memRequest_bits_data_lo_347};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_hi, memRequest_bits_data_hi_346, memRequest_bits_data_lo_346};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_lo_hi_8, memRequest_bits_data_hi_hi_hi_lo_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_hi = {memRequest_bits_data_hi_351, memRequest_bits_data_lo_351, memRequest_bits_data_hi_350, memRequest_bits_data_lo_350};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_hi, memRequest_bits_data_hi_349, memRequest_bits_data_lo_349};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_hi = {memRequest_bits_data_hi_354, memRequest_bits_data_lo_354, memRequest_bits_data_hi_353, memRequest_bits_data_lo_353};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_hi, memRequest_bits_data_hi_352, memRequest_bits_data_lo_352};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_lo_hi_8, memRequest_bits_data_hi_hi_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_hi = {memRequest_bits_data_hi_357, memRequest_bits_data_lo_357, memRequest_bits_data_hi_356, memRequest_bits_data_lo_356};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_hi, memRequest_bits_data_hi_355, memRequest_bits_data_lo_355};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_hi = {memRequest_bits_data_hi_360, memRequest_bits_data_lo_360, memRequest_bits_data_hi_359, memRequest_bits_data_lo_359};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_hi, memRequest_bits_data_hi_358, memRequest_bits_data_lo_358};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_lo_hi_8, memRequest_bits_data_hi_hi_hi_lo_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_hi = {memRequest_bits_data_hi_363, memRequest_bits_data_lo_363, memRequest_bits_data_hi_362, memRequest_bits_data_lo_362};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_hi, memRequest_bits_data_hi_361, memRequest_bits_data_lo_361};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_hi = {memRequest_bits_data_hi_366, memRequest_bits_data_lo_366, memRequest_bits_data_hi_365, memRequest_bits_data_lo_365};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_hi, memRequest_bits_data_hi_364, memRequest_bits_data_lo_364};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_hi = {memRequest_bits_data_hi_369, memRequest_bits_data_lo_369, memRequest_bits_data_hi_368, memRequest_bits_data_lo_368};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_hi, memRequest_bits_data_hi_367, memRequest_bits_data_lo_367};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_hi = {memRequest_bits_data_hi_372, memRequest_bits_data_lo_372, memRequest_bits_data_hi_371, memRequest_bits_data_lo_371};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_hi, memRequest_bits_data_hi_370, memRequest_bits_data_lo_370};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_lo_hi_8, memRequest_bits_data_hi_hi_hi_hi_lo_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_hi = {memRequest_bits_data_hi_375, memRequest_bits_data_lo_375, memRequest_bits_data_hi_374, memRequest_bits_data_lo_374};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_hi, memRequest_bits_data_hi_373, memRequest_bits_data_lo_373};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_hi = {memRequest_bits_data_hi_378, memRequest_bits_data_lo_378, memRequest_bits_data_hi_377, memRequest_bits_data_lo_377};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_hi, memRequest_bits_data_hi_376, memRequest_bits_data_lo_376};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_hi_8, memRequest_bits_data_hi_hi_hi_hi_lo_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_hi = {memRequest_bits_data_hi_381, memRequest_bits_data_lo_381, memRequest_bits_data_hi_380, memRequest_bits_data_lo_380};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_hi, memRequest_bits_data_hi_379, memRequest_bits_data_lo_379};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_hi = {memRequest_bits_data_hi_384, memRequest_bits_data_lo_384, memRequest_bits_data_hi_383, memRequest_bits_data_lo_383};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_hi, memRequest_bits_data_hi_382, memRequest_bits_data_lo_382};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_lo_hi_8, memRequest_bits_data_hi_hi_hi_hi_hi_lo_lo_8};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_hi = {memRequest_bits_data_hi_387, memRequest_bits_data_lo_387, memRequest_bits_data_hi_386, memRequest_bits_data_lo_386};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_hi, memRequest_bits_data_hi_385, memRequest_bits_data_lo_385};
  wire [15:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_hi = {memRequest_bits_data_hi_390, memRequest_bits_data_lo_390, memRequest_bits_data_hi_389, memRequest_bits_data_lo_389};
  wire [23:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_hi, memRequest_bits_data_hi_388, memRequest_bits_data_lo_388};
  wire [47:0]       memRequest_bits_data_hi_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_hi_hi_hi_lo_8};
  wire [95:0]       memRequest_bits_data_hi_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_hi_hi_lo_8};
  wire [191:0]      memRequest_bits_data_hi_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_hi_lo_8};
  wire [383:0]      memRequest_bits_data_hi_hi_hi_8 = {memRequest_bits_data_hi_hi_hi_hi_8, memRequest_bits_data_hi_hi_hi_lo_8};
  wire [767:0]      memRequest_bits_data_hi_hi_391 = {memRequest_bits_data_hi_hi_hi_8, memRequest_bits_data_hi_hi_lo_8};
  wire [1535:0]     memRequest_bits_data_hi_391 = {memRequest_bits_data_hi_hi_391, memRequest_bits_data_hi_lo_391};
  wire [1023:0]     memRequest_bits_data_0 = {memRequest_bits_data_hi_391[519:0], memRequest_bits_data_lo_391[1527:1024]};
  wire [127:0]      selectMaskForTail = bufferValid ? _GEN_1129 : 128'h0;
  wire [382:0]      _memRequest_bits_mask_T_1 = {127'h0, selectMaskForTail, maskTemp} << _GEN_1130;
  wire [127:0]      memRequest_bits_mask_0 = _memRequest_bits_mask_T_1[255:128];
  assign alignedDequeueAddress = {lsuRequestReg_rs1Data[31:7] + {21'h0, bufferBaseCacheLineIndex}, 7'h0};
  wire [31:0]       memRequest_bits_address_0 = alignedDequeueAddress;
  wire [31:0]       addressQueue_enq_bits = alignedDequeueAddress;
  assign addressQueueFree = addressQueue_enq_ready;
  wire              addressQueue_deq_valid;
  assign addressQueue_deq_valid = ~_addressQueue_fifo_empty;
  assign addressQueue_enq_ready = ~_addressQueue_fifo_full;
  wire              _status_idle_output = ~bufferValid & ~readStageValid & readQueueClear & ~bufferFull & ~addressQueue_deq_valid;
  reg               idleNext;
  wire [31:0]       addressQueue_deq_bits;
  always @(posedge clock) begin
    if (reset) begin
      lsuRequestReg_instructionInformation_nf <= 3'h0;
      lsuRequestReg_instructionInformation_mew <= 1'h0;
      lsuRequestReg_instructionInformation_mop <= 2'h0;
      lsuRequestReg_instructionInformation_lumop <= 5'h0;
      lsuRequestReg_instructionInformation_eew <= 2'h0;
      lsuRequestReg_instructionInformation_vs3 <= 5'h0;
      lsuRequestReg_instructionInformation_isStore <= 1'h0;
      lsuRequestReg_instructionInformation_maskedLoadStore <= 1'h0;
      lsuRequestReg_rs1Data <= 32'h0;
      lsuRequestReg_rs2Data <= 32'h0;
      lsuRequestReg_instructionIndex <= 3'h0;
      csrInterfaceReg_vl <= 11'h0;
      csrInterfaceReg_vStart <= 11'h0;
      csrInterfaceReg_vlmul <= 3'h0;
      csrInterfaceReg_vSew <= 2'h0;
      csrInterfaceReg_vxrm <= 2'h0;
      csrInterfaceReg_vta <= 1'h0;
      csrInterfaceReg_vma <= 1'h0;
      requestFireNext <= 1'h0;
      dataEEW <= 2'h0;
      maskReg <= 128'h0;
      needAmend <= 1'h0;
      lastMaskAmendReg <= 127'h0;
      maskGroupCounter <= 3'h0;
      maskCounterInGroup <= 2'h0;
      isLastMaskGroup <= 1'h0;
      accessData_0 <= 1024'h0;
      accessData_1 <= 1024'h0;
      accessData_2 <= 1024'h0;
      accessData_3 <= 1024'h0;
      accessData_4 <= 1024'h0;
      accessData_5 <= 1024'h0;
      accessData_6 <= 1024'h0;
      accessData_7 <= 1024'h0;
      accessPtr <= 3'h0;
      dataGroup <= 3'h0;
      dataBuffer_0 <= 1024'h0;
      dataBuffer_1 <= 1024'h0;
      dataBuffer_2 <= 1024'h0;
      dataBuffer_3 <= 1024'h0;
      dataBuffer_4 <= 1024'h0;
      dataBuffer_5 <= 1024'h0;
      dataBuffer_6 <= 1024'h0;
      dataBuffer_7 <= 1024'h0;
      bufferBaseCacheLineIndex <= 4'h0;
      cacheLineIndexInBuffer <= 3'h0;
      segmentInstructionIndexInterval <= 4'h0;
      lastWriteVrfIndexReg <= 11'h0;
      lastCacheNeedPush <= 1'h0;
      cacheLineNumberReg <= 11'h0;
      lastDataGroupReg <= 7'h0;
      hazardCheck <= 1'h0;
      readStageValid_segPtr <= 3'h0;
      readStageValid_readCount <= 3'h0;
      readStageValid_stageValid <= 1'h0;
      readStageValid_readCounter <= 4'h0;
      readStageValid_segPtr_1 <= 3'h0;
      readStageValid_readCount_1 <= 3'h0;
      readStageValid_stageValid_1 <= 1'h0;
      readStageValid_readCounter_1 <= 4'h0;
      readStageValid_segPtr_2 <= 3'h0;
      readStageValid_readCount_2 <= 3'h0;
      readStageValid_stageValid_2 <= 1'h0;
      readStageValid_readCounter_2 <= 4'h0;
      readStageValid_segPtr_3 <= 3'h0;
      readStageValid_readCount_3 <= 3'h0;
      readStageValid_stageValid_3 <= 1'h0;
      readStageValid_readCounter_3 <= 4'h0;
      readStageValid_segPtr_4 <= 3'h0;
      readStageValid_readCount_4 <= 3'h0;
      readStageValid_stageValid_4 <= 1'h0;
      readStageValid_readCounter_4 <= 4'h0;
      readStageValid_segPtr_5 <= 3'h0;
      readStageValid_readCount_5 <= 3'h0;
      readStageValid_stageValid_5 <= 1'h0;
      readStageValid_readCounter_5 <= 4'h0;
      readStageValid_segPtr_6 <= 3'h0;
      readStageValid_readCount_6 <= 3'h0;
      readStageValid_stageValid_6 <= 1'h0;
      readStageValid_readCounter_6 <= 4'h0;
      readStageValid_segPtr_7 <= 3'h0;
      readStageValid_readCount_7 <= 3'h0;
      readStageValid_stageValid_7 <= 1'h0;
      readStageValid_readCounter_7 <= 4'h0;
      readStageValid_segPtr_8 <= 3'h0;
      readStageValid_readCount_8 <= 3'h0;
      readStageValid_stageValid_8 <= 1'h0;
      readStageValid_readCounter_8 <= 4'h0;
      readStageValid_segPtr_9 <= 3'h0;
      readStageValid_readCount_9 <= 3'h0;
      readStageValid_stageValid_9 <= 1'h0;
      readStageValid_readCounter_9 <= 4'h0;
      readStageValid_segPtr_10 <= 3'h0;
      readStageValid_readCount_10 <= 3'h0;
      readStageValid_stageValid_10 <= 1'h0;
      readStageValid_readCounter_10 <= 4'h0;
      readStageValid_segPtr_11 <= 3'h0;
      readStageValid_readCount_11 <= 3'h0;
      readStageValid_stageValid_11 <= 1'h0;
      readStageValid_readCounter_11 <= 4'h0;
      readStageValid_segPtr_12 <= 3'h0;
      readStageValid_readCount_12 <= 3'h0;
      readStageValid_stageValid_12 <= 1'h0;
      readStageValid_readCounter_12 <= 4'h0;
      readStageValid_segPtr_13 <= 3'h0;
      readStageValid_readCount_13 <= 3'h0;
      readStageValid_stageValid_13 <= 1'h0;
      readStageValid_readCounter_13 <= 4'h0;
      readStageValid_segPtr_14 <= 3'h0;
      readStageValid_readCount_14 <= 3'h0;
      readStageValid_stageValid_14 <= 1'h0;
      readStageValid_readCounter_14 <= 4'h0;
      readStageValid_segPtr_15 <= 3'h0;
      readStageValid_readCount_15 <= 3'h0;
      readStageValid_stageValid_15 <= 1'h0;
      readStageValid_readCounter_15 <= 4'h0;
      readStageValid_segPtr_16 <= 3'h0;
      readStageValid_readCount_16 <= 3'h0;
      readStageValid_stageValid_16 <= 1'h0;
      readStageValid_readCounter_16 <= 4'h0;
      readStageValid_segPtr_17 <= 3'h0;
      readStageValid_readCount_17 <= 3'h0;
      readStageValid_stageValid_17 <= 1'h0;
      readStageValid_readCounter_17 <= 4'h0;
      readStageValid_segPtr_18 <= 3'h0;
      readStageValid_readCount_18 <= 3'h0;
      readStageValid_stageValid_18 <= 1'h0;
      readStageValid_readCounter_18 <= 4'h0;
      readStageValid_segPtr_19 <= 3'h0;
      readStageValid_readCount_19 <= 3'h0;
      readStageValid_stageValid_19 <= 1'h0;
      readStageValid_readCounter_19 <= 4'h0;
      readStageValid_segPtr_20 <= 3'h0;
      readStageValid_readCount_20 <= 3'h0;
      readStageValid_stageValid_20 <= 1'h0;
      readStageValid_readCounter_20 <= 4'h0;
      readStageValid_segPtr_21 <= 3'h0;
      readStageValid_readCount_21 <= 3'h0;
      readStageValid_stageValid_21 <= 1'h0;
      readStageValid_readCounter_21 <= 4'h0;
      readStageValid_segPtr_22 <= 3'h0;
      readStageValid_readCount_22 <= 3'h0;
      readStageValid_stageValid_22 <= 1'h0;
      readStageValid_readCounter_22 <= 4'h0;
      readStageValid_segPtr_23 <= 3'h0;
      readStageValid_readCount_23 <= 3'h0;
      readStageValid_stageValid_23 <= 1'h0;
      readStageValid_readCounter_23 <= 4'h0;
      readStageValid_segPtr_24 <= 3'h0;
      readStageValid_readCount_24 <= 3'h0;
      readStageValid_stageValid_24 <= 1'h0;
      readStageValid_readCounter_24 <= 4'h0;
      readStageValid_segPtr_25 <= 3'h0;
      readStageValid_readCount_25 <= 3'h0;
      readStageValid_stageValid_25 <= 1'h0;
      readStageValid_readCounter_25 <= 4'h0;
      readStageValid_segPtr_26 <= 3'h0;
      readStageValid_readCount_26 <= 3'h0;
      readStageValid_stageValid_26 <= 1'h0;
      readStageValid_readCounter_26 <= 4'h0;
      readStageValid_segPtr_27 <= 3'h0;
      readStageValid_readCount_27 <= 3'h0;
      readStageValid_stageValid_27 <= 1'h0;
      readStageValid_readCounter_27 <= 4'h0;
      readStageValid_segPtr_28 <= 3'h0;
      readStageValid_readCount_28 <= 3'h0;
      readStageValid_stageValid_28 <= 1'h0;
      readStageValid_readCounter_28 <= 4'h0;
      readStageValid_segPtr_29 <= 3'h0;
      readStageValid_readCount_29 <= 3'h0;
      readStageValid_stageValid_29 <= 1'h0;
      readStageValid_readCounter_29 <= 4'h0;
      readStageValid_segPtr_30 <= 3'h0;
      readStageValid_readCount_30 <= 3'h0;
      readStageValid_stageValid_30 <= 1'h0;
      readStageValid_readCounter_30 <= 4'h0;
      readStageValid_segPtr_31 <= 3'h0;
      readStageValid_readCount_31 <= 3'h0;
      readStageValid_stageValid_31 <= 1'h0;
      readStageValid_readCounter_31 <= 4'h0;
      bufferFull <= 1'h0;
      bufferValid <= 1'h0;
      maskForBufferData_0 <= 128'h0;
      maskForBufferData_1 <= 128'h0;
      maskForBufferData_2 <= 128'h0;
      maskForBufferData_3 <= 128'h0;
      maskForBufferData_4 <= 128'h0;
      maskForBufferData_5 <= 128'h0;
      maskForBufferData_6 <= 128'h0;
      maskForBufferData_7 <= 128'h0;
      lastDataGroupInDataBuffer <= 1'h0;
      cacheLineTemp <= 1024'h0;
      maskTemp <= 128'h0;
      canSendTail <= 1'h0;
      idleNext <= 1'h1;
    end
    else begin
      if (lsuRequest_valid) begin
        lsuRequestReg_instructionInformation_nf <= nfCorrection;
        lsuRequestReg_instructionInformation_mew <= ~invalidInstruction & lsuRequest_bits_instructionInformation_mew;
        lsuRequestReg_instructionInformation_mop <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_mop;
        lsuRequestReg_instructionInformation_lumop <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_lumop;
        lsuRequestReg_instructionInformation_eew <= invalidInstruction ? 2'h0 : lsuRequest_bits_instructionInformation_eew;
        lsuRequestReg_instructionInformation_vs3 <= invalidInstruction ? 5'h0 : lsuRequest_bits_instructionInformation_vs3;
        lsuRequestReg_instructionInformation_isStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_isStore;
        lsuRequestReg_instructionInformation_maskedLoadStore <= ~invalidInstruction & lsuRequest_bits_instructionInformation_maskedLoadStore;
        lsuRequestReg_rs1Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs1Data;
        lsuRequestReg_rs2Data <= invalidInstruction ? 32'h0 : lsuRequest_bits_rs2Data;
        lsuRequestReg_instructionIndex <= lsuRequest_bits_instructionIndex;
        csrInterfaceReg_vl <= csrInterface_vl;
        csrInterfaceReg_vStart <= csrInterface_vStart;
        csrInterfaceReg_vlmul <= csrInterface_vlmul;
        csrInterfaceReg_vSew <= csrInterface_vSew;
        csrInterfaceReg_vxrm <= csrInterface_vxrm;
        csrInterfaceReg_vta <= csrInterface_vta;
        csrInterfaceReg_vma <= csrInterface_vma;
        dataEEW <= lsuRequest_bits_instructionInformation_eew;
        needAmend <= |(csrInterface_vl[6:0]);
        lastMaskAmendReg <= lastMaskAmend;
        segmentInstructionIndexInterval <= csrInterface_vlmul[2] ? 4'h1 : 4'h1 << csrInterface_vlmul[1:0];
        lastWriteVrfIndexReg <= lastWriteVrfIndex;
        lastCacheNeedPush <= lastCacheLineIndex == lastWriteVrfIndex;
        cacheLineNumberReg <= lastCacheLineIndex;
        lastDataGroupReg <= lastDataGroupForInstruction;
      end
      requestFireNext <= lsuRequest_valid;
      if (_maskSelect_valid_output | lsuRequest_valid) begin
        maskReg <= maskAmend;
        isLastMaskGroup <= lsuRequest_valid ? csrInterface_vl[10:7] == 4'h0 : {1'h0, _maskSelect_bits_output} == csrInterfaceReg_vl[10:7];
      end
      if (_GEN_1126 & (_GEN_1127 | lsuRequest_valid))
        maskGroupCounter <= _maskSelect_bits_output;
      if (_GEN_1126) begin
        maskCounterInGroup <= isLastDataGroup | lsuRequest_valid ? 2'h0 : nextMaskCount;
        dataGroup <= nextDataGroup;
      end
      if (accessBufferDequeueFire | accessBufferEnqueueFire | requestFireNext) begin
        accessData_0 <= accessDataUpdate_0;
        accessData_1 <= accessDataUpdate_1;
        accessData_2 <= accessDataUpdate_2;
        accessData_3 <= accessDataUpdate_3;
        accessData_4 <= accessDataUpdate_4;
        accessData_5 <= accessDataUpdate_5;
        accessData_6 <= accessDataUpdate_6;
        accessData_7 <= accessDataUpdate_7;
        accessPtr <= accessBufferDequeueFire | lastPtr | requestFireNext ? lsuRequestReg_instructionInformation_nf - {2'h0, accessBufferEnqueueFire & ~lastPtr} : accessPtr - 3'h1;
      end
      if (accessBufferDequeueFire) begin
        automatic logic [8191:0] _GEN_1131 =
          (dataEEWOH[0]
             ? (_fillBySeg_T[0] ? regroupLoadData_0_0 : 8192'h0) | (_fillBySeg_T[1] ? regroupLoadData_0_1 : 8192'h0) | (_fillBySeg_T[2] ? regroupLoadData_0_2 : 8192'h0) | (_fillBySeg_T[3] ? regroupLoadData_0_3 : 8192'h0)
               | (_fillBySeg_T[4] ? regroupLoadData_0_4 : 8192'h0) | (_fillBySeg_T[5] ? regroupLoadData_0_5 : 8192'h0) | (_fillBySeg_T[6] ? regroupLoadData_0_6 : 8192'h0) | (_fillBySeg_T[7] ? regroupLoadData_0_7 : 8192'h0)
             : 8192'h0)
          | (dataEEWOH[1]
               ? (_fillBySeg_T[0] ? regroupLoadData_1_0 : 8192'h0) | (_fillBySeg_T[1] ? regroupLoadData_1_1 : 8192'h0) | (_fillBySeg_T[2] ? regroupLoadData_1_2 : 8192'h0) | (_fillBySeg_T[3] ? regroupLoadData_1_3 : 8192'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_1_4 : 8192'h0) | (_fillBySeg_T[5] ? regroupLoadData_1_5 : 8192'h0) | (_fillBySeg_T[6] ? regroupLoadData_1_6 : 8192'h0) | (_fillBySeg_T[7] ? regroupLoadData_1_7 : 8192'h0)
               : 8192'h0)
          | (dataEEWOH[2]
               ? (_fillBySeg_T[0] ? regroupLoadData_2_0 : 8192'h0) | (_fillBySeg_T[1] ? regroupLoadData_2_1 : 8192'h0) | (_fillBySeg_T[2] ? regroupLoadData_2_2 : 8192'h0) | (_fillBySeg_T[3] ? regroupLoadData_2_3 : 8192'h0)
                 | (_fillBySeg_T[4] ? regroupLoadData_2_4 : 8192'h0) | (_fillBySeg_T[5] ? regroupLoadData_2_5 : 8192'h0) | (_fillBySeg_T[6] ? regroupLoadData_2_6 : 8192'h0) | (_fillBySeg_T[7] ? regroupLoadData_2_7 : 8192'h0)
               : 8192'h0);
        dataBuffer_0 <= _GEN_1131[1023:0];
        dataBuffer_1 <= _GEN_1131[2047:1024];
        dataBuffer_2 <= _GEN_1131[3071:2048];
        dataBuffer_3 <= _GEN_1131[4095:3072];
        dataBuffer_4 <= _GEN_1131[5119:4096];
        dataBuffer_5 <= _GEN_1131[6143:5120];
        dataBuffer_6 <= _GEN_1131[7167:6144];
        dataBuffer_7 <= _GEN_1131[8191:7168];
        maskForBufferData_0 <= fillBySeg[127:0];
        maskForBufferData_1 <= fillBySeg[255:128];
        maskForBufferData_2 <= fillBySeg[383:256];
        maskForBufferData_3 <= fillBySeg[511:384];
        maskForBufferData_4 <= fillBySeg[639:512];
        maskForBufferData_5 <= fillBySeg[767:640];
        maskForBufferData_6 <= fillBySeg[895:768];
        maskForBufferData_7 <= fillBySeg[1023:896];
        lastDataGroupInDataBuffer <= isLastRead;
      end
      else if (alignedDequeueFire) begin
        dataBuffer_0 <= dataBuffer_1;
        dataBuffer_1 <= dataBuffer_2;
        dataBuffer_2 <= dataBuffer_3;
        dataBuffer_3 <= dataBuffer_4;
        dataBuffer_4 <= dataBuffer_5;
        dataBuffer_5 <= dataBuffer_6;
        dataBuffer_6 <= dataBuffer_7;
        dataBuffer_7 <= 1024'h0;
      end
      if (lsuRequest_valid | alignedDequeueFire) begin
        bufferBaseCacheLineIndex <= lsuRequest_valid ? 4'h0 : bufferBaseCacheLineIndex + 4'h1;
        maskTemp <= lsuRequest_valid ? 128'h0 : _GEN_1129;
        canSendTail <= ~lsuRequest_valid & bufferValid & isLastCacheLineInBuffer & lastDataGroupInDataBuffer;
      end
      if (accessBufferDequeueFire | alignedDequeueFire)
        cacheLineIndexInBuffer <= accessBufferDequeueFire ? 3'h0 : cacheLineIndexInBuffer + 3'h1;
      hazardCheck <= ~lsuRequest_valid;
      if (lsuRequest_valid | _readStageValid_T_11)
        readStageValid_segPtr <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_11 & readStageValid_lastReadPtr)
        readStageValid_readCount <= readStageValid_nextReadCount;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup & readStageValid_lastReadPtr & _readStageValid_T_11)
        readStageValid_stageValid <= lsuRequest_valid;
      if (_readStageValid_T_11 ^ vrfReadQueueVec_0_deq_ready & vrfReadQueueVec_0_deq_valid)
        readStageValid_readCounter <= readStageValid_readCounter + readStageValid_counterChange;
      if (lsuRequest_valid | _readStageValid_T_30)
        readStageValid_segPtr_1 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_1 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_1 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_30 & readStageValid_lastReadPtr_1)
        readStageValid_readCount_1 <= readStageValid_nextReadCount_1;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_1 & readStageValid_lastReadPtr_1 & _readStageValid_T_30)
        readStageValid_stageValid_1 <= lsuRequest_valid;
      if (_readStageValid_T_30 ^ vrfReadQueueVec_1_deq_ready & vrfReadQueueVec_1_deq_valid)
        readStageValid_readCounter_1 <= readStageValid_readCounter_1 + readStageValid_counterChange_1;
      if (lsuRequest_valid | _readStageValid_T_49)
        readStageValid_segPtr_2 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_2 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_2 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_49 & readStageValid_lastReadPtr_2)
        readStageValid_readCount_2 <= readStageValid_nextReadCount_2;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_2 & readStageValid_lastReadPtr_2 & _readStageValid_T_49)
        readStageValid_stageValid_2 <= lsuRequest_valid;
      if (_readStageValid_T_49 ^ vrfReadQueueVec_2_deq_ready & vrfReadQueueVec_2_deq_valid)
        readStageValid_readCounter_2 <= readStageValid_readCounter_2 + readStageValid_counterChange_2;
      if (lsuRequest_valid | _readStageValid_T_68)
        readStageValid_segPtr_3 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_3 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_3 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_68 & readStageValid_lastReadPtr_3)
        readStageValid_readCount_3 <= readStageValid_nextReadCount_3;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_3 & readStageValid_lastReadPtr_3 & _readStageValid_T_68)
        readStageValid_stageValid_3 <= lsuRequest_valid;
      if (_readStageValid_T_68 ^ vrfReadQueueVec_3_deq_ready & vrfReadQueueVec_3_deq_valid)
        readStageValid_readCounter_3 <= readStageValid_readCounter_3 + readStageValid_counterChange_3;
      if (lsuRequest_valid | _readStageValid_T_87)
        readStageValid_segPtr_4 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_4 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_4 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_87 & readStageValid_lastReadPtr_4)
        readStageValid_readCount_4 <= readStageValid_nextReadCount_4;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_4 & readStageValid_lastReadPtr_4 & _readStageValid_T_87)
        readStageValid_stageValid_4 <= lsuRequest_valid;
      if (_readStageValid_T_87 ^ vrfReadQueueVec_4_deq_ready & vrfReadQueueVec_4_deq_valid)
        readStageValid_readCounter_4 <= readStageValid_readCounter_4 + readStageValid_counterChange_4;
      if (lsuRequest_valid | _readStageValid_T_106)
        readStageValid_segPtr_5 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_5 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_5 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_106 & readStageValid_lastReadPtr_5)
        readStageValid_readCount_5 <= readStageValid_nextReadCount_5;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_5 & readStageValid_lastReadPtr_5 & _readStageValid_T_106)
        readStageValid_stageValid_5 <= lsuRequest_valid;
      if (_readStageValid_T_106 ^ vrfReadQueueVec_5_deq_ready & vrfReadQueueVec_5_deq_valid)
        readStageValid_readCounter_5 <= readStageValid_readCounter_5 + readStageValid_counterChange_5;
      if (lsuRequest_valid | _readStageValid_T_125)
        readStageValid_segPtr_6 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_6 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_6 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_125 & readStageValid_lastReadPtr_6)
        readStageValid_readCount_6 <= readStageValid_nextReadCount_6;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_6 & readStageValid_lastReadPtr_6 & _readStageValid_T_125)
        readStageValid_stageValid_6 <= lsuRequest_valid;
      if (_readStageValid_T_125 ^ vrfReadQueueVec_6_deq_ready & vrfReadQueueVec_6_deq_valid)
        readStageValid_readCounter_6 <= readStageValid_readCounter_6 + readStageValid_counterChange_6;
      if (lsuRequest_valid | _readStageValid_T_144)
        readStageValid_segPtr_7 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_7 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_7 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_144 & readStageValid_lastReadPtr_7)
        readStageValid_readCount_7 <= readStageValid_nextReadCount_7;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_7 & readStageValid_lastReadPtr_7 & _readStageValid_T_144)
        readStageValid_stageValid_7 <= lsuRequest_valid;
      if (_readStageValid_T_144 ^ vrfReadQueueVec_7_deq_ready & vrfReadQueueVec_7_deq_valid)
        readStageValid_readCounter_7 <= readStageValid_readCounter_7 + readStageValid_counterChange_7;
      if (lsuRequest_valid | _readStageValid_T_163)
        readStageValid_segPtr_8 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_8 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_8 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_163 & readStageValid_lastReadPtr_8)
        readStageValid_readCount_8 <= readStageValid_nextReadCount_8;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_8 & readStageValid_lastReadPtr_8 & _readStageValid_T_163)
        readStageValid_stageValid_8 <= lsuRequest_valid;
      if (_readStageValid_T_163 ^ vrfReadQueueVec_8_deq_ready & vrfReadQueueVec_8_deq_valid)
        readStageValid_readCounter_8 <= readStageValid_readCounter_8 + readStageValid_counterChange_8;
      if (lsuRequest_valid | _readStageValid_T_182)
        readStageValid_segPtr_9 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_9 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_9 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_182 & readStageValid_lastReadPtr_9)
        readStageValid_readCount_9 <= readStageValid_nextReadCount_9;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_9 & readStageValid_lastReadPtr_9 & _readStageValid_T_182)
        readStageValid_stageValid_9 <= lsuRequest_valid;
      if (_readStageValid_T_182 ^ vrfReadQueueVec_9_deq_ready & vrfReadQueueVec_9_deq_valid)
        readStageValid_readCounter_9 <= readStageValid_readCounter_9 + readStageValid_counterChange_9;
      if (lsuRequest_valid | _readStageValid_T_201)
        readStageValid_segPtr_10 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_10 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_10 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_201 & readStageValid_lastReadPtr_10)
        readStageValid_readCount_10 <= readStageValid_nextReadCount_10;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_10 & readStageValid_lastReadPtr_10 & _readStageValid_T_201)
        readStageValid_stageValid_10 <= lsuRequest_valid;
      if (_readStageValid_T_201 ^ vrfReadQueueVec_10_deq_ready & vrfReadQueueVec_10_deq_valid)
        readStageValid_readCounter_10 <= readStageValid_readCounter_10 + readStageValid_counterChange_10;
      if (lsuRequest_valid | _readStageValid_T_220)
        readStageValid_segPtr_11 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_11 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_11 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_220 & readStageValid_lastReadPtr_11)
        readStageValid_readCount_11 <= readStageValid_nextReadCount_11;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_11 & readStageValid_lastReadPtr_11 & _readStageValid_T_220)
        readStageValid_stageValid_11 <= lsuRequest_valid;
      if (_readStageValid_T_220 ^ vrfReadQueueVec_11_deq_ready & vrfReadQueueVec_11_deq_valid)
        readStageValid_readCounter_11 <= readStageValid_readCounter_11 + readStageValid_counterChange_11;
      if (lsuRequest_valid | _readStageValid_T_239)
        readStageValid_segPtr_12 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_12 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_12 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_239 & readStageValid_lastReadPtr_12)
        readStageValid_readCount_12 <= readStageValid_nextReadCount_12;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_12 & readStageValid_lastReadPtr_12 & _readStageValid_T_239)
        readStageValid_stageValid_12 <= lsuRequest_valid;
      if (_readStageValid_T_239 ^ vrfReadQueueVec_12_deq_ready & vrfReadQueueVec_12_deq_valid)
        readStageValid_readCounter_12 <= readStageValid_readCounter_12 + readStageValid_counterChange_12;
      if (lsuRequest_valid | _readStageValid_T_258)
        readStageValid_segPtr_13 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_13 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_13 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_258 & readStageValid_lastReadPtr_13)
        readStageValid_readCount_13 <= readStageValid_nextReadCount_13;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_13 & readStageValid_lastReadPtr_13 & _readStageValid_T_258)
        readStageValid_stageValid_13 <= lsuRequest_valid;
      if (_readStageValid_T_258 ^ vrfReadQueueVec_13_deq_ready & vrfReadQueueVec_13_deq_valid)
        readStageValid_readCounter_13 <= readStageValid_readCounter_13 + readStageValid_counterChange_13;
      if (lsuRequest_valid | _readStageValid_T_277)
        readStageValid_segPtr_14 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_14 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_14 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_277 & readStageValid_lastReadPtr_14)
        readStageValid_readCount_14 <= readStageValid_nextReadCount_14;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_14 & readStageValid_lastReadPtr_14 & _readStageValid_T_277)
        readStageValid_stageValid_14 <= lsuRequest_valid;
      if (_readStageValid_T_277 ^ vrfReadQueueVec_14_deq_ready & vrfReadQueueVec_14_deq_valid)
        readStageValid_readCounter_14 <= readStageValid_readCounter_14 + readStageValid_counterChange_14;
      if (lsuRequest_valid | _readStageValid_T_296)
        readStageValid_segPtr_15 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_15 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_15 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_296 & readStageValid_lastReadPtr_15)
        readStageValid_readCount_15 <= readStageValid_nextReadCount_15;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_15 & readStageValid_lastReadPtr_15 & _readStageValid_T_296)
        readStageValid_stageValid_15 <= lsuRequest_valid;
      if (_readStageValid_T_296 ^ vrfReadQueueVec_15_deq_ready & vrfReadQueueVec_15_deq_valid)
        readStageValid_readCounter_15 <= readStageValid_readCounter_15 + readStageValid_counterChange_15;
      if (lsuRequest_valid | _readStageValid_T_315)
        readStageValid_segPtr_16 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_16 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_16 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_315 & readStageValid_lastReadPtr_16)
        readStageValid_readCount_16 <= readStageValid_nextReadCount_16;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_16 & readStageValid_lastReadPtr_16 & _readStageValid_T_315)
        readStageValid_stageValid_16 <= lsuRequest_valid;
      if (_readStageValid_T_315 ^ vrfReadQueueVec_16_deq_ready & vrfReadQueueVec_16_deq_valid)
        readStageValid_readCounter_16 <= readStageValid_readCounter_16 + readStageValid_counterChange_16;
      if (lsuRequest_valid | _readStageValid_T_334)
        readStageValid_segPtr_17 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_17 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_17 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_334 & readStageValid_lastReadPtr_17)
        readStageValid_readCount_17 <= readStageValid_nextReadCount_17;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_17 & readStageValid_lastReadPtr_17 & _readStageValid_T_334)
        readStageValid_stageValid_17 <= lsuRequest_valid;
      if (_readStageValid_T_334 ^ vrfReadQueueVec_17_deq_ready & vrfReadQueueVec_17_deq_valid)
        readStageValid_readCounter_17 <= readStageValid_readCounter_17 + readStageValid_counterChange_17;
      if (lsuRequest_valid | _readStageValid_T_353)
        readStageValid_segPtr_18 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_18 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_18 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_353 & readStageValid_lastReadPtr_18)
        readStageValid_readCount_18 <= readStageValid_nextReadCount_18;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_18 & readStageValid_lastReadPtr_18 & _readStageValid_T_353)
        readStageValid_stageValid_18 <= lsuRequest_valid;
      if (_readStageValid_T_353 ^ vrfReadQueueVec_18_deq_ready & vrfReadQueueVec_18_deq_valid)
        readStageValid_readCounter_18 <= readStageValid_readCounter_18 + readStageValid_counterChange_18;
      if (lsuRequest_valid | _readStageValid_T_372)
        readStageValid_segPtr_19 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_19 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_19 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_372 & readStageValid_lastReadPtr_19)
        readStageValid_readCount_19 <= readStageValid_nextReadCount_19;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_19 & readStageValid_lastReadPtr_19 & _readStageValid_T_372)
        readStageValid_stageValid_19 <= lsuRequest_valid;
      if (_readStageValid_T_372 ^ vrfReadQueueVec_19_deq_ready & vrfReadQueueVec_19_deq_valid)
        readStageValid_readCounter_19 <= readStageValid_readCounter_19 + readStageValid_counterChange_19;
      if (lsuRequest_valid | _readStageValid_T_391)
        readStageValid_segPtr_20 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_20 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_20 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_391 & readStageValid_lastReadPtr_20)
        readStageValid_readCount_20 <= readStageValid_nextReadCount_20;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_20 & readStageValid_lastReadPtr_20 & _readStageValid_T_391)
        readStageValid_stageValid_20 <= lsuRequest_valid;
      if (_readStageValid_T_391 ^ vrfReadQueueVec_20_deq_ready & vrfReadQueueVec_20_deq_valid)
        readStageValid_readCounter_20 <= readStageValid_readCounter_20 + readStageValid_counterChange_20;
      if (lsuRequest_valid | _readStageValid_T_410)
        readStageValid_segPtr_21 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_21 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_21 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_410 & readStageValid_lastReadPtr_21)
        readStageValid_readCount_21 <= readStageValid_nextReadCount_21;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_21 & readStageValid_lastReadPtr_21 & _readStageValid_T_410)
        readStageValid_stageValid_21 <= lsuRequest_valid;
      if (_readStageValid_T_410 ^ vrfReadQueueVec_21_deq_ready & vrfReadQueueVec_21_deq_valid)
        readStageValid_readCounter_21 <= readStageValid_readCounter_21 + readStageValid_counterChange_21;
      if (lsuRequest_valid | _readStageValid_T_429)
        readStageValid_segPtr_22 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_22 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_22 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_429 & readStageValid_lastReadPtr_22)
        readStageValid_readCount_22 <= readStageValid_nextReadCount_22;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_22 & readStageValid_lastReadPtr_22 & _readStageValid_T_429)
        readStageValid_stageValid_22 <= lsuRequest_valid;
      if (_readStageValid_T_429 ^ vrfReadQueueVec_22_deq_ready & vrfReadQueueVec_22_deq_valid)
        readStageValid_readCounter_22 <= readStageValid_readCounter_22 + readStageValid_counterChange_22;
      if (lsuRequest_valid | _readStageValid_T_448)
        readStageValid_segPtr_23 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_23 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_23 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_448 & readStageValid_lastReadPtr_23)
        readStageValid_readCount_23 <= readStageValid_nextReadCount_23;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_23 & readStageValid_lastReadPtr_23 & _readStageValid_T_448)
        readStageValid_stageValid_23 <= lsuRequest_valid;
      if (_readStageValid_T_448 ^ vrfReadQueueVec_23_deq_ready & vrfReadQueueVec_23_deq_valid)
        readStageValid_readCounter_23 <= readStageValid_readCounter_23 + readStageValid_counterChange_23;
      if (lsuRequest_valid | _readStageValid_T_467)
        readStageValid_segPtr_24 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_24 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_24 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_467 & readStageValid_lastReadPtr_24)
        readStageValid_readCount_24 <= readStageValid_nextReadCount_24;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_24 & readStageValid_lastReadPtr_24 & _readStageValid_T_467)
        readStageValid_stageValid_24 <= lsuRequest_valid;
      if (_readStageValid_T_467 ^ vrfReadQueueVec_24_deq_ready & vrfReadQueueVec_24_deq_valid)
        readStageValid_readCounter_24 <= readStageValid_readCounter_24 + readStageValid_counterChange_24;
      if (lsuRequest_valid | _readStageValid_T_486)
        readStageValid_segPtr_25 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_25 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_25 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_486 & readStageValid_lastReadPtr_25)
        readStageValid_readCount_25 <= readStageValid_nextReadCount_25;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_25 & readStageValid_lastReadPtr_25 & _readStageValid_T_486)
        readStageValid_stageValid_25 <= lsuRequest_valid;
      if (_readStageValid_T_486 ^ vrfReadQueueVec_25_deq_ready & vrfReadQueueVec_25_deq_valid)
        readStageValid_readCounter_25 <= readStageValid_readCounter_25 + readStageValid_counterChange_25;
      if (lsuRequest_valid | _readStageValid_T_505)
        readStageValid_segPtr_26 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_26 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_26 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_505 & readStageValid_lastReadPtr_26)
        readStageValid_readCount_26 <= readStageValid_nextReadCount_26;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_26 & readStageValid_lastReadPtr_26 & _readStageValid_T_505)
        readStageValid_stageValid_26 <= lsuRequest_valid;
      if (_readStageValid_T_505 ^ vrfReadQueueVec_26_deq_ready & vrfReadQueueVec_26_deq_valid)
        readStageValid_readCounter_26 <= readStageValid_readCounter_26 + readStageValid_counterChange_26;
      if (lsuRequest_valid | _readStageValid_T_524)
        readStageValid_segPtr_27 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_27 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_27 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_524 & readStageValid_lastReadPtr_27)
        readStageValid_readCount_27 <= readStageValid_nextReadCount_27;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_27 & readStageValid_lastReadPtr_27 & _readStageValid_T_524)
        readStageValid_stageValid_27 <= lsuRequest_valid;
      if (_readStageValid_T_524 ^ vrfReadQueueVec_27_deq_ready & vrfReadQueueVec_27_deq_valid)
        readStageValid_readCounter_27 <= readStageValid_readCounter_27 + readStageValid_counterChange_27;
      if (lsuRequest_valid | _readStageValid_T_543)
        readStageValid_segPtr_28 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_28 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_28 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_543 & readStageValid_lastReadPtr_28)
        readStageValid_readCount_28 <= readStageValid_nextReadCount_28;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_28 & readStageValid_lastReadPtr_28 & _readStageValid_T_543)
        readStageValid_stageValid_28 <= lsuRequest_valid;
      if (_readStageValid_T_543 ^ vrfReadQueueVec_28_deq_ready & vrfReadQueueVec_28_deq_valid)
        readStageValid_readCounter_28 <= readStageValid_readCounter_28 + readStageValid_counterChange_28;
      if (lsuRequest_valid | _readStageValid_T_562)
        readStageValid_segPtr_29 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_29 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_29 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_562 & readStageValid_lastReadPtr_29)
        readStageValid_readCount_29 <= readStageValid_nextReadCount_29;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_29 & readStageValid_lastReadPtr_29 & _readStageValid_T_562)
        readStageValid_stageValid_29 <= lsuRequest_valid;
      if (_readStageValid_T_562 ^ vrfReadQueueVec_29_deq_ready & vrfReadQueueVec_29_deq_valid)
        readStageValid_readCounter_29 <= readStageValid_readCounter_29 + readStageValid_counterChange_29;
      if (lsuRequest_valid | _readStageValid_T_581)
        readStageValid_segPtr_30 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_30 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_30 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_581 & readStageValid_lastReadPtr_30)
        readStageValid_readCount_30 <= readStageValid_nextReadCount_30;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_30 & readStageValid_lastReadPtr_30 & _readStageValid_T_581)
        readStageValid_stageValid_30 <= lsuRequest_valid;
      if (_readStageValid_T_581 ^ vrfReadQueueVec_30_deq_ready & vrfReadQueueVec_30_deq_valid)
        readStageValid_readCounter_30 <= readStageValid_readCounter_30 + readStageValid_counterChange_30;
      if (lsuRequest_valid | _readStageValid_T_600)
        readStageValid_segPtr_31 <= lsuRequest_valid ? nfCorrection : readStageValid_lastReadPtr_31 ? lsuRequestReg_instructionInformation_nf : readStageValid_segPtr_31 - 3'h1;
      if (lsuRequest_valid | _readStageValid_T_600 & readStageValid_lastReadPtr_31)
        readStageValid_readCount_31 <= readStageValid_nextReadCount_31;
      if (lsuRequest_valid & ~invalidInstruction | readStageValid_lastReadGroup_31 & readStageValid_lastReadPtr_31 & _readStageValid_T_600)
        readStageValid_stageValid_31 <= lsuRequest_valid;
      if (_readStageValid_T_600 ^ vrfReadQueueVec_31_deq_ready & vrfReadQueueVec_31_deq_valid)
        readStageValid_readCounter_31 <= readStageValid_readCounter_31 + readStageValid_counterChange_31;
      if (lastPtrEnq ^ accessBufferDequeueFire)
        bufferFull <= lastPtrEnq;
      if (accessBufferDequeueFire ^ bufferWillClear)
        bufferValid <= accessBufferDequeueFire;
      if (alignedDequeueFire)
        cacheLineTemp <= dataBuffer_0;
      idleNext <= _status_idle_output;
    end
    invalidInstructionNext <= invalidInstruction & lsuRequest_valid;
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:609];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [9:0] i = 10'h0; i < 10'h262; i += 10'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        lsuRequestReg_instructionInformation_nf = _RANDOM[10'h0][2:0];
        lsuRequestReg_instructionInformation_mew = _RANDOM[10'h0][3];
        lsuRequestReg_instructionInformation_mop = _RANDOM[10'h0][5:4];
        lsuRequestReg_instructionInformation_lumop = _RANDOM[10'h0][10:6];
        lsuRequestReg_instructionInformation_eew = _RANDOM[10'h0][12:11];
        lsuRequestReg_instructionInformation_vs3 = _RANDOM[10'h0][17:13];
        lsuRequestReg_instructionInformation_isStore = _RANDOM[10'h0][18];
        lsuRequestReg_instructionInformation_maskedLoadStore = _RANDOM[10'h0][19];
        lsuRequestReg_rs1Data = {_RANDOM[10'h0][31:20], _RANDOM[10'h1][19:0]};
        lsuRequestReg_rs2Data = {_RANDOM[10'h1][31:20], _RANDOM[10'h2][19:0]};
        lsuRequestReg_instructionIndex = _RANDOM[10'h2][22:20];
        csrInterfaceReg_vl = {_RANDOM[10'h2][31:23], _RANDOM[10'h3][1:0]};
        csrInterfaceReg_vStart = _RANDOM[10'h3][12:2];
        csrInterfaceReg_vlmul = _RANDOM[10'h3][15:13];
        csrInterfaceReg_vSew = _RANDOM[10'h3][17:16];
        csrInterfaceReg_vxrm = _RANDOM[10'h3][19:18];
        csrInterfaceReg_vta = _RANDOM[10'h3][20];
        csrInterfaceReg_vma = _RANDOM[10'h3][21];
        requestFireNext = _RANDOM[10'h3][22];
        dataEEW = _RANDOM[10'h3][24:23];
        maskReg = {_RANDOM[10'h3][31:25], _RANDOM[10'h4], _RANDOM[10'h5], _RANDOM[10'h6], _RANDOM[10'h7][24:0]};
        needAmend = _RANDOM[10'h7][25];
        lastMaskAmendReg = {_RANDOM[10'h7][31:26], _RANDOM[10'h8], _RANDOM[10'h9], _RANDOM[10'hA], _RANDOM[10'hB][24:0]};
        maskGroupCounter = _RANDOM[10'hB][27:25];
        maskCounterInGroup = _RANDOM[10'hB][29:28];
        isLastMaskGroup = _RANDOM[10'hF][30];
        accessData_0 =
          {_RANDOM[10'hF][31],
           _RANDOM[10'h10],
           _RANDOM[10'h11],
           _RANDOM[10'h12],
           _RANDOM[10'h13],
           _RANDOM[10'h14],
           _RANDOM[10'h15],
           _RANDOM[10'h16],
           _RANDOM[10'h17],
           _RANDOM[10'h18],
           _RANDOM[10'h19],
           _RANDOM[10'h1A],
           _RANDOM[10'h1B],
           _RANDOM[10'h1C],
           _RANDOM[10'h1D],
           _RANDOM[10'h1E],
           _RANDOM[10'h1F],
           _RANDOM[10'h20],
           _RANDOM[10'h21],
           _RANDOM[10'h22],
           _RANDOM[10'h23],
           _RANDOM[10'h24],
           _RANDOM[10'h25],
           _RANDOM[10'h26],
           _RANDOM[10'h27],
           _RANDOM[10'h28],
           _RANDOM[10'h29],
           _RANDOM[10'h2A],
           _RANDOM[10'h2B],
           _RANDOM[10'h2C],
           _RANDOM[10'h2D],
           _RANDOM[10'h2E],
           _RANDOM[10'h2F][30:0]};
        accessData_1 =
          {_RANDOM[10'h2F][31],
           _RANDOM[10'h30],
           _RANDOM[10'h31],
           _RANDOM[10'h32],
           _RANDOM[10'h33],
           _RANDOM[10'h34],
           _RANDOM[10'h35],
           _RANDOM[10'h36],
           _RANDOM[10'h37],
           _RANDOM[10'h38],
           _RANDOM[10'h39],
           _RANDOM[10'h3A],
           _RANDOM[10'h3B],
           _RANDOM[10'h3C],
           _RANDOM[10'h3D],
           _RANDOM[10'h3E],
           _RANDOM[10'h3F],
           _RANDOM[10'h40],
           _RANDOM[10'h41],
           _RANDOM[10'h42],
           _RANDOM[10'h43],
           _RANDOM[10'h44],
           _RANDOM[10'h45],
           _RANDOM[10'h46],
           _RANDOM[10'h47],
           _RANDOM[10'h48],
           _RANDOM[10'h49],
           _RANDOM[10'h4A],
           _RANDOM[10'h4B],
           _RANDOM[10'h4C],
           _RANDOM[10'h4D],
           _RANDOM[10'h4E],
           _RANDOM[10'h4F][30:0]};
        accessData_2 =
          {_RANDOM[10'h4F][31],
           _RANDOM[10'h50],
           _RANDOM[10'h51],
           _RANDOM[10'h52],
           _RANDOM[10'h53],
           _RANDOM[10'h54],
           _RANDOM[10'h55],
           _RANDOM[10'h56],
           _RANDOM[10'h57],
           _RANDOM[10'h58],
           _RANDOM[10'h59],
           _RANDOM[10'h5A],
           _RANDOM[10'h5B],
           _RANDOM[10'h5C],
           _RANDOM[10'h5D],
           _RANDOM[10'h5E],
           _RANDOM[10'h5F],
           _RANDOM[10'h60],
           _RANDOM[10'h61],
           _RANDOM[10'h62],
           _RANDOM[10'h63],
           _RANDOM[10'h64],
           _RANDOM[10'h65],
           _RANDOM[10'h66],
           _RANDOM[10'h67],
           _RANDOM[10'h68],
           _RANDOM[10'h69],
           _RANDOM[10'h6A],
           _RANDOM[10'h6B],
           _RANDOM[10'h6C],
           _RANDOM[10'h6D],
           _RANDOM[10'h6E],
           _RANDOM[10'h6F][30:0]};
        accessData_3 =
          {_RANDOM[10'h6F][31],
           _RANDOM[10'h70],
           _RANDOM[10'h71],
           _RANDOM[10'h72],
           _RANDOM[10'h73],
           _RANDOM[10'h74],
           _RANDOM[10'h75],
           _RANDOM[10'h76],
           _RANDOM[10'h77],
           _RANDOM[10'h78],
           _RANDOM[10'h79],
           _RANDOM[10'h7A],
           _RANDOM[10'h7B],
           _RANDOM[10'h7C],
           _RANDOM[10'h7D],
           _RANDOM[10'h7E],
           _RANDOM[10'h7F],
           _RANDOM[10'h80],
           _RANDOM[10'h81],
           _RANDOM[10'h82],
           _RANDOM[10'h83],
           _RANDOM[10'h84],
           _RANDOM[10'h85],
           _RANDOM[10'h86],
           _RANDOM[10'h87],
           _RANDOM[10'h88],
           _RANDOM[10'h89],
           _RANDOM[10'h8A],
           _RANDOM[10'h8B],
           _RANDOM[10'h8C],
           _RANDOM[10'h8D],
           _RANDOM[10'h8E],
           _RANDOM[10'h8F][30:0]};
        accessData_4 =
          {_RANDOM[10'h8F][31],
           _RANDOM[10'h90],
           _RANDOM[10'h91],
           _RANDOM[10'h92],
           _RANDOM[10'h93],
           _RANDOM[10'h94],
           _RANDOM[10'h95],
           _RANDOM[10'h96],
           _RANDOM[10'h97],
           _RANDOM[10'h98],
           _RANDOM[10'h99],
           _RANDOM[10'h9A],
           _RANDOM[10'h9B],
           _RANDOM[10'h9C],
           _RANDOM[10'h9D],
           _RANDOM[10'h9E],
           _RANDOM[10'h9F],
           _RANDOM[10'hA0],
           _RANDOM[10'hA1],
           _RANDOM[10'hA2],
           _RANDOM[10'hA3],
           _RANDOM[10'hA4],
           _RANDOM[10'hA5],
           _RANDOM[10'hA6],
           _RANDOM[10'hA7],
           _RANDOM[10'hA8],
           _RANDOM[10'hA9],
           _RANDOM[10'hAA],
           _RANDOM[10'hAB],
           _RANDOM[10'hAC],
           _RANDOM[10'hAD],
           _RANDOM[10'hAE],
           _RANDOM[10'hAF][30:0]};
        accessData_5 =
          {_RANDOM[10'hAF][31],
           _RANDOM[10'hB0],
           _RANDOM[10'hB1],
           _RANDOM[10'hB2],
           _RANDOM[10'hB3],
           _RANDOM[10'hB4],
           _RANDOM[10'hB5],
           _RANDOM[10'hB6],
           _RANDOM[10'hB7],
           _RANDOM[10'hB8],
           _RANDOM[10'hB9],
           _RANDOM[10'hBA],
           _RANDOM[10'hBB],
           _RANDOM[10'hBC],
           _RANDOM[10'hBD],
           _RANDOM[10'hBE],
           _RANDOM[10'hBF],
           _RANDOM[10'hC0],
           _RANDOM[10'hC1],
           _RANDOM[10'hC2],
           _RANDOM[10'hC3],
           _RANDOM[10'hC4],
           _RANDOM[10'hC5],
           _RANDOM[10'hC6],
           _RANDOM[10'hC7],
           _RANDOM[10'hC8],
           _RANDOM[10'hC9],
           _RANDOM[10'hCA],
           _RANDOM[10'hCB],
           _RANDOM[10'hCC],
           _RANDOM[10'hCD],
           _RANDOM[10'hCE],
           _RANDOM[10'hCF][30:0]};
        accessData_6 =
          {_RANDOM[10'hCF][31],
           _RANDOM[10'hD0],
           _RANDOM[10'hD1],
           _RANDOM[10'hD2],
           _RANDOM[10'hD3],
           _RANDOM[10'hD4],
           _RANDOM[10'hD5],
           _RANDOM[10'hD6],
           _RANDOM[10'hD7],
           _RANDOM[10'hD8],
           _RANDOM[10'hD9],
           _RANDOM[10'hDA],
           _RANDOM[10'hDB],
           _RANDOM[10'hDC],
           _RANDOM[10'hDD],
           _RANDOM[10'hDE],
           _RANDOM[10'hDF],
           _RANDOM[10'hE0],
           _RANDOM[10'hE1],
           _RANDOM[10'hE2],
           _RANDOM[10'hE3],
           _RANDOM[10'hE4],
           _RANDOM[10'hE5],
           _RANDOM[10'hE6],
           _RANDOM[10'hE7],
           _RANDOM[10'hE8],
           _RANDOM[10'hE9],
           _RANDOM[10'hEA],
           _RANDOM[10'hEB],
           _RANDOM[10'hEC],
           _RANDOM[10'hED],
           _RANDOM[10'hEE],
           _RANDOM[10'hEF][30:0]};
        accessData_7 =
          {_RANDOM[10'hEF][31],
           _RANDOM[10'hF0],
           _RANDOM[10'hF1],
           _RANDOM[10'hF2],
           _RANDOM[10'hF3],
           _RANDOM[10'hF4],
           _RANDOM[10'hF5],
           _RANDOM[10'hF6],
           _RANDOM[10'hF7],
           _RANDOM[10'hF8],
           _RANDOM[10'hF9],
           _RANDOM[10'hFA],
           _RANDOM[10'hFB],
           _RANDOM[10'hFC],
           _RANDOM[10'hFD],
           _RANDOM[10'hFE],
           _RANDOM[10'hFF],
           _RANDOM[10'h100],
           _RANDOM[10'h101],
           _RANDOM[10'h102],
           _RANDOM[10'h103],
           _RANDOM[10'h104],
           _RANDOM[10'h105],
           _RANDOM[10'h106],
           _RANDOM[10'h107],
           _RANDOM[10'h108],
           _RANDOM[10'h109],
           _RANDOM[10'h10A],
           _RANDOM[10'h10B],
           _RANDOM[10'h10C],
           _RANDOM[10'h10D],
           _RANDOM[10'h10E],
           _RANDOM[10'h10F][30:0]};
        accessPtr = {_RANDOM[10'h10F][31], _RANDOM[10'h110][1:0]};
        dataGroup = _RANDOM[10'h111][4:2];
        dataBuffer_0 =
          {_RANDOM[10'h111][31:5],
           _RANDOM[10'h112],
           _RANDOM[10'h113],
           _RANDOM[10'h114],
           _RANDOM[10'h115],
           _RANDOM[10'h116],
           _RANDOM[10'h117],
           _RANDOM[10'h118],
           _RANDOM[10'h119],
           _RANDOM[10'h11A],
           _RANDOM[10'h11B],
           _RANDOM[10'h11C],
           _RANDOM[10'h11D],
           _RANDOM[10'h11E],
           _RANDOM[10'h11F],
           _RANDOM[10'h120],
           _RANDOM[10'h121],
           _RANDOM[10'h122],
           _RANDOM[10'h123],
           _RANDOM[10'h124],
           _RANDOM[10'h125],
           _RANDOM[10'h126],
           _RANDOM[10'h127],
           _RANDOM[10'h128],
           _RANDOM[10'h129],
           _RANDOM[10'h12A],
           _RANDOM[10'h12B],
           _RANDOM[10'h12C],
           _RANDOM[10'h12D],
           _RANDOM[10'h12E],
           _RANDOM[10'h12F],
           _RANDOM[10'h130],
           _RANDOM[10'h131][4:0]};
        dataBuffer_1 =
          {_RANDOM[10'h131][31:5],
           _RANDOM[10'h132],
           _RANDOM[10'h133],
           _RANDOM[10'h134],
           _RANDOM[10'h135],
           _RANDOM[10'h136],
           _RANDOM[10'h137],
           _RANDOM[10'h138],
           _RANDOM[10'h139],
           _RANDOM[10'h13A],
           _RANDOM[10'h13B],
           _RANDOM[10'h13C],
           _RANDOM[10'h13D],
           _RANDOM[10'h13E],
           _RANDOM[10'h13F],
           _RANDOM[10'h140],
           _RANDOM[10'h141],
           _RANDOM[10'h142],
           _RANDOM[10'h143],
           _RANDOM[10'h144],
           _RANDOM[10'h145],
           _RANDOM[10'h146],
           _RANDOM[10'h147],
           _RANDOM[10'h148],
           _RANDOM[10'h149],
           _RANDOM[10'h14A],
           _RANDOM[10'h14B],
           _RANDOM[10'h14C],
           _RANDOM[10'h14D],
           _RANDOM[10'h14E],
           _RANDOM[10'h14F],
           _RANDOM[10'h150],
           _RANDOM[10'h151][4:0]};
        dataBuffer_2 =
          {_RANDOM[10'h151][31:5],
           _RANDOM[10'h152],
           _RANDOM[10'h153],
           _RANDOM[10'h154],
           _RANDOM[10'h155],
           _RANDOM[10'h156],
           _RANDOM[10'h157],
           _RANDOM[10'h158],
           _RANDOM[10'h159],
           _RANDOM[10'h15A],
           _RANDOM[10'h15B],
           _RANDOM[10'h15C],
           _RANDOM[10'h15D],
           _RANDOM[10'h15E],
           _RANDOM[10'h15F],
           _RANDOM[10'h160],
           _RANDOM[10'h161],
           _RANDOM[10'h162],
           _RANDOM[10'h163],
           _RANDOM[10'h164],
           _RANDOM[10'h165],
           _RANDOM[10'h166],
           _RANDOM[10'h167],
           _RANDOM[10'h168],
           _RANDOM[10'h169],
           _RANDOM[10'h16A],
           _RANDOM[10'h16B],
           _RANDOM[10'h16C],
           _RANDOM[10'h16D],
           _RANDOM[10'h16E],
           _RANDOM[10'h16F],
           _RANDOM[10'h170],
           _RANDOM[10'h171][4:0]};
        dataBuffer_3 =
          {_RANDOM[10'h171][31:5],
           _RANDOM[10'h172],
           _RANDOM[10'h173],
           _RANDOM[10'h174],
           _RANDOM[10'h175],
           _RANDOM[10'h176],
           _RANDOM[10'h177],
           _RANDOM[10'h178],
           _RANDOM[10'h179],
           _RANDOM[10'h17A],
           _RANDOM[10'h17B],
           _RANDOM[10'h17C],
           _RANDOM[10'h17D],
           _RANDOM[10'h17E],
           _RANDOM[10'h17F],
           _RANDOM[10'h180],
           _RANDOM[10'h181],
           _RANDOM[10'h182],
           _RANDOM[10'h183],
           _RANDOM[10'h184],
           _RANDOM[10'h185],
           _RANDOM[10'h186],
           _RANDOM[10'h187],
           _RANDOM[10'h188],
           _RANDOM[10'h189],
           _RANDOM[10'h18A],
           _RANDOM[10'h18B],
           _RANDOM[10'h18C],
           _RANDOM[10'h18D],
           _RANDOM[10'h18E],
           _RANDOM[10'h18F],
           _RANDOM[10'h190],
           _RANDOM[10'h191][4:0]};
        dataBuffer_4 =
          {_RANDOM[10'h191][31:5],
           _RANDOM[10'h192],
           _RANDOM[10'h193],
           _RANDOM[10'h194],
           _RANDOM[10'h195],
           _RANDOM[10'h196],
           _RANDOM[10'h197],
           _RANDOM[10'h198],
           _RANDOM[10'h199],
           _RANDOM[10'h19A],
           _RANDOM[10'h19B],
           _RANDOM[10'h19C],
           _RANDOM[10'h19D],
           _RANDOM[10'h19E],
           _RANDOM[10'h19F],
           _RANDOM[10'h1A0],
           _RANDOM[10'h1A1],
           _RANDOM[10'h1A2],
           _RANDOM[10'h1A3],
           _RANDOM[10'h1A4],
           _RANDOM[10'h1A5],
           _RANDOM[10'h1A6],
           _RANDOM[10'h1A7],
           _RANDOM[10'h1A8],
           _RANDOM[10'h1A9],
           _RANDOM[10'h1AA],
           _RANDOM[10'h1AB],
           _RANDOM[10'h1AC],
           _RANDOM[10'h1AD],
           _RANDOM[10'h1AE],
           _RANDOM[10'h1AF],
           _RANDOM[10'h1B0],
           _RANDOM[10'h1B1][4:0]};
        dataBuffer_5 =
          {_RANDOM[10'h1B1][31:5],
           _RANDOM[10'h1B2],
           _RANDOM[10'h1B3],
           _RANDOM[10'h1B4],
           _RANDOM[10'h1B5],
           _RANDOM[10'h1B6],
           _RANDOM[10'h1B7],
           _RANDOM[10'h1B8],
           _RANDOM[10'h1B9],
           _RANDOM[10'h1BA],
           _RANDOM[10'h1BB],
           _RANDOM[10'h1BC],
           _RANDOM[10'h1BD],
           _RANDOM[10'h1BE],
           _RANDOM[10'h1BF],
           _RANDOM[10'h1C0],
           _RANDOM[10'h1C1],
           _RANDOM[10'h1C2],
           _RANDOM[10'h1C3],
           _RANDOM[10'h1C4],
           _RANDOM[10'h1C5],
           _RANDOM[10'h1C6],
           _RANDOM[10'h1C7],
           _RANDOM[10'h1C8],
           _RANDOM[10'h1C9],
           _RANDOM[10'h1CA],
           _RANDOM[10'h1CB],
           _RANDOM[10'h1CC],
           _RANDOM[10'h1CD],
           _RANDOM[10'h1CE],
           _RANDOM[10'h1CF],
           _RANDOM[10'h1D0],
           _RANDOM[10'h1D1][4:0]};
        dataBuffer_6 =
          {_RANDOM[10'h1D1][31:5],
           _RANDOM[10'h1D2],
           _RANDOM[10'h1D3],
           _RANDOM[10'h1D4],
           _RANDOM[10'h1D5],
           _RANDOM[10'h1D6],
           _RANDOM[10'h1D7],
           _RANDOM[10'h1D8],
           _RANDOM[10'h1D9],
           _RANDOM[10'h1DA],
           _RANDOM[10'h1DB],
           _RANDOM[10'h1DC],
           _RANDOM[10'h1DD],
           _RANDOM[10'h1DE],
           _RANDOM[10'h1DF],
           _RANDOM[10'h1E0],
           _RANDOM[10'h1E1],
           _RANDOM[10'h1E2],
           _RANDOM[10'h1E3],
           _RANDOM[10'h1E4],
           _RANDOM[10'h1E5],
           _RANDOM[10'h1E6],
           _RANDOM[10'h1E7],
           _RANDOM[10'h1E8],
           _RANDOM[10'h1E9],
           _RANDOM[10'h1EA],
           _RANDOM[10'h1EB],
           _RANDOM[10'h1EC],
           _RANDOM[10'h1ED],
           _RANDOM[10'h1EE],
           _RANDOM[10'h1EF],
           _RANDOM[10'h1F0],
           _RANDOM[10'h1F1][4:0]};
        dataBuffer_7 =
          {_RANDOM[10'h1F1][31:5],
           _RANDOM[10'h1F2],
           _RANDOM[10'h1F3],
           _RANDOM[10'h1F4],
           _RANDOM[10'h1F5],
           _RANDOM[10'h1F6],
           _RANDOM[10'h1F7],
           _RANDOM[10'h1F8],
           _RANDOM[10'h1F9],
           _RANDOM[10'h1FA],
           _RANDOM[10'h1FB],
           _RANDOM[10'h1FC],
           _RANDOM[10'h1FD],
           _RANDOM[10'h1FE],
           _RANDOM[10'h1FF],
           _RANDOM[10'h200],
           _RANDOM[10'h201],
           _RANDOM[10'h202],
           _RANDOM[10'h203],
           _RANDOM[10'h204],
           _RANDOM[10'h205],
           _RANDOM[10'h206],
           _RANDOM[10'h207],
           _RANDOM[10'h208],
           _RANDOM[10'h209],
           _RANDOM[10'h20A],
           _RANDOM[10'h20B],
           _RANDOM[10'h20C],
           _RANDOM[10'h20D],
           _RANDOM[10'h20E],
           _RANDOM[10'h20F],
           _RANDOM[10'h210],
           _RANDOM[10'h211][4:0]};
        bufferBaseCacheLineIndex = _RANDOM[10'h211][8:5];
        cacheLineIndexInBuffer = _RANDOM[10'h211][11:9];
        invalidInstructionNext = _RANDOM[10'h211][12];
        segmentInstructionIndexInterval = _RANDOM[10'h211][16:13];
        lastWriteVrfIndexReg = _RANDOM[10'h211][27:17];
        lastCacheNeedPush = _RANDOM[10'h211][28];
        cacheLineNumberReg = {_RANDOM[10'h211][31:29], _RANDOM[10'h212][7:0]};
        lastDataGroupReg = _RANDOM[10'h212][14:8];
        hazardCheck = _RANDOM[10'h212][15];
        readStageValid_segPtr = _RANDOM[10'h212][18:16];
        readStageValid_readCount = _RANDOM[10'h212][21:19];
        readStageValid_stageValid = _RANDOM[10'h212][22];
        readStageValid_readCounter = _RANDOM[10'h212][26:23];
        readStageValid_segPtr_1 = _RANDOM[10'h212][29:27];
        readStageValid_readCount_1 = {_RANDOM[10'h212][31:30], _RANDOM[10'h213][0]};
        readStageValid_stageValid_1 = _RANDOM[10'h213][1];
        readStageValid_readCounter_1 = _RANDOM[10'h213][5:2];
        readStageValid_segPtr_2 = _RANDOM[10'h213][8:6];
        readStageValid_readCount_2 = _RANDOM[10'h213][11:9];
        readStageValid_stageValid_2 = _RANDOM[10'h213][12];
        readStageValid_readCounter_2 = _RANDOM[10'h213][16:13];
        readStageValid_segPtr_3 = _RANDOM[10'h213][19:17];
        readStageValid_readCount_3 = _RANDOM[10'h213][22:20];
        readStageValid_stageValid_3 = _RANDOM[10'h213][23];
        readStageValid_readCounter_3 = _RANDOM[10'h213][27:24];
        readStageValid_segPtr_4 = _RANDOM[10'h213][30:28];
        readStageValid_readCount_4 = {_RANDOM[10'h213][31], _RANDOM[10'h214][1:0]};
        readStageValid_stageValid_4 = _RANDOM[10'h214][2];
        readStageValid_readCounter_4 = _RANDOM[10'h214][6:3];
        readStageValid_segPtr_5 = _RANDOM[10'h214][9:7];
        readStageValid_readCount_5 = _RANDOM[10'h214][12:10];
        readStageValid_stageValid_5 = _RANDOM[10'h214][13];
        readStageValid_readCounter_5 = _RANDOM[10'h214][17:14];
        readStageValid_segPtr_6 = _RANDOM[10'h214][20:18];
        readStageValid_readCount_6 = _RANDOM[10'h214][23:21];
        readStageValid_stageValid_6 = _RANDOM[10'h214][24];
        readStageValid_readCounter_6 = _RANDOM[10'h214][28:25];
        readStageValid_segPtr_7 = _RANDOM[10'h214][31:29];
        readStageValid_readCount_7 = _RANDOM[10'h215][2:0];
        readStageValid_stageValid_7 = _RANDOM[10'h215][3];
        readStageValid_readCounter_7 = _RANDOM[10'h215][7:4];
        readStageValid_segPtr_8 = _RANDOM[10'h215][10:8];
        readStageValid_readCount_8 = _RANDOM[10'h215][13:11];
        readStageValid_stageValid_8 = _RANDOM[10'h215][14];
        readStageValid_readCounter_8 = _RANDOM[10'h215][18:15];
        readStageValid_segPtr_9 = _RANDOM[10'h215][21:19];
        readStageValid_readCount_9 = _RANDOM[10'h215][24:22];
        readStageValid_stageValid_9 = _RANDOM[10'h215][25];
        readStageValid_readCounter_9 = _RANDOM[10'h215][29:26];
        readStageValid_segPtr_10 = {_RANDOM[10'h215][31:30], _RANDOM[10'h216][0]};
        readStageValid_readCount_10 = _RANDOM[10'h216][3:1];
        readStageValid_stageValid_10 = _RANDOM[10'h216][4];
        readStageValid_readCounter_10 = _RANDOM[10'h216][8:5];
        readStageValid_segPtr_11 = _RANDOM[10'h216][11:9];
        readStageValid_readCount_11 = _RANDOM[10'h216][14:12];
        readStageValid_stageValid_11 = _RANDOM[10'h216][15];
        readStageValid_readCounter_11 = _RANDOM[10'h216][19:16];
        readStageValid_segPtr_12 = _RANDOM[10'h216][22:20];
        readStageValid_readCount_12 = _RANDOM[10'h216][25:23];
        readStageValid_stageValid_12 = _RANDOM[10'h216][26];
        readStageValid_readCounter_12 = _RANDOM[10'h216][30:27];
        readStageValid_segPtr_13 = {_RANDOM[10'h216][31], _RANDOM[10'h217][1:0]};
        readStageValid_readCount_13 = _RANDOM[10'h217][4:2];
        readStageValid_stageValid_13 = _RANDOM[10'h217][5];
        readStageValid_readCounter_13 = _RANDOM[10'h217][9:6];
        readStageValid_segPtr_14 = _RANDOM[10'h217][12:10];
        readStageValid_readCount_14 = _RANDOM[10'h217][15:13];
        readStageValid_stageValid_14 = _RANDOM[10'h217][16];
        readStageValid_readCounter_14 = _RANDOM[10'h217][20:17];
        readStageValid_segPtr_15 = _RANDOM[10'h217][23:21];
        readStageValid_readCount_15 = _RANDOM[10'h217][26:24];
        readStageValid_stageValid_15 = _RANDOM[10'h217][27];
        readStageValid_readCounter_15 = _RANDOM[10'h217][31:28];
        readStageValid_segPtr_16 = _RANDOM[10'h218][2:0];
        readStageValid_readCount_16 = _RANDOM[10'h218][5:3];
        readStageValid_stageValid_16 = _RANDOM[10'h218][6];
        readStageValid_readCounter_16 = _RANDOM[10'h218][10:7];
        readStageValid_segPtr_17 = _RANDOM[10'h218][13:11];
        readStageValid_readCount_17 = _RANDOM[10'h218][16:14];
        readStageValid_stageValid_17 = _RANDOM[10'h218][17];
        readStageValid_readCounter_17 = _RANDOM[10'h218][21:18];
        readStageValid_segPtr_18 = _RANDOM[10'h218][24:22];
        readStageValid_readCount_18 = _RANDOM[10'h218][27:25];
        readStageValid_stageValid_18 = _RANDOM[10'h218][28];
        readStageValid_readCounter_18 = {_RANDOM[10'h218][31:29], _RANDOM[10'h219][0]};
        readStageValid_segPtr_19 = _RANDOM[10'h219][3:1];
        readStageValid_readCount_19 = _RANDOM[10'h219][6:4];
        readStageValid_stageValid_19 = _RANDOM[10'h219][7];
        readStageValid_readCounter_19 = _RANDOM[10'h219][11:8];
        readStageValid_segPtr_20 = _RANDOM[10'h219][14:12];
        readStageValid_readCount_20 = _RANDOM[10'h219][17:15];
        readStageValid_stageValid_20 = _RANDOM[10'h219][18];
        readStageValid_readCounter_20 = _RANDOM[10'h219][22:19];
        readStageValid_segPtr_21 = _RANDOM[10'h219][25:23];
        readStageValid_readCount_21 = _RANDOM[10'h219][28:26];
        readStageValid_stageValid_21 = _RANDOM[10'h219][29];
        readStageValid_readCounter_21 = {_RANDOM[10'h219][31:30], _RANDOM[10'h21A][1:0]};
        readStageValid_segPtr_22 = _RANDOM[10'h21A][4:2];
        readStageValid_readCount_22 = _RANDOM[10'h21A][7:5];
        readStageValid_stageValid_22 = _RANDOM[10'h21A][8];
        readStageValid_readCounter_22 = _RANDOM[10'h21A][12:9];
        readStageValid_segPtr_23 = _RANDOM[10'h21A][15:13];
        readStageValid_readCount_23 = _RANDOM[10'h21A][18:16];
        readStageValid_stageValid_23 = _RANDOM[10'h21A][19];
        readStageValid_readCounter_23 = _RANDOM[10'h21A][23:20];
        readStageValid_segPtr_24 = _RANDOM[10'h21A][26:24];
        readStageValid_readCount_24 = _RANDOM[10'h21A][29:27];
        readStageValid_stageValid_24 = _RANDOM[10'h21A][30];
        readStageValid_readCounter_24 = {_RANDOM[10'h21A][31], _RANDOM[10'h21B][2:0]};
        readStageValid_segPtr_25 = _RANDOM[10'h21B][5:3];
        readStageValid_readCount_25 = _RANDOM[10'h21B][8:6];
        readStageValid_stageValid_25 = _RANDOM[10'h21B][9];
        readStageValid_readCounter_25 = _RANDOM[10'h21B][13:10];
        readStageValid_segPtr_26 = _RANDOM[10'h21B][16:14];
        readStageValid_readCount_26 = _RANDOM[10'h21B][19:17];
        readStageValid_stageValid_26 = _RANDOM[10'h21B][20];
        readStageValid_readCounter_26 = _RANDOM[10'h21B][24:21];
        readStageValid_segPtr_27 = _RANDOM[10'h21B][27:25];
        readStageValid_readCount_27 = _RANDOM[10'h21B][30:28];
        readStageValid_stageValid_27 = _RANDOM[10'h21B][31];
        readStageValid_readCounter_27 = _RANDOM[10'h21C][3:0];
        readStageValid_segPtr_28 = _RANDOM[10'h21C][6:4];
        readStageValid_readCount_28 = _RANDOM[10'h21C][9:7];
        readStageValid_stageValid_28 = _RANDOM[10'h21C][10];
        readStageValid_readCounter_28 = _RANDOM[10'h21C][14:11];
        readStageValid_segPtr_29 = _RANDOM[10'h21C][17:15];
        readStageValid_readCount_29 = _RANDOM[10'h21C][20:18];
        readStageValid_stageValid_29 = _RANDOM[10'h21C][21];
        readStageValid_readCounter_29 = _RANDOM[10'h21C][25:22];
        readStageValid_segPtr_30 = _RANDOM[10'h21C][28:26];
        readStageValid_readCount_30 = _RANDOM[10'h21C][31:29];
        readStageValid_stageValid_30 = _RANDOM[10'h21D][0];
        readStageValid_readCounter_30 = _RANDOM[10'h21D][4:1];
        readStageValid_segPtr_31 = _RANDOM[10'h21D][7:5];
        readStageValid_readCount_31 = _RANDOM[10'h21D][10:8];
        readStageValid_stageValid_31 = _RANDOM[10'h21D][11];
        readStageValid_readCounter_31 = _RANDOM[10'h21D][15:12];
        bufferFull = _RANDOM[10'h21D][16];
        bufferValid = _RANDOM[10'h21D][17];
        maskForBufferData_0 = {_RANDOM[10'h21D][31:18], _RANDOM[10'h21E], _RANDOM[10'h21F], _RANDOM[10'h220], _RANDOM[10'h221][17:0]};
        maskForBufferData_1 = {_RANDOM[10'h221][31:18], _RANDOM[10'h222], _RANDOM[10'h223], _RANDOM[10'h224], _RANDOM[10'h225][17:0]};
        maskForBufferData_2 = {_RANDOM[10'h225][31:18], _RANDOM[10'h226], _RANDOM[10'h227], _RANDOM[10'h228], _RANDOM[10'h229][17:0]};
        maskForBufferData_3 = {_RANDOM[10'h229][31:18], _RANDOM[10'h22A], _RANDOM[10'h22B], _RANDOM[10'h22C], _RANDOM[10'h22D][17:0]};
        maskForBufferData_4 = {_RANDOM[10'h22D][31:18], _RANDOM[10'h22E], _RANDOM[10'h22F], _RANDOM[10'h230], _RANDOM[10'h231][17:0]};
        maskForBufferData_5 = {_RANDOM[10'h231][31:18], _RANDOM[10'h232], _RANDOM[10'h233], _RANDOM[10'h234], _RANDOM[10'h235][17:0]};
        maskForBufferData_6 = {_RANDOM[10'h235][31:18], _RANDOM[10'h236], _RANDOM[10'h237], _RANDOM[10'h238], _RANDOM[10'h239][17:0]};
        maskForBufferData_7 = {_RANDOM[10'h239][31:18], _RANDOM[10'h23A], _RANDOM[10'h23B], _RANDOM[10'h23C], _RANDOM[10'h23D][17:0]};
        lastDataGroupInDataBuffer = _RANDOM[10'h23D][18];
        cacheLineTemp =
          {_RANDOM[10'h23D][31:19],
           _RANDOM[10'h23E],
           _RANDOM[10'h23F],
           _RANDOM[10'h240],
           _RANDOM[10'h241],
           _RANDOM[10'h242],
           _RANDOM[10'h243],
           _RANDOM[10'h244],
           _RANDOM[10'h245],
           _RANDOM[10'h246],
           _RANDOM[10'h247],
           _RANDOM[10'h248],
           _RANDOM[10'h249],
           _RANDOM[10'h24A],
           _RANDOM[10'h24B],
           _RANDOM[10'h24C],
           _RANDOM[10'h24D],
           _RANDOM[10'h24E],
           _RANDOM[10'h24F],
           _RANDOM[10'h250],
           _RANDOM[10'h251],
           _RANDOM[10'h252],
           _RANDOM[10'h253],
           _RANDOM[10'h254],
           _RANDOM[10'h255],
           _RANDOM[10'h256],
           _RANDOM[10'h257],
           _RANDOM[10'h258],
           _RANDOM[10'h259],
           _RANDOM[10'h25A],
           _RANDOM[10'h25B],
           _RANDOM[10'h25C],
           _RANDOM[10'h25D][18:0]};
        maskTemp = {_RANDOM[10'h25D][31:19], _RANDOM[10'h25E], _RANDOM[10'h25F], _RANDOM[10'h260], _RANDOM[10'h261][18:0]};
        canSendTail = _RANDOM[10'h261][19];
        idleNext = _RANDOM[10'h261][20];
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  wire              vrfReadQueueVec_0_empty;
  assign vrfReadQueueVec_0_empty = _vrfReadQueueVec_fifo_empty;
  wire              vrfReadQueueVec_0_full;
  assign vrfReadQueueVec_0_full = _vrfReadQueueVec_fifo_full;
  wire              vrfReadQueueVec_1_empty;
  assign vrfReadQueueVec_1_empty = _vrfReadQueueVec_fifo_1_empty;
  wire              vrfReadQueueVec_1_full;
  assign vrfReadQueueVec_1_full = _vrfReadQueueVec_fifo_1_full;
  wire              vrfReadQueueVec_2_empty;
  assign vrfReadQueueVec_2_empty = _vrfReadQueueVec_fifo_2_empty;
  wire              vrfReadQueueVec_2_full;
  assign vrfReadQueueVec_2_full = _vrfReadQueueVec_fifo_2_full;
  wire              vrfReadQueueVec_3_empty;
  assign vrfReadQueueVec_3_empty = _vrfReadQueueVec_fifo_3_empty;
  wire              vrfReadQueueVec_3_full;
  assign vrfReadQueueVec_3_full = _vrfReadQueueVec_fifo_3_full;
  wire              vrfReadQueueVec_4_empty;
  assign vrfReadQueueVec_4_empty = _vrfReadQueueVec_fifo_4_empty;
  wire              vrfReadQueueVec_4_full;
  assign vrfReadQueueVec_4_full = _vrfReadQueueVec_fifo_4_full;
  wire              vrfReadQueueVec_5_empty;
  assign vrfReadQueueVec_5_empty = _vrfReadQueueVec_fifo_5_empty;
  wire              vrfReadQueueVec_5_full;
  assign vrfReadQueueVec_5_full = _vrfReadQueueVec_fifo_5_full;
  wire              vrfReadQueueVec_6_empty;
  assign vrfReadQueueVec_6_empty = _vrfReadQueueVec_fifo_6_empty;
  wire              vrfReadQueueVec_6_full;
  assign vrfReadQueueVec_6_full = _vrfReadQueueVec_fifo_6_full;
  wire              vrfReadQueueVec_7_empty;
  assign vrfReadQueueVec_7_empty = _vrfReadQueueVec_fifo_7_empty;
  wire              vrfReadQueueVec_7_full;
  assign vrfReadQueueVec_7_full = _vrfReadQueueVec_fifo_7_full;
  wire              vrfReadQueueVec_8_empty;
  assign vrfReadQueueVec_8_empty = _vrfReadQueueVec_fifo_8_empty;
  wire              vrfReadQueueVec_8_full;
  assign vrfReadQueueVec_8_full = _vrfReadQueueVec_fifo_8_full;
  wire              vrfReadQueueVec_9_empty;
  assign vrfReadQueueVec_9_empty = _vrfReadQueueVec_fifo_9_empty;
  wire              vrfReadQueueVec_9_full;
  assign vrfReadQueueVec_9_full = _vrfReadQueueVec_fifo_9_full;
  wire              vrfReadQueueVec_10_empty;
  assign vrfReadQueueVec_10_empty = _vrfReadQueueVec_fifo_10_empty;
  wire              vrfReadQueueVec_10_full;
  assign vrfReadQueueVec_10_full = _vrfReadQueueVec_fifo_10_full;
  wire              vrfReadQueueVec_11_empty;
  assign vrfReadQueueVec_11_empty = _vrfReadQueueVec_fifo_11_empty;
  wire              vrfReadQueueVec_11_full;
  assign vrfReadQueueVec_11_full = _vrfReadQueueVec_fifo_11_full;
  wire              vrfReadQueueVec_12_empty;
  assign vrfReadQueueVec_12_empty = _vrfReadQueueVec_fifo_12_empty;
  wire              vrfReadQueueVec_12_full;
  assign vrfReadQueueVec_12_full = _vrfReadQueueVec_fifo_12_full;
  wire              vrfReadQueueVec_13_empty;
  assign vrfReadQueueVec_13_empty = _vrfReadQueueVec_fifo_13_empty;
  wire              vrfReadQueueVec_13_full;
  assign vrfReadQueueVec_13_full = _vrfReadQueueVec_fifo_13_full;
  wire              vrfReadQueueVec_14_empty;
  assign vrfReadQueueVec_14_empty = _vrfReadQueueVec_fifo_14_empty;
  wire              vrfReadQueueVec_14_full;
  assign vrfReadQueueVec_14_full = _vrfReadQueueVec_fifo_14_full;
  wire              vrfReadQueueVec_15_empty;
  assign vrfReadQueueVec_15_empty = _vrfReadQueueVec_fifo_15_empty;
  wire              vrfReadQueueVec_15_full;
  assign vrfReadQueueVec_15_full = _vrfReadQueueVec_fifo_15_full;
  wire              vrfReadQueueVec_16_empty;
  assign vrfReadQueueVec_16_empty = _vrfReadQueueVec_fifo_16_empty;
  wire              vrfReadQueueVec_16_full;
  assign vrfReadQueueVec_16_full = _vrfReadQueueVec_fifo_16_full;
  wire              vrfReadQueueVec_17_empty;
  assign vrfReadQueueVec_17_empty = _vrfReadQueueVec_fifo_17_empty;
  wire              vrfReadQueueVec_17_full;
  assign vrfReadQueueVec_17_full = _vrfReadQueueVec_fifo_17_full;
  wire              vrfReadQueueVec_18_empty;
  assign vrfReadQueueVec_18_empty = _vrfReadQueueVec_fifo_18_empty;
  wire              vrfReadQueueVec_18_full;
  assign vrfReadQueueVec_18_full = _vrfReadQueueVec_fifo_18_full;
  wire              vrfReadQueueVec_19_empty;
  assign vrfReadQueueVec_19_empty = _vrfReadQueueVec_fifo_19_empty;
  wire              vrfReadQueueVec_19_full;
  assign vrfReadQueueVec_19_full = _vrfReadQueueVec_fifo_19_full;
  wire              vrfReadQueueVec_20_empty;
  assign vrfReadQueueVec_20_empty = _vrfReadQueueVec_fifo_20_empty;
  wire              vrfReadQueueVec_20_full;
  assign vrfReadQueueVec_20_full = _vrfReadQueueVec_fifo_20_full;
  wire              vrfReadQueueVec_21_empty;
  assign vrfReadQueueVec_21_empty = _vrfReadQueueVec_fifo_21_empty;
  wire              vrfReadQueueVec_21_full;
  assign vrfReadQueueVec_21_full = _vrfReadQueueVec_fifo_21_full;
  wire              vrfReadQueueVec_22_empty;
  assign vrfReadQueueVec_22_empty = _vrfReadQueueVec_fifo_22_empty;
  wire              vrfReadQueueVec_22_full;
  assign vrfReadQueueVec_22_full = _vrfReadQueueVec_fifo_22_full;
  wire              vrfReadQueueVec_23_empty;
  assign vrfReadQueueVec_23_empty = _vrfReadQueueVec_fifo_23_empty;
  wire              vrfReadQueueVec_23_full;
  assign vrfReadQueueVec_23_full = _vrfReadQueueVec_fifo_23_full;
  wire              vrfReadQueueVec_24_empty;
  assign vrfReadQueueVec_24_empty = _vrfReadQueueVec_fifo_24_empty;
  wire              vrfReadQueueVec_24_full;
  assign vrfReadQueueVec_24_full = _vrfReadQueueVec_fifo_24_full;
  wire              vrfReadQueueVec_25_empty;
  assign vrfReadQueueVec_25_empty = _vrfReadQueueVec_fifo_25_empty;
  wire              vrfReadQueueVec_25_full;
  assign vrfReadQueueVec_25_full = _vrfReadQueueVec_fifo_25_full;
  wire              vrfReadQueueVec_26_empty;
  assign vrfReadQueueVec_26_empty = _vrfReadQueueVec_fifo_26_empty;
  wire              vrfReadQueueVec_26_full;
  assign vrfReadQueueVec_26_full = _vrfReadQueueVec_fifo_26_full;
  wire              vrfReadQueueVec_27_empty;
  assign vrfReadQueueVec_27_empty = _vrfReadQueueVec_fifo_27_empty;
  wire              vrfReadQueueVec_27_full;
  assign vrfReadQueueVec_27_full = _vrfReadQueueVec_fifo_27_full;
  wire              vrfReadQueueVec_28_empty;
  assign vrfReadQueueVec_28_empty = _vrfReadQueueVec_fifo_28_empty;
  wire              vrfReadQueueVec_28_full;
  assign vrfReadQueueVec_28_full = _vrfReadQueueVec_fifo_28_full;
  wire              vrfReadQueueVec_29_empty;
  assign vrfReadQueueVec_29_empty = _vrfReadQueueVec_fifo_29_empty;
  wire              vrfReadQueueVec_29_full;
  assign vrfReadQueueVec_29_full = _vrfReadQueueVec_fifo_29_full;
  wire              vrfReadQueueVec_30_empty;
  assign vrfReadQueueVec_30_empty = _vrfReadQueueVec_fifo_30_empty;
  wire              vrfReadQueueVec_30_full;
  assign vrfReadQueueVec_30_full = _vrfReadQueueVec_fifo_30_full;
  wire              vrfReadQueueVec_31_empty;
  assign vrfReadQueueVec_31_empty = _vrfReadQueueVec_fifo_31_empty;
  wire              vrfReadQueueVec_31_full;
  assign vrfReadQueueVec_31_full = _vrfReadQueueVec_fifo_31_full;
  wire              addressQueue_empty;
  assign addressQueue_empty = _addressQueue_fifo_empty;
  wire              addressQueue_full;
  assign addressQueue_full = _addressQueue_fifo_full;
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_0_enq_ready & vrfReadQueueVec_0_enq_valid & ~(_vrfReadQueueVec_fifo_empty & vrfReadQueueVec_0_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_0_deq_ready & ~_vrfReadQueueVec_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_0_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_empty),
    .almost_empty (vrfReadQueueVec_0_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_0_almostFull),
    .full         (_vrfReadQueueVec_fifo_full),
    .error        (_vrfReadQueueVec_fifo_error),
    .data_out     (_vrfReadQueueVec_fifo_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_1 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_1_enq_ready & vrfReadQueueVec_1_enq_valid & ~(_vrfReadQueueVec_fifo_1_empty & vrfReadQueueVec_1_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_1_deq_ready & ~_vrfReadQueueVec_fifo_1_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_1_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_1_empty),
    .almost_empty (vrfReadQueueVec_1_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_1_almostFull),
    .full         (_vrfReadQueueVec_fifo_1_full),
    .error        (_vrfReadQueueVec_fifo_1_error),
    .data_out     (_vrfReadQueueVec_fifo_1_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_2 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_2_enq_ready & vrfReadQueueVec_2_enq_valid & ~(_vrfReadQueueVec_fifo_2_empty & vrfReadQueueVec_2_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_2_deq_ready & ~_vrfReadQueueVec_fifo_2_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_2_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_2_empty),
    .almost_empty (vrfReadQueueVec_2_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_2_almostFull),
    .full         (_vrfReadQueueVec_fifo_2_full),
    .error        (_vrfReadQueueVec_fifo_2_error),
    .data_out     (_vrfReadQueueVec_fifo_2_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_3 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_3_enq_ready & vrfReadQueueVec_3_enq_valid & ~(_vrfReadQueueVec_fifo_3_empty & vrfReadQueueVec_3_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_3_deq_ready & ~_vrfReadQueueVec_fifo_3_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_3_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_3_empty),
    .almost_empty (vrfReadQueueVec_3_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_3_almostFull),
    .full         (_vrfReadQueueVec_fifo_3_full),
    .error        (_vrfReadQueueVec_fifo_3_error),
    .data_out     (_vrfReadQueueVec_fifo_3_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_4 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_4_enq_ready & vrfReadQueueVec_4_enq_valid & ~(_vrfReadQueueVec_fifo_4_empty & vrfReadQueueVec_4_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_4_deq_ready & ~_vrfReadQueueVec_fifo_4_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_4_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_4_empty),
    .almost_empty (vrfReadQueueVec_4_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_4_almostFull),
    .full         (_vrfReadQueueVec_fifo_4_full),
    .error        (_vrfReadQueueVec_fifo_4_error),
    .data_out     (_vrfReadQueueVec_fifo_4_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_5 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_5_enq_ready & vrfReadQueueVec_5_enq_valid & ~(_vrfReadQueueVec_fifo_5_empty & vrfReadQueueVec_5_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_5_deq_ready & ~_vrfReadQueueVec_fifo_5_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_5_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_5_empty),
    .almost_empty (vrfReadQueueVec_5_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_5_almostFull),
    .full         (_vrfReadQueueVec_fifo_5_full),
    .error        (_vrfReadQueueVec_fifo_5_error),
    .data_out     (_vrfReadQueueVec_fifo_5_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_6 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_6_enq_ready & vrfReadQueueVec_6_enq_valid & ~(_vrfReadQueueVec_fifo_6_empty & vrfReadQueueVec_6_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_6_deq_ready & ~_vrfReadQueueVec_fifo_6_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_6_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_6_empty),
    .almost_empty (vrfReadQueueVec_6_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_6_almostFull),
    .full         (_vrfReadQueueVec_fifo_6_full),
    .error        (_vrfReadQueueVec_fifo_6_error),
    .data_out     (_vrfReadQueueVec_fifo_6_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_7 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_7_enq_ready & vrfReadQueueVec_7_enq_valid & ~(_vrfReadQueueVec_fifo_7_empty & vrfReadQueueVec_7_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_7_deq_ready & ~_vrfReadQueueVec_fifo_7_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_7_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_7_empty),
    .almost_empty (vrfReadQueueVec_7_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_7_almostFull),
    .full         (_vrfReadQueueVec_fifo_7_full),
    .error        (_vrfReadQueueVec_fifo_7_error),
    .data_out     (_vrfReadQueueVec_fifo_7_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_8 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_8_enq_ready & vrfReadQueueVec_8_enq_valid & ~(_vrfReadQueueVec_fifo_8_empty & vrfReadQueueVec_8_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_8_deq_ready & ~_vrfReadQueueVec_fifo_8_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_8_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_8_empty),
    .almost_empty (vrfReadQueueVec_8_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_8_almostFull),
    .full         (_vrfReadQueueVec_fifo_8_full),
    .error        (_vrfReadQueueVec_fifo_8_error),
    .data_out     (_vrfReadQueueVec_fifo_8_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_9 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_9_enq_ready & vrfReadQueueVec_9_enq_valid & ~(_vrfReadQueueVec_fifo_9_empty & vrfReadQueueVec_9_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_9_deq_ready & ~_vrfReadQueueVec_fifo_9_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_9_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_9_empty),
    .almost_empty (vrfReadQueueVec_9_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_9_almostFull),
    .full         (_vrfReadQueueVec_fifo_9_full),
    .error        (_vrfReadQueueVec_fifo_9_error),
    .data_out     (_vrfReadQueueVec_fifo_9_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_10 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_10_enq_ready & vrfReadQueueVec_10_enq_valid & ~(_vrfReadQueueVec_fifo_10_empty & vrfReadQueueVec_10_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_10_deq_ready & ~_vrfReadQueueVec_fifo_10_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_10_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_10_empty),
    .almost_empty (vrfReadQueueVec_10_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_10_almostFull),
    .full         (_vrfReadQueueVec_fifo_10_full),
    .error        (_vrfReadQueueVec_fifo_10_error),
    .data_out     (_vrfReadQueueVec_fifo_10_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_11 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_11_enq_ready & vrfReadQueueVec_11_enq_valid & ~(_vrfReadQueueVec_fifo_11_empty & vrfReadQueueVec_11_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_11_deq_ready & ~_vrfReadQueueVec_fifo_11_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_11_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_11_empty),
    .almost_empty (vrfReadQueueVec_11_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_11_almostFull),
    .full         (_vrfReadQueueVec_fifo_11_full),
    .error        (_vrfReadQueueVec_fifo_11_error),
    .data_out     (_vrfReadQueueVec_fifo_11_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_12 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_12_enq_ready & vrfReadQueueVec_12_enq_valid & ~(_vrfReadQueueVec_fifo_12_empty & vrfReadQueueVec_12_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_12_deq_ready & ~_vrfReadQueueVec_fifo_12_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_12_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_12_empty),
    .almost_empty (vrfReadQueueVec_12_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_12_almostFull),
    .full         (_vrfReadQueueVec_fifo_12_full),
    .error        (_vrfReadQueueVec_fifo_12_error),
    .data_out     (_vrfReadQueueVec_fifo_12_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_13 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_13_enq_ready & vrfReadQueueVec_13_enq_valid & ~(_vrfReadQueueVec_fifo_13_empty & vrfReadQueueVec_13_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_13_deq_ready & ~_vrfReadQueueVec_fifo_13_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_13_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_13_empty),
    .almost_empty (vrfReadQueueVec_13_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_13_almostFull),
    .full         (_vrfReadQueueVec_fifo_13_full),
    .error        (_vrfReadQueueVec_fifo_13_error),
    .data_out     (_vrfReadQueueVec_fifo_13_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_14 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_14_enq_ready & vrfReadQueueVec_14_enq_valid & ~(_vrfReadQueueVec_fifo_14_empty & vrfReadQueueVec_14_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_14_deq_ready & ~_vrfReadQueueVec_fifo_14_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_14_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_14_empty),
    .almost_empty (vrfReadQueueVec_14_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_14_almostFull),
    .full         (_vrfReadQueueVec_fifo_14_full),
    .error        (_vrfReadQueueVec_fifo_14_error),
    .data_out     (_vrfReadQueueVec_fifo_14_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_15 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_15_enq_ready & vrfReadQueueVec_15_enq_valid & ~(_vrfReadQueueVec_fifo_15_empty & vrfReadQueueVec_15_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_15_deq_ready & ~_vrfReadQueueVec_fifo_15_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_15_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_15_empty),
    .almost_empty (vrfReadQueueVec_15_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_15_almostFull),
    .full         (_vrfReadQueueVec_fifo_15_full),
    .error        (_vrfReadQueueVec_fifo_15_error),
    .data_out     (_vrfReadQueueVec_fifo_15_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_16 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_16_enq_ready & vrfReadQueueVec_16_enq_valid & ~(_vrfReadQueueVec_fifo_16_empty & vrfReadQueueVec_16_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_16_deq_ready & ~_vrfReadQueueVec_fifo_16_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_16_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_16_empty),
    .almost_empty (vrfReadQueueVec_16_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_16_almostFull),
    .full         (_vrfReadQueueVec_fifo_16_full),
    .error        (_vrfReadQueueVec_fifo_16_error),
    .data_out     (_vrfReadQueueVec_fifo_16_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_17 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_17_enq_ready & vrfReadQueueVec_17_enq_valid & ~(_vrfReadQueueVec_fifo_17_empty & vrfReadQueueVec_17_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_17_deq_ready & ~_vrfReadQueueVec_fifo_17_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_17_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_17_empty),
    .almost_empty (vrfReadQueueVec_17_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_17_almostFull),
    .full         (_vrfReadQueueVec_fifo_17_full),
    .error        (_vrfReadQueueVec_fifo_17_error),
    .data_out     (_vrfReadQueueVec_fifo_17_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_18 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_18_enq_ready & vrfReadQueueVec_18_enq_valid & ~(_vrfReadQueueVec_fifo_18_empty & vrfReadQueueVec_18_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_18_deq_ready & ~_vrfReadQueueVec_fifo_18_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_18_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_18_empty),
    .almost_empty (vrfReadQueueVec_18_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_18_almostFull),
    .full         (_vrfReadQueueVec_fifo_18_full),
    .error        (_vrfReadQueueVec_fifo_18_error),
    .data_out     (_vrfReadQueueVec_fifo_18_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_19 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_19_enq_ready & vrfReadQueueVec_19_enq_valid & ~(_vrfReadQueueVec_fifo_19_empty & vrfReadQueueVec_19_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_19_deq_ready & ~_vrfReadQueueVec_fifo_19_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_19_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_19_empty),
    .almost_empty (vrfReadQueueVec_19_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_19_almostFull),
    .full         (_vrfReadQueueVec_fifo_19_full),
    .error        (_vrfReadQueueVec_fifo_19_error),
    .data_out     (_vrfReadQueueVec_fifo_19_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_20 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_20_enq_ready & vrfReadQueueVec_20_enq_valid & ~(_vrfReadQueueVec_fifo_20_empty & vrfReadQueueVec_20_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_20_deq_ready & ~_vrfReadQueueVec_fifo_20_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_20_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_20_empty),
    .almost_empty (vrfReadQueueVec_20_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_20_almostFull),
    .full         (_vrfReadQueueVec_fifo_20_full),
    .error        (_vrfReadQueueVec_fifo_20_error),
    .data_out     (_vrfReadQueueVec_fifo_20_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_21 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_21_enq_ready & vrfReadQueueVec_21_enq_valid & ~(_vrfReadQueueVec_fifo_21_empty & vrfReadQueueVec_21_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_21_deq_ready & ~_vrfReadQueueVec_fifo_21_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_21_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_21_empty),
    .almost_empty (vrfReadQueueVec_21_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_21_almostFull),
    .full         (_vrfReadQueueVec_fifo_21_full),
    .error        (_vrfReadQueueVec_fifo_21_error),
    .data_out     (_vrfReadQueueVec_fifo_21_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_22 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_22_enq_ready & vrfReadQueueVec_22_enq_valid & ~(_vrfReadQueueVec_fifo_22_empty & vrfReadQueueVec_22_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_22_deq_ready & ~_vrfReadQueueVec_fifo_22_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_22_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_22_empty),
    .almost_empty (vrfReadQueueVec_22_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_22_almostFull),
    .full         (_vrfReadQueueVec_fifo_22_full),
    .error        (_vrfReadQueueVec_fifo_22_error),
    .data_out     (_vrfReadQueueVec_fifo_22_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_23 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_23_enq_ready & vrfReadQueueVec_23_enq_valid & ~(_vrfReadQueueVec_fifo_23_empty & vrfReadQueueVec_23_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_23_deq_ready & ~_vrfReadQueueVec_fifo_23_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_23_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_23_empty),
    .almost_empty (vrfReadQueueVec_23_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_23_almostFull),
    .full         (_vrfReadQueueVec_fifo_23_full),
    .error        (_vrfReadQueueVec_fifo_23_error),
    .data_out     (_vrfReadQueueVec_fifo_23_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_24 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_24_enq_ready & vrfReadQueueVec_24_enq_valid & ~(_vrfReadQueueVec_fifo_24_empty & vrfReadQueueVec_24_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_24_deq_ready & ~_vrfReadQueueVec_fifo_24_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_24_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_24_empty),
    .almost_empty (vrfReadQueueVec_24_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_24_almostFull),
    .full         (_vrfReadQueueVec_fifo_24_full),
    .error        (_vrfReadQueueVec_fifo_24_error),
    .data_out     (_vrfReadQueueVec_fifo_24_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_25 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_25_enq_ready & vrfReadQueueVec_25_enq_valid & ~(_vrfReadQueueVec_fifo_25_empty & vrfReadQueueVec_25_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_25_deq_ready & ~_vrfReadQueueVec_fifo_25_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_25_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_25_empty),
    .almost_empty (vrfReadQueueVec_25_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_25_almostFull),
    .full         (_vrfReadQueueVec_fifo_25_full),
    .error        (_vrfReadQueueVec_fifo_25_error),
    .data_out     (_vrfReadQueueVec_fifo_25_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_26 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_26_enq_ready & vrfReadQueueVec_26_enq_valid & ~(_vrfReadQueueVec_fifo_26_empty & vrfReadQueueVec_26_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_26_deq_ready & ~_vrfReadQueueVec_fifo_26_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_26_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_26_empty),
    .almost_empty (vrfReadQueueVec_26_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_26_almostFull),
    .full         (_vrfReadQueueVec_fifo_26_full),
    .error        (_vrfReadQueueVec_fifo_26_error),
    .data_out     (_vrfReadQueueVec_fifo_26_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_27 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_27_enq_ready & vrfReadQueueVec_27_enq_valid & ~(_vrfReadQueueVec_fifo_27_empty & vrfReadQueueVec_27_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_27_deq_ready & ~_vrfReadQueueVec_fifo_27_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_27_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_27_empty),
    .almost_empty (vrfReadQueueVec_27_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_27_almostFull),
    .full         (_vrfReadQueueVec_fifo_27_full),
    .error        (_vrfReadQueueVec_fifo_27_error),
    .data_out     (_vrfReadQueueVec_fifo_27_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_28 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_28_enq_ready & vrfReadQueueVec_28_enq_valid & ~(_vrfReadQueueVec_fifo_28_empty & vrfReadQueueVec_28_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_28_deq_ready & ~_vrfReadQueueVec_fifo_28_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_28_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_28_empty),
    .almost_empty (vrfReadQueueVec_28_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_28_almostFull),
    .full         (_vrfReadQueueVec_fifo_28_full),
    .error        (_vrfReadQueueVec_fifo_28_error),
    .data_out     (_vrfReadQueueVec_fifo_28_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_29 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_29_enq_ready & vrfReadQueueVec_29_enq_valid & ~(_vrfReadQueueVec_fifo_29_empty & vrfReadQueueVec_29_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_29_deq_ready & ~_vrfReadQueueVec_fifo_29_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_29_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_29_empty),
    .almost_empty (vrfReadQueueVec_29_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_29_almostFull),
    .full         (_vrfReadQueueVec_fifo_29_full),
    .error        (_vrfReadQueueVec_fifo_29_error),
    .data_out     (_vrfReadQueueVec_fifo_29_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_30 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_30_enq_ready & vrfReadQueueVec_30_enq_valid & ~(_vrfReadQueueVec_fifo_30_empty & vrfReadQueueVec_30_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_30_deq_ready & ~_vrfReadQueueVec_fifo_30_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_30_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_30_empty),
    .almost_empty (vrfReadQueueVec_30_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_30_almostFull),
    .full         (_vrfReadQueueVec_fifo_30_full),
    .error        (_vrfReadQueueVec_fifo_30_error),
    .data_out     (_vrfReadQueueVec_fifo_30_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(8),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) vrfReadQueueVec_fifo_31 (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(vrfReadQueueVec_31_enq_ready & vrfReadQueueVec_31_enq_valid & ~(_vrfReadQueueVec_fifo_31_empty & vrfReadQueueVec_31_deq_ready))),
    .pop_req_n    (~(vrfReadQueueVec_31_deq_ready & ~_vrfReadQueueVec_fifo_31_empty)),
    .diag_n       (1'h1),
    .data_in      (vrfReadQueueVec_31_enq_bits),
    .empty        (_vrfReadQueueVec_fifo_31_empty),
    .almost_empty (vrfReadQueueVec_31_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (vrfReadQueueVec_31_almostFull),
    .full         (_vrfReadQueueVec_fifo_31_full),
    .error        (_vrfReadQueueVec_fifo_31_error),
    .data_out     (_vrfReadQueueVec_fifo_31_data_out)
  );
  DW_fifo_s1_sf #(
    .ae_level(1),
    .af_level(1),
    .depth(9),
    .err_mode(2),
    .rst_mode(3),
    .width(32)
  ) addressQueue_fifo (
    .clk          (clock),
    .rst_n        (~reset),
    .push_req_n   (~(addressQueue_enq_ready & addressQueue_enq_valid)),
    .pop_req_n    (~(addressQueue_deq_ready & ~_addressQueue_fifo_empty)),
    .diag_n       (1'h1),
    .data_in      (addressQueue_enq_bits),
    .empty        (_addressQueue_fifo_empty),
    .almost_empty (addressQueue_almostEmpty),
    .half_full    (/* unused */),
    .almost_full  (addressQueue_almostFull),
    .full         (_addressQueue_fifo_full),
    .error        (_addressQueue_fifo_error),
    .data_out     (addressQueue_deq_bits)
  );
  assign maskSelect_valid = _maskSelect_valid_output;
  assign maskSelect_bits = _maskSelect_bits_output;
  assign memRequest_valid = memRequest_valid_0;
  assign memRequest_bits_data = memRequest_bits_data_0;
  assign memRequest_bits_mask = memRequest_bits_mask_0;
  assign memRequest_bits_index = memRequest_bits_index_0;
  assign memRequest_bits_address = memRequest_bits_address_0;
  assign status_idle = _status_idle_output;
  assign status_last = ~idleNext & _status_idle_output | invalidInstructionNext;
  assign status_instructionIndex = lsuRequestReg_instructionIndex;
  assign status_changeMaskGroup = _maskSelect_valid_output & ~lsuRequest_valid;
  assign status_startAddress = addressQueue_deq_valid ? addressQueue_deq_bits : alignedDequeueAddress;
  assign status_endAddress = {lsuRequestReg_rs1Data[31:7] + {14'h0, cacheLineNumberReg}, 7'h0};
  assign vrfReadDataPorts_0_valid = vrfReadDataPorts_0_valid_0;
  assign vrfReadDataPorts_0_bits_vs = vrfReadDataPorts_0_bits_vs_0;
  assign vrfReadDataPorts_0_bits_instructionIndex = vrfReadDataPorts_0_bits_instructionIndex_0;
  assign vrfReadDataPorts_1_valid = vrfReadDataPorts_1_valid_0;
  assign vrfReadDataPorts_1_bits_vs = vrfReadDataPorts_1_bits_vs_0;
  assign vrfReadDataPorts_1_bits_instructionIndex = vrfReadDataPorts_1_bits_instructionIndex_0;
  assign vrfReadDataPorts_2_valid = vrfReadDataPorts_2_valid_0;
  assign vrfReadDataPorts_2_bits_vs = vrfReadDataPorts_2_bits_vs_0;
  assign vrfReadDataPorts_2_bits_instructionIndex = vrfReadDataPorts_2_bits_instructionIndex_0;
  assign vrfReadDataPorts_3_valid = vrfReadDataPorts_3_valid_0;
  assign vrfReadDataPorts_3_bits_vs = vrfReadDataPorts_3_bits_vs_0;
  assign vrfReadDataPorts_3_bits_instructionIndex = vrfReadDataPorts_3_bits_instructionIndex_0;
  assign vrfReadDataPorts_4_valid = vrfReadDataPorts_4_valid_0;
  assign vrfReadDataPorts_4_bits_vs = vrfReadDataPorts_4_bits_vs_0;
  assign vrfReadDataPorts_4_bits_instructionIndex = vrfReadDataPorts_4_bits_instructionIndex_0;
  assign vrfReadDataPorts_5_valid = vrfReadDataPorts_5_valid_0;
  assign vrfReadDataPorts_5_bits_vs = vrfReadDataPorts_5_bits_vs_0;
  assign vrfReadDataPorts_5_bits_instructionIndex = vrfReadDataPorts_5_bits_instructionIndex_0;
  assign vrfReadDataPorts_6_valid = vrfReadDataPorts_6_valid_0;
  assign vrfReadDataPorts_6_bits_vs = vrfReadDataPorts_6_bits_vs_0;
  assign vrfReadDataPorts_6_bits_instructionIndex = vrfReadDataPorts_6_bits_instructionIndex_0;
  assign vrfReadDataPorts_7_valid = vrfReadDataPorts_7_valid_0;
  assign vrfReadDataPorts_7_bits_vs = vrfReadDataPorts_7_bits_vs_0;
  assign vrfReadDataPorts_7_bits_instructionIndex = vrfReadDataPorts_7_bits_instructionIndex_0;
  assign vrfReadDataPorts_8_valid = vrfReadDataPorts_8_valid_0;
  assign vrfReadDataPorts_8_bits_vs = vrfReadDataPorts_8_bits_vs_0;
  assign vrfReadDataPorts_8_bits_instructionIndex = vrfReadDataPorts_8_bits_instructionIndex_0;
  assign vrfReadDataPorts_9_valid = vrfReadDataPorts_9_valid_0;
  assign vrfReadDataPorts_9_bits_vs = vrfReadDataPorts_9_bits_vs_0;
  assign vrfReadDataPorts_9_bits_instructionIndex = vrfReadDataPorts_9_bits_instructionIndex_0;
  assign vrfReadDataPorts_10_valid = vrfReadDataPorts_10_valid_0;
  assign vrfReadDataPorts_10_bits_vs = vrfReadDataPorts_10_bits_vs_0;
  assign vrfReadDataPorts_10_bits_instructionIndex = vrfReadDataPorts_10_bits_instructionIndex_0;
  assign vrfReadDataPorts_11_valid = vrfReadDataPorts_11_valid_0;
  assign vrfReadDataPorts_11_bits_vs = vrfReadDataPorts_11_bits_vs_0;
  assign vrfReadDataPorts_11_bits_instructionIndex = vrfReadDataPorts_11_bits_instructionIndex_0;
  assign vrfReadDataPorts_12_valid = vrfReadDataPorts_12_valid_0;
  assign vrfReadDataPorts_12_bits_vs = vrfReadDataPorts_12_bits_vs_0;
  assign vrfReadDataPorts_12_bits_instructionIndex = vrfReadDataPorts_12_bits_instructionIndex_0;
  assign vrfReadDataPorts_13_valid = vrfReadDataPorts_13_valid_0;
  assign vrfReadDataPorts_13_bits_vs = vrfReadDataPorts_13_bits_vs_0;
  assign vrfReadDataPorts_13_bits_instructionIndex = vrfReadDataPorts_13_bits_instructionIndex_0;
  assign vrfReadDataPorts_14_valid = vrfReadDataPorts_14_valid_0;
  assign vrfReadDataPorts_14_bits_vs = vrfReadDataPorts_14_bits_vs_0;
  assign vrfReadDataPorts_14_bits_instructionIndex = vrfReadDataPorts_14_bits_instructionIndex_0;
  assign vrfReadDataPorts_15_valid = vrfReadDataPorts_15_valid_0;
  assign vrfReadDataPorts_15_bits_vs = vrfReadDataPorts_15_bits_vs_0;
  assign vrfReadDataPorts_15_bits_instructionIndex = vrfReadDataPorts_15_bits_instructionIndex_0;
  assign vrfReadDataPorts_16_valid = vrfReadDataPorts_16_valid_0;
  assign vrfReadDataPorts_16_bits_vs = vrfReadDataPorts_16_bits_vs_0;
  assign vrfReadDataPorts_16_bits_instructionIndex = vrfReadDataPorts_16_bits_instructionIndex_0;
  assign vrfReadDataPorts_17_valid = vrfReadDataPorts_17_valid_0;
  assign vrfReadDataPorts_17_bits_vs = vrfReadDataPorts_17_bits_vs_0;
  assign vrfReadDataPorts_17_bits_instructionIndex = vrfReadDataPorts_17_bits_instructionIndex_0;
  assign vrfReadDataPorts_18_valid = vrfReadDataPorts_18_valid_0;
  assign vrfReadDataPorts_18_bits_vs = vrfReadDataPorts_18_bits_vs_0;
  assign vrfReadDataPorts_18_bits_instructionIndex = vrfReadDataPorts_18_bits_instructionIndex_0;
  assign vrfReadDataPorts_19_valid = vrfReadDataPorts_19_valid_0;
  assign vrfReadDataPorts_19_bits_vs = vrfReadDataPorts_19_bits_vs_0;
  assign vrfReadDataPorts_19_bits_instructionIndex = vrfReadDataPorts_19_bits_instructionIndex_0;
  assign vrfReadDataPorts_20_valid = vrfReadDataPorts_20_valid_0;
  assign vrfReadDataPorts_20_bits_vs = vrfReadDataPorts_20_bits_vs_0;
  assign vrfReadDataPorts_20_bits_instructionIndex = vrfReadDataPorts_20_bits_instructionIndex_0;
  assign vrfReadDataPorts_21_valid = vrfReadDataPorts_21_valid_0;
  assign vrfReadDataPorts_21_bits_vs = vrfReadDataPorts_21_bits_vs_0;
  assign vrfReadDataPorts_21_bits_instructionIndex = vrfReadDataPorts_21_bits_instructionIndex_0;
  assign vrfReadDataPorts_22_valid = vrfReadDataPorts_22_valid_0;
  assign vrfReadDataPorts_22_bits_vs = vrfReadDataPorts_22_bits_vs_0;
  assign vrfReadDataPorts_22_bits_instructionIndex = vrfReadDataPorts_22_bits_instructionIndex_0;
  assign vrfReadDataPorts_23_valid = vrfReadDataPorts_23_valid_0;
  assign vrfReadDataPorts_23_bits_vs = vrfReadDataPorts_23_bits_vs_0;
  assign vrfReadDataPorts_23_bits_instructionIndex = vrfReadDataPorts_23_bits_instructionIndex_0;
  assign vrfReadDataPorts_24_valid = vrfReadDataPorts_24_valid_0;
  assign vrfReadDataPorts_24_bits_vs = vrfReadDataPorts_24_bits_vs_0;
  assign vrfReadDataPorts_24_bits_instructionIndex = vrfReadDataPorts_24_bits_instructionIndex_0;
  assign vrfReadDataPorts_25_valid = vrfReadDataPorts_25_valid_0;
  assign vrfReadDataPorts_25_bits_vs = vrfReadDataPorts_25_bits_vs_0;
  assign vrfReadDataPorts_25_bits_instructionIndex = vrfReadDataPorts_25_bits_instructionIndex_0;
  assign vrfReadDataPorts_26_valid = vrfReadDataPorts_26_valid_0;
  assign vrfReadDataPorts_26_bits_vs = vrfReadDataPorts_26_bits_vs_0;
  assign vrfReadDataPorts_26_bits_instructionIndex = vrfReadDataPorts_26_bits_instructionIndex_0;
  assign vrfReadDataPorts_27_valid = vrfReadDataPorts_27_valid_0;
  assign vrfReadDataPorts_27_bits_vs = vrfReadDataPorts_27_bits_vs_0;
  assign vrfReadDataPorts_27_bits_instructionIndex = vrfReadDataPorts_27_bits_instructionIndex_0;
  assign vrfReadDataPorts_28_valid = vrfReadDataPorts_28_valid_0;
  assign vrfReadDataPorts_28_bits_vs = vrfReadDataPorts_28_bits_vs_0;
  assign vrfReadDataPorts_28_bits_instructionIndex = vrfReadDataPorts_28_bits_instructionIndex_0;
  assign vrfReadDataPorts_29_valid = vrfReadDataPorts_29_valid_0;
  assign vrfReadDataPorts_29_bits_vs = vrfReadDataPorts_29_bits_vs_0;
  assign vrfReadDataPorts_29_bits_instructionIndex = vrfReadDataPorts_29_bits_instructionIndex_0;
  assign vrfReadDataPorts_30_valid = vrfReadDataPorts_30_valid_0;
  assign vrfReadDataPorts_30_bits_vs = vrfReadDataPorts_30_bits_vs_0;
  assign vrfReadDataPorts_30_bits_instructionIndex = vrfReadDataPorts_30_bits_instructionIndex_0;
  assign vrfReadDataPorts_31_valid = vrfReadDataPorts_31_valid_0;
  assign vrfReadDataPorts_31_bits_vs = vrfReadDataPorts_31_bits_vs_0;
  assign vrfReadDataPorts_31_bits_instructionIndex = vrfReadDataPorts_31_bits_instructionIndex_0;
endmodule

